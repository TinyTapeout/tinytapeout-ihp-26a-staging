module tt_um_andreasp00 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire miso;
 wire pdm;
 wire \tt6581_inst.accum_en ;
 wire \tt6581_inst.accum_in_mux ;
 wire \tt6581_inst.accum_rst ;
 wire \tt6581_inst.ad_pack[0] ;
 wire \tt6581_inst.ad_pack[10] ;
 wire \tt6581_inst.ad_pack[11] ;
 wire \tt6581_inst.ad_pack[12] ;
 wire \tt6581_inst.ad_pack[13] ;
 wire \tt6581_inst.ad_pack[14] ;
 wire \tt6581_inst.ad_pack[15] ;
 wire \tt6581_inst.ad_pack[16] ;
 wire \tt6581_inst.ad_pack[17] ;
 wire \tt6581_inst.ad_pack[18] ;
 wire \tt6581_inst.ad_pack[19] ;
 wire \tt6581_inst.ad_pack[1] ;
 wire \tt6581_inst.ad_pack[20] ;
 wire \tt6581_inst.ad_pack[21] ;
 wire \tt6581_inst.ad_pack[22] ;
 wire \tt6581_inst.ad_pack[23] ;
 wire \tt6581_inst.ad_pack[2] ;
 wire \tt6581_inst.ad_pack[3] ;
 wire \tt6581_inst.ad_pack[4] ;
 wire \tt6581_inst.ad_pack[5] ;
 wire \tt6581_inst.ad_pack[6] ;
 wire \tt6581_inst.ad_pack[7] ;
 wire \tt6581_inst.ad_pack[8] ;
 wire \tt6581_inst.ad_pack[9] ;
 wire \tt6581_inst.audio_valid ;
 wire \tt6581_inst.bypass_accum[0] ;
 wire \tt6581_inst.bypass_accum[10] ;
 wire \tt6581_inst.bypass_accum[11] ;
 wire \tt6581_inst.bypass_accum[12] ;
 wire \tt6581_inst.bypass_accum[13] ;
 wire \tt6581_inst.bypass_accum[1] ;
 wire \tt6581_inst.bypass_accum[2] ;
 wire \tt6581_inst.bypass_accum[3] ;
 wire \tt6581_inst.bypass_accum[4] ;
 wire \tt6581_inst.bypass_accum[5] ;
 wire \tt6581_inst.bypass_accum[6] ;
 wire \tt6581_inst.bypass_accum[7] ;
 wire \tt6581_inst.bypass_accum[8] ;
 wire \tt6581_inst.bypass_accum[9] ;
 wire \tt6581_inst.control_pack[0] ;
 wire \tt6581_inst.control_pack[10] ;
 wire \tt6581_inst.control_pack[11] ;
 wire \tt6581_inst.control_pack[12] ;
 wire \tt6581_inst.control_pack[13] ;
 wire \tt6581_inst.control_pack[14] ;
 wire \tt6581_inst.control_pack[15] ;
 wire \tt6581_inst.control_pack[16] ;
 wire \tt6581_inst.control_pack[17] ;
 wire \tt6581_inst.control_pack[18] ;
 wire \tt6581_inst.control_pack[19] ;
 wire \tt6581_inst.control_pack[1] ;
 wire \tt6581_inst.control_pack[20] ;
 wire \tt6581_inst.control_pack[21] ;
 wire \tt6581_inst.control_pack[22] ;
 wire \tt6581_inst.control_pack[23] ;
 wire \tt6581_inst.control_pack[2] ;
 wire \tt6581_inst.control_pack[3] ;
 wire \tt6581_inst.control_pack[4] ;
 wire \tt6581_inst.control_pack[5] ;
 wire \tt6581_inst.control_pack[6] ;
 wire \tt6581_inst.control_pack[7] ;
 wire \tt6581_inst.control_pack[8] ;
 wire \tt6581_inst.control_pack[9] ;
 wire \tt6581_inst.controller_inst.cur_state[0] ;
 wire \tt6581_inst.controller_inst.cur_state[10] ;
 wire \tt6581_inst.controller_inst.cur_state[1] ;
 wire \tt6581_inst.controller_inst.cur_state[2] ;
 wire \tt6581_inst.controller_inst.cur_state[3] ;
 wire \tt6581_inst.controller_inst.cur_state[4] ;
 wire \tt6581_inst.controller_inst.cur_state[5] ;
 wire \tt6581_inst.controller_inst.cur_state[6] ;
 wire \tt6581_inst.controller_inst.cur_state[7] ;
 wire \tt6581_inst.controller_inst.cur_state[8] ;
 wire \tt6581_inst.controller_inst.cur_state[9] ;
 wire \tt6581_inst.controller_inst.cur_voice[0] ;
 wire \tt6581_inst.controller_inst.cur_voice[1] ;
 wire \tt6581_inst.controller_inst.env_start_o ;
 wire \tt6581_inst.controller_inst.filt_en_i[0] ;
 wire \tt6581_inst.controller_inst.filt_en_i[1] ;
 wire \tt6581_inst.controller_inst.filt_en_i[2] ;
 wire \tt6581_inst.controller_inst.filt_ready_i ;
 wire \tt6581_inst.controller_inst.filt_start_o ;
 wire \tt6581_inst.controller_inst.freq_hi_i[0] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[10] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[11] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[12] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[13] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[14] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[15] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[16] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[17] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[18] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[19] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[1] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[20] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[21] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[22] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[23] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[2] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[3] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[4] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[5] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[6] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[7] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[8] ;
 wire \tt6581_inst.controller_inst.freq_hi_i[9] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[0] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[10] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[11] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[12] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[13] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[14] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[15] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[16] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[17] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[18] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[19] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[1] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[20] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[21] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[22] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[23] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[2] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[3] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[4] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[5] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[6] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[7] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[8] ;
 wire \tt6581_inst.controller_inst.freq_lo_i[9] ;
 wire \tt6581_inst.controller_inst.mult_in_mux_o[1] ;
 wire \tt6581_inst.controller_inst.mult_in_mux_o[2] ;
 wire \tt6581_inst.controller_inst.mult_start_o ;
 wire \tt6581_inst.controller_inst.pw_hi_i[0] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[10] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[11] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[12] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[13] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[14] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[15] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[16] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[17] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[18] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[19] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[1] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[20] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[21] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[22] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[23] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[2] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[3] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[4] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[5] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[6] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[7] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[8] ;
 wire \tt6581_inst.controller_inst.pw_hi_i[9] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[0] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[10] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[11] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[12] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[13] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[14] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[15] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[16] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[17] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[18] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[19] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[1] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[20] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[21] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[22] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[23] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[2] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[3] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[4] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[5] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[6] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[7] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[8] ;
 wire \tt6581_inst.controller_inst.pw_lo_i[9] ;
 wire \tt6581_inst.controller_inst.sample_tick_i ;
 wire \tt6581_inst.controller_inst.sr_i[0] ;
 wire \tt6581_inst.controller_inst.sr_i[10] ;
 wire \tt6581_inst.controller_inst.sr_i[11] ;
 wire \tt6581_inst.controller_inst.sr_i[12] ;
 wire \tt6581_inst.controller_inst.sr_i[13] ;
 wire \tt6581_inst.controller_inst.sr_i[14] ;
 wire \tt6581_inst.controller_inst.sr_i[15] ;
 wire \tt6581_inst.controller_inst.sr_i[16] ;
 wire \tt6581_inst.controller_inst.sr_i[17] ;
 wire \tt6581_inst.controller_inst.sr_i[18] ;
 wire \tt6581_inst.controller_inst.sr_i[19] ;
 wire \tt6581_inst.controller_inst.sr_i[1] ;
 wire \tt6581_inst.controller_inst.sr_i[20] ;
 wire \tt6581_inst.controller_inst.sr_i[21] ;
 wire \tt6581_inst.controller_inst.sr_i[22] ;
 wire \tt6581_inst.controller_inst.sr_i[23] ;
 wire \tt6581_inst.controller_inst.sr_i[2] ;
 wire \tt6581_inst.controller_inst.sr_i[3] ;
 wire \tt6581_inst.controller_inst.sr_i[4] ;
 wire \tt6581_inst.controller_inst.sr_i[5] ;
 wire \tt6581_inst.controller_inst.sr_i[6] ;
 wire \tt6581_inst.controller_inst.sr_i[7] ;
 wire \tt6581_inst.controller_inst.sr_i[8] ;
 wire \tt6581_inst.controller_inst.sr_i[9] ;
 wire \tt6581_inst.controller_inst.voice_ready_i ;
 wire \tt6581_inst.controller_inst.voice_start_o ;
 wire \tt6581_inst.delta_sigma_inst.audio[10] ;
 wire \tt6581_inst.delta_sigma_inst.audio[11] ;
 wire \tt6581_inst.delta_sigma_inst.audio[12] ;
 wire \tt6581_inst.delta_sigma_inst.audio[13] ;
 wire \tt6581_inst.delta_sigma_inst.audio[14] ;
 wire \tt6581_inst.delta_sigma_inst.audio[15] ;
 wire \tt6581_inst.delta_sigma_inst.audio[16] ;
 wire \tt6581_inst.delta_sigma_inst.audio[17] ;
 wire \tt6581_inst.delta_sigma_inst.audio[4] ;
 wire \tt6581_inst.delta_sigma_inst.audio[5] ;
 wire \tt6581_inst.delta_sigma_inst.audio[6] ;
 wire \tt6581_inst.delta_sigma_inst.audio[7] ;
 wire \tt6581_inst.delta_sigma_inst.audio[8] ;
 wire \tt6581_inst.delta_sigma_inst.audio[9] ;
 wire \tt6581_inst.delta_sigma_inst.cnt[0] ;
 wire \tt6581_inst.delta_sigma_inst.cnt[1] ;
 wire \tt6581_inst.delta_sigma_inst.cnt[2] ;
 wire \tt6581_inst.delta_sigma_inst.e1[0] ;
 wire \tt6581_inst.delta_sigma_inst.e1[10] ;
 wire \tt6581_inst.delta_sigma_inst.e1[11] ;
 wire \tt6581_inst.delta_sigma_inst.e1[12] ;
 wire \tt6581_inst.delta_sigma_inst.e1[13] ;
 wire \tt6581_inst.delta_sigma_inst.e1[14] ;
 wire \tt6581_inst.delta_sigma_inst.e1[15] ;
 wire \tt6581_inst.delta_sigma_inst.e1[16] ;
 wire \tt6581_inst.delta_sigma_inst.e1[17] ;
 wire \tt6581_inst.delta_sigma_inst.e1[18] ;
 wire \tt6581_inst.delta_sigma_inst.e1[1] ;
 wire \tt6581_inst.delta_sigma_inst.e1[2] ;
 wire \tt6581_inst.delta_sigma_inst.e1[3] ;
 wire \tt6581_inst.delta_sigma_inst.e1[4] ;
 wire \tt6581_inst.delta_sigma_inst.e1[5] ;
 wire \tt6581_inst.delta_sigma_inst.e1[6] ;
 wire \tt6581_inst.delta_sigma_inst.e1[7] ;
 wire \tt6581_inst.delta_sigma_inst.e1[8] ;
 wire \tt6581_inst.delta_sigma_inst.e1[9] ;
 wire \tt6581_inst.delta_sigma_inst.e2[0] ;
 wire \tt6581_inst.delta_sigma_inst.e2[10] ;
 wire \tt6581_inst.delta_sigma_inst.e2[11] ;
 wire \tt6581_inst.delta_sigma_inst.e2[12] ;
 wire \tt6581_inst.delta_sigma_inst.e2[13] ;
 wire \tt6581_inst.delta_sigma_inst.e2[14] ;
 wire \tt6581_inst.delta_sigma_inst.e2[15] ;
 wire \tt6581_inst.delta_sigma_inst.e2[16] ;
 wire \tt6581_inst.delta_sigma_inst.e2[17] ;
 wire \tt6581_inst.delta_sigma_inst.e2[18] ;
 wire \tt6581_inst.delta_sigma_inst.e2[1] ;
 wire \tt6581_inst.delta_sigma_inst.e2[2] ;
 wire \tt6581_inst.delta_sigma_inst.e2[3] ;
 wire \tt6581_inst.delta_sigma_inst.e2[4] ;
 wire \tt6581_inst.delta_sigma_inst.e2[5] ;
 wire \tt6581_inst.delta_sigma_inst.e2[6] ;
 wire \tt6581_inst.delta_sigma_inst.e2[7] ;
 wire \tt6581_inst.delta_sigma_inst.e2[8] ;
 wire \tt6581_inst.delta_sigma_inst.e2[9] ;
 wire \tt6581_inst.delta_sigma_inst.en ;
 wire \tt6581_inst.envelope_inst.cur_state[0] ;
 wire \tt6581_inst.envelope_inst.cur_state[1] ;
 wire \tt6581_inst.envelope_inst.nxt_state[0] ;
 wire \tt6581_inst.envelope_inst.nxt_state[1] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][0] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][10] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][11] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][12] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][13] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][14] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][15] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][16] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][17] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][18] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][19] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][1] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][20] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][21] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][22] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][23] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][2] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][3] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][4] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][5] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][6] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][7] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][8] ;
 wire \tt6581_inst.envelope_inst.vol_regs[0][9] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][0] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][10] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][11] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][12] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][13] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][14] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][15] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][16] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][17] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][18] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][19] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][1] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][20] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][21] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][22] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][23] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][2] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][3] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][4] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][5] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][6] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][7] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][8] ;
 wire \tt6581_inst.envelope_inst.vol_regs[1][9] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][0] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][10] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][11] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][12] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][13] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][14] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][15] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][16] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][17] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][18] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][19] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][1] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][20] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][21] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][22] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][23] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][2] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][3] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][4] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][5] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][6] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][7] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][8] ;
 wire \tt6581_inst.envelope_inst.vol_regs[2][9] ;
 wire \tt6581_inst.filt_en_mode[0] ;
 wire \tt6581_inst.filt_en_mode[1] ;
 wire \tt6581_inst.filt_en_mode[2] ;
 wire \tt6581_inst.filt_en_mode[6] ;
 wire \tt6581_inst.filt_en_mode[7] ;
 wire \tt6581_inst.filt_f_hi[0] ;
 wire \tt6581_inst.filt_f_hi[1] ;
 wire \tt6581_inst.filt_f_hi[2] ;
 wire \tt6581_inst.filt_f_hi[3] ;
 wire \tt6581_inst.filt_f_hi[4] ;
 wire \tt6581_inst.filt_f_hi[5] ;
 wire \tt6581_inst.filt_f_hi[6] ;
 wire \tt6581_inst.filt_f_hi[7] ;
 wire \tt6581_inst.filt_f_lo[0] ;
 wire \tt6581_inst.filt_f_lo[1] ;
 wire \tt6581_inst.filt_f_lo[2] ;
 wire \tt6581_inst.filt_f_lo[3] ;
 wire \tt6581_inst.filt_f_lo[4] ;
 wire \tt6581_inst.filt_f_lo[5] ;
 wire \tt6581_inst.filt_f_lo[6] ;
 wire \tt6581_inst.filt_f_lo[7] ;
 wire \tt6581_inst.filt_q_hi[0] ;
 wire \tt6581_inst.filt_q_hi[1] ;
 wire \tt6581_inst.filt_q_hi[2] ;
 wire \tt6581_inst.filt_q_hi[3] ;
 wire \tt6581_inst.filt_q_hi[4] ;
 wire \tt6581_inst.filt_q_hi[5] ;
 wire \tt6581_inst.filt_q_hi[6] ;
 wire \tt6581_inst.filt_q_hi[7] ;
 wire \tt6581_inst.filt_q_lo[0] ;
 wire \tt6581_inst.filt_q_lo[1] ;
 wire \tt6581_inst.filt_q_lo[2] ;
 wire \tt6581_inst.filt_q_lo[3] ;
 wire \tt6581_inst.filt_q_lo[4] ;
 wire \tt6581_inst.filt_q_lo[5] ;
 wire \tt6581_inst.filt_q_lo[6] ;
 wire \tt6581_inst.filt_q_lo[7] ;
 wire \tt6581_inst.filt_volume[0] ;
 wire \tt6581_inst.filt_volume[1] ;
 wire \tt6581_inst.filt_volume[2] ;
 wire \tt6581_inst.filt_volume[3] ;
 wire \tt6581_inst.filt_volume[4] ;
 wire \tt6581_inst.filt_volume[5] ;
 wire \tt6581_inst.filt_volume[6] ;
 wire \tt6581_inst.filt_volume[7] ;
 wire \tt6581_inst.filter_accum[0] ;
 wire \tt6581_inst.filter_accum[10] ;
 wire \tt6581_inst.filter_accum[11] ;
 wire \tt6581_inst.filter_accum[12] ;
 wire \tt6581_inst.filter_accum[13] ;
 wire \tt6581_inst.filter_accum[1] ;
 wire \tt6581_inst.filter_accum[2] ;
 wire \tt6581_inst.filter_accum[3] ;
 wire \tt6581_inst.filter_accum[4] ;
 wire \tt6581_inst.filter_accum[5] ;
 wire \tt6581_inst.filter_accum[6] ;
 wire \tt6581_inst.filter_accum[7] ;
 wire \tt6581_inst.filter_accum[8] ;
 wire \tt6581_inst.filter_accum[9] ;
 wire \tt6581_inst.mult_inst.a_reg[0] ;
 wire \tt6581_inst.mult_inst.a_reg[10] ;
 wire \tt6581_inst.mult_inst.a_reg[11] ;
 wire \tt6581_inst.mult_inst.a_reg[12] ;
 wire \tt6581_inst.mult_inst.a_reg[13] ;
 wire \tt6581_inst.mult_inst.a_reg[14] ;
 wire \tt6581_inst.mult_inst.a_reg[15] ;
 wire \tt6581_inst.mult_inst.a_reg[16] ;
 wire \tt6581_inst.mult_inst.a_reg[17] ;
 wire \tt6581_inst.mult_inst.a_reg[18] ;
 wire \tt6581_inst.mult_inst.a_reg[19] ;
 wire \tt6581_inst.mult_inst.a_reg[1] ;
 wire \tt6581_inst.mult_inst.a_reg[20] ;
 wire \tt6581_inst.mult_inst.a_reg[21] ;
 wire \tt6581_inst.mult_inst.a_reg[22] ;
 wire \tt6581_inst.mult_inst.a_reg[23] ;
 wire \tt6581_inst.mult_inst.a_reg[24] ;
 wire \tt6581_inst.mult_inst.a_reg[25] ;
 wire \tt6581_inst.mult_inst.a_reg[26] ;
 wire \tt6581_inst.mult_inst.a_reg[27] ;
 wire \tt6581_inst.mult_inst.a_reg[28] ;
 wire \tt6581_inst.mult_inst.a_reg[29] ;
 wire \tt6581_inst.mult_inst.a_reg[2] ;
 wire \tt6581_inst.mult_inst.a_reg[30] ;
 wire \tt6581_inst.mult_inst.a_reg[31] ;
 wire \tt6581_inst.mult_inst.a_reg[32] ;
 wire \tt6581_inst.mult_inst.a_reg[33] ;
 wire \tt6581_inst.mult_inst.a_reg[34] ;
 wire \tt6581_inst.mult_inst.a_reg[35] ;
 wire \tt6581_inst.mult_inst.a_reg[36] ;
 wire \tt6581_inst.mult_inst.a_reg[37] ;
 wire \tt6581_inst.mult_inst.a_reg[38] ;
 wire \tt6581_inst.mult_inst.a_reg[3] ;
 wire \tt6581_inst.mult_inst.a_reg[4] ;
 wire \tt6581_inst.mult_inst.a_reg[5] ;
 wire \tt6581_inst.mult_inst.a_reg[6] ;
 wire \tt6581_inst.mult_inst.a_reg[7] ;
 wire \tt6581_inst.mult_inst.a_reg[8] ;
 wire \tt6581_inst.mult_inst.a_reg[9] ;
 wire \tt6581_inst.mult_inst.accum[0] ;
 wire \tt6581_inst.mult_inst.accum[10] ;
 wire \tt6581_inst.mult_inst.accum[11] ;
 wire \tt6581_inst.mult_inst.accum[12] ;
 wire \tt6581_inst.mult_inst.accum[13] ;
 wire \tt6581_inst.mult_inst.accum[14] ;
 wire \tt6581_inst.mult_inst.accum[15] ;
 wire \tt6581_inst.mult_inst.accum[16] ;
 wire \tt6581_inst.mult_inst.accum[17] ;
 wire \tt6581_inst.mult_inst.accum[18] ;
 wire \tt6581_inst.mult_inst.accum[19] ;
 wire \tt6581_inst.mult_inst.accum[1] ;
 wire \tt6581_inst.mult_inst.accum[20] ;
 wire \tt6581_inst.mult_inst.accum[21] ;
 wire \tt6581_inst.mult_inst.accum[22] ;
 wire \tt6581_inst.mult_inst.accum[23] ;
 wire \tt6581_inst.mult_inst.accum[24] ;
 wire \tt6581_inst.mult_inst.accum[25] ;
 wire \tt6581_inst.mult_inst.accum[26] ;
 wire \tt6581_inst.mult_inst.accum[27] ;
 wire \tt6581_inst.mult_inst.accum[28] ;
 wire \tt6581_inst.mult_inst.accum[29] ;
 wire \tt6581_inst.mult_inst.accum[2] ;
 wire \tt6581_inst.mult_inst.accum[30] ;
 wire \tt6581_inst.mult_inst.accum[31] ;
 wire \tt6581_inst.mult_inst.accum[32] ;
 wire \tt6581_inst.mult_inst.accum[33] ;
 wire \tt6581_inst.mult_inst.accum[34] ;
 wire \tt6581_inst.mult_inst.accum[35] ;
 wire \tt6581_inst.mult_inst.accum[36] ;
 wire \tt6581_inst.mult_inst.accum[37] ;
 wire \tt6581_inst.mult_inst.accum[38] ;
 wire \tt6581_inst.mult_inst.accum[3] ;
 wire \tt6581_inst.mult_inst.accum[4] ;
 wire \tt6581_inst.mult_inst.accum[5] ;
 wire \tt6581_inst.mult_inst.accum[6] ;
 wire \tt6581_inst.mult_inst.accum[7] ;
 wire \tt6581_inst.mult_inst.accum[8] ;
 wire \tt6581_inst.mult_inst.accum[9] ;
 wire \tt6581_inst.mult_inst.b_reg[0] ;
 wire \tt6581_inst.mult_inst.b_reg[10] ;
 wire \tt6581_inst.mult_inst.b_reg[11] ;
 wire \tt6581_inst.mult_inst.b_reg[12] ;
 wire \tt6581_inst.mult_inst.b_reg[13] ;
 wire \tt6581_inst.mult_inst.b_reg[14] ;
 wire \tt6581_inst.mult_inst.b_reg[15] ;
 wire \tt6581_inst.mult_inst.b_reg[1] ;
 wire \tt6581_inst.mult_inst.b_reg[2] ;
 wire \tt6581_inst.mult_inst.b_reg[3] ;
 wire \tt6581_inst.mult_inst.b_reg[4] ;
 wire \tt6581_inst.mult_inst.b_reg[5] ;
 wire \tt6581_inst.mult_inst.b_reg[6] ;
 wire \tt6581_inst.mult_inst.b_reg[7] ;
 wire \tt6581_inst.mult_inst.b_reg[8] ;
 wire \tt6581_inst.mult_inst.b_reg[9] ;
 wire \tt6581_inst.mult_inst.cur_state ;
 wire \tt6581_inst.mult_inst.iter[0] ;
 wire \tt6581_inst.mult_inst.iter[1] ;
 wire \tt6581_inst.mult_inst.iter[2] ;
 wire \tt6581_inst.mult_inst.iter[3] ;
 wire \tt6581_inst.mult_inst.iter[4] ;
 wire \tt6581_inst.mult_inst.neg_result ;
 wire \tt6581_inst.mult_inst.nxt_state ;
 wire \tt6581_inst.multi_voice_inst.cur_state[0] ;
 wire \tt6581_inst.multi_voice_inst.cur_state[1] ;
 wire \tt6581_inst.multi_voice_inst.nxt_state[0] ;
 wire \tt6581_inst.multi_voice_inst.nxt_state[1] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[0][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[0][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[1][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[1][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[2][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_last_msb[2][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][10] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][11] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][12] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][13] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][14] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][15] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][16] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][17] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][2] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][3] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][4] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][5] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][6] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][7] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][8] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[0][9] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][10] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][11] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][12] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][13] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][14] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][15] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][16] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][17] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][2] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][3] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][4] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][5] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][6] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][7] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][8] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[1][9] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][0] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][10] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][11] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][12] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][13] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][14] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][15] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][16] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][17] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][1] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][2] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][3] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][4] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][5] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][6] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][7] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][8] ;
 wire \tt6581_inst.multi_voice_inst.phase_regs[2][9] ;
 wire \tt6581_inst.reg_addr[0] ;
 wire \tt6581_inst.reg_addr[1] ;
 wire \tt6581_inst.reg_addr[2] ;
 wire \tt6581_inst.reg_addr[3] ;
 wire \tt6581_inst.reg_addr[4] ;
 wire \tt6581_inst.reg_addr[5] ;
 wire \tt6581_inst.reg_addr[6] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[0] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[1] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[2] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[3] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[4] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[5] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[6] ;
 wire \tt6581_inst.reg_file_inst.wdata_i[7] ;
 wire \tt6581_inst.reg_file_inst.we_i ;
 wire \tt6581_inst.spi_inst.bit_cnt[0] ;
 wire \tt6581_inst.spi_inst.bit_cnt[1] ;
 wire \tt6581_inst.spi_inst.bit_cnt[2] ;
 wire \tt6581_inst.spi_inst.bit_cnt[3] ;
 wire \tt6581_inst.spi_inst.cs_sync[0] ;
 wire \tt6581_inst.spi_inst.cs_sync[1] ;
 wire \tt6581_inst.spi_inst.data_out_reg[0] ;
 wire \tt6581_inst.spi_inst.data_out_reg[1] ;
 wire \tt6581_inst.spi_inst.data_out_reg[2] ;
 wire \tt6581_inst.spi_inst.data_out_reg[3] ;
 wire \tt6581_inst.spi_inst.data_out_reg[4] ;
 wire \tt6581_inst.spi_inst.data_out_reg[5] ;
 wire \tt6581_inst.spi_inst.data_out_reg[6] ;
 wire \tt6581_inst.spi_inst.data_out_reg[7] ;
 wire \tt6581_inst.spi_inst.is_write_cmd ;
 wire \tt6581_inst.spi_inst.mosi_sync[0] ;
 wire \tt6581_inst.spi_inst.mosi_sync[1] ;
 wire \tt6581_inst.spi_inst.sclk_sync[0] ;
 wire \tt6581_inst.spi_inst.sclk_sync[1] ;
 wire \tt6581_inst.spi_inst.sclk_sync[2] ;
 wire \tt6581_inst.spi_inst.shift_reg[0] ;
 wire \tt6581_inst.spi_inst.shift_reg[1] ;
 wire \tt6581_inst.spi_inst.shift_reg[2] ;
 wire \tt6581_inst.spi_inst.shift_reg[3] ;
 wire \tt6581_inst.spi_inst.shift_reg[4] ;
 wire \tt6581_inst.spi_inst.shift_reg[5] ;
 wire \tt6581_inst.spi_inst.shift_reg[6] ;
 wire \tt6581_inst.svf_inst.cur_state[10] ;
 wire \tt6581_inst.svf_inst.cur_state[1] ;
 wire \tt6581_inst.svf_inst.cur_state[2] ;
 wire \tt6581_inst.svf_inst.cur_state[3] ;
 wire \tt6581_inst.svf_inst.cur_state[5] ;
 wire \tt6581_inst.svf_inst.cur_state[6] ;
 wire \tt6581_inst.svf_inst.cur_state[7] ;
 wire \tt6581_inst.svf_inst.cur_state[8] ;
 wire \tt6581_inst.svf_inst.cur_state[9] ;
 wire \tt6581_inst.svf_inst.hp_node[0] ;
 wire \tt6581_inst.svf_inst.hp_node[10] ;
 wire \tt6581_inst.svf_inst.hp_node[11] ;
 wire \tt6581_inst.svf_inst.hp_node[12] ;
 wire \tt6581_inst.svf_inst.hp_node[13] ;
 wire \tt6581_inst.svf_inst.hp_node[14] ;
 wire \tt6581_inst.svf_inst.hp_node[15] ;
 wire \tt6581_inst.svf_inst.hp_node[16] ;
 wire \tt6581_inst.svf_inst.hp_node[17] ;
 wire \tt6581_inst.svf_inst.hp_node[18] ;
 wire \tt6581_inst.svf_inst.hp_node[19] ;
 wire \tt6581_inst.svf_inst.hp_node[1] ;
 wire \tt6581_inst.svf_inst.hp_node[20] ;
 wire \tt6581_inst.svf_inst.hp_node[21] ;
 wire \tt6581_inst.svf_inst.hp_node[22] ;
 wire \tt6581_inst.svf_inst.hp_node[23] ;
 wire \tt6581_inst.svf_inst.hp_node[2] ;
 wire \tt6581_inst.svf_inst.hp_node[3] ;
 wire \tt6581_inst.svf_inst.hp_node[4] ;
 wire \tt6581_inst.svf_inst.hp_node[5] ;
 wire \tt6581_inst.svf_inst.hp_node[6] ;
 wire \tt6581_inst.svf_inst.hp_node[7] ;
 wire \tt6581_inst.svf_inst.hp_node[8] ;
 wire \tt6581_inst.svf_inst.hp_node[9] ;
 wire \tt6581_inst.svf_inst.reg_band[0] ;
 wire \tt6581_inst.svf_inst.reg_band[10] ;
 wire \tt6581_inst.svf_inst.reg_band[11] ;
 wire \tt6581_inst.svf_inst.reg_band[12] ;
 wire \tt6581_inst.svf_inst.reg_band[13] ;
 wire \tt6581_inst.svf_inst.reg_band[14] ;
 wire \tt6581_inst.svf_inst.reg_band[15] ;
 wire \tt6581_inst.svf_inst.reg_band[16] ;
 wire \tt6581_inst.svf_inst.reg_band[17] ;
 wire \tt6581_inst.svf_inst.reg_band[18] ;
 wire \tt6581_inst.svf_inst.reg_band[19] ;
 wire \tt6581_inst.svf_inst.reg_band[1] ;
 wire \tt6581_inst.svf_inst.reg_band[20] ;
 wire \tt6581_inst.svf_inst.reg_band[21] ;
 wire \tt6581_inst.svf_inst.reg_band[22] ;
 wire \tt6581_inst.svf_inst.reg_band[23] ;
 wire \tt6581_inst.svf_inst.reg_band[2] ;
 wire \tt6581_inst.svf_inst.reg_band[3] ;
 wire \tt6581_inst.svf_inst.reg_band[4] ;
 wire \tt6581_inst.svf_inst.reg_band[5] ;
 wire \tt6581_inst.svf_inst.reg_band[6] ;
 wire \tt6581_inst.svf_inst.reg_band[7] ;
 wire \tt6581_inst.svf_inst.reg_band[8] ;
 wire \tt6581_inst.svf_inst.reg_band[9] ;
 wire \tt6581_inst.svf_inst.reg_low[0] ;
 wire \tt6581_inst.svf_inst.reg_low[10] ;
 wire \tt6581_inst.svf_inst.reg_low[11] ;
 wire \tt6581_inst.svf_inst.reg_low[12] ;
 wire \tt6581_inst.svf_inst.reg_low[13] ;
 wire \tt6581_inst.svf_inst.reg_low[14] ;
 wire \tt6581_inst.svf_inst.reg_low[15] ;
 wire \tt6581_inst.svf_inst.reg_low[16] ;
 wire \tt6581_inst.svf_inst.reg_low[17] ;
 wire \tt6581_inst.svf_inst.reg_low[18] ;
 wire \tt6581_inst.svf_inst.reg_low[19] ;
 wire \tt6581_inst.svf_inst.reg_low[1] ;
 wire \tt6581_inst.svf_inst.reg_low[20] ;
 wire \tt6581_inst.svf_inst.reg_low[21] ;
 wire \tt6581_inst.svf_inst.reg_low[22] ;
 wire \tt6581_inst.svf_inst.reg_low[23] ;
 wire \tt6581_inst.svf_inst.reg_low[2] ;
 wire \tt6581_inst.svf_inst.reg_low[3] ;
 wire \tt6581_inst.svf_inst.reg_low[4] ;
 wire \tt6581_inst.svf_inst.reg_low[5] ;
 wire \tt6581_inst.svf_inst.reg_low[6] ;
 wire \tt6581_inst.svf_inst.reg_low[7] ;
 wire \tt6581_inst.svf_inst.reg_low[8] ;
 wire \tt6581_inst.svf_inst.reg_low[9] ;
 wire \tt6581_inst.tick_gen_inst.cnt[0] ;
 wire \tt6581_inst.tick_gen_inst.cnt[1] ;
 wire \tt6581_inst.tick_gen_inst.cnt[2] ;
 wire \tt6581_inst.tick_gen_inst.cnt[3] ;
 wire \tt6581_inst.tick_gen_inst.cnt[4] ;
 wire \tt6581_inst.tick_gen_inst.cnt[5] ;
 wire \tt6581_inst.tick_gen_inst.cnt[6] ;
 wire \tt6581_inst.tick_gen_inst.cnt[7] ;
 wire \tt6581_inst.tick_gen_inst.cnt[8] ;
 wire \tt6581_inst.tick_gen_inst.cnt[9] ;
 wire net5;
 wire net6;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;

 sg13g2_inv_1 _4451_ (.Y(_0831_),
    .A(net198));
 sg13g2_inv_1 _4452_ (.Y(_0832_),
    .A(net181));
 sg13g2_inv_1 _4453_ (.Y(_0833_),
    .A(net172));
 sg13g2_inv_1 _4454_ (.Y(_0834_),
    .A(net254));
 sg13g2_inv_1 _4455_ (.Y(_0835_),
    .A(net200));
 sg13g2_inv_1 _4456_ (.Y(_0836_),
    .A(net241));
 sg13g2_inv_1 _4457_ (.Y(_0837_),
    .A(net203));
 sg13g2_inv_1 _4458_ (.Y(_0838_),
    .A(_0042_));
 sg13g2_inv_1 _4459_ (.Y(_0839_),
    .A(\tt6581_inst.envelope_inst.vol_regs[0][17] ));
 sg13g2_inv_1 _4460_ (.Y(_0840_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][17] ));
 sg13g2_inv_1 _4461_ (.Y(_0841_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][18] ));
 sg13g2_inv_1 _4462_ (.Y(_0842_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][18] ));
 sg13g2_inv_1 _4463_ (.Y(_0843_),
    .A(\tt6581_inst.envelope_inst.vol_regs[0][23] ));
 sg13g2_inv_1 _4464_ (.Y(_0844_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][23] ));
 sg13g2_inv_1 _4465_ (.Y(_0845_),
    .A(\tt6581_inst.envelope_inst.vol_regs[0][22] ));
 sg13g2_inv_1 _4466_ (.Y(_0846_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][22] ));
 sg13g2_inv_1 _4467_ (.Y(_0847_),
    .A(\tt6581_inst.envelope_inst.vol_regs[0][21] ));
 sg13g2_inv_1 _4468_ (.Y(_0848_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][21] ));
 sg13g2_inv_1 _4469_ (.Y(_0849_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][20] ));
 sg13g2_inv_1 _4470_ (.Y(_0850_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][20] ));
 sg13g2_inv_1 _4471_ (.Y(_0851_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][1] ));
 sg13g2_inv_1 _4472_ (.Y(_0852_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][1] ));
 sg13g2_inv_1 _4473_ (.Y(_0853_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][5] ));
 sg13g2_inv_1 _4474_ (.Y(_0854_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][5] ));
 sg13g2_inv_1 _4475_ (.Y(_0855_),
    .A(net223));
 sg13g2_inv_1 _4476_ (.Y(_0856_),
    .A(net249));
 sg13g2_inv_1 _4477_ (.Y(_0857_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][7] ));
 sg13g2_inv_1 _4478_ (.Y(_0858_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][7] ));
 sg13g2_inv_1 _4479_ (.Y(_0859_),
    .A(net233));
 sg13g2_inv_1 _4480_ (.Y(_0860_),
    .A(net258));
 sg13g2_inv_1 _4481_ (.Y(_0861_),
    .A(net154));
 sg13g2_inv_1 _4482_ (.Y(_0862_),
    .A(net184));
 sg13g2_inv_1 _4483_ (.Y(_0863_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][8] ));
 sg13g2_inv_1 _4484_ (.Y(_0864_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][8] ));
 sg13g2_inv_1 _4485_ (.Y(_0865_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][11] ));
 sg13g2_inv_1 _4486_ (.Y(_0866_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][11] ));
 sg13g2_inv_1 _4487_ (.Y(_0867_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][10] ));
 sg13g2_inv_1 _4488_ (.Y(_0868_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][10] ));
 sg13g2_inv_1 _4489_ (.Y(_0869_),
    .A(net264));
 sg13g2_inv_1 _4490_ (.Y(_0870_),
    .A(net193));
 sg13g2_inv_1 _4491_ (.Y(_0871_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][15] ));
 sg13g2_inv_1 _4492_ (.Y(_0872_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][15] ));
 sg13g2_inv_1 _4493_ (.Y(_0873_),
    .A(\tt6581_inst.envelope_inst.vol_regs[2][14] ));
 sg13g2_inv_1 _4494_ (.Y(_0874_),
    .A(\tt6581_inst.envelope_inst.vol_regs[1][14] ));
 sg13g2_inv_1 _4495_ (.Y(_0875_),
    .A(net777));
 sg13g2_inv_2 _4496_ (.Y(_0876_),
    .A(net488));
 sg13g2_inv_2 _4497_ (.Y(_0877_),
    .A(net823));
 sg13g2_inv_1 _4498_ (.Y(_0878_),
    .A(net989));
 sg13g2_inv_2 _4499_ (.Y(_0879_),
    .A(\tt6581_inst.reg_addr[4] ));
 sg13g2_inv_1 _4500_ (.Y(_0880_),
    .A(\tt6581_inst.mult_inst.iter[3] ));
 sg13g2_inv_1 _4501_ (.Y(_0881_),
    .A(net77));
 sg13g2_inv_1 _4502_ (.Y(_0882_),
    .A(net514));
 sg13g2_inv_1 _4503_ (.Y(_0883_),
    .A(\tt6581_inst.delta_sigma_inst.e2[17] ));
 sg13g2_inv_1 _4504_ (.Y(_0884_),
    .A(\tt6581_inst.controller_inst.voice_ready_i ));
 sg13g2_inv_1 _4505_ (.Y(_0885_),
    .A(\tt6581_inst.controller_inst.sample_tick_i ));
 sg13g2_inv_2 _4506_ (.Y(_0886_),
    .A(net34));
 sg13g2_inv_1 _4507_ (.Y(_0887_),
    .A(net42));
 sg13g2_inv_4 _4508_ (.A(net1538),
    .Y(_0888_));
 sg13g2_inv_1 _4509_ (.Y(_0025_),
    .A(net46));
 sg13g2_inv_1 _4510_ (.Y(_0889_),
    .A(net67));
 sg13g2_inv_1 _4511_ (.Y(_0890_),
    .A(net454));
 sg13g2_inv_1 _4512_ (.Y(_0891_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][9] ));
 sg13g2_inv_1 _4513_ (.Y(_0892_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][9] ));
 sg13g2_inv_1 _4514_ (.Y(_0893_),
    .A(net493));
 sg13g2_inv_1 _4515_ (.Y(_0894_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][8] ));
 sg13g2_inv_1 _4516_ (.Y(_0895_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][8] ));
 sg13g2_inv_1 _4517_ (.Y(_0896_),
    .A(net718));
 sg13g2_inv_1 _4518_ (.Y(_0897_),
    .A(net521));
 sg13g2_inv_1 _4519_ (.Y(_0898_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][6] ));
 sg13g2_inv_1 _4520_ (.Y(_0899_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][6] ));
 sg13g2_inv_1 _4521_ (.Y(_0900_),
    .A(net669));
 sg13g2_inv_1 _4522_ (.Y(_0901_),
    .A(net527));
 sg13g2_inv_1 _4523_ (.Y(_0902_),
    .A(net1017));
 sg13g2_inv_1 _4524_ (.Y(_0903_),
    .A(net546));
 sg13g2_inv_1 _4525_ (.Y(_0904_),
    .A(net563));
 sg13g2_inv_1 _4526_ (.Y(_0905_),
    .A(net242));
 sg13g2_inv_1 _4527_ (.Y(_0906_),
    .A(net175));
 sg13g2_inv_1 _4528_ (.Y(_0907_),
    .A(net262));
 sg13g2_inv_1 _4529_ (.Y(_0908_),
    .A(\tt6581_inst.mult_inst.accum[8] ));
 sg13g2_inv_8 _4530_ (.Y(_0909_),
    .A(net1500));
 sg13g2_inv_2 _4531_ (.Y(_0910_),
    .A(net1705));
 sg13g2_inv_1 _4532_ (.Y(_0911_),
    .A(net1536));
 sg13g2_inv_1 _4533_ (.Y(_0912_),
    .A(\tt6581_inst.mult_inst.accum[12] ));
 sg13g2_inv_1 _4534_ (.Y(_0913_),
    .A(\tt6581_inst.mult_inst.accum[14] ));
 sg13g2_inv_1 _4535_ (.Y(_0914_),
    .A(\tt6581_inst.mult_inst.accum[15] ));
 sg13g2_inv_1 _4536_ (.Y(_0915_),
    .A(\tt6581_inst.mult_inst.accum[16] ));
 sg13g2_inv_4 _4537_ (.A(net1492),
    .Y(_0916_));
 sg13g2_inv_1 _4538_ (.Y(_0917_),
    .A(net1491));
 sg13g2_inv_1 _4539_ (.Y(_0918_),
    .A(\tt6581_inst.svf_inst.reg_low[23] ));
 sg13g2_inv_1 _4540_ (.Y(_0919_),
    .A(net1053));
 sg13g2_inv_4 _4541_ (.A(net1081),
    .Y(_0920_));
 sg13g2_inv_1 _4542_ (.Y(_0921_),
    .A(net802));
 sg13g2_inv_2 _4543_ (.Y(_0922_),
    .A(\tt6581_inst.svf_inst.reg_low[21] ));
 sg13g2_inv_2 _4544_ (.Y(_0923_),
    .A(net1113));
 sg13g2_inv_2 _4545_ (.Y(_0924_),
    .A(\tt6581_inst.svf_inst.reg_low[19] ));
 sg13g2_inv_2 _4546_ (.Y(_0925_),
    .A(\tt6581_inst.svf_inst.reg_low[18] ));
 sg13g2_inv_1 _4547_ (.Y(_0926_),
    .A(\tt6581_inst.svf_inst.hp_node[17] ));
 sg13g2_inv_2 _4548_ (.Y(_0927_),
    .A(\tt6581_inst.svf_inst.reg_low[17] ));
 sg13g2_inv_2 _4549_ (.Y(_0928_),
    .A(\tt6581_inst.svf_inst.reg_low[16] ));
 sg13g2_inv_1 _4550_ (.Y(_0929_),
    .A(net1094));
 sg13g2_inv_2 _4551_ (.Y(_0930_),
    .A(\tt6581_inst.svf_inst.reg_low[15] ));
 sg13g2_inv_1 _4552_ (.Y(_0931_),
    .A(net516));
 sg13g2_inv_1 _4553_ (.Y(_0932_),
    .A(net1132));
 sg13g2_inv_1 _4554_ (.Y(_0933_),
    .A(net892));
 sg13g2_inv_2 _4555_ (.Y(_0934_),
    .A(net1116));
 sg13g2_inv_1 _4556_ (.Y(_0935_),
    .A(net1002));
 sg13g2_inv_1 _4557_ (.Y(_0936_),
    .A(\tt6581_inst.svf_inst.reg_low[11] ));
 sg13g2_inv_2 _4558_ (.Y(_0937_),
    .A(net1118));
 sg13g2_inv_2 _4559_ (.Y(_0938_),
    .A(net1128));
 sg13g2_inv_2 _4560_ (.Y(_0939_),
    .A(net1115));
 sg13g2_inv_2 _4561_ (.Y(_0940_),
    .A(net1698));
 sg13g2_inv_1 _4562_ (.Y(_0941_),
    .A(\tt6581_inst.svf_inst.reg_low[4] ));
 sg13g2_inv_1 _4563_ (.Y(_0942_),
    .A(\tt6581_inst.svf_inst.reg_low[2] ));
 sg13g2_inv_1 _4564_ (.Y(_0943_),
    .A(net1508));
 sg13g2_inv_1 _4565_ (.Y(_0944_),
    .A(\tt6581_inst.svf_inst.reg_band[21] ));
 sg13g2_inv_1 _4566_ (.Y(_0945_),
    .A(net1049));
 sg13g2_inv_1 _4567_ (.Y(_0946_),
    .A(net818));
 sg13g2_inv_1 _4568_ (.Y(_0947_),
    .A(net880));
 sg13g2_inv_1 _4569_ (.Y(_0948_),
    .A(net430));
 sg13g2_inv_1 _4570_ (.Y(_0949_),
    .A(net337));
 sg13g2_inv_1 _4571_ (.Y(_0950_),
    .A(\tt6581_inst.bypass_accum[0] ));
 sg13g2_inv_1 _4572_ (.Y(_0951_),
    .A(net539));
 sg13g2_inv_1 _4573_ (.Y(_0952_),
    .A(net439));
 sg13g2_inv_1 _4574_ (.Y(_0953_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][13] ));
 sg13g2_inv_1 _4575_ (.Y(_0954_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][13] ));
 sg13g2_inv_1 _4576_ (.Y(_0955_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][12] ));
 sg13g2_inv_1 _4577_ (.Y(_0956_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][12] ));
 sg13g2_inv_1 _4578_ (.Y(_0957_),
    .A(net447));
 sg13g2_inv_1 _4579_ (.Y(_0958_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[0][11] ));
 sg13g2_inv_1 _4580_ (.Y(_0959_),
    .A(\tt6581_inst.multi_voice_inst.phase_regs[1][11] ));
 sg13g2_inv_1 _4581_ (.Y(_0960_),
    .A(net394));
 sg13g2_inv_1 _4582_ (.Y(_0961_),
    .A(net166));
 sg13g2_inv_1 _4583_ (.Y(_0962_),
    .A(net161));
 sg13g2_inv_1 _4584_ (.Y(_0963_),
    .A(net234));
 sg13g2_inv_1 _4585_ (.Y(_0964_),
    .A(net269));
 sg13g2_inv_1 _4586_ (.Y(_0965_),
    .A(net600));
 sg13g2_inv_1 _4587_ (.Y(_0966_),
    .A(net366));
 sg13g2_inv_1 _4588_ (.Y(_0967_),
    .A(net512));
 sg13g2_inv_1 _4589_ (.Y(_0968_),
    .A(net548));
 sg13g2_inv_1 _4590_ (.Y(_0969_),
    .A(net614));
 sg13g2_inv_1 _4591_ (.Y(_0970_),
    .A(net167));
 sg13g2_inv_1 _4592_ (.Y(_0971_),
    .A(net230));
 sg13g2_inv_1 _4593_ (.Y(_0972_),
    .A(net460));
 sg13g2_inv_2 _4594_ (.Y(_0973_),
    .A(net631));
 sg13g2_inv_1 _4595_ (.Y(_0974_),
    .A(net571));
 sg13g2_inv_1 _4596_ (.Y(_0975_),
    .A(net1072));
 sg13g2_inv_1 _4597_ (.Y(_0976_),
    .A(net1068));
 sg13g2_inv_1 _4598_ (.Y(_0977_),
    .A(net1026));
 sg13g2_inv_1 _4599_ (.Y(_0978_),
    .A(net972));
 sg13g2_inv_1 _4600_ (.Y(_0979_),
    .A(net803));
 sg13g2_inv_1 _4601_ (.Y(_0980_),
    .A(net871));
 sg13g2_inv_1 _4602_ (.Y(_0981_),
    .A(net553));
 sg13g2_inv_1 _4603_ (.Y(_0982_),
    .A(net529));
 sg13g2_inv_1 _4604_ (.Y(_0983_),
    .A(net674));
 sg13g2_inv_1 _4605_ (.Y(_0984_),
    .A(net579));
 sg13g2_inv_1 _4606_ (.Y(_0985_),
    .A(net963));
 sg13g2_inv_1 _4607_ (.Y(_0986_),
    .A(net1015));
 sg13g2_inv_1 _4608_ (.Y(_0987_),
    .A(\tt6581_inst.mult_inst.accum[29] ));
 sg13g2_inv_1 _4609_ (.Y(_0988_),
    .A(\tt6581_inst.mult_inst.accum[31] ));
 sg13g2_inv_1 _4610_ (.Y(_0989_),
    .A(net290));
 sg13g2_inv_2 _4611_ (.Y(_0990_),
    .A(net955));
 sg13g2_inv_1 _4612_ (.Y(_0991_),
    .A(net1054));
 sg13g2_inv_1 _4613_ (.Y(_0992_),
    .A(net1120));
 sg13g2_inv_2 _4614_ (.Y(_0993_),
    .A(net1108));
 sg13g2_inv_2 _4615_ (.Y(_0994_),
    .A(net1019));
 sg13g2_inv_8 _4616_ (.Y(_0995_),
    .A(net1130));
 sg13g2_inv_1 _4617_ (.Y(_0996_),
    .A(net40));
 sg13g2_inv_4 _4618_ (.A(net1513),
    .Y(_0997_));
 sg13g2_inv_2 _4619_ (.Y(\tt6581_inst.controller_inst.cur_state[0] ),
    .A(net36));
 sg13g2_inv_2 _4620_ (.Y(_0998_),
    .A(net1550));
 sg13g2_inv_1 _4621_ (.Y(_0999_),
    .A(net187));
 sg13g2_inv_2 _4622_ (.Y(_1000_),
    .A(net1516));
 sg13g2_inv_2 _4623_ (.Y(_1001_),
    .A(net1527));
 sg13g2_inv_1 _4624_ (.Y(_1002_),
    .A(net1494));
 sg13g2_or2_1 _4625_ (.X(_0014_),
    .B(net33),
    .A(net60));
 sg13g2_or2_1 _4626_ (.X(_0015_),
    .B(net32),
    .A(net64));
 sg13g2_or2_1 _4627_ (.X(_0116_),
    .B(_0015_),
    .A(_0014_));
 sg13g2_nor2_1 _4628_ (.A(\tt6581_inst.controller_inst.filt_start_o ),
    .B(net38),
    .Y(_1003_));
 sg13g2_nor2_1 _4629_ (.A(net42),
    .B(_1003_),
    .Y(_0115_));
 sg13g2_a21oi_1 _4630_ (.A1(_0885_),
    .A2(\tt6581_inst.controller_inst.cur_state[0] ),
    .Y(_0114_),
    .B1(net31));
 sg13g2_or2_1 _4631_ (.X(_1004_),
    .B(\tt6581_inst.svf_inst.cur_state[10] ),
    .A(net1526));
 sg13g2_nand2b_2 _4632_ (.Y(_1005_),
    .B(\tt6581_inst.envelope_inst.cur_state[0] ),
    .A_N(\tt6581_inst.envelope_inst.cur_state[1] ));
 sg13g2_nor3_1 _4633_ (.A(net72),
    .B(net1534),
    .C(net1429),
    .Y(_1006_));
 sg13g2_nand2_1 _4634_ (.Y(_1007_),
    .A(_1005_),
    .B(_1006_));
 sg13g2_nor3_1 _4635_ (.A(\tt6581_inst.mult_inst.iter[1] ),
    .B(\tt6581_inst.mult_inst.iter[0] ),
    .C(\tt6581_inst.mult_inst.iter[3] ),
    .Y(_1008_));
 sg13g2_nand3b_1 _4636_ (.B(_1008_),
    .C(\tt6581_inst.mult_inst.iter[4] ),
    .Y(_1009_),
    .A_N(\tt6581_inst.mult_inst.iter[2] ));
 sg13g2_nor2_2 _4637_ (.A(_1007_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_or2_1 _4638_ (.X(_1011_),
    .B(_1009_),
    .A(_1007_));
 sg13g2_a21o_1 _4639_ (.A2(_1011_),
    .A1(net49),
    .B1(net1526),
    .X(_0017_));
 sg13g2_a21o_1 _4640_ (.A2(_1011_),
    .A1(net51),
    .B1(net1534),
    .X(_0018_));
 sg13g2_a21o_1 _4641_ (.A2(_0884_),
    .A1(net57),
    .B1(net29),
    .X(_0011_));
 sg13g2_nand2_1 _4642_ (.Y(_1012_),
    .A(\tt6581_inst.envelope_inst.cur_state[0] ),
    .B(\tt6581_inst.envelope_inst.cur_state[1] ));
 sg13g2_a21o_1 _4643_ (.A2(_1012_),
    .A1(net55),
    .B1(net30),
    .X(_0010_));
 sg13g2_nand2_1 _4644_ (.Y(_1013_),
    .A(net759),
    .B(\tt6581_inst.controller_inst.cur_state[0] ));
 sg13g2_a21oi_1 _4645_ (.A1(net759),
    .A2(\tt6581_inst.controller_inst.cur_state[0] ),
    .Y(_1014_),
    .B1(net34));
 sg13g2_nor2b_1 _4646_ (.A(net1545),
    .B_N(net1544),
    .Y(_1015_));
 sg13g2_nand2b_2 _4647_ (.Y(_1016_),
    .B(net1544),
    .A_N(net1545));
 sg13g2_o21ai_1 _4648_ (.B1(_1013_),
    .Y(_0012_),
    .A1(_0886_),
    .A2(net1423));
 sg13g2_a21o_1 _4649_ (.A2(_1011_),
    .A1(net53),
    .B1(net213),
    .X(_0016_));
 sg13g2_nand2b_2 _4650_ (.Y(_1017_),
    .B(net47),
    .A_N(net1086));
 sg13g2_inv_1 _4651_ (.Y(_0024_),
    .A(_1017_));
 sg13g2_a21oi_2 _4652_ (.B1(net1542),
    .Y(_1018_),
    .A2(_1006_),
    .A1(_1005_));
 sg13g2_inv_1 _4653_ (.Y(_1019_),
    .A(_1018_));
 sg13g2_and2_1 _4654_ (.A(net1537),
    .B(_1009_),
    .X(_1020_));
 sg13g2_nor2_2 _4655_ (.A(_1018_),
    .B(net1290),
    .Y(_1021_));
 sg13g2_inv_1 _4656_ (.Y(\tt6581_inst.mult_inst.nxt_state ),
    .A(net1229));
 sg13g2_a21o_1 _4657_ (.A2(net64),
    .A1(_0887_),
    .B1(net32),
    .X(_0009_));
 sg13g2_a21o_1 _4658_ (.A2(_1011_),
    .A1(net60),
    .B1(net33),
    .X(_0013_));
 sg13g2_nor2_1 _4659_ (.A(net636),
    .B(net44),
    .Y(_1022_));
 sg13g2_and2_1 _4660_ (.A(net112),
    .B(_1022_),
    .X(_0023_));
 sg13g2_nand3_1 _4661_ (.B(net46),
    .C(net1040),
    .A(net81),
    .Y(_1023_));
 sg13g2_nand4_1 _4662_ (.B(\tt6581_inst.tick_gen_inst.cnt[6] ),
    .C(\tt6581_inst.tick_gen_inst.cnt[8] ),
    .A(\tt6581_inst.tick_gen_inst.cnt[7] ),
    .Y(_1024_),
    .D(\tt6581_inst.tick_gen_inst.cnt[9] ));
 sg13g2_nand2_1 _4663_ (.Y(_1025_),
    .A(_0889_),
    .B(\tt6581_inst.tick_gen_inst.cnt[5] ));
 sg13g2_nor4_2 _4664_ (.A(net266),
    .B(_1023_),
    .C(_1024_),
    .Y(_0035_),
    .D(_1025_));
 sg13g2_nor2_1 _4665_ (.A(net44),
    .B(_0023_),
    .Y(_0020_));
 sg13g2_and2_1 _4666_ (.A(net636),
    .B(net44),
    .X(_1026_));
 sg13g2_nor2_1 _4667_ (.A(_1022_),
    .B(_1026_),
    .Y(_0021_));
 sg13g2_mux2_1 _4668_ (.A0(_1026_),
    .A1(_0021_),
    .S(net112),
    .X(_0022_));
 sg13g2_nor2b_1 _4669_ (.A(\tt6581_inst.spi_inst.cs_sync[1] ),
    .B_N(\tt6581_inst.spi_inst.data_out_reg[7] ),
    .Y(miso));
 sg13g2_xor2_1 _4670_ (.B(net46),
    .A(net81),
    .X(_0026_));
 sg13g2_a21o_1 _4671_ (.A2(net46),
    .A1(net81),
    .B1(net1040),
    .X(_1027_));
 sg13g2_and2_1 _4672_ (.A(_1023_),
    .B(_1027_),
    .X(_0027_));
 sg13g2_xor2_1 _4673_ (.B(_1023_),
    .A(net266),
    .X(_1028_));
 sg13g2_nor2_1 _4674_ (.A(net267),
    .B(_1028_),
    .Y(_0028_));
 sg13g2_nand4_1 _4675_ (.B(net46),
    .C(net266),
    .A(net81),
    .Y(_1029_),
    .D(net1107));
 sg13g2_nor2_1 _4676_ (.A(_0889_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_xnor2_1 _4677_ (.Y(_0029_),
    .A(net67),
    .B(_1029_));
 sg13g2_nor2_1 _4678_ (.A(net468),
    .B(_1030_),
    .Y(_1031_));
 sg13g2_and2_1 _4679_ (.A(net468),
    .B(_1030_),
    .X(_1032_));
 sg13g2_nor3_1 _4680_ (.A(net267),
    .B(net469),
    .C(_1032_),
    .Y(_0030_));
 sg13g2_nor2_1 _4681_ (.A(net502),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_and2_1 _4682_ (.A(net502),
    .B(_1032_),
    .X(_1034_));
 sg13g2_nor3_1 _4683_ (.A(net267),
    .B(net503),
    .C(_1034_),
    .Y(_0031_));
 sg13g2_nor2_1 _4684_ (.A(net526),
    .B(_1034_),
    .Y(_1035_));
 sg13g2_and2_1 _4685_ (.A(net526),
    .B(_1034_),
    .X(_1036_));
 sg13g2_nor3_1 _4686_ (.A(net267),
    .B(_1035_),
    .C(_1036_),
    .Y(_0032_));
 sg13g2_nor2_1 _4687_ (.A(net545),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_and2_1 _4688_ (.A(net545),
    .B(_1036_),
    .X(_1038_));
 sg13g2_nor3_1 _4689_ (.A(net267),
    .B(_1037_),
    .C(_1038_),
    .Y(_0033_));
 sg13g2_a21oi_1 _4690_ (.A1(net825),
    .A2(_1038_),
    .Y(_1039_),
    .B1(net267));
 sg13g2_o21ai_1 _4691_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net825),
    .A2(_1038_));
 sg13g2_inv_1 _4692_ (.Y(_0034_),
    .A(_1040_));
 sg13g2_o21ai_1 _4693_ (.B1(_0881_),
    .Y(_1041_),
    .A1(net114),
    .A2(net120));
 sg13g2_a21oi_1 _4694_ (.A1(net114),
    .A2(_1011_),
    .Y(\tt6581_inst.envelope_inst.nxt_state[0] ),
    .B1(_1041_));
 sg13g2_xor2_1 _4695_ (.B(net114),
    .A(net77),
    .X(\tt6581_inst.envelope_inst.nxt_state[1] ));
 sg13g2_nor3_1 _4696_ (.A(\tt6581_inst.multi_voice_inst.cur_state[1] ),
    .B(\tt6581_inst.multi_voice_inst.cur_state[0] ),
    .C(_0996_),
    .Y(\tt6581_inst.multi_voice_inst.nxt_state[0] ));
 sg13g2_nor2b_1 _4697_ (.A(net47),
    .B_N(\tt6581_inst.multi_voice_inst.cur_state[0] ),
    .Y(\tt6581_inst.multi_voice_inst.nxt_state[1] ));
 sg13g2_and2_1 _4698_ (.A(net51),
    .B(_1010_),
    .X(_0005_));
 sg13g2_nor2b_1 _4699_ (.A(net38),
    .B_N(\tt6581_inst.controller_inst.filt_start_o ),
    .Y(_0006_));
 sg13g2_and2_1 _4700_ (.A(net53),
    .B(_1010_),
    .X(_0007_));
 sg13g2_and2_1 _4701_ (.A(net49),
    .B(_1010_),
    .X(_0008_));
 sg13g2_and2_1 _4702_ (.A(net60),
    .B(_1010_),
    .X(_0001_));
 sg13g2_nor2_1 _4703_ (.A(_0886_),
    .B(net1416),
    .Y(_0002_));
 sg13g2_and2_1 _4704_ (.A(net42),
    .B(net64),
    .X(_0000_));
 sg13g2_nor2b_2 _4705_ (.A(net1544),
    .B_N(net1545),
    .Y(_1042_));
 sg13g2_nand2b_2 _4706_ (.Y(_1043_),
    .B(net1545),
    .A_N(net1544));
 sg13g2_nor2_1 _4707_ (.A(\tt6581_inst.controller_inst.cur_voice[1] ),
    .B(\tt6581_inst.controller_inst.cur_voice[0] ),
    .Y(_1044_));
 sg13g2_nand2_1 _4708_ (.Y(_1045_),
    .A(net764),
    .B(net1419));
 sg13g2_a22oi_1 _4709_ (.Y(_1046_),
    .B1(net1383),
    .B2(net593),
    .A2(net1398),
    .A1(net873));
 sg13g2_a21oi_1 _4710_ (.A1(_1045_),
    .A2(_1046_),
    .Y(_0019_),
    .B1(_0886_));
 sg13g2_and2_1 _4711_ (.A(net57),
    .B(net59),
    .X(_0004_));
 sg13g2_and3_1 _4712_ (.X(_0003_),
    .A(net77),
    .B(\tt6581_inst.envelope_inst.cur_state[1] ),
    .C(net55));
 sg13g2_nand2b_2 _4713_ (.Y(_1047_),
    .B(net1451),
    .A_N(net1449));
 sg13g2_nor2_2 _4714_ (.A(\tt6581_inst.reg_addr[5] ),
    .B(\tt6581_inst.reg_addr[6] ),
    .Y(_1048_));
 sg13g2_nand2_2 _4715_ (.Y(_1049_),
    .A(_0879_),
    .B(_1048_));
 sg13g2_nor2b_1 _4716_ (.A(\tt6581_inst.reg_addr[2] ),
    .B_N(\tt6581_inst.reg_addr[3] ),
    .Y(_1050_));
 sg13g2_nand3_1 _4717_ (.B(_1048_),
    .C(_1050_),
    .A(_0879_),
    .Y(_1051_));
 sg13g2_nor2_1 _4718_ (.A(_1047_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_nand2_2 _4719_ (.Y(_1053_),
    .A(net1445),
    .B(net1286));
 sg13g2_mux2_1 _4720_ (.A0(net1485),
    .A1(net1046),
    .S(net1220),
    .X(_0117_));
 sg13g2_mux2_1 _4721_ (.A0(net1481),
    .A1(net744),
    .S(net1220),
    .X(_0118_));
 sg13g2_mux2_1 _4722_ (.A0(net1476),
    .A1(net830),
    .S(net1220),
    .X(_0119_));
 sg13g2_mux2_1 _4723_ (.A0(net1471),
    .A1(net595),
    .S(_1053_),
    .X(_0120_));
 sg13g2_mux2_1 _4724_ (.A0(net1467),
    .A1(net700),
    .S(net1220),
    .X(_0121_));
 sg13g2_nor2_1 _4725_ (.A(net1463),
    .B(net1220),
    .Y(_1054_));
 sg13g2_a21oi_1 _4726_ (.A1(_0967_),
    .A2(net1220),
    .Y(_0122_),
    .B1(_1054_));
 sg13g2_mux2_1 _4727_ (.A0(net1457),
    .A1(net639),
    .S(_1053_),
    .X(_0123_));
 sg13g2_nor2_1 _4728_ (.A(net1453),
    .B(net1220),
    .Y(_1055_));
 sg13g2_a21oi_1 _4729_ (.A1(_0965_),
    .A2(net1220),
    .Y(_0124_),
    .B1(_1055_));
 sg13g2_or2_1 _4730_ (.X(_1056_),
    .B(\tt6581_inst.reg_addr[2] ),
    .A(\tt6581_inst.reg_addr[3] ));
 sg13g2_nand2b_2 _4731_ (.Y(_1057_),
    .B(net1449),
    .A_N(net1451));
 sg13g2_nor3_1 _4732_ (.A(_1049_),
    .B(_1056_),
    .C(_1057_),
    .Y(_1058_));
 sg13g2_nand2_2 _4733_ (.Y(_1059_),
    .A(net1445),
    .B(net1285));
 sg13g2_mux2_1 _4734_ (.A0(net1486),
    .A1(net1028),
    .S(_1059_),
    .X(_0125_));
 sg13g2_mux2_1 _4735_ (.A0(net1481),
    .A1(net990),
    .S(_1059_),
    .X(_0126_));
 sg13g2_mux2_1 _4736_ (.A0(net1478),
    .A1(net936),
    .S(_1059_),
    .X(_0127_));
 sg13g2_mux2_1 _4737_ (.A0(net1473),
    .A1(net558),
    .S(_1059_),
    .X(_0128_));
 sg13g2_mux2_1 _4738_ (.A0(net1466),
    .A1(net994),
    .S(_1059_),
    .X(_0129_));
 sg13g2_mux2_1 _4739_ (.A0(net1462),
    .A1(net952),
    .S(_1059_),
    .X(_0130_));
 sg13g2_mux2_1 _4740_ (.A0(net1457),
    .A1(net768),
    .S(_1059_),
    .X(_0131_));
 sg13g2_mux2_1 _4741_ (.A0(net1453),
    .A1(net523),
    .S(_1059_),
    .X(_0132_));
 sg13g2_nor3_2 _4742_ (.A(net1451),
    .B(net1449),
    .C(_1051_),
    .Y(_1060_));
 sg13g2_nand2_2 _4743_ (.Y(_1061_),
    .A(net1445),
    .B(net1284));
 sg13g2_mux2_1 _4744_ (.A0(net1485),
    .A1(net785),
    .S(net1219),
    .X(_0133_));
 sg13g2_mux2_1 _4745_ (.A0(net1481),
    .A1(net739),
    .S(net1219),
    .X(_0134_));
 sg13g2_mux2_1 _4746_ (.A0(net1476),
    .A1(net671),
    .S(_1061_),
    .X(_0135_));
 sg13g2_mux2_1 _4747_ (.A0(net1471),
    .A1(net581),
    .S(_1061_),
    .X(_0136_));
 sg13g2_mux2_1 _4748_ (.A0(net1467),
    .A1(net987),
    .S(net1219),
    .X(_0137_));
 sg13g2_mux2_1 _4749_ (.A0(net1463),
    .A1(net619),
    .S(net1219),
    .X(_0138_));
 sg13g2_nor2_1 _4750_ (.A(net1457),
    .B(net1219),
    .Y(_1062_));
 sg13g2_a21oi_1 _4751_ (.A1(_0952_),
    .A2(net1219),
    .Y(_0139_),
    .B1(_1062_));
 sg13g2_nor2_1 _4752_ (.A(net1453),
    .B(net1219),
    .Y(_1063_));
 sg13g2_a21oi_1 _4753_ (.A1(_0951_),
    .A2(net1219),
    .Y(_0140_),
    .B1(_1063_));
 sg13g2_nor3_2 _4754_ (.A(_1047_),
    .B(_1049_),
    .C(_1056_),
    .Y(_1064_));
 sg13g2_nand2_2 _4755_ (.Y(_1065_),
    .A(net1445),
    .B(net1283));
 sg13g2_mux2_1 _4756_ (.A0(net1485),
    .A1(net708),
    .S(_1065_),
    .X(_0141_));
 sg13g2_mux2_1 _4757_ (.A0(net1481),
    .A1(net621),
    .S(_1065_),
    .X(_0142_));
 sg13g2_mux2_1 _4758_ (.A0(net1476),
    .A1(net618),
    .S(_1065_),
    .X(_0143_));
 sg13g2_mux2_1 _4759_ (.A0(net1471),
    .A1(net628),
    .S(_1065_),
    .X(_0144_));
 sg13g2_mux2_1 _4760_ (.A0(net1467),
    .A1(net835),
    .S(_1065_),
    .X(_0145_));
 sg13g2_mux2_1 _4761_ (.A0(net1463),
    .A1(net926),
    .S(_1065_),
    .X(_0146_));
 sg13g2_mux2_1 _4762_ (.A0(net1458),
    .A1(net551),
    .S(_1065_),
    .X(_0147_));
 sg13g2_mux2_1 _4763_ (.A0(net1453),
    .A1(net575),
    .S(_1065_),
    .X(_0148_));
 sg13g2_nand2_2 _4764_ (.Y(_1066_),
    .A(net1451),
    .B(net1449));
 sg13g2_nand2b_2 _4765_ (.Y(_1067_),
    .B(\tt6581_inst.reg_addr[2] ),
    .A_N(\tt6581_inst.reg_addr[3] ));
 sg13g2_nor3_1 _4766_ (.A(_1049_),
    .B(_1066_),
    .C(_1067_),
    .Y(_1068_));
 sg13g2_nand2_2 _4767_ (.Y(_1069_),
    .A(net1446),
    .B(net1282));
 sg13g2_nor2_1 _4768_ (.A(net1486),
    .B(net1218),
    .Y(_1070_));
 sg13g2_a21oi_1 _4769_ (.A1(_0907_),
    .A2(net1218),
    .Y(_0149_),
    .B1(_1070_));
 sg13g2_mux2_1 _4770_ (.A0(net1482),
    .A1(net999),
    .S(net1218),
    .X(_0150_));
 sg13g2_mux2_1 _4771_ (.A0(net1478),
    .A1(net808),
    .S(_1069_),
    .X(_0151_));
 sg13g2_mux2_1 _4772_ (.A0(net1473),
    .A1(net746),
    .S(net1218),
    .X(_0152_));
 sg13g2_mux2_1 _4773_ (.A0(net1466),
    .A1(net929),
    .S(net1218),
    .X(_0153_));
 sg13g2_mux2_1 _4774_ (.A0(net1462),
    .A1(net734),
    .S(net1218),
    .X(_0154_));
 sg13g2_mux2_1 _4775_ (.A0(net1458),
    .A1(net697),
    .S(net1218),
    .X(_0155_));
 sg13g2_mux2_1 _4776_ (.A0(net1454),
    .A1(net753),
    .S(net1218),
    .X(_0156_));
 sg13g2_nor4_1 _4777_ (.A(net1452),
    .B(net1450),
    .C(_1049_),
    .D(_1056_),
    .Y(_1071_));
 sg13g2_nand2_2 _4778_ (.Y(_1072_),
    .A(net1446),
    .B(net1281));
 sg13g2_mux2_1 _4779_ (.A0(net1486),
    .A1(net799),
    .S(_1072_),
    .X(_0157_));
 sg13g2_mux2_1 _4780_ (.A0(net1484),
    .A1(net756),
    .S(_1072_),
    .X(_0158_));
 sg13g2_mux2_1 _4781_ (.A0(net1478),
    .A1(net696),
    .S(_1072_),
    .X(_0159_));
 sg13g2_mux2_1 _4782_ (.A0(net1473),
    .A1(net814),
    .S(_1072_),
    .X(_0160_));
 sg13g2_mux2_1 _4783_ (.A0(net1466),
    .A1(net633),
    .S(_1072_),
    .X(_0161_));
 sg13g2_mux2_1 _4784_ (.A0(net1462),
    .A1(net797),
    .S(_1072_),
    .X(_0162_));
 sg13g2_mux2_1 _4785_ (.A0(net1458),
    .A1(net676),
    .S(_1072_),
    .X(_0163_));
 sg13g2_mux2_1 _4786_ (.A0(net1454),
    .A1(net1070),
    .S(_1072_),
    .X(_0164_));
 sg13g2_nor4_2 _4787_ (.A(\tt6581_inst.mult_inst.accum[3] ),
    .B(\tt6581_inst.mult_inst.accum[2] ),
    .C(\tt6581_inst.mult_inst.accum[1] ),
    .Y(_1073_),
    .D(\tt6581_inst.mult_inst.accum[0] ));
 sg13g2_nor4_2 _4788_ (.A(\tt6581_inst.mult_inst.accum[7] ),
    .B(\tt6581_inst.mult_inst.accum[6] ),
    .C(\tt6581_inst.mult_inst.accum[5] ),
    .Y(_1074_),
    .D(\tt6581_inst.mult_inst.accum[4] ));
 sg13g2_nand2_1 _4789_ (.Y(_1075_),
    .A(_1073_),
    .B(_1074_));
 sg13g2_nand4_1 _4790_ (.B(_0910_),
    .C(_1073_),
    .A(_0908_),
    .Y(_1076_),
    .D(_1074_));
 sg13g2_or3_1 _4791_ (.A(net1536),
    .B(\tt6581_inst.mult_inst.accum[11] ),
    .C(_1076_),
    .X(_1077_));
 sg13g2_a21oi_2 _4792_ (.B1(_0912_),
    .Y(_1078_),
    .A2(_1077_),
    .A1(net1501));
 sg13g2_and3_2 _4793_ (.X(_1079_),
    .A(net1501),
    .B(_0912_),
    .C(_1077_));
 sg13g2_or2_1 _4794_ (.X(_1080_),
    .B(_1079_),
    .A(_1078_));
 sg13g2_nor3_1 _4795_ (.A(\tt6581_inst.svf_inst.reg_low[0] ),
    .B(_1078_),
    .C(_1079_),
    .Y(_1081_));
 sg13g2_o21ai_1 _4796_ (.B1(\tt6581_inst.svf_inst.reg_low[0] ),
    .Y(_1082_),
    .A1(_1078_),
    .A2(_1079_));
 sg13g2_nor2b_1 _4797_ (.A(_1081_),
    .B_N(_1082_),
    .Y(_1083_));
 sg13g2_o21ai_1 _4798_ (.B1(net1513),
    .Y(_1084_),
    .A1(\tt6581_inst.filter_accum[0] ),
    .A2(_1083_));
 sg13g2_a21oi_1 _4799_ (.A1(\tt6581_inst.filter_accum[0] ),
    .A2(_1083_),
    .Y(_1085_),
    .B1(_1084_));
 sg13g2_a21o_1 _4800_ (.A2(_0997_),
    .A1(net640),
    .B1(_1085_),
    .X(_0165_));
 sg13g2_nor2_1 _4801_ (.A(net996),
    .B(net1514),
    .Y(_1086_));
 sg13g2_a21oi_1 _4802_ (.A1(\tt6581_inst.filter_accum[0] ),
    .A2(_1082_),
    .Y(_1087_),
    .B1(_1081_));
 sg13g2_or4_1 _4803_ (.A(net1536),
    .B(\tt6581_inst.mult_inst.accum[11] ),
    .C(\tt6581_inst.mult_inst.accum[12] ),
    .D(_1076_),
    .X(_1088_));
 sg13g2_nand2_1 _4804_ (.Y(_1089_),
    .A(net1501),
    .B(_1088_));
 sg13g2_xnor2_1 _4805_ (.Y(_1090_),
    .A(\tt6581_inst.mult_inst.accum[13] ),
    .B(_1089_));
 sg13g2_xnor2_1 _4806_ (.Y(_1091_),
    .A(\tt6581_inst.svf_inst.reg_low[1] ),
    .B(net1191));
 sg13g2_nand2b_1 _4807_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_1087_));
 sg13g2_xor2_1 _4808_ (.B(_1091_),
    .A(_1087_),
    .X(_1093_));
 sg13g2_xnor2_1 _4809_ (.Y(_1094_),
    .A(_0990_),
    .B(_1093_));
 sg13g2_a21oi_1 _4810_ (.A1(net1514),
    .A2(_1094_),
    .Y(_0166_),
    .B1(_1086_));
 sg13g2_o21ai_1 _4811_ (.B1(_1092_),
    .Y(_1095_),
    .A1(_0990_),
    .A2(_1093_));
 sg13g2_o21ai_1 _4812_ (.B1(net1501),
    .Y(_1096_),
    .A1(\tt6581_inst.mult_inst.accum[13] ),
    .A2(_1088_));
 sg13g2_xnor2_1 _4813_ (.Y(_1097_),
    .A(\tt6581_inst.mult_inst.accum[14] ),
    .B(_1096_));
 sg13g2_nor2_1 _4814_ (.A(\tt6581_inst.svf_inst.reg_low[2] ),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_xnor2_1 _4815_ (.Y(_1099_),
    .A(_0942_),
    .B(_1097_));
 sg13g2_xnor2_1 _4816_ (.Y(_1100_),
    .A(\tt6581_inst.filter_accum[2] ),
    .B(_1099_));
 sg13g2_a21oi_1 _4817_ (.A1(\tt6581_inst.svf_inst.reg_low[1] ),
    .A2(net1191),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_nand3_1 _4818_ (.B(net1191),
    .C(_1100_),
    .A(\tt6581_inst.svf_inst.reg_low[1] ),
    .Y(_1102_));
 sg13g2_nand2b_1 _4819_ (.Y(_1103_),
    .B(_1102_),
    .A_N(_1101_));
 sg13g2_xor2_1 _4820_ (.B(_1103_),
    .A(_1095_),
    .X(_1104_));
 sg13g2_nor2_1 _4821_ (.A(net597),
    .B(net1514),
    .Y(_1105_));
 sg13g2_a21oi_1 _4822_ (.A1(net1514),
    .A2(_1104_),
    .Y(_0167_),
    .B1(_1105_));
 sg13g2_a21oi_1 _4823_ (.A1(_1095_),
    .A2(_1102_),
    .Y(_1106_),
    .B1(_1101_));
 sg13g2_or3_1 _4824_ (.A(\tt6581_inst.mult_inst.accum[13] ),
    .B(\tt6581_inst.mult_inst.accum[14] ),
    .C(_1088_),
    .X(_1107_));
 sg13g2_a21oi_2 _4825_ (.B1(_0914_),
    .Y(_1108_),
    .A2(_1107_),
    .A1(net1501));
 sg13g2_and3_2 _4826_ (.X(_1109_),
    .A(net1501),
    .B(_0914_),
    .C(_1107_));
 sg13g2_or2_1 _4827_ (.X(_1110_),
    .B(_1109_),
    .A(_1108_));
 sg13g2_nor2_1 _4828_ (.A(net1507),
    .B(net1185),
    .Y(_1111_));
 sg13g2_xor2_1 _4829_ (.B(net1185),
    .A(\tt6581_inst.svf_inst.reg_low[3] ),
    .X(_1112_));
 sg13g2_xnor2_1 _4830_ (.Y(_1113_),
    .A(\tt6581_inst.filter_accum[3] ),
    .B(_1112_));
 sg13g2_a21oi_1 _4831_ (.A1(\tt6581_inst.filter_accum[2] ),
    .A2(_1099_),
    .Y(_1114_),
    .B1(_1098_));
 sg13g2_or2_1 _4832_ (.X(_1115_),
    .B(_1114_),
    .A(_1113_));
 sg13g2_xnor2_1 _4833_ (.Y(_1116_),
    .A(_1113_),
    .B(_1114_));
 sg13g2_xor2_1 _4834_ (.B(_1116_),
    .A(_1106_),
    .X(_1117_));
 sg13g2_mux2_1 _4835_ (.A0(net1105),
    .A1(_1117_),
    .S(net1514),
    .X(_0168_));
 sg13g2_nor2_1 _4836_ (.A(net747),
    .B(net1513),
    .Y(_1118_));
 sg13g2_o21ai_1 _4837_ (.B1(_1115_),
    .Y(_1119_),
    .A1(_1106_),
    .A2(_1116_));
 sg13g2_nor4_1 _4838_ (.A(\tt6581_inst.mult_inst.accum[13] ),
    .B(\tt6581_inst.mult_inst.accum[14] ),
    .C(\tt6581_inst.mult_inst.accum[15] ),
    .D(_1088_),
    .Y(_1120_));
 sg13g2_or4_1 _4839_ (.A(\tt6581_inst.mult_inst.accum[13] ),
    .B(\tt6581_inst.mult_inst.accum[14] ),
    .C(\tt6581_inst.mult_inst.accum[15] ),
    .D(_1088_),
    .X(_1121_));
 sg13g2_a21oi_2 _4840_ (.B1(_0915_),
    .Y(_1122_),
    .A2(_1121_),
    .A1(net1501));
 sg13g2_nor3_2 _4841_ (.A(_0909_),
    .B(\tt6581_inst.mult_inst.accum[16] ),
    .C(_1120_),
    .Y(_1123_));
 sg13g2_or2_1 _4842_ (.X(_1124_),
    .B(_1123_),
    .A(_1122_));
 sg13g2_nor2_1 _4843_ (.A(\tt6581_inst.svf_inst.reg_low[4] ),
    .B(net1184),
    .Y(_1125_));
 sg13g2_xnor2_1 _4844_ (.Y(_1126_),
    .A(_0941_),
    .B(net1184));
 sg13g2_xnor2_1 _4845_ (.Y(_1127_),
    .A(\tt6581_inst.filter_accum[4] ),
    .B(_1126_));
 sg13g2_a21oi_1 _4846_ (.A1(\tt6581_inst.filter_accum[3] ),
    .A2(_1112_),
    .Y(_1128_),
    .B1(_1111_));
 sg13g2_nor2_1 _4847_ (.A(_1127_),
    .B(_1128_),
    .Y(_1129_));
 sg13g2_nand2_1 _4848_ (.Y(_1130_),
    .A(_1127_),
    .B(_1128_));
 sg13g2_nand2b_1 _4849_ (.Y(_1131_),
    .B(_1130_),
    .A_N(_1129_));
 sg13g2_xor2_1 _4850_ (.B(_1131_),
    .A(_1119_),
    .X(_1132_));
 sg13g2_a21oi_1 _4851_ (.A1(net1513),
    .A2(_1132_),
    .Y(_0169_),
    .B1(net748));
 sg13g2_a21oi_1 _4852_ (.A1(_1119_),
    .A2(_1130_),
    .Y(_1133_),
    .B1(_1129_));
 sg13g2_nand2_1 _4853_ (.Y(_1134_),
    .A(_0915_),
    .B(_1120_));
 sg13g2_o21ai_1 _4854_ (.B1(net1502),
    .Y(_1135_),
    .A1(\tt6581_inst.mult_inst.accum[16] ),
    .A2(_1121_));
 sg13g2_xnor2_1 _4855_ (.Y(_1136_),
    .A(\tt6581_inst.mult_inst.accum[17] ),
    .B(_1135_));
 sg13g2_nor2_1 _4856_ (.A(net1506),
    .B(net1182),
    .Y(_1137_));
 sg13g2_xor2_1 _4857_ (.B(net1182),
    .A(net1506),
    .X(_1138_));
 sg13g2_xnor2_1 _4858_ (.Y(_1139_),
    .A(\tt6581_inst.filter_accum[5] ),
    .B(_1138_));
 sg13g2_a21oi_1 _4859_ (.A1(\tt6581_inst.filter_accum[4] ),
    .A2(_1126_),
    .Y(_1140_),
    .B1(_1125_));
 sg13g2_or2_1 _4860_ (.X(_1141_),
    .B(_1140_),
    .A(_1139_));
 sg13g2_xnor2_1 _4861_ (.Y(_1142_),
    .A(_1139_),
    .B(_1140_));
 sg13g2_nor2_1 _4862_ (.A(_1133_),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_nand2_1 _4863_ (.Y(_1144_),
    .A(net710),
    .B(_0997_));
 sg13g2_a21o_1 _4864_ (.A2(_1142_),
    .A1(_1133_),
    .B1(_0997_),
    .X(_1145_));
 sg13g2_o21ai_1 _4865_ (.B1(_1144_),
    .Y(_0170_),
    .A1(_1143_),
    .A2(_1145_));
 sg13g2_nor2_1 _4866_ (.A(net715),
    .B(net1513),
    .Y(_1146_));
 sg13g2_o21ai_1 _4867_ (.B1(_1141_),
    .Y(_1147_),
    .A1(_1133_),
    .A2(_1142_));
 sg13g2_o21ai_1 _4868_ (.B1(net1503),
    .Y(_1148_),
    .A1(\tt6581_inst.mult_inst.accum[17] ),
    .A2(_1134_));
 sg13g2_xnor2_1 _4869_ (.Y(_1149_),
    .A(\tt6581_inst.mult_inst.accum[18] ),
    .B(_1148_));
 sg13g2_nor2_1 _4870_ (.A(\tt6581_inst.svf_inst.reg_low[6] ),
    .B(net1173),
    .Y(_1150_));
 sg13g2_xnor2_1 _4871_ (.Y(_1151_),
    .A(_0940_),
    .B(net1173));
 sg13g2_xnor2_1 _4872_ (.Y(_1152_),
    .A(\tt6581_inst.filter_accum[6] ),
    .B(_1151_));
 sg13g2_a21oi_1 _4873_ (.A1(\tt6581_inst.filter_accum[5] ),
    .A2(_1138_),
    .Y(_1153_),
    .B1(_1137_));
 sg13g2_nor2_1 _4874_ (.A(_1152_),
    .B(_1153_),
    .Y(_1154_));
 sg13g2_nand2_1 _4875_ (.Y(_1155_),
    .A(_1152_),
    .B(_1153_));
 sg13g2_nand2b_1 _4876_ (.Y(_1156_),
    .B(_1155_),
    .A_N(_1154_));
 sg13g2_xor2_1 _4877_ (.B(_1156_),
    .A(_1147_),
    .X(_1157_));
 sg13g2_a21oi_1 _4878_ (.A1(net1513),
    .A2(_1157_),
    .Y(_0171_),
    .B1(net716));
 sg13g2_nor2_1 _4879_ (.A(net847),
    .B(net1513),
    .Y(_1158_));
 sg13g2_a21oi_1 _4880_ (.A1(_1147_),
    .A2(_1155_),
    .Y(_1159_),
    .B1(_1154_));
 sg13g2_nor3_1 _4881_ (.A(\tt6581_inst.mult_inst.accum[17] ),
    .B(\tt6581_inst.mult_inst.accum[18] ),
    .C(_1134_),
    .Y(_1160_));
 sg13g2_nor2_1 _4882_ (.A(_0909_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_xor2_1 _4883_ (.B(_1161_),
    .A(\tt6581_inst.mult_inst.accum[19] ),
    .X(_1162_));
 sg13g2_nor2_1 _4884_ (.A(\tt6581_inst.svf_inst.reg_low[7] ),
    .B(net1166),
    .Y(_1163_));
 sg13g2_xnor2_1 _4885_ (.Y(_1164_),
    .A(_0939_),
    .B(net1166));
 sg13g2_xnor2_1 _4886_ (.Y(_1165_),
    .A(\tt6581_inst.filter_accum[7] ),
    .B(_1164_));
 sg13g2_a21oi_1 _4887_ (.A1(\tt6581_inst.filter_accum[6] ),
    .A2(_1151_),
    .Y(_1166_),
    .B1(_1150_));
 sg13g2_nor2_1 _4888_ (.A(_1165_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_inv_1 _4889_ (.Y(_1168_),
    .A(_1167_));
 sg13g2_xor2_1 _4890_ (.B(_1166_),
    .A(_1165_),
    .X(_1169_));
 sg13g2_inv_1 _4891_ (.Y(_1170_),
    .A(_1169_));
 sg13g2_xnor2_1 _4892_ (.Y(_1171_),
    .A(_1159_),
    .B(_1170_));
 sg13g2_a21oi_1 _4893_ (.A1(net1513),
    .A2(_1171_),
    .Y(_0172_),
    .B1(net848));
 sg13g2_nor2_1 _4894_ (.A(net864),
    .B(net1515),
    .Y(_1172_));
 sg13g2_o21ai_1 _4895_ (.B1(_1168_),
    .Y(_1173_),
    .A1(_1159_),
    .A2(_1170_));
 sg13g2_or4_1 _4896_ (.A(\tt6581_inst.mult_inst.accum[17] ),
    .B(\tt6581_inst.mult_inst.accum[18] ),
    .C(\tt6581_inst.mult_inst.accum[19] ),
    .D(_1134_),
    .X(_1174_));
 sg13g2_nand2_1 _4897_ (.Y(_1175_),
    .A(net1503),
    .B(_1174_));
 sg13g2_xnor2_1 _4898_ (.Y(_1176_),
    .A(\tt6581_inst.mult_inst.accum[20] ),
    .B(_1175_));
 sg13g2_nor2_1 _4899_ (.A(\tt6581_inst.svf_inst.reg_low[8] ),
    .B(net1164),
    .Y(_1177_));
 sg13g2_xnor2_1 _4900_ (.Y(_1178_),
    .A(_0938_),
    .B(net1164));
 sg13g2_xnor2_1 _4901_ (.Y(_1179_),
    .A(\tt6581_inst.filter_accum[8] ),
    .B(_1178_));
 sg13g2_a21oi_1 _4902_ (.A1(\tt6581_inst.filter_accum[7] ),
    .A2(_1164_),
    .Y(_1180_),
    .B1(_1163_));
 sg13g2_nor2_1 _4903_ (.A(_1179_),
    .B(_1180_),
    .Y(_1181_));
 sg13g2_xor2_1 _4904_ (.B(_1180_),
    .A(_1179_),
    .X(_1182_));
 sg13g2_xnor2_1 _4905_ (.Y(_1183_),
    .A(_1173_),
    .B(_1182_));
 sg13g2_a21oi_1 _4906_ (.A1(net1515),
    .A2(_1183_),
    .Y(_0173_),
    .B1(net865));
 sg13g2_nor2_1 _4907_ (.A(net1008),
    .B(net1515),
    .Y(_1184_));
 sg13g2_a21o_1 _4908_ (.A2(_1182_),
    .A1(_1173_),
    .B1(_1181_),
    .X(_1185_));
 sg13g2_o21ai_1 _4909_ (.B1(net1503),
    .Y(_1186_),
    .A1(\tt6581_inst.mult_inst.accum[20] ),
    .A2(_1174_));
 sg13g2_xnor2_1 _4910_ (.Y(_1187_),
    .A(\tt6581_inst.mult_inst.accum[21] ),
    .B(_1186_));
 sg13g2_xor2_1 _4911_ (.B(_1186_),
    .A(\tt6581_inst.mult_inst.accum[21] ),
    .X(_1188_));
 sg13g2_nor2_1 _4912_ (.A(net1505),
    .B(_1187_),
    .Y(_1189_));
 sg13g2_xnor2_1 _4913_ (.Y(_1190_),
    .A(net1505),
    .B(_1188_));
 sg13g2_xnor2_1 _4914_ (.Y(_1191_),
    .A(\tt6581_inst.filter_accum[9] ),
    .B(_1190_));
 sg13g2_a21oi_1 _4915_ (.A1(\tt6581_inst.filter_accum[8] ),
    .A2(_1178_),
    .Y(_1192_),
    .B1(_1177_));
 sg13g2_nor2_1 _4916_ (.A(_1191_),
    .B(_1192_),
    .Y(_1193_));
 sg13g2_xor2_1 _4917_ (.B(_1192_),
    .A(_1191_),
    .X(_1194_));
 sg13g2_xnor2_1 _4918_ (.Y(_1195_),
    .A(_1185_),
    .B(_1194_));
 sg13g2_a21oi_1 _4919_ (.A1(net1515),
    .A2(_1195_),
    .Y(_0174_),
    .B1(net1009));
 sg13g2_nor2_1 _4920_ (.A(net957),
    .B(net1515),
    .Y(_1196_));
 sg13g2_a21o_2 _4921_ (.A2(_1194_),
    .A1(_1185_),
    .B1(_1193_),
    .X(_1197_));
 sg13g2_nor3_1 _4922_ (.A(\tt6581_inst.mult_inst.accum[20] ),
    .B(\tt6581_inst.mult_inst.accum[21] ),
    .C(_1174_),
    .Y(_1198_));
 sg13g2_nor2_1 _4923_ (.A(_0909_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_xor2_1 _4924_ (.B(_1199_),
    .A(\tt6581_inst.mult_inst.accum[22] ),
    .X(_1200_));
 sg13g2_xnor2_1 _4925_ (.Y(_1201_),
    .A(_0937_),
    .B(_1200_));
 sg13g2_nand2_1 _4926_ (.Y(_1202_),
    .A(\tt6581_inst.filter_accum[10] ),
    .B(_1201_));
 sg13g2_xnor2_1 _4927_ (.Y(_1203_),
    .A(\tt6581_inst.filter_accum[10] ),
    .B(_1201_));
 sg13g2_a21oi_1 _4928_ (.A1(\tt6581_inst.filter_accum[9] ),
    .A2(_1190_),
    .Y(_1204_),
    .B1(_1189_));
 sg13g2_nor2_1 _4929_ (.A(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_xor2_1 _4930_ (.B(_1204_),
    .A(_1203_),
    .X(_1206_));
 sg13g2_xnor2_1 _4931_ (.Y(_1207_),
    .A(_1197_),
    .B(_1206_));
 sg13g2_a21oi_1 _4932_ (.A1(net1515),
    .A2(_1207_),
    .Y(_0175_),
    .B1(net958));
 sg13g2_a21oi_1 _4933_ (.A1(_1197_),
    .A2(_1206_),
    .Y(_1208_),
    .B1(_1205_));
 sg13g2_nand2b_2 _4934_ (.Y(_1209_),
    .B(_1198_),
    .A_N(\tt6581_inst.mult_inst.accum[22] ));
 sg13g2_nand2_1 _4935_ (.Y(_1210_),
    .A(net1503),
    .B(_1209_));
 sg13g2_xnor2_1 _4936_ (.Y(_1211_),
    .A(\tt6581_inst.mult_inst.accum[23] ),
    .B(_1210_));
 sg13g2_xor2_1 _4937_ (.B(_1210_),
    .A(\tt6581_inst.mult_inst.accum[23] ),
    .X(_1212_));
 sg13g2_xnor2_1 _4938_ (.Y(_1213_),
    .A(\tt6581_inst.svf_inst.reg_low[11] ),
    .B(_1211_));
 sg13g2_nor2_1 _4939_ (.A(_0993_),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_xnor2_1 _4940_ (.Y(_1215_),
    .A(_0993_),
    .B(_1213_));
 sg13g2_inv_1 _4941_ (.Y(_1216_),
    .A(_1215_));
 sg13g2_o21ai_1 _4942_ (.B1(_1202_),
    .Y(_1217_),
    .A1(\tt6581_inst.svf_inst.reg_low[10] ),
    .A2(_1200_));
 sg13g2_nand2b_1 _4943_ (.Y(_1218_),
    .B(_1215_),
    .A_N(_1217_));
 sg13g2_inv_1 _4944_ (.Y(_1219_),
    .A(_1218_));
 sg13g2_xor2_1 _4945_ (.B(_1217_),
    .A(_1215_),
    .X(_1220_));
 sg13g2_xor2_1 _4946_ (.B(_1220_),
    .A(_1208_),
    .X(_1221_));
 sg13g2_nor2_1 _4947_ (.A(_0997_),
    .B(_1221_),
    .Y(_1222_));
 sg13g2_a21oi_1 _4948_ (.A1(_0935_),
    .A2(_0997_),
    .Y(_0176_),
    .B1(_1222_));
 sg13g2_o21ai_1 _4949_ (.B1(net1503),
    .Y(_1223_),
    .A1(\tt6581_inst.mult_inst.accum[23] ),
    .A2(_1209_));
 sg13g2_xor2_1 _4950_ (.B(_1223_),
    .A(\tt6581_inst.mult_inst.accum[24] ),
    .X(_1224_));
 sg13g2_inv_1 _4951_ (.Y(_1225_),
    .A(_1224_));
 sg13g2_xnor2_1 _4952_ (.Y(_1226_),
    .A(_0934_),
    .B(_1224_));
 sg13g2_nor2_1 _4953_ (.A(_0994_),
    .B(_1226_),
    .Y(_1227_));
 sg13g2_xnor2_1 _4954_ (.Y(_1228_),
    .A(_0994_),
    .B(_1226_));
 sg13g2_a21oi_1 _4955_ (.A1(_0936_),
    .A2(_1212_),
    .Y(_1229_),
    .B1(_1214_));
 sg13g2_nor2_1 _4956_ (.A(_1228_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_xnor2_1 _4957_ (.Y(_1231_),
    .A(_1228_),
    .B(_1229_));
 sg13g2_a221oi_1 _4958_ (.B2(_1217_),
    .C1(_1205_),
    .B1(_1216_),
    .A1(_1197_),
    .Y(_1232_),
    .A2(_1206_));
 sg13g2_nor3_1 _4959_ (.A(_1219_),
    .B(_1231_),
    .C(_1232_),
    .Y(_1233_));
 sg13g2_o21ai_1 _4960_ (.B1(_1231_),
    .Y(_1234_),
    .A1(_1219_),
    .A2(_1232_));
 sg13g2_nand2b_1 _4961_ (.Y(_1235_),
    .B(_1234_),
    .A_N(_1233_));
 sg13g2_nor2_1 _4962_ (.A(net720),
    .B(net1512),
    .Y(_1236_));
 sg13g2_a21oi_1 _4963_ (.A1(net1512),
    .A2(_1235_),
    .Y(_0177_),
    .B1(net721));
 sg13g2_nor3_1 _4964_ (.A(\tt6581_inst.mult_inst.accum[23] ),
    .B(\tt6581_inst.mult_inst.accum[24] ),
    .C(_1209_),
    .Y(_1237_));
 sg13g2_nor2_1 _4965_ (.A(_0909_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_xor2_1 _4966_ (.B(_1238_),
    .A(\tt6581_inst.mult_inst.accum[25] ),
    .X(_1239_));
 sg13g2_nor2_1 _4967_ (.A(\tt6581_inst.svf_inst.reg_low[13] ),
    .B(_1239_),
    .Y(_1240_));
 sg13g2_xor2_1 _4968_ (.B(_1239_),
    .A(\tt6581_inst.svf_inst.reg_low[13] ),
    .X(_1241_));
 sg13g2_xnor2_1 _4969_ (.Y(_1242_),
    .A(net1497),
    .B(_1241_));
 sg13g2_a21oi_1 _4970_ (.A1(_0934_),
    .A2(_1224_),
    .Y(_1243_),
    .B1(_1227_));
 sg13g2_nor2_1 _4971_ (.A(_1242_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_inv_1 _4972_ (.Y(_1245_),
    .A(_1244_));
 sg13g2_xnor2_1 _4973_ (.Y(_1246_),
    .A(_1242_),
    .B(_1243_));
 sg13g2_inv_1 _4974_ (.Y(_1247_),
    .A(_1246_));
 sg13g2_o21ai_1 _4975_ (.B1(_1247_),
    .Y(_1248_),
    .A1(_1230_),
    .A2(_1233_));
 sg13g2_or3_1 _4976_ (.A(_1230_),
    .B(_1233_),
    .C(_1247_),
    .X(_1249_));
 sg13g2_nand3_1 _4977_ (.B(_1248_),
    .C(_1249_),
    .A(net1512),
    .Y(_1250_));
 sg13g2_o21ai_1 _4978_ (.B1(_1250_),
    .Y(_0178_),
    .A1(_0933_),
    .A2(net1512));
 sg13g2_nand2b_2 _4979_ (.Y(_1251_),
    .B(_1237_),
    .A_N(\tt6581_inst.mult_inst.accum[25] ));
 sg13g2_nand2_1 _4980_ (.Y(_1252_),
    .A(net1504),
    .B(_1251_));
 sg13g2_xnor2_1 _4981_ (.Y(_1253_),
    .A(\tt6581_inst.mult_inst.accum[26] ),
    .B(_1252_));
 sg13g2_xor2_1 _4982_ (.B(_1252_),
    .A(\tt6581_inst.mult_inst.accum[26] ),
    .X(_1254_));
 sg13g2_xnor2_1 _4983_ (.Y(_1255_),
    .A(\tt6581_inst.svf_inst.reg_low[14] ),
    .B(_1253_));
 sg13g2_nor2_1 _4984_ (.A(_0995_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_xnor2_1 _4985_ (.Y(_1257_),
    .A(_0995_),
    .B(_1255_));
 sg13g2_a21oi_1 _4986_ (.A1(net1497),
    .A2(_1241_),
    .Y(_1258_),
    .B1(_1240_));
 sg13g2_nor2_1 _4987_ (.A(_1257_),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_inv_1 _4988_ (.Y(_1260_),
    .A(_1259_));
 sg13g2_xnor2_1 _4989_ (.Y(_1261_),
    .A(_1257_),
    .B(_1258_));
 sg13g2_a21o_1 _4990_ (.A2(_1248_),
    .A1(_1245_),
    .B1(_1261_),
    .X(_1262_));
 sg13g2_nand3_1 _4991_ (.B(_1248_),
    .C(_1261_),
    .A(_1245_),
    .Y(_1263_));
 sg13g2_a21oi_1 _4992_ (.A1(_1262_),
    .A2(_1263_),
    .Y(_1264_),
    .B1(_0997_));
 sg13g2_a21oi_1 _4993_ (.A1(_0931_),
    .A2(_0997_),
    .Y(_0179_),
    .B1(_1264_));
 sg13g2_o21ai_1 _4994_ (.B1(net1500),
    .Y(_1265_),
    .A1(\tt6581_inst.mult_inst.accum[26] ),
    .A2(_1251_));
 sg13g2_inv_1 _4995_ (.Y(_1266_),
    .A(_1265_));
 sg13g2_xnor2_1 _4996_ (.Y(_1267_),
    .A(\tt6581_inst.mult_inst.accum[27] ),
    .B(_1265_));
 sg13g2_nor2_1 _4997_ (.A(\tt6581_inst.svf_inst.reg_low[15] ),
    .B(_1267_),
    .Y(_1268_));
 sg13g2_xnor2_1 _4998_ (.Y(_1269_),
    .A(\tt6581_inst.svf_inst.reg_low[15] ),
    .B(_1267_));
 sg13g2_nor2_1 _4999_ (.A(_0995_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_xnor2_1 _5000_ (.Y(_1271_),
    .A(_0995_),
    .B(_1269_));
 sg13g2_a21oi_1 _5001_ (.A1(_0932_),
    .A2(_1254_),
    .Y(_1272_),
    .B1(_1256_));
 sg13g2_nor2_1 _5002_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_inv_1 _5003_ (.Y(_1274_),
    .A(_1273_));
 sg13g2_xnor2_1 _5004_ (.Y(_1275_),
    .A(_1271_),
    .B(_1272_));
 sg13g2_a21o_1 _5005_ (.A2(_1262_),
    .A1(_1260_),
    .B1(_1275_),
    .X(_1276_));
 sg13g2_nand3_1 _5006_ (.B(_1262_),
    .C(_1275_),
    .A(_1260_),
    .Y(_1277_));
 sg13g2_nand3_1 _5007_ (.B(_1276_),
    .C(_1277_),
    .A(net1509),
    .Y(_1278_));
 sg13g2_o21ai_1 _5008_ (.B1(_1278_),
    .Y(_0180_),
    .A1(_0929_),
    .A2(net1511));
 sg13g2_a21oi_1 _5009_ (.A1(net1500),
    .A2(\tt6581_inst.mult_inst.accum[27] ),
    .Y(_1279_),
    .B1(_1266_));
 sg13g2_xnor2_1 _5010_ (.Y(_1280_),
    .A(\tt6581_inst.mult_inst.accum[28] ),
    .B(_1279_));
 sg13g2_nand2b_1 _5011_ (.Y(_1281_),
    .B(_0928_),
    .A_N(_1280_));
 sg13g2_xnor2_1 _5012_ (.Y(_1282_),
    .A(_0928_),
    .B(_1280_));
 sg13g2_nand2_1 _5013_ (.Y(_1283_),
    .A(net1495),
    .B(_1282_));
 sg13g2_xnor2_1 _5014_ (.Y(_1284_),
    .A(net1495),
    .B(_1282_));
 sg13g2_nor2_1 _5015_ (.A(_1268_),
    .B(_1270_),
    .Y(_1285_));
 sg13g2_nor2_1 _5016_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_xnor2_1 _5017_ (.Y(_1287_),
    .A(_1284_),
    .B(_1285_));
 sg13g2_a21oi_1 _5018_ (.A1(_1274_),
    .A2(_1276_),
    .Y(_1288_),
    .B1(_1287_));
 sg13g2_nand3_1 _5019_ (.B(_1276_),
    .C(_1287_),
    .A(_1274_),
    .Y(_1289_));
 sg13g2_nand2b_1 _5020_ (.Y(_1290_),
    .B(net499),
    .A_N(net1509));
 sg13g2_nand2_1 _5021_ (.Y(_1291_),
    .A(net1509),
    .B(_1289_));
 sg13g2_o21ai_1 _5022_ (.B1(_1290_),
    .Y(_0181_),
    .A1(_1288_),
    .A2(_1291_));
 sg13g2_nor2_1 _5023_ (.A(net851),
    .B(net1509),
    .Y(_1292_));
 sg13g2_nor2_1 _5024_ (.A(_1286_),
    .B(_1288_),
    .Y(_1293_));
 sg13g2_nor4_1 _5025_ (.A(\tt6581_inst.mult_inst.accum[26] ),
    .B(\tt6581_inst.mult_inst.accum[27] ),
    .C(\tt6581_inst.mult_inst.accum[28] ),
    .D(_1251_),
    .Y(_1294_));
 sg13g2_nor2_1 _5026_ (.A(_0909_),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_xnor2_1 _5027_ (.Y(_1296_),
    .A(_0987_),
    .B(_1295_));
 sg13g2_xnor2_1 _5028_ (.Y(_1297_),
    .A(_0927_),
    .B(_1296_));
 sg13g2_nand2_1 _5029_ (.Y(_1298_),
    .A(net1495),
    .B(_1297_));
 sg13g2_xnor2_1 _5030_ (.Y(_1299_),
    .A(net1495),
    .B(_1297_));
 sg13g2_nand3_1 _5031_ (.B(_1283_),
    .C(_1299_),
    .A(_1281_),
    .Y(_1300_));
 sg13g2_a21o_1 _5032_ (.A2(_1283_),
    .A1(_1281_),
    .B1(_1299_),
    .X(_1301_));
 sg13g2_nand2_1 _5033_ (.Y(_1302_),
    .A(_1300_),
    .B(_1301_));
 sg13g2_xnor2_1 _5034_ (.Y(_1303_),
    .A(_1293_),
    .B(_1302_));
 sg13g2_a21oi_1 _5035_ (.A1(net1509),
    .A2(_1303_),
    .Y(_0182_),
    .B1(_1292_));
 sg13g2_a21oi_2 _5036_ (.B1(_0909_),
    .Y(_1304_),
    .A2(_1294_),
    .A1(_0987_));
 sg13g2_xor2_1 _5037_ (.B(_1304_),
    .A(\tt6581_inst.mult_inst.accum[30] ),
    .X(_1305_));
 sg13g2_xnor2_1 _5038_ (.Y(_1306_),
    .A(\tt6581_inst.mult_inst.accum[30] ),
    .B(_1304_));
 sg13g2_nand2_1 _5039_ (.Y(_1307_),
    .A(_0925_),
    .B(_1306_));
 sg13g2_xnor2_1 _5040_ (.Y(_1308_),
    .A(_0925_),
    .B(_1305_));
 sg13g2_nand2_1 _5041_ (.Y(_1309_),
    .A(net1495),
    .B(_1308_));
 sg13g2_xnor2_1 _5042_ (.Y(_1310_),
    .A(net1495),
    .B(_1308_));
 sg13g2_o21ai_1 _5043_ (.B1(_1298_),
    .Y(_1311_),
    .A1(\tt6581_inst.svf_inst.reg_low[17] ),
    .A2(_1296_));
 sg13g2_nor2b_1 _5044_ (.A(_1310_),
    .B_N(_1311_),
    .Y(_1312_));
 sg13g2_xor2_1 _5045_ (.B(_1311_),
    .A(_1310_),
    .X(_1313_));
 sg13g2_o21ai_1 _5046_ (.B1(_1300_),
    .Y(_1314_),
    .A1(_1286_),
    .A2(_1288_));
 sg13g2_a21oi_1 _5047_ (.A1(_1301_),
    .A2(_1314_),
    .Y(_1315_),
    .B1(_1313_));
 sg13g2_nand3_1 _5048_ (.B(_1313_),
    .C(_1314_),
    .A(_1301_),
    .Y(_1316_));
 sg13g2_nand2b_1 _5049_ (.Y(_1317_),
    .B(net694),
    .A_N(net1509));
 sg13g2_nand2_1 _5050_ (.Y(_1318_),
    .A(net1509),
    .B(_1316_));
 sg13g2_o21ai_1 _5051_ (.B1(_1317_),
    .Y(_0183_),
    .A1(_1315_),
    .A2(_1318_));
 sg13g2_a21oi_1 _5052_ (.A1(net1500),
    .A2(\tt6581_inst.mult_inst.accum[30] ),
    .Y(_1319_),
    .B1(_1304_));
 sg13g2_xnor2_1 _5053_ (.Y(_1320_),
    .A(\tt6581_inst.mult_inst.accum[31] ),
    .B(_1319_));
 sg13g2_nor2_1 _5054_ (.A(\tt6581_inst.svf_inst.reg_low[19] ),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_xnor2_1 _5055_ (.Y(_1322_),
    .A(_0924_),
    .B(_1320_));
 sg13g2_xnor2_1 _5056_ (.Y(_1323_),
    .A(net1495),
    .B(_1322_));
 sg13g2_a21oi_1 _5057_ (.A1(_1307_),
    .A2(_1309_),
    .Y(_1324_),
    .B1(_1323_));
 sg13g2_nand3_1 _5058_ (.B(_1309_),
    .C(_1323_),
    .A(_1307_),
    .Y(_1325_));
 sg13g2_nor2b_1 _5059_ (.A(_1324_),
    .B_N(_1325_),
    .Y(_1326_));
 sg13g2_nor2_1 _5060_ (.A(_1312_),
    .B(_1315_),
    .Y(_1327_));
 sg13g2_xnor2_1 _5061_ (.Y(_1328_),
    .A(_1326_),
    .B(_1327_));
 sg13g2_mux2_1 _5062_ (.A0(net1106),
    .A1(_1328_),
    .S(net1509),
    .X(_0184_));
 sg13g2_nor2_1 _5063_ (.A(net559),
    .B(net1510),
    .Y(_1329_));
 sg13g2_o21ai_1 _5064_ (.B1(_1319_),
    .Y(_1330_),
    .A1(_0909_),
    .A2(_0988_));
 sg13g2_xnor2_1 _5065_ (.Y(_1331_),
    .A(\tt6581_inst.mult_inst.accum[32] ),
    .B(_1330_));
 sg13g2_and2_1 _5066_ (.A(_0923_),
    .B(_1331_),
    .X(_1332_));
 sg13g2_xnor2_1 _5067_ (.Y(_1333_),
    .A(\tt6581_inst.svf_inst.reg_low[20] ),
    .B(_1331_));
 sg13g2_xnor2_1 _5068_ (.Y(_1334_),
    .A(net1496),
    .B(_1333_));
 sg13g2_a21oi_1 _5069_ (.A1(net1496),
    .A2(_1322_),
    .Y(_1335_),
    .B1(_1321_));
 sg13g2_nor2_1 _5070_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_xnor2_1 _5071_ (.Y(_1337_),
    .A(_1334_),
    .B(_1335_));
 sg13g2_or2_1 _5072_ (.X(_1338_),
    .B(_1324_),
    .A(_1312_));
 sg13g2_o21ai_1 _5073_ (.B1(_1325_),
    .Y(_1339_),
    .A1(_1315_),
    .A2(_1338_));
 sg13g2_nor2_1 _5074_ (.A(_1337_),
    .B(_1339_),
    .Y(_1340_));
 sg13g2_xnor2_1 _5075_ (.Y(_1341_),
    .A(_1337_),
    .B(_1339_));
 sg13g2_a21oi_1 _5076_ (.A1(net1510),
    .A2(_1341_),
    .Y(_0185_),
    .B1(_1329_));
 sg13g2_a21o_1 _5077_ (.A2(\tt6581_inst.mult_inst.accum[32] ),
    .A1(net1500),
    .B1(_1330_),
    .X(_1342_));
 sg13g2_xor2_1 _5078_ (.B(_1342_),
    .A(\tt6581_inst.mult_inst.accum[33] ),
    .X(_1343_));
 sg13g2_nor2_1 _5079_ (.A(\tt6581_inst.svf_inst.reg_low[21] ),
    .B(_1343_),
    .Y(_1344_));
 sg13g2_xnor2_1 _5080_ (.Y(_1345_),
    .A(_0922_),
    .B(_1343_));
 sg13g2_xnor2_1 _5081_ (.Y(_1346_),
    .A(net1496),
    .B(_1345_));
 sg13g2_a21oi_1 _5082_ (.A1(net1496),
    .A2(_1333_),
    .Y(_1347_),
    .B1(_1332_));
 sg13g2_nor2_1 _5083_ (.A(_1346_),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_inv_1 _5084_ (.Y(_1349_),
    .A(_1348_));
 sg13g2_xor2_1 _5085_ (.B(_1347_),
    .A(_1346_),
    .X(_1350_));
 sg13g2_o21ai_1 _5086_ (.B1(_1350_),
    .Y(_1351_),
    .A1(_1336_),
    .A2(_1340_));
 sg13g2_or3_1 _5087_ (.A(_1336_),
    .B(_1340_),
    .C(_1350_),
    .X(_1352_));
 sg13g2_nand3_1 _5088_ (.B(_1351_),
    .C(_1352_),
    .A(net1510),
    .Y(_1353_));
 sg13g2_o21ai_1 _5089_ (.B1(_1353_),
    .Y(_0186_),
    .A1(_0921_),
    .A2(net1510));
 sg13g2_a21oi_1 _5090_ (.A1(net1500),
    .A2(\tt6581_inst.mult_inst.accum[33] ),
    .Y(_1354_),
    .B1(_1342_));
 sg13g2_xor2_1 _5091_ (.B(_1354_),
    .A(\tt6581_inst.mult_inst.accum[34] ),
    .X(_1355_));
 sg13g2_inv_2 _5092_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_xnor2_1 _5093_ (.Y(_1357_),
    .A(_0920_),
    .B(_1355_));
 sg13g2_nor2_1 _5094_ (.A(_0995_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_xnor2_1 _5095_ (.Y(_1359_),
    .A(_0995_),
    .B(_1357_));
 sg13g2_a21oi_1 _5096_ (.A1(net1495),
    .A2(_1345_),
    .Y(_1360_),
    .B1(_1344_));
 sg13g2_nor2_1 _5097_ (.A(_1359_),
    .B(_1360_),
    .Y(_1361_));
 sg13g2_xnor2_1 _5098_ (.Y(_1362_),
    .A(_1359_),
    .B(_1360_));
 sg13g2_a21oi_1 _5099_ (.A1(_1349_),
    .A2(_1351_),
    .Y(_1363_),
    .B1(_1362_));
 sg13g2_nand3_1 _5100_ (.B(_1351_),
    .C(_1362_),
    .A(_1349_),
    .Y(_1364_));
 sg13g2_nand2b_1 _5101_ (.Y(_1365_),
    .B(net500),
    .A_N(net1510));
 sg13g2_nand2_1 _5102_ (.Y(_1366_),
    .A(net1511),
    .B(_1364_));
 sg13g2_o21ai_1 _5103_ (.B1(_1365_),
    .Y(_0187_),
    .A1(_1363_),
    .A2(_1366_));
 sg13g2_nor2_1 _5104_ (.A(net535),
    .B(net1510),
    .Y(_1367_));
 sg13g2_nor2_1 _5105_ (.A(_1361_),
    .B(_1363_),
    .Y(_1368_));
 sg13g2_a21oi_1 _5106_ (.A1(_0920_),
    .A2(_1355_),
    .Y(_1369_),
    .B1(_1358_));
 sg13g2_nor3_1 _5107_ (.A(\tt6581_inst.mult_inst.accum[33] ),
    .B(\tt6581_inst.mult_inst.accum[34] ),
    .C(_1342_),
    .Y(_1370_));
 sg13g2_nor2_1 _5108_ (.A(_0909_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_xor2_1 _5109_ (.B(_1371_),
    .A(\tt6581_inst.mult_inst.accum[35] ),
    .X(_1372_));
 sg13g2_xor2_1 _5110_ (.B(net1496),
    .A(\tt6581_inst.svf_inst.reg_low[23] ),
    .X(_1373_));
 sg13g2_xnor2_1 _5111_ (.Y(_1374_),
    .A(_1372_),
    .B(_1373_));
 sg13g2_xnor2_1 _5112_ (.Y(_1375_),
    .A(_1369_),
    .B(_1374_));
 sg13g2_xnor2_1 _5113_ (.Y(_1376_),
    .A(_1368_),
    .B(_1375_));
 sg13g2_a21oi_1 _5114_ (.A1(net1510),
    .A2(_1376_),
    .Y(_0188_),
    .B1(_1367_));
 sg13g2_nor3_1 _5115_ (.A(_1049_),
    .B(_1057_),
    .C(_1067_),
    .Y(_1377_));
 sg13g2_nand2_2 _5116_ (.Y(_1378_),
    .A(net1448),
    .B(net1280));
 sg13g2_mux2_1 _5117_ (.A0(net1487),
    .A1(net933),
    .S(_1378_),
    .X(_0189_));
 sg13g2_mux2_1 _5118_ (.A0(net1483),
    .A1(net1037),
    .S(_1378_),
    .X(_0190_));
 sg13g2_mux2_1 _5119_ (.A0(net1479),
    .A1(net1066),
    .S(_1378_),
    .X(_0191_));
 sg13g2_mux2_1 _5120_ (.A0(net1474),
    .A1(net1092),
    .S(_1378_),
    .X(_0192_));
 sg13g2_mux2_1 _5121_ (.A0(net1470),
    .A1(net1085),
    .S(_1378_),
    .X(_0193_));
 sg13g2_mux2_1 _5122_ (.A0(net1464),
    .A1(net860),
    .S(_1378_),
    .X(_0194_));
 sg13g2_mux2_1 _5123_ (.A0(net1460),
    .A1(net954),
    .S(_1378_),
    .X(_0195_));
 sg13g2_mux2_1 _5124_ (.A0(net1456),
    .A1(net948),
    .S(_1378_),
    .X(_0196_));
 sg13g2_nand4_1 _5125_ (.B(\tt6581_inst.reg_addr[2] ),
    .C(_0879_),
    .A(\tt6581_inst.reg_addr[3] ),
    .Y(_1379_),
    .D(_1048_));
 sg13g2_nor2_2 _5126_ (.A(_1047_),
    .B(_1379_),
    .Y(_1380_));
 sg13g2_nand2_2 _5127_ (.Y(_1381_),
    .A(net1447),
    .B(net1279));
 sg13g2_mux2_1 _5128_ (.A0(net1487),
    .A1(net741),
    .S(_1381_),
    .X(_0197_));
 sg13g2_mux2_1 _5129_ (.A0(net1484),
    .A1(net805),
    .S(_1381_),
    .X(_0198_));
 sg13g2_mux2_1 _5130_ (.A0(net1479),
    .A1(net1013),
    .S(_1381_),
    .X(_0199_));
 sg13g2_mux2_1 _5131_ (.A0(net1474),
    .A1(net906),
    .S(_1381_),
    .X(_0200_));
 sg13g2_mux2_1 _5132_ (.A0(net1468),
    .A1(net678),
    .S(_1381_),
    .X(_0201_));
 sg13g2_mux2_1 _5133_ (.A0(net1464),
    .A1(net1007),
    .S(_1381_),
    .X(_0202_));
 sg13g2_mux2_1 _5134_ (.A0(net1459),
    .A1(net962),
    .S(_1381_),
    .X(_0203_));
 sg13g2_mux2_1 _5135_ (.A0(net1455),
    .A1(net940),
    .S(_1381_),
    .X(_0204_));
 sg13g2_nor3_2 _5136_ (.A(net1452),
    .B(net1450),
    .C(_1379_),
    .Y(_1382_));
 sg13g2_nand2_2 _5137_ (.Y(_1383_),
    .A(net1448),
    .B(net1278));
 sg13g2_mux2_1 _5138_ (.A0(net1487),
    .A1(net680),
    .S(_1383_),
    .X(_0205_));
 sg13g2_mux2_1 _5139_ (.A0(net1483),
    .A1(net844),
    .S(_1383_),
    .X(_0206_));
 sg13g2_mux2_1 _5140_ (.A0(net1479),
    .A1(net931),
    .S(_1383_),
    .X(_0207_));
 sg13g2_mux2_1 _5141_ (.A0(net1474),
    .A1(net760),
    .S(_1383_),
    .X(_0208_));
 sg13g2_mux2_1 _5142_ (.A0(net1468),
    .A1(net751),
    .S(_1383_),
    .X(_0209_));
 sg13g2_mux2_1 _5143_ (.A0(net1465),
    .A1(net950),
    .S(_1383_),
    .X(_0210_));
 sg13g2_mux2_1 _5144_ (.A0(net1459),
    .A1(net1058),
    .S(_1383_),
    .X(_0211_));
 sg13g2_mux2_1 _5145_ (.A0(net1456),
    .A1(net1033),
    .S(_1383_),
    .X(_0212_));
 sg13g2_nor3_1 _5146_ (.A(_1047_),
    .B(_1049_),
    .C(_1067_),
    .Y(_1384_));
 sg13g2_nand2_2 _5147_ (.Y(_1385_),
    .A(net1447),
    .B(net1277));
 sg13g2_mux2_1 _5148_ (.A0(net1487),
    .A1(net911),
    .S(_1385_),
    .X(_0213_));
 sg13g2_mux2_1 _5149_ (.A0(net1484),
    .A1(net966),
    .S(_1385_),
    .X(_0214_));
 sg13g2_mux2_1 _5150_ (.A0(net1479),
    .A1(net1056),
    .S(_1385_),
    .X(_0215_));
 sg13g2_mux2_1 _5151_ (.A0(net1475),
    .A1(net1051),
    .S(_1385_),
    .X(_0216_));
 sg13g2_mux2_1 _5152_ (.A0(net1468),
    .A1(net664),
    .S(_1385_),
    .X(_0217_));
 sg13g2_mux2_1 _5153_ (.A0(net1465),
    .A1(net692),
    .S(_1385_),
    .X(_0218_));
 sg13g2_mux2_1 _5154_ (.A0(net1459),
    .A1(net534),
    .S(_1385_),
    .X(_0219_));
 sg13g2_mux2_1 _5155_ (.A0(net1456),
    .A1(net637),
    .S(_1385_),
    .X(_0220_));
 sg13g2_nor2_1 _5156_ (.A(_1051_),
    .B(_1066_),
    .Y(_1386_));
 sg13g2_nand2_2 _5157_ (.Y(_1387_),
    .A(net1448),
    .B(net1276));
 sg13g2_mux2_1 _5158_ (.A0(net1488),
    .A1(net774),
    .S(net1217),
    .X(_0221_));
 sg13g2_mux2_1 _5159_ (.A0(net1481),
    .A1(net787),
    .S(net1217),
    .X(_0222_));
 sg13g2_nor2_1 _5160_ (.A(net1478),
    .B(_1387_),
    .Y(_1388_));
 sg13g2_a21oi_1 _5161_ (.A1(_0972_),
    .A2(_1387_),
    .Y(_0223_),
    .B1(_1388_));
 sg13g2_mux2_1 _5162_ (.A0(net1474),
    .A1(net406),
    .S(_1387_),
    .X(_0224_));
 sg13g2_mux2_1 _5163_ (.A0(net1466),
    .A1(net867),
    .S(net1217),
    .X(_0225_));
 sg13g2_mux2_1 _5164_ (.A0(net1463),
    .A1(net934),
    .S(net1217),
    .X(_0226_));
 sg13g2_nor2_1 _5165_ (.A(net1457),
    .B(net1217),
    .Y(_1389_));
 sg13g2_a21oi_1 _5166_ (.A1(_0970_),
    .A2(net1217),
    .Y(_0227_),
    .B1(_1389_));
 sg13g2_nor2_1 _5167_ (.A(net1453),
    .B(net1217),
    .Y(_1390_));
 sg13g2_a21oi_1 _5168_ (.A1(_0971_),
    .A2(net1217),
    .Y(_0228_),
    .B1(_1390_));
 sg13g2_nor4_2 _5169_ (.A(net1451),
    .B(net1449),
    .C(_1049_),
    .Y(_1391_),
    .D(_1067_));
 sg13g2_nand2_2 _5170_ (.Y(_1392_),
    .A(net1446),
    .B(net1275));
 sg13g2_mux2_1 _5171_ (.A0(net1487),
    .A1(net852),
    .S(_1392_),
    .X(_0229_));
 sg13g2_mux2_1 _5172_ (.A0(net1482),
    .A1(net737),
    .S(_1392_),
    .X(_0230_));
 sg13g2_mux2_1 _5173_ (.A0(net1478),
    .A1(net602),
    .S(_1392_),
    .X(_0231_));
 sg13g2_mux2_1 _5174_ (.A0(net1473),
    .A1(net386),
    .S(_1392_),
    .X(_0232_));
 sg13g2_mux2_1 _5175_ (.A0(net1466),
    .A1(net688),
    .S(_1392_),
    .X(_0233_));
 sg13g2_mux2_1 _5176_ (.A0(net1462),
    .A1(net591),
    .S(_1392_),
    .X(_0234_));
 sg13g2_mux2_1 _5177_ (.A0(net1461),
    .A1(net585),
    .S(_1392_),
    .X(_0235_));
 sg13g2_mux2_1 _5178_ (.A0(net1453),
    .A1(net625),
    .S(_1392_),
    .X(_0236_));
 sg13g2_nor2_1 _5179_ (.A(_1051_),
    .B(_1057_),
    .Y(_1393_));
 sg13g2_nand2_2 _5180_ (.Y(_1394_),
    .A(net1445),
    .B(net1274));
 sg13g2_nor2_1 _5181_ (.A(net1485),
    .B(net1216),
    .Y(_1395_));
 sg13g2_a21oi_1 _5182_ (.A1(_0964_),
    .A2(net1216),
    .Y(_0237_),
    .B1(_1395_));
 sg13g2_mux2_1 _5183_ (.A0(net1482),
    .A1(net567),
    .S(net1216),
    .X(_0238_));
 sg13g2_nor2_1 _5184_ (.A(net1477),
    .B(net1216),
    .Y(_1396_));
 sg13g2_a21oi_1 _5185_ (.A1(_0963_),
    .A2(net1216),
    .Y(_0239_),
    .B1(_1396_));
 sg13g2_mux2_1 _5186_ (.A0(net1471),
    .A1(net903),
    .S(net1216),
    .X(_0240_));
 sg13g2_mux2_1 _5187_ (.A0(net1468),
    .A1(net374),
    .S(net1216),
    .X(_0241_));
 sg13g2_mux2_1 _5188_ (.A0(net1464),
    .A1(net335),
    .S(_1394_),
    .X(_0242_));
 sg13g2_mux2_1 _5189_ (.A0(net1457),
    .A1(net506),
    .S(_1394_),
    .X(_0243_));
 sg13g2_mux2_1 _5190_ (.A0(net1455),
    .A1(net313),
    .S(net1216),
    .X(_0244_));
 sg13g2_nor3_1 _5191_ (.A(_1049_),
    .B(_1056_),
    .C(_1066_),
    .Y(_1397_));
 sg13g2_nand2_2 _5192_ (.Y(_1398_),
    .A(net1446),
    .B(net1273));
 sg13g2_mux2_1 _5193_ (.A0(net1486),
    .A1(net878),
    .S(_1398_),
    .X(_0245_));
 sg13g2_mux2_1 _5194_ (.A0(net1482),
    .A1(net504),
    .S(_1398_),
    .X(_0246_));
 sg13g2_mux2_1 _5195_ (.A0(net1478),
    .A1(net946),
    .S(_1398_),
    .X(_0247_));
 sg13g2_mux2_1 _5196_ (.A0(net1473),
    .A1(net831),
    .S(_1398_),
    .X(_0248_));
 sg13g2_mux2_1 _5197_ (.A0(net1466),
    .A1(net489),
    .S(_1398_),
    .X(_0249_));
 sg13g2_mux2_1 _5198_ (.A0(net1462),
    .A1(net451),
    .S(_1398_),
    .X(_0250_));
 sg13g2_mux2_1 _5199_ (.A0(net1458),
    .A1(net288),
    .S(_1398_),
    .X(_0251_));
 sg13g2_mux2_1 _5200_ (.A0(net1454),
    .A1(net391),
    .S(_1398_),
    .X(_0252_));
 sg13g2_xor2_1 _5201_ (.B(\tt6581_inst.delta_sigma_inst.audio[16] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[15] ),
    .X(_1399_));
 sg13g2_nor2b_1 _5202_ (.A(\tt6581_inst.delta_sigma_inst.e2[16] ),
    .B_N(_1399_),
    .Y(_1400_));
 sg13g2_a21oi_1 _5203_ (.A1(\tt6581_inst.delta_sigma_inst.e1[15] ),
    .A2(\tt6581_inst.delta_sigma_inst.audio[16] ),
    .Y(_1401_),
    .B1(_1400_));
 sg13g2_xnor2_1 _5204_ (.Y(_1402_),
    .A(\tt6581_inst.delta_sigma_inst.e1[16] ),
    .B(\tt6581_inst.delta_sigma_inst.e2[17] ));
 sg13g2_xnor2_1 _5205_ (.Y(_1403_),
    .A(\tt6581_inst.delta_sigma_inst.audio[17] ),
    .B(_1402_));
 sg13g2_nor2_1 _5206_ (.A(_1401_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_xnor2_1 _5207_ (.Y(_1405_),
    .A(_1401_),
    .B(_1403_));
 sg13g2_nand2_1 _5208_ (.Y(_1406_),
    .A(\tt6581_inst.delta_sigma_inst.e1[14] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[15] ));
 sg13g2_nor2_1 _5209_ (.A(\tt6581_inst.delta_sigma_inst.e1[14] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[15] ),
    .Y(_1407_));
 sg13g2_xor2_1 _5210_ (.B(\tt6581_inst.delta_sigma_inst.audio[15] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[14] ),
    .X(_1408_));
 sg13g2_o21ai_1 _5211_ (.B1(_1406_),
    .Y(_1409_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[15] ),
    .A2(_1407_));
 sg13g2_xnor2_1 _5212_ (.Y(_1410_),
    .A(\tt6581_inst.delta_sigma_inst.e2[16] ),
    .B(_1399_));
 sg13g2_nand2_1 _5213_ (.Y(_1411_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_xnor2_1 _5214_ (.Y(_1412_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_xnor2_1 _5215_ (.Y(_1413_),
    .A(\tt6581_inst.delta_sigma_inst.e2[15] ),
    .B(_1408_));
 sg13g2_and2_1 _5216_ (.A(\tt6581_inst.delta_sigma_inst.e1[13] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[14] ),
    .X(_1414_));
 sg13g2_xor2_1 _5217_ (.B(\tt6581_inst.delta_sigma_inst.audio[14] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[13] ),
    .X(_1415_));
 sg13g2_nor2b_1 _5218_ (.A(\tt6581_inst.delta_sigma_inst.e2[14] ),
    .B_N(_1415_),
    .Y(_1416_));
 sg13g2_or3_1 _5219_ (.A(_1413_),
    .B(_1414_),
    .C(_1416_),
    .X(_1417_));
 sg13g2_o21ai_1 _5220_ (.B1(_1413_),
    .Y(_1418_),
    .A1(_1414_),
    .A2(_1416_));
 sg13g2_inv_1 _5221_ (.Y(_1419_),
    .A(_1418_));
 sg13g2_xnor2_1 _5222_ (.Y(_1420_),
    .A(\tt6581_inst.delta_sigma_inst.e2[14] ),
    .B(_1415_));
 sg13g2_nand2_1 _5223_ (.Y(_1421_),
    .A(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[13] ));
 sg13g2_nor2_1 _5224_ (.A(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[13] ),
    .Y(_1422_));
 sg13g2_xor2_1 _5225_ (.B(\tt6581_inst.delta_sigma_inst.audio[13] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .X(_1423_));
 sg13g2_o21ai_1 _5226_ (.B1(_1421_),
    .Y(_1424_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[13] ),
    .A2(_1422_));
 sg13g2_and2_1 _5227_ (.A(_1420_),
    .B(_1424_),
    .X(_1425_));
 sg13g2_xor2_1 _5228_ (.B(_1424_),
    .A(_1420_),
    .X(_1426_));
 sg13g2_and2_1 _5229_ (.A(\tt6581_inst.delta_sigma_inst.e1[11] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[12] ),
    .X(_1427_));
 sg13g2_xor2_1 _5230_ (.B(\tt6581_inst.delta_sigma_inst.audio[12] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[11] ),
    .X(_1428_));
 sg13g2_nor2b_1 _5231_ (.A(\tt6581_inst.delta_sigma_inst.e2[12] ),
    .B_N(_1428_),
    .Y(_1429_));
 sg13g2_xnor2_1 _5232_ (.Y(_1430_),
    .A(\tt6581_inst.delta_sigma_inst.e2[13] ),
    .B(_1423_));
 sg13g2_nor3_1 _5233_ (.A(_1427_),
    .B(_1429_),
    .C(_1430_),
    .Y(_1431_));
 sg13g2_o21ai_1 _5234_ (.B1(_1430_),
    .Y(_1432_),
    .A1(_1427_),
    .A2(_1429_));
 sg13g2_xnor2_1 _5235_ (.Y(_1433_),
    .A(\tt6581_inst.delta_sigma_inst.e2[12] ),
    .B(_1428_));
 sg13g2_nand2_1 _5236_ (.Y(_1434_),
    .A(\tt6581_inst.delta_sigma_inst.e1[10] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[11] ));
 sg13g2_nor2_1 _5237_ (.A(\tt6581_inst.delta_sigma_inst.e1[10] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[11] ),
    .Y(_1435_));
 sg13g2_xor2_1 _5238_ (.B(\tt6581_inst.delta_sigma_inst.audio[11] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[10] ),
    .X(_1436_));
 sg13g2_o21ai_1 _5239_ (.B1(_1434_),
    .Y(_1437_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[11] ),
    .A2(_1435_));
 sg13g2_xnor2_1 _5240_ (.Y(_1438_),
    .A(\tt6581_inst.delta_sigma_inst.e2[11] ),
    .B(_1436_));
 sg13g2_nand2_1 _5241_ (.Y(_1439_),
    .A(\tt6581_inst.delta_sigma_inst.e1[9] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[10] ));
 sg13g2_nor2_1 _5242_ (.A(\tt6581_inst.delta_sigma_inst.e1[9] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[10] ),
    .Y(_1440_));
 sg13g2_xor2_1 _5243_ (.B(\tt6581_inst.delta_sigma_inst.audio[10] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[9] ),
    .X(_1441_));
 sg13g2_o21ai_1 _5244_ (.B1(_1439_),
    .Y(_1442_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[10] ),
    .A2(_1440_));
 sg13g2_nand2_1 _5245_ (.Y(_1443_),
    .A(_1438_),
    .B(_1442_));
 sg13g2_xnor2_1 _5246_ (.Y(_1444_),
    .A(\tt6581_inst.delta_sigma_inst.e2[10] ),
    .B(_1441_));
 sg13g2_nand2_1 _5247_ (.Y(_1445_),
    .A(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[9] ));
 sg13g2_nor2_1 _5248_ (.A(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[9] ),
    .Y(_1446_));
 sg13g2_xor2_1 _5249_ (.B(\tt6581_inst.delta_sigma_inst.audio[9] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .X(_1447_));
 sg13g2_o21ai_1 _5250_ (.B1(_1445_),
    .Y(_1448_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[9] ),
    .A2(_1446_));
 sg13g2_and2_1 _5251_ (.A(_1444_),
    .B(_1448_),
    .X(_1449_));
 sg13g2_xnor2_1 _5252_ (.Y(_1450_),
    .A(\tt6581_inst.delta_sigma_inst.e2[9] ),
    .B(_1447_));
 sg13g2_nand2_1 _5253_ (.Y(_1451_),
    .A(\tt6581_inst.delta_sigma_inst.e1[7] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[8] ));
 sg13g2_nor2_1 _5254_ (.A(\tt6581_inst.delta_sigma_inst.e1[7] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[8] ),
    .Y(_1452_));
 sg13g2_xor2_1 _5255_ (.B(\tt6581_inst.delta_sigma_inst.audio[8] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[7] ),
    .X(_1453_));
 sg13g2_o21ai_1 _5256_ (.B1(_1451_),
    .Y(_1454_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[8] ),
    .A2(_1452_));
 sg13g2_nand2_1 _5257_ (.Y(_1455_),
    .A(_1450_),
    .B(_1454_));
 sg13g2_xnor2_1 _5258_ (.Y(_1456_),
    .A(\tt6581_inst.delta_sigma_inst.e2[8] ),
    .B(_1453_));
 sg13g2_nand2_1 _5259_ (.Y(_1457_),
    .A(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[7] ));
 sg13g2_nor2_1 _5260_ (.A(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[7] ),
    .Y(_1458_));
 sg13g2_xor2_1 _5261_ (.B(\tt6581_inst.delta_sigma_inst.audio[7] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .X(_1459_));
 sg13g2_o21ai_1 _5262_ (.B1(_1457_),
    .Y(_1460_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[7] ),
    .A2(_1458_));
 sg13g2_and2_1 _5263_ (.A(_1456_),
    .B(_1460_),
    .X(_1461_));
 sg13g2_xnor2_1 _5264_ (.Y(_1462_),
    .A(\tt6581_inst.delta_sigma_inst.e2[7] ),
    .B(_1459_));
 sg13g2_nand2_1 _5265_ (.Y(_1463_),
    .A(\tt6581_inst.delta_sigma_inst.e1[5] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[6] ));
 sg13g2_nor2_1 _5266_ (.A(\tt6581_inst.delta_sigma_inst.e1[5] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[6] ),
    .Y(_1464_));
 sg13g2_xor2_1 _5267_ (.B(\tt6581_inst.delta_sigma_inst.audio[6] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[5] ),
    .X(_1465_));
 sg13g2_o21ai_1 _5268_ (.B1(_1463_),
    .Y(_1466_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[6] ),
    .A2(_1464_));
 sg13g2_nand2_1 _5269_ (.Y(_1467_),
    .A(_1462_),
    .B(_1466_));
 sg13g2_xnor2_1 _5270_ (.Y(_1468_),
    .A(\tt6581_inst.delta_sigma_inst.e2[6] ),
    .B(_1465_));
 sg13g2_nand2_1 _5271_ (.Y(_1469_),
    .A(\tt6581_inst.delta_sigma_inst.e1[4] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[5] ));
 sg13g2_nor2_1 _5272_ (.A(\tt6581_inst.delta_sigma_inst.e1[4] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[5] ),
    .Y(_1470_));
 sg13g2_xor2_1 _5273_ (.B(\tt6581_inst.delta_sigma_inst.audio[5] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[4] ),
    .X(_1471_));
 sg13g2_o21ai_1 _5274_ (.B1(_1469_),
    .Y(_1472_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[5] ),
    .A2(_1470_));
 sg13g2_and2_1 _5275_ (.A(_1468_),
    .B(_1472_),
    .X(_1473_));
 sg13g2_xnor2_1 _5276_ (.Y(_1474_),
    .A(\tt6581_inst.delta_sigma_inst.e2[5] ),
    .B(_1471_));
 sg13g2_nand2_1 _5277_ (.Y(_1475_),
    .A(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[4] ));
 sg13g2_nor2_1 _5278_ (.A(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .B(\tt6581_inst.delta_sigma_inst.audio[4] ),
    .Y(_1476_));
 sg13g2_xor2_1 _5279_ (.B(\tt6581_inst.delta_sigma_inst.audio[4] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .X(_1477_));
 sg13g2_o21ai_1 _5280_ (.B1(_1475_),
    .Y(_1478_),
    .A1(\tt6581_inst.delta_sigma_inst.e2[4] ),
    .A2(_1476_));
 sg13g2_nand2_1 _5281_ (.Y(_1479_),
    .A(_1474_),
    .B(_1478_));
 sg13g2_nor2b_1 _5282_ (.A(\tt6581_inst.delta_sigma_inst.e2[3] ),
    .B_N(\tt6581_inst.delta_sigma_inst.e1[2] ),
    .Y(_1480_));
 sg13g2_xnor2_1 _5283_ (.Y(_1481_),
    .A(\tt6581_inst.delta_sigma_inst.e2[4] ),
    .B(_1477_));
 sg13g2_and2_1 _5284_ (.A(_1480_),
    .B(_1481_),
    .X(_1482_));
 sg13g2_nor2_1 _5285_ (.A(_0876_),
    .B(\tt6581_inst.delta_sigma_inst.e2[1] ),
    .Y(_1483_));
 sg13g2_xor2_1 _5286_ (.B(\tt6581_inst.delta_sigma_inst.e2[1] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[0] ),
    .X(_1484_));
 sg13g2_nor2_1 _5287_ (.A(net216),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_nand2b_1 _5288_ (.Y(_1486_),
    .B(\tt6581_inst.delta_sigma_inst.e1[1] ),
    .A_N(\tt6581_inst.delta_sigma_inst.e2[2] ));
 sg13g2_xor2_1 _5289_ (.B(\tt6581_inst.delta_sigma_inst.e2[2] ),
    .A(\tt6581_inst.delta_sigma_inst.e1[1] ),
    .X(_1487_));
 sg13g2_nor3_1 _5290_ (.A(_0876_),
    .B(\tt6581_inst.delta_sigma_inst.e2[1] ),
    .C(_1487_),
    .Y(_1488_));
 sg13g2_xnor2_1 _5291_ (.Y(_1489_),
    .A(_1483_),
    .B(_1487_));
 sg13g2_and2_1 _5292_ (.A(_1485_),
    .B(_1489_),
    .X(_1490_));
 sg13g2_xnor2_1 _5293_ (.Y(_1491_),
    .A(\tt6581_inst.delta_sigma_inst.e1[2] ),
    .B(\tt6581_inst.delta_sigma_inst.e2[3] ));
 sg13g2_inv_1 _5294_ (.Y(_1492_),
    .A(_1491_));
 sg13g2_nor2_1 _5295_ (.A(_1486_),
    .B(_1492_),
    .Y(_1493_));
 sg13g2_nand2_1 _5296_ (.Y(_1494_),
    .A(_1486_),
    .B(_1492_));
 sg13g2_nand2b_1 _5297_ (.Y(_1495_),
    .B(_1494_),
    .A_N(_1493_));
 sg13g2_a221oi_1 _5298_ (.B2(_1490_),
    .C1(_1493_),
    .B1(_1494_),
    .A1(_1488_),
    .Y(_1496_),
    .A2(_1491_));
 sg13g2_xnor2_1 _5299_ (.Y(_1497_),
    .A(_1480_),
    .B(_1481_));
 sg13g2_nor2_1 _5300_ (.A(_1496_),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_xor2_1 _5301_ (.B(_1478_),
    .A(_1474_),
    .X(_1499_));
 sg13g2_o21ai_1 _5302_ (.B1(_1499_),
    .Y(_1500_),
    .A1(_1482_),
    .A2(_1498_));
 sg13g2_xnor2_1 _5303_ (.Y(_1501_),
    .A(_1468_),
    .B(_1472_));
 sg13g2_a21oi_1 _5304_ (.A1(_1479_),
    .A2(_1500_),
    .Y(_1502_),
    .B1(_1501_));
 sg13g2_xor2_1 _5305_ (.B(_1466_),
    .A(_1462_),
    .X(_1503_));
 sg13g2_o21ai_1 _5306_ (.B1(_1503_),
    .Y(_1504_),
    .A1(_1473_),
    .A2(_1502_));
 sg13g2_xnor2_1 _5307_ (.Y(_1505_),
    .A(_1456_),
    .B(_1460_));
 sg13g2_a21oi_1 _5308_ (.A1(_1467_),
    .A2(_1504_),
    .Y(_1506_),
    .B1(_1505_));
 sg13g2_xor2_1 _5309_ (.B(_1454_),
    .A(_1450_),
    .X(_1507_));
 sg13g2_o21ai_1 _5310_ (.B1(_1507_),
    .Y(_1508_),
    .A1(_1461_),
    .A2(_1506_));
 sg13g2_xnor2_1 _5311_ (.Y(_1509_),
    .A(_1444_),
    .B(_1448_));
 sg13g2_a21oi_1 _5312_ (.A1(_1455_),
    .A2(_1508_),
    .Y(_1510_),
    .B1(_1509_));
 sg13g2_xor2_1 _5313_ (.B(_1442_),
    .A(_1438_),
    .X(_1511_));
 sg13g2_o21ai_1 _5314_ (.B1(_1511_),
    .Y(_1512_),
    .A1(_1449_),
    .A2(_1510_));
 sg13g2_xnor2_1 _5315_ (.Y(_1513_),
    .A(_1433_),
    .B(_1437_));
 sg13g2_a21oi_1 _5316_ (.A1(_1443_),
    .A2(_1512_),
    .Y(_1514_),
    .B1(_1513_));
 sg13g2_a21o_1 _5317_ (.A2(_1437_),
    .A1(_1433_),
    .B1(_1514_),
    .X(_1515_));
 sg13g2_inv_1 _5318_ (.Y(_1516_),
    .A(_1515_));
 sg13g2_o21ai_1 _5319_ (.B1(_1432_),
    .Y(_1517_),
    .A1(_1431_),
    .A2(_1516_));
 sg13g2_a21o_1 _5320_ (.A2(_1517_),
    .A1(_1426_),
    .B1(_1425_),
    .X(_1518_));
 sg13g2_a21oi_1 _5321_ (.A1(_1417_),
    .A2(_1518_),
    .Y(_1519_),
    .B1(_1419_));
 sg13g2_or2_1 _5322_ (.X(_1520_),
    .B(_1519_),
    .A(_1412_));
 sg13g2_a21oi_1 _5323_ (.A1(_1411_),
    .A2(_1520_),
    .Y(_1521_),
    .B1(_1405_));
 sg13g2_nor2_1 _5324_ (.A(_1404_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_xnor2_1 _5325_ (.Y(_1523_),
    .A(\tt6581_inst.delta_sigma_inst.e1[17] ),
    .B(\tt6581_inst.delta_sigma_inst.e2[18] ));
 sg13g2_a21oi_1 _5326_ (.A1(\tt6581_inst.delta_sigma_inst.e1[16] ),
    .A2(_0883_),
    .Y(_1524_),
    .B1(\tt6581_inst.delta_sigma_inst.audio[17] ));
 sg13g2_o21ai_1 _5327_ (.B1(\tt6581_inst.delta_sigma_inst.audio[17] ),
    .Y(_1525_),
    .A1(\tt6581_inst.delta_sigma_inst.e1[16] ),
    .A2(_0883_));
 sg13g2_nor2b_1 _5328_ (.A(_1524_),
    .B_N(_1525_),
    .Y(_1526_));
 sg13g2_xnor2_1 _5329_ (.Y(_1527_),
    .A(_1523_),
    .B(_1526_));
 sg13g2_xnor2_1 _5330_ (.Y(_1528_),
    .A(_1522_),
    .B(_1527_));
 sg13g2_mux2_1 _5331_ (.A0(net758),
    .A1(_1528_),
    .S(net1549),
    .X(_0253_));
 sg13g2_nand2_1 _5332_ (.Y(_1529_),
    .A(net34),
    .B(_1013_));
 sg13g2_nand2_1 _5333_ (.Y(_1530_),
    .A(net1545),
    .B(_1014_));
 sg13g2_o21ai_1 _5334_ (.B1(_1530_),
    .Y(_0254_),
    .A1(net1545),
    .A2(_1529_));
 sg13g2_nand2_1 _5335_ (.Y(_1531_),
    .A(net1544),
    .B(_1014_));
 sg13g2_xnor2_1 _5336_ (.Y(_1532_),
    .A(net1544),
    .B(\tt6581_inst.controller_inst.cur_voice[0] ));
 sg13g2_xor2_1 _5337_ (.B(net1545),
    .A(net1544),
    .X(_1533_));
 sg13g2_o21ai_1 _5338_ (.B1(_1531_),
    .Y(_0255_),
    .A1(_1529_),
    .A2(net1373));
 sg13g2_nand2_1 _5339_ (.Y(_1534_),
    .A(net216),
    .B(net1546));
 sg13g2_o21ai_1 _5340_ (.B1(_1534_),
    .Y(_0256_),
    .A1(_0876_),
    .A2(net1546));
 sg13g2_nor2_1 _5341_ (.A(net471),
    .B(net1546),
    .Y(_1535_));
 sg13g2_xnor2_1 _5342_ (.Y(_1536_),
    .A(net216),
    .B(_1484_));
 sg13g2_a21oi_1 _5343_ (.A1(net1546),
    .A2(_1536_),
    .Y(_0257_),
    .B1(_1535_));
 sg13g2_nor2_1 _5344_ (.A(_1485_),
    .B(_1489_),
    .Y(_1537_));
 sg13g2_nor3_1 _5345_ (.A(net1432),
    .B(_1490_),
    .C(_1537_),
    .Y(_1538_));
 sg13g2_a21o_1 _5346_ (.A2(net1432),
    .A1(net566),
    .B1(_1538_),
    .X(_0258_));
 sg13g2_nor2_1 _5347_ (.A(net762),
    .B(net1547),
    .Y(_1539_));
 sg13g2_nor2_1 _5348_ (.A(_1488_),
    .B(_1490_),
    .Y(_1540_));
 sg13g2_xnor2_1 _5349_ (.Y(_1541_),
    .A(_1495_),
    .B(_1540_));
 sg13g2_a21oi_1 _5350_ (.A1(net1547),
    .A2(_1541_),
    .Y(_0259_),
    .B1(_1539_));
 sg13g2_and2_1 _5351_ (.A(_1496_),
    .B(_1497_),
    .X(_1542_));
 sg13g2_nor3_1 _5352_ (.A(net1432),
    .B(_1498_),
    .C(_1542_),
    .Y(_1543_));
 sg13g2_a21o_1 _5353_ (.A2(net1432),
    .A1(net960),
    .B1(_1543_),
    .X(_0260_));
 sg13g2_nor3_1 _5354_ (.A(_1482_),
    .B(_1498_),
    .C(_1499_),
    .Y(_1544_));
 sg13g2_nand2_1 _5355_ (.Y(_1545_),
    .A(net479),
    .B(net1432));
 sg13g2_nand2_1 _5356_ (.Y(_1546_),
    .A(net1547),
    .B(_1500_));
 sg13g2_o21ai_1 _5357_ (.B1(_1545_),
    .Y(_0261_),
    .A1(_1544_),
    .A2(_1546_));
 sg13g2_and3_1 _5358_ (.X(_1547_),
    .A(_1479_),
    .B(_1500_),
    .C(_1501_));
 sg13g2_nor3_1 _5359_ (.A(net1432),
    .B(_1502_),
    .C(_1547_),
    .Y(_1548_));
 sg13g2_a21o_1 _5360_ (.A2(net1432),
    .A1(net869),
    .B1(_1548_),
    .X(_0262_));
 sg13g2_nor3_1 _5361_ (.A(_1473_),
    .B(_1502_),
    .C(_1503_),
    .Y(_1549_));
 sg13g2_nand2_1 _5362_ (.Y(_1550_),
    .A(net464),
    .B(net1433));
 sg13g2_nand2_1 _5363_ (.Y(_1551_),
    .A(net1548),
    .B(_1504_));
 sg13g2_o21ai_1 _5364_ (.B1(_1550_),
    .Y(_0263_),
    .A1(_1549_),
    .A2(_1551_));
 sg13g2_and3_1 _5365_ (.X(_1552_),
    .A(_1467_),
    .B(_1504_),
    .C(_1505_));
 sg13g2_nor3_1 _5366_ (.A(net1432),
    .B(_1506_),
    .C(_1552_),
    .Y(_1553_));
 sg13g2_a21o_1 _5367_ (.A2(net1433),
    .A1(net901),
    .B1(_1553_),
    .X(_0264_));
 sg13g2_nor3_1 _5368_ (.A(_1461_),
    .B(_1506_),
    .C(_1507_),
    .Y(_1554_));
 sg13g2_nand2_1 _5369_ (.Y(_1555_),
    .A(net280),
    .B(net1433));
 sg13g2_nand2_1 _5370_ (.Y(_1556_),
    .A(net1548),
    .B(_1508_));
 sg13g2_o21ai_1 _5371_ (.B1(_1555_),
    .Y(_0265_),
    .A1(_1554_),
    .A2(_1556_));
 sg13g2_and3_1 _5372_ (.X(_1557_),
    .A(_1455_),
    .B(_1508_),
    .C(_1509_));
 sg13g2_nor3_1 _5373_ (.A(_0998_),
    .B(_1510_),
    .C(_1557_),
    .Y(_1558_));
 sg13g2_a21o_1 _5374_ (.A2(_0998_),
    .A1(net838),
    .B1(_1558_),
    .X(_0266_));
 sg13g2_nor3_1 _5375_ (.A(_1449_),
    .B(_1510_),
    .C(_1511_),
    .Y(_1559_));
 sg13g2_nand2_1 _5376_ (.Y(_1560_),
    .A(net285),
    .B(net1433));
 sg13g2_nand2_1 _5377_ (.Y(_1561_),
    .A(net1551),
    .B(_1512_));
 sg13g2_o21ai_1 _5378_ (.B1(_1560_),
    .Y(_0267_),
    .A1(_1559_),
    .A2(_1561_));
 sg13g2_and3_1 _5379_ (.X(_1562_),
    .A(_1443_),
    .B(_1512_),
    .C(_1513_));
 sg13g2_nor3_1 _5380_ (.A(net1433),
    .B(_1514_),
    .C(_1562_),
    .Y(_1563_));
 sg13g2_a21o_1 _5381_ (.A2(net1433),
    .A1(net979),
    .B1(_1563_),
    .X(_0268_));
 sg13g2_nor2_1 _5382_ (.A(net515),
    .B(net1551),
    .Y(_1564_));
 sg13g2_nor2b_1 _5383_ (.A(_1431_),
    .B_N(_1432_),
    .Y(_1565_));
 sg13g2_xnor2_1 _5384_ (.Y(_1566_),
    .A(_1515_),
    .B(_1565_));
 sg13g2_a21oi_1 _5385_ (.A1(net1551),
    .A2(_1566_),
    .Y(_0269_),
    .B1(_1564_));
 sg13g2_xnor2_1 _5386_ (.Y(_1567_),
    .A(_1426_),
    .B(_1517_));
 sg13g2_nor2_1 _5387_ (.A(net656),
    .B(net1551),
    .Y(_1568_));
 sg13g2_a21oi_1 _5388_ (.A1(net1551),
    .A2(_1567_),
    .Y(_0270_),
    .B1(_1568_));
 sg13g2_nand2_1 _5389_ (.Y(_1569_),
    .A(_1417_),
    .B(_1418_));
 sg13g2_xnor2_1 _5390_ (.Y(_1570_),
    .A(_1518_),
    .B(_1569_));
 sg13g2_nor2_1 _5391_ (.A(net470),
    .B(net1549),
    .Y(_1571_));
 sg13g2_a21oi_1 _5392_ (.A1(net1549),
    .A2(_1570_),
    .Y(_0271_),
    .B1(_1571_));
 sg13g2_xor2_1 _5393_ (.B(_1519_),
    .A(_1412_),
    .X(_1572_));
 sg13g2_xnor2_1 _5394_ (.Y(_1573_),
    .A(_1528_),
    .B(_1572_));
 sg13g2_nor2b_1 _5395_ (.A(_1573_),
    .B_N(_1570_),
    .Y(_1574_));
 sg13g2_xor2_1 _5396_ (.B(_1573_),
    .A(_1570_),
    .X(_1575_));
 sg13g2_nor2_1 _5397_ (.A(net791),
    .B(net1549),
    .Y(_1576_));
 sg13g2_a21oi_1 _5398_ (.A1(net1549),
    .A2(_1575_),
    .Y(_0272_),
    .B1(_1576_));
 sg13g2_a21o_1 _5399_ (.A2(_1572_),
    .A1(_1528_),
    .B1(_1574_),
    .X(_1577_));
 sg13g2_nand3_1 _5400_ (.B(_1411_),
    .C(_1520_),
    .A(_1405_),
    .Y(_1578_));
 sg13g2_nand2b_1 _5401_ (.Y(_1579_),
    .B(_1578_),
    .A_N(_1521_));
 sg13g2_nand2b_1 _5402_ (.Y(_1580_),
    .B(_1528_),
    .A_N(_1579_));
 sg13g2_xnor2_1 _5403_ (.Y(_1581_),
    .A(_1528_),
    .B(_1579_));
 sg13g2_a21oi_1 _5404_ (.A1(_1577_),
    .A2(_1581_),
    .Y(_1582_),
    .B1(net1433));
 sg13g2_o21ai_1 _5405_ (.B1(_1582_),
    .Y(_1583_),
    .A1(_1577_),
    .A2(_1581_));
 sg13g2_o21ai_1 _5406_ (.B1(_1583_),
    .Y(_0273_),
    .A1(_0882_),
    .A2(net1550));
 sg13g2_nand2_1 _5407_ (.Y(_1584_),
    .A(_1580_),
    .B(_1582_));
 sg13g2_o21ai_1 _5408_ (.B1(_1584_),
    .Y(_0274_),
    .A1(net1550),
    .A2(_0999_));
 sg13g2_nor2_1 _5409_ (.A(net216),
    .B(net1546),
    .Y(_1585_));
 sg13g2_a21oi_1 _5410_ (.A1(_0876_),
    .A2(net1546),
    .Y(_0275_),
    .B1(_1585_));
 sg13g2_mux2_1 _5411_ (.A0(net781),
    .A1(net471),
    .S(net1547),
    .X(_0276_));
 sg13g2_mux2_1 _5412_ (.A0(net657),
    .A1(net566),
    .S(net1546),
    .X(_0277_));
 sg13g2_mux2_1 _5413_ (.A0(net711),
    .A1(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .S(net1546),
    .X(_0278_));
 sg13g2_mux2_1 _5414_ (.A0(net970),
    .A1(net960),
    .S(net1547),
    .X(_0279_));
 sg13g2_mux2_1 _5415_ (.A0(net945),
    .A1(net479),
    .S(net1548),
    .X(_0280_));
 sg13g2_mux2_1 _5416_ (.A0(net667),
    .A1(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .S(net1548),
    .X(_0281_));
 sg13g2_mux2_1 _5417_ (.A0(net603),
    .A1(net464),
    .S(net1548),
    .X(_0282_));
 sg13g2_mux2_1 _5418_ (.A0(net686),
    .A1(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .S(net1548),
    .X(_0283_));
 sg13g2_mux2_1 _5419_ (.A0(net801),
    .A1(net280),
    .S(net1548),
    .X(_0284_));
 sg13g2_mux2_1 _5420_ (.A0(net910),
    .A1(net838),
    .S(net1551),
    .X(_0285_));
 sg13g2_mux2_1 _5421_ (.A0(net675),
    .A1(net285),
    .S(net1551),
    .X(_0286_));
 sg13g2_mux2_1 _5422_ (.A0(net672),
    .A1(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .S(net1550),
    .X(_0287_));
 sg13g2_mux2_1 _5423_ (.A0(net947),
    .A1(net515),
    .S(net1550),
    .X(_0288_));
 sg13g2_mux2_1 _5424_ (.A0(net870),
    .A1(net656),
    .S(net1551),
    .X(_0289_));
 sg13g2_mux2_1 _5425_ (.A0(net875),
    .A1(net470),
    .S(net1549),
    .X(_0290_));
 sg13g2_mux2_1 _5426_ (.A0(net889),
    .A1(net791),
    .S(net1549),
    .X(_0291_));
 sg13g2_nor2_1 _5427_ (.A(net424),
    .B(net1549),
    .Y(_1586_));
 sg13g2_a21oi_1 _5428_ (.A1(_0882_),
    .A2(net1550),
    .Y(_0292_),
    .B1(_1586_));
 sg13g2_nor2_1 _5429_ (.A(\tt6581_inst.delta_sigma_inst.e2[18] ),
    .B(net1550),
    .Y(_1587_));
 sg13g2_a21oi_1 _5430_ (.A1(net1550),
    .A2(_0999_),
    .Y(_0293_),
    .B1(_1587_));
 sg13g2_nor2_1 _5431_ (.A(net169),
    .B(net1290),
    .Y(_1588_));
 sg13g2_a21oi_1 _5432_ (.A1(net169),
    .A2(net1192),
    .Y(_0294_),
    .B1(_1588_));
 sg13g2_xor2_1 _5433_ (.B(net169),
    .A(net1069),
    .X(_1589_));
 sg13g2_a22oi_1 _5434_ (.Y(_1590_),
    .B1(_1589_),
    .B2(net1537),
    .A2(net1224),
    .A1(net1069));
 sg13g2_inv_1 _5435_ (.Y(_0295_),
    .A(_1590_));
 sg13g2_a21oi_1 _5436_ (.A1(\tt6581_inst.mult_inst.iter[1] ),
    .A2(net169),
    .Y(_1591_),
    .B1(net881));
 sg13g2_nand3_1 _5437_ (.B(net169),
    .C(net881),
    .A(\tt6581_inst.mult_inst.iter[1] ),
    .Y(_1592_));
 sg13g2_nor2b_1 _5438_ (.A(_1591_),
    .B_N(_1592_),
    .Y(_1593_));
 sg13g2_a22oi_1 _5439_ (.Y(_1594_),
    .B1(_1593_),
    .B2(net1290),
    .A2(net1224),
    .A1(net881));
 sg13g2_inv_1 _5440_ (.Y(_0296_),
    .A(net882));
 sg13g2_xnor2_1 _5441_ (.Y(_1595_),
    .A(net967),
    .B(_1592_));
 sg13g2_a22oi_1 _5442_ (.Y(_1596_),
    .B1(_1595_),
    .B2(net1290),
    .A2(net1224),
    .A1(net967));
 sg13g2_inv_1 _5443_ (.Y(_0297_),
    .A(net968));
 sg13g2_nor3_1 _5444_ (.A(_0880_),
    .B(net1225),
    .C(_1592_),
    .Y(_1597_));
 sg13g2_o21ai_1 _5445_ (.B1(_1019_),
    .Y(_1598_),
    .A1(net65),
    .A2(_1597_));
 sg13g2_a21oi_1 _5446_ (.A1(net65),
    .A2(_1597_),
    .Y(_0298_),
    .B1(_1598_));
 sg13g2_nand2_1 _5447_ (.Y(_1599_),
    .A(\tt6581_inst.control_pack[13] ),
    .B(net1397));
 sg13g2_a22oi_1 _5448_ (.Y(_1600_),
    .B1(net1376),
    .B2(\tt6581_inst.control_pack[5] ),
    .A2(net1420),
    .A1(\tt6581_inst.control_pack[21] ));
 sg13g2_and2_1 _5449_ (.A(_1599_),
    .B(_1600_),
    .X(_1601_));
 sg13g2_nand2_1 _5450_ (.Y(_1602_),
    .A(_1599_),
    .B(_1600_));
 sg13g2_and2_1 _5451_ (.A(\tt6581_inst.control_pack[12] ),
    .B(net1399),
    .X(_1603_));
 sg13g2_a221oi_1 _5452_ (.B2(\tt6581_inst.control_pack[4] ),
    .C1(_1603_),
    .B1(net1376),
    .A1(\tt6581_inst.control_pack[20] ),
    .Y(_1604_),
    .A2(net1420));
 sg13g2_a22oi_1 _5453_ (.Y(_1605_),
    .B1(net1376),
    .B2(\tt6581_inst.control_pack[7] ),
    .A2(net1418),
    .A1(\tt6581_inst.control_pack[23] ));
 sg13g2_o21ai_1 _5454_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_0971_),
    .A2(net1391));
 sg13g2_a22oi_1 _5455_ (.Y(_1607_),
    .B1(net1376),
    .B2(\tt6581_inst.control_pack[6] ),
    .A2(net1420),
    .A1(\tt6581_inst.control_pack[22] ));
 sg13g2_o21ai_1 _5456_ (.B1(_1607_),
    .Y(_1608_),
    .A1(_0970_),
    .A2(net1390));
 sg13g2_nand3_1 _5457_ (.B(_1604_),
    .C(_1606_),
    .A(_1601_),
    .Y(_1609_));
 sg13g2_nor2_2 _5458_ (.A(_1608_),
    .B(_1609_),
    .Y(_1610_));
 sg13g2_nor2_1 _5459_ (.A(_1606_),
    .B(_1608_),
    .Y(_1611_));
 sg13g2_and3_2 _5460_ (.X(_1612_),
    .A(_1602_),
    .B(_1604_),
    .C(_1611_));
 sg13g2_nand3_1 _5461_ (.B(_1604_),
    .C(_1611_),
    .A(_1602_),
    .Y(_1613_));
 sg13g2_nor2b_1 _5462_ (.A(_1606_),
    .B_N(_1608_),
    .Y(_1614_));
 sg13g2_nand3_1 _5463_ (.B(_1604_),
    .C(_1614_),
    .A(_1601_),
    .Y(_1615_));
 sg13g2_inv_1 _5464_ (.Y(_1616_),
    .A(net1190));
 sg13g2_nor4_2 _5465_ (.A(_1602_),
    .B(_1604_),
    .C(_1606_),
    .Y(_1617_),
    .D(_1608_));
 sg13g2_nor3_1 _5466_ (.A(_1610_),
    .B(_1612_),
    .C(net1215),
    .Y(_1618_));
 sg13g2_a21oi_2 _5467_ (.B1(net1494),
    .Y(_1619_),
    .A2(_1618_),
    .A1(net1190));
 sg13g2_a21o_2 _5468_ (.A2(_1618_),
    .A1(net1190),
    .B1(net1494),
    .X(_1620_));
 sg13g2_nor2_1 _5469_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][16] ),
    .B(net1369),
    .Y(_1621_));
 sg13g2_nor2_1 _5470_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][16] ),
    .B(net1413),
    .Y(_1622_));
 sg13g2_nor2_1 _5471_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][16] ),
    .B(net1390),
    .Y(_1623_));
 sg13g2_nor3_1 _5472_ (.A(_1621_),
    .B(_1622_),
    .C(_1623_),
    .Y(_1624_));
 sg13g2_a22oi_1 _5473_ (.Y(_1625_),
    .B1(net1377),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[7] ),
    .A2(net1419),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[23] ));
 sg13g2_o21ai_1 _5474_ (.B1(_1625_),
    .Y(_1626_),
    .A1(_0951_),
    .A2(net1390));
 sg13g2_nor2_1 _5475_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][15] ),
    .B(net1369),
    .Y(_1627_));
 sg13g2_nor2_1 _5476_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][15] ),
    .B(net1413),
    .Y(_1628_));
 sg13g2_nor2_1 _5477_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][15] ),
    .B(net1390),
    .Y(_1629_));
 sg13g2_nor3_1 _5478_ (.A(_1627_),
    .B(_1628_),
    .C(_1629_),
    .Y(_1630_));
 sg13g2_nor2_1 _5479_ (.A(_1626_),
    .B(_1630_),
    .Y(_1631_));
 sg13g2_a22oi_1 _5480_ (.Y(_1632_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[6] ),
    .A2(net1419),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[22] ));
 sg13g2_o21ai_1 _5481_ (.B1(_1632_),
    .Y(_1633_),
    .A1(_0952_),
    .A2(net1390));
 sg13g2_nor2_1 _5482_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][14] ),
    .B(net1369),
    .Y(_1634_));
 sg13g2_nor2_1 _5483_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][14] ),
    .B(net1413),
    .Y(_1635_));
 sg13g2_nor2_1 _5484_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][14] ),
    .B(net1390),
    .Y(_1636_));
 sg13g2_nor3_1 _5485_ (.A(_1634_),
    .B(_1635_),
    .C(_1636_),
    .Y(_1637_));
 sg13g2_and2_1 _5486_ (.A(_1633_),
    .B(_1637_),
    .X(_1638_));
 sg13g2_nand2_1 _5487_ (.Y(_1639_),
    .A(_1633_),
    .B(_1637_));
 sg13g2_nand2_1 _5488_ (.Y(_1640_),
    .A(_1626_),
    .B(_1630_));
 sg13g2_and2_1 _5489_ (.A(\tt6581_inst.controller_inst.freq_hi_i[5] ),
    .B(net1378),
    .X(_1641_));
 sg13g2_a221oi_1 _5490_ (.B2(\tt6581_inst.controller_inst.freq_hi_i[13] ),
    .C1(_1641_),
    .B1(net1397),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[21] ),
    .Y(_1642_),
    .A2(net1419));
 sg13g2_a22oi_1 _5491_ (.Y(_1643_),
    .B1(net1374),
    .B2(_0953_),
    .A2(net1393),
    .A1(_0954_));
 sg13g2_o21ai_1 _5492_ (.B1(_1643_),
    .Y(_1644_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][13] ),
    .A2(net1408));
 sg13g2_nor2_1 _5493_ (.A(_1642_),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_nand2_1 _5494_ (.Y(_1646_),
    .A(_1642_),
    .B(_1644_));
 sg13g2_and2_1 _5495_ (.A(\tt6581_inst.controller_inst.freq_hi_i[4] ),
    .B(net1378),
    .X(_1647_));
 sg13g2_a221oi_1 _5496_ (.B2(\tt6581_inst.controller_inst.freq_hi_i[12] ),
    .C1(_1647_),
    .B1(net1398),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[20] ),
    .Y(_1648_),
    .A2(net1420));
 sg13g2_a22oi_1 _5497_ (.Y(_1649_),
    .B1(net1374),
    .B2(_0955_),
    .A2(net1394),
    .A1(_0956_));
 sg13g2_o21ai_1 _5498_ (.B1(_1649_),
    .Y(_1650_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][12] ),
    .A2(net1408));
 sg13g2_nor2_1 _5499_ (.A(_1648_),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_inv_1 _5500_ (.Y(_1652_),
    .A(_1651_));
 sg13g2_a22oi_1 _5501_ (.Y(_1653_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[3] ),
    .A2(net1398),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[11] ));
 sg13g2_o21ai_1 _5502_ (.B1(_1653_),
    .Y(_1654_),
    .A1(_0957_),
    .A2(net1413));
 sg13g2_a22oi_1 _5503_ (.Y(_1655_),
    .B1(net1374),
    .B2(_0958_),
    .A2(net1394),
    .A1(_0959_));
 sg13g2_o21ai_1 _5504_ (.B1(_1655_),
    .Y(_1656_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][11] ),
    .A2(net1408));
 sg13g2_nand2b_1 _5505_ (.Y(_1657_),
    .B(_1654_),
    .A_N(_1656_));
 sg13g2_a22oi_1 _5506_ (.Y(_1658_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[2] ),
    .A2(net1397),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[10] ));
 sg13g2_o21ai_1 _5507_ (.B1(_1658_),
    .Y(_1659_),
    .A1(_0960_),
    .A2(net1413));
 sg13g2_a22oi_1 _5508_ (.Y(_1660_),
    .B1(net1393),
    .B2(_0962_),
    .A2(net1417),
    .A1(_0961_));
 sg13g2_o21ai_1 _5509_ (.B1(_1660_),
    .Y(_1661_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[0][10] ),
    .A2(net1365));
 sg13g2_nor2b_1 _5510_ (.A(_1661_),
    .B_N(_1659_),
    .Y(_1662_));
 sg13g2_inv_1 _5511_ (.Y(_1663_),
    .A(_1662_));
 sg13g2_nand2b_1 _5512_ (.Y(_1664_),
    .B(_1661_),
    .A_N(_1659_));
 sg13g2_nand2_1 _5513_ (.Y(_1665_),
    .A(_1663_),
    .B(_1664_));
 sg13g2_a22oi_1 _5514_ (.Y(_1666_),
    .B1(net1377),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[1] ),
    .A2(net1394),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[9] ));
 sg13g2_o21ai_1 _5515_ (.B1(_1666_),
    .Y(_1667_),
    .A1(_0890_),
    .A2(net1408));
 sg13g2_a22oi_1 _5516_ (.Y(_1668_),
    .B1(net1374),
    .B2(_0891_),
    .A2(net1393),
    .A1(_0892_));
 sg13g2_o21ai_1 _5517_ (.B1(_1668_),
    .Y(_1669_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][9] ),
    .A2(net1407));
 sg13g2_inv_1 _5518_ (.Y(_1670_),
    .A(_1669_));
 sg13g2_nand2b_2 _5519_ (.Y(_1671_),
    .B(_1669_),
    .A_N(_1667_));
 sg13g2_inv_1 _5520_ (.Y(_1672_),
    .A(_1671_));
 sg13g2_a22oi_1 _5521_ (.Y(_1673_),
    .B1(net1377),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[0] ),
    .A2(net1398),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[8] ));
 sg13g2_o21ai_1 _5522_ (.B1(_1673_),
    .Y(_1674_),
    .A1(_0893_),
    .A2(net1409));
 sg13g2_a22oi_1 _5523_ (.Y(_1675_),
    .B1(net1374),
    .B2(_0894_),
    .A2(net1393),
    .A1(_0895_));
 sg13g2_o21ai_1 _5524_ (.B1(_1675_),
    .Y(_1676_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][8] ),
    .A2(net1407));
 sg13g2_nor2b_1 _5525_ (.A(_1676_),
    .B_N(_1674_),
    .Y(_1677_));
 sg13g2_a22oi_1 _5526_ (.Y(_1678_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[7] ),
    .A2(net1395),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[15] ));
 sg13g2_o21ai_1 _5527_ (.B1(_1678_),
    .Y(_1679_),
    .A1(_0896_),
    .A2(net1411));
 sg13g2_nor2_1 _5528_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][7] ),
    .B(net1367),
    .Y(_1680_));
 sg13g2_nor2_1 _5529_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][7] ),
    .B(net1410),
    .Y(_1681_));
 sg13g2_nor2_1 _5530_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][7] ),
    .B(net1388),
    .Y(_1682_));
 sg13g2_nor3_1 _5531_ (.A(_1680_),
    .B(_1681_),
    .C(_1682_),
    .Y(_1683_));
 sg13g2_and2_1 _5532_ (.A(_1679_),
    .B(_1683_),
    .X(_1684_));
 sg13g2_a22oi_1 _5533_ (.Y(_1685_),
    .B1(net1376),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[6] ),
    .A2(net1399),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[14] ));
 sg13g2_o21ai_1 _5534_ (.B1(_1685_),
    .Y(_1686_),
    .A1(_0897_),
    .A2(net1413));
 sg13g2_a22oi_1 _5535_ (.Y(_1687_),
    .B1(net1374),
    .B2(_0898_),
    .A2(net1395),
    .A1(_0899_));
 sg13g2_o21ai_1 _5536_ (.B1(_1687_),
    .Y(_1688_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[2][6] ),
    .A2(net1410));
 sg13g2_nor2b_1 _5537_ (.A(_1688_),
    .B_N(_1686_),
    .Y(_1689_));
 sg13g2_a22oi_1 _5538_ (.Y(_1690_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[5] ),
    .A2(net1395),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[13] ));
 sg13g2_o21ai_1 _5539_ (.B1(_1690_),
    .Y(_1691_),
    .A1(_0900_),
    .A2(net1411));
 sg13g2_nor2_1 _5540_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][5] ),
    .B(net1367),
    .Y(_1692_));
 sg13g2_nor2_1 _5541_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][5] ),
    .B(net1410),
    .Y(_1693_));
 sg13g2_nor2_1 _5542_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][5] ),
    .B(net1388),
    .Y(_1694_));
 sg13g2_nor3_1 _5543_ (.A(_1692_),
    .B(_1693_),
    .C(_1694_),
    .Y(_1695_));
 sg13g2_nand2_1 _5544_ (.Y(_1696_),
    .A(_1691_),
    .B(_1695_));
 sg13g2_a22oi_1 _5545_ (.Y(_1697_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[4] ),
    .A2(net1395),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[12] ));
 sg13g2_o21ai_1 _5546_ (.B1(_1697_),
    .Y(_1698_),
    .A1(_0901_),
    .A2(net1411));
 sg13g2_nor2_1 _5547_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][4] ),
    .B(net1367),
    .Y(_1699_));
 sg13g2_nor2_1 _5548_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][4] ),
    .B(net1410),
    .Y(_1700_));
 sg13g2_nor2_1 _5549_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][4] ),
    .B(net1388),
    .Y(_1701_));
 sg13g2_nor3_1 _5550_ (.A(_1699_),
    .B(_1700_),
    .C(_1701_),
    .Y(_1702_));
 sg13g2_and2_1 _5551_ (.A(_1698_),
    .B(_1702_),
    .X(_1703_));
 sg13g2_nor2_1 _5552_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][3] ),
    .B(net1367),
    .Y(_1704_));
 sg13g2_nor2_1 _5553_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][3] ),
    .B(net1410),
    .Y(_1705_));
 sg13g2_nor2_1 _5554_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][3] ),
    .B(net1388),
    .Y(_1706_));
 sg13g2_nor3_1 _5555_ (.A(_1704_),
    .B(_1705_),
    .C(_1706_),
    .Y(_1707_));
 sg13g2_a22oi_1 _5556_ (.Y(_1708_),
    .B1(net1379),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[3] ),
    .A2(net1399),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[11] ));
 sg13g2_o21ai_1 _5557_ (.B1(_1708_),
    .Y(_1709_),
    .A1(_0902_),
    .A2(net1414));
 sg13g2_nand2_1 _5558_ (.Y(_1710_),
    .A(_1707_),
    .B(_1709_));
 sg13g2_a22oi_1 _5559_ (.Y(_1711_),
    .B1(net1379),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[2] ),
    .A2(net1399),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[10] ));
 sg13g2_o21ai_1 _5560_ (.B1(_1711_),
    .Y(_1712_),
    .A1(_0903_),
    .A2(net1414));
 sg13g2_nor2_1 _5561_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][2] ),
    .B(net1368),
    .Y(_1713_));
 sg13g2_nor2_1 _5562_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][2] ),
    .B(net1412),
    .Y(_1714_));
 sg13g2_nor2_1 _5563_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][2] ),
    .B(net1389),
    .Y(_1715_));
 sg13g2_nor3_1 _5564_ (.A(_1713_),
    .B(_1714_),
    .C(_1715_),
    .Y(_1716_));
 sg13g2_and2_1 _5565_ (.A(_1712_),
    .B(_1716_),
    .X(_1717_));
 sg13g2_a22oi_1 _5566_ (.Y(_1718_),
    .B1(net1379),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[1] ),
    .A2(net1399),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[9] ));
 sg13g2_o21ai_1 _5567_ (.B1(_1718_),
    .Y(_1719_),
    .A1(_0904_),
    .A2(net1411));
 sg13g2_a22oi_1 _5568_ (.Y(_1720_),
    .B1(net1396),
    .B2(_0906_),
    .A2(net1418),
    .A1(_0905_));
 sg13g2_o21ai_1 _5569_ (.B1(_1720_),
    .Y(_1721_),
    .A1(\tt6581_inst.multi_voice_inst.phase_regs[0][1] ),
    .A2(net1368));
 sg13g2_nand2b_1 _5570_ (.Y(_1722_),
    .B(_1719_),
    .A_N(_1721_));
 sg13g2_a22oi_1 _5571_ (.Y(_1723_),
    .B1(net1376),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[0] ),
    .A2(net1418),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[16] ));
 sg13g2_o21ai_1 _5572_ (.B1(_1723_),
    .Y(_1724_),
    .A1(_0907_),
    .A2(net1389));
 sg13g2_nor2_1 _5573_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][0] ),
    .B(net1368),
    .Y(_1725_));
 sg13g2_nor2_1 _5574_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][0] ),
    .B(net1412),
    .Y(_1726_));
 sg13g2_nor2_1 _5575_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][0] ),
    .B(net1389),
    .Y(_1727_));
 sg13g2_nor3_1 _5576_ (.A(_1725_),
    .B(_1726_),
    .C(_1727_),
    .Y(_1728_));
 sg13g2_nand2_1 _5577_ (.Y(_1729_),
    .A(_1724_),
    .B(_1728_));
 sg13g2_xor2_1 _5578_ (.B(_1721_),
    .A(_1719_),
    .X(_1730_));
 sg13g2_o21ai_1 _5579_ (.B1(_1722_),
    .Y(_1731_),
    .A1(_1729_),
    .A2(_1730_));
 sg13g2_or2_1 _5580_ (.X(_1732_),
    .B(_1716_),
    .A(_1712_));
 sg13g2_nand2b_1 _5581_ (.Y(_1733_),
    .B(_1732_),
    .A_N(_1717_));
 sg13g2_a21oi_1 _5582_ (.A1(_1731_),
    .A2(_1732_),
    .Y(_1734_),
    .B1(_1717_));
 sg13g2_nor2_1 _5583_ (.A(_1707_),
    .B(_1709_),
    .Y(_1735_));
 sg13g2_xor2_1 _5584_ (.B(_1709_),
    .A(_1707_),
    .X(_1736_));
 sg13g2_nand2b_1 _5585_ (.Y(_1737_),
    .B(_1736_),
    .A_N(_1734_));
 sg13g2_o21ai_1 _5586_ (.B1(_1710_),
    .Y(_1738_),
    .A1(_1734_),
    .A2(_1735_));
 sg13g2_or2_1 _5587_ (.X(_1739_),
    .B(_1702_),
    .A(_1698_));
 sg13g2_nand2b_1 _5588_ (.Y(_1740_),
    .B(_1739_),
    .A_N(_1703_));
 sg13g2_a21oi_1 _5589_ (.A1(_1738_),
    .A2(_1739_),
    .Y(_1741_),
    .B1(_1703_));
 sg13g2_nor2_1 _5590_ (.A(_1691_),
    .B(_1695_),
    .Y(_1742_));
 sg13g2_xor2_1 _5591_ (.B(_1695_),
    .A(_1691_),
    .X(_1743_));
 sg13g2_nand2b_1 _5592_ (.Y(_1744_),
    .B(_1743_),
    .A_N(_1741_));
 sg13g2_o21ai_1 _5593_ (.B1(_1696_),
    .Y(_1745_),
    .A1(_1741_),
    .A2(_1742_));
 sg13g2_xor2_1 _5594_ (.B(_1688_),
    .A(_1686_),
    .X(_1746_));
 sg13g2_inv_1 _5595_ (.Y(_1747_),
    .A(_1746_));
 sg13g2_a21o_2 _5596_ (.A2(_1747_),
    .A1(_1745_),
    .B1(_1689_),
    .X(_1748_));
 sg13g2_or2_1 _5597_ (.X(_1749_),
    .B(_1683_),
    .A(_1679_));
 sg13g2_nor2b_1 _5598_ (.A(_1684_),
    .B_N(_1749_),
    .Y(_1750_));
 sg13g2_a21o_2 _5599_ (.A2(_1749_),
    .A1(_1748_),
    .B1(_1684_),
    .X(_1751_));
 sg13g2_xnor2_1 _5600_ (.Y(_1752_),
    .A(_1674_),
    .B(_1676_));
 sg13g2_a21o_1 _5601_ (.A2(_1752_),
    .A1(_1751_),
    .B1(_1677_),
    .X(_1753_));
 sg13g2_nand2_1 _5602_ (.Y(_1754_),
    .A(_1667_),
    .B(_1670_));
 sg13g2_inv_1 _5603_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_a221oi_1 _5604_ (.B2(_1752_),
    .C1(_1677_),
    .B1(_1751_),
    .A1(_1667_),
    .Y(_1756_),
    .A2(_1670_));
 sg13g2_nor3_1 _5605_ (.A(_1665_),
    .B(_1672_),
    .C(_1756_),
    .Y(_1757_));
 sg13g2_xnor2_1 _5606_ (.Y(_1758_),
    .A(_1654_),
    .B(_1656_));
 sg13g2_o21ai_1 _5607_ (.B1(_1758_),
    .Y(_1759_),
    .A1(_1662_),
    .A2(_1757_));
 sg13g2_xnor2_1 _5608_ (.Y(_1760_),
    .A(_1648_),
    .B(_1650_));
 sg13g2_a21o_2 _5609_ (.A2(_1759_),
    .A1(_1657_),
    .B1(_1760_),
    .X(_1761_));
 sg13g2_nor2_1 _5610_ (.A(_1645_),
    .B(_1651_),
    .Y(_1762_));
 sg13g2_a22oi_1 _5611_ (.Y(_1763_),
    .B1(_1761_),
    .B2(_1762_),
    .A2(_1644_),
    .A1(_1642_));
 sg13g2_xnor2_1 _5612_ (.Y(_1764_),
    .A(_1633_),
    .B(_1637_));
 sg13g2_a221oi_1 _5613_ (.B2(_1762_),
    .C1(_1764_),
    .B1(_1761_),
    .A1(_1642_),
    .Y(_1765_),
    .A2(_1644_));
 sg13g2_a21oi_1 _5614_ (.A1(_1639_),
    .A2(_1640_),
    .Y(_1766_),
    .B1(_1631_));
 sg13g2_nand2b_1 _5615_ (.Y(_1767_),
    .B(_1640_),
    .A_N(_1631_));
 sg13g2_inv_1 _5616_ (.Y(_1768_),
    .A(_1767_));
 sg13g2_or2_1 _5617_ (.X(_1769_),
    .B(_1767_),
    .A(_1764_));
 sg13g2_a221oi_1 _5618_ (.B2(_1762_),
    .C1(_1769_),
    .B1(_1761_),
    .A1(_1642_),
    .Y(_1770_),
    .A2(_1644_));
 sg13g2_nor3_1 _5619_ (.A(_1624_),
    .B(_1766_),
    .C(_1770_),
    .Y(_1771_));
 sg13g2_nor2_1 _5620_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[2][0] ),
    .B(net1365),
    .Y(_1772_));
 sg13g2_nor2_1 _5621_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[1][0] ),
    .B(net1407),
    .Y(_1773_));
 sg13g2_nor2_1 _5622_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[0][0] ),
    .B(net1386),
    .Y(_1774_));
 sg13g2_nor3_2 _5623_ (.A(_1772_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1775_));
 sg13g2_a22oi_1 _5624_ (.Y(_1776_),
    .B1(net1374),
    .B2(\tt6581_inst.multi_voice_inst.phase_last_msb[2][1] ),
    .A2(net1393),
    .A1(\tt6581_inst.multi_voice_inst.phase_last_msb[0][1] ));
 sg13g2_inv_1 _5625_ (.Y(_1777_),
    .A(_1776_));
 sg13g2_nand2_1 _5626_ (.Y(_1778_),
    .A(\tt6581_inst.control_pack[9] ),
    .B(net1394));
 sg13g2_a22oi_1 _5627_ (.Y(_1779_),
    .B1(net1375),
    .B2(\tt6581_inst.control_pack[1] ),
    .A2(net1418),
    .A1(\tt6581_inst.control_pack[17] ));
 sg13g2_a221oi_1 _5628_ (.B2(_1779_),
    .C1(_1777_),
    .B1(_1778_),
    .A1(\tt6581_inst.multi_voice_inst.phase_last_msb[1][1] ),
    .Y(_1780_),
    .A2(net1417));
 sg13g2_and2_1 _5629_ (.A(_1775_),
    .B(_1780_),
    .X(_1781_));
 sg13g2_nand2_2 _5630_ (.Y(_1782_),
    .A(_1775_),
    .B(_1780_));
 sg13g2_o21ai_1 _5631_ (.B1(_1624_),
    .Y(_1783_),
    .A1(_1766_),
    .A2(_1770_));
 sg13g2_nand2_1 _5632_ (.Y(_1784_),
    .A(net1188),
    .B(_1783_));
 sg13g2_nor2_2 _5633_ (.A(_1771_),
    .B(_1784_),
    .Y(_1785_));
 sg13g2_and2_1 _5634_ (.A(\tt6581_inst.controller_inst.pw_hi_i[1] ),
    .B(net1376),
    .X(_1786_));
 sg13g2_a221oi_1 _5635_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[9] ),
    .C1(_1786_),
    .B1(net1397),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[17] ),
    .Y(_1787_),
    .A2(net1419));
 sg13g2_nand2_1 _5636_ (.Y(_1788_),
    .A(_1785_),
    .B(_1787_));
 sg13g2_a22oi_1 _5637_ (.Y(_1789_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[0] ),
    .A2(net1419),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[16] ));
 sg13g2_o21ai_1 _5638_ (.B1(_1789_),
    .Y(_1790_),
    .A1(_0964_),
    .A2(net1391));
 sg13g2_or3_1 _5639_ (.A(_1638_),
    .B(_1765_),
    .C(_1768_),
    .X(_1791_));
 sg13g2_o21ai_1 _5640_ (.B1(_1768_),
    .Y(_1792_),
    .A1(_1638_),
    .A2(_1765_));
 sg13g2_and3_1 _5641_ (.X(_1793_),
    .A(net1189),
    .B(_1791_),
    .C(_1792_));
 sg13g2_nand3_1 _5642_ (.B(_1791_),
    .C(_1792_),
    .A(net1188),
    .Y(_1794_));
 sg13g2_nor2_1 _5643_ (.A(_1790_),
    .B(_1794_),
    .Y(_1795_));
 sg13g2_nand2b_1 _5644_ (.Y(_1796_),
    .B(_1764_),
    .A_N(_1763_));
 sg13g2_nand3b_1 _5645_ (.B(net1188),
    .C(_1796_),
    .Y(_1797_),
    .A_N(_1765_));
 sg13g2_a22oi_1 _5646_ (.Y(_1798_),
    .B1(net1377),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[7] ),
    .A2(net1417),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[23] ));
 sg13g2_o21ai_1 _5647_ (.B1(_1798_),
    .Y(_1799_),
    .A1(_0965_),
    .A2(net1391));
 sg13g2_nor2_1 _5648_ (.A(_1797_),
    .B(_1799_),
    .Y(_1800_));
 sg13g2_nand2b_1 _5649_ (.Y(_1801_),
    .B(_1646_),
    .A_N(_1645_));
 sg13g2_a21o_1 _5650_ (.A2(_1761_),
    .A1(_1652_),
    .B1(_1801_),
    .X(_1802_));
 sg13g2_nand3_1 _5651_ (.B(_1761_),
    .C(_1801_),
    .A(_1652_),
    .Y(_1803_));
 sg13g2_nand3_1 _5652_ (.B(_1802_),
    .C(_1803_),
    .A(net1188),
    .Y(_1804_));
 sg13g2_a22oi_1 _5653_ (.Y(_1805_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[6] ),
    .A2(net1397),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[14] ));
 sg13g2_o21ai_1 _5654_ (.B1(_1805_),
    .Y(_1806_),
    .A1(_0966_),
    .A2(net1413));
 sg13g2_and2_1 _5655_ (.A(_1804_),
    .B(_1806_),
    .X(_1807_));
 sg13g2_or2_1 _5656_ (.X(_1808_),
    .B(_1806_),
    .A(_1804_));
 sg13g2_nand3_1 _5657_ (.B(_1759_),
    .C(_1760_),
    .A(_1657_),
    .Y(_1809_));
 sg13g2_nand3_1 _5658_ (.B(net1188),
    .C(_1809_),
    .A(_1761_),
    .Y(_1810_));
 sg13g2_a22oi_1 _5659_ (.Y(_1811_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[5] ),
    .A2(net1418),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[21] ));
 sg13g2_o21ai_1 _5660_ (.B1(_1811_),
    .Y(_1812_),
    .A1(_0967_),
    .A2(net1387));
 sg13g2_nor2_1 _5661_ (.A(_1810_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_nand2_1 _5662_ (.Y(_1814_),
    .A(_1810_),
    .B(_1812_));
 sg13g2_or3_1 _5663_ (.A(_1662_),
    .B(_1757_),
    .C(_1758_),
    .X(_1815_));
 sg13g2_nand3_1 _5664_ (.B(net1188),
    .C(_1815_),
    .A(_1759_),
    .Y(_1816_));
 sg13g2_a22oi_1 _5665_ (.Y(_1817_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[4] ),
    .A2(net1393),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[12] ));
 sg13g2_o21ai_1 _5666_ (.B1(_1817_),
    .Y(_1818_),
    .A1(_0968_),
    .A2(net1411));
 sg13g2_nand2_1 _5667_ (.Y(_1819_),
    .A(_1816_),
    .B(_1818_));
 sg13g2_nor2_1 _5668_ (.A(_1816_),
    .B(_1818_),
    .Y(_1820_));
 sg13g2_a221oi_1 _5669_ (.B2(_1753_),
    .C1(_1755_),
    .B1(_1671_),
    .A1(_1663_),
    .Y(_1821_),
    .A2(_1664_));
 sg13g2_nor3_2 _5670_ (.A(_1757_),
    .B(_1781_),
    .C(_1821_),
    .Y(_1822_));
 sg13g2_and2_1 _5671_ (.A(\tt6581_inst.controller_inst.pw_lo_i[3] ),
    .B(net1379),
    .X(_1823_));
 sg13g2_a221oi_1 _5672_ (.B2(\tt6581_inst.controller_inst.pw_lo_i[11] ),
    .C1(_1823_),
    .B1(net1397),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[19] ),
    .Y(_1824_),
    .A2(net1420));
 sg13g2_and2_1 _5673_ (.A(_1822_),
    .B(_1824_),
    .X(_1825_));
 sg13g2_or2_1 _5674_ (.X(_1826_),
    .B(_1824_),
    .A(_1822_));
 sg13g2_a21oi_1 _5675_ (.A1(_1751_),
    .A2(_1752_),
    .Y(_1827_),
    .B1(_1781_));
 sg13g2_o21ai_1 _5676_ (.B1(_1827_),
    .Y(_1828_),
    .A1(_1751_),
    .A2(_1752_));
 sg13g2_and2_1 _5677_ (.A(\tt6581_inst.controller_inst.pw_lo_i[9] ),
    .B(net1394),
    .X(_1829_));
 sg13g2_a221oi_1 _5678_ (.B2(\tt6581_inst.controller_inst.pw_lo_i[1] ),
    .C1(_1829_),
    .B1(net1375),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[17] ),
    .Y(_1830_),
    .A2(net1417));
 sg13g2_inv_1 _5679_ (.Y(_1831_),
    .A(_1830_));
 sg13g2_a21oi_1 _5680_ (.A1(_1748_),
    .A2(_1750_),
    .Y(_1832_),
    .B1(_1781_));
 sg13g2_o21ai_1 _5681_ (.B1(_1832_),
    .Y(_1833_),
    .A1(_1748_),
    .A2(_1750_));
 sg13g2_a22oi_1 _5682_ (.Y(_1834_),
    .B1(net1375),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[0] ),
    .A2(net1395),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[8] ));
 sg13g2_o21ai_1 _5683_ (.B1(_1834_),
    .Y(_1835_),
    .A1(_0969_),
    .A2(net1411));
 sg13g2_a21o_1 _5684_ (.A2(_1835_),
    .A1(_1833_),
    .B1(_1831_),
    .X(_1836_));
 sg13g2_and3_1 _5685_ (.X(_1837_),
    .A(_1831_),
    .B(_1833_),
    .C(_1835_));
 sg13g2_a21o_1 _5686_ (.A2(_1836_),
    .A1(_1828_),
    .B1(_1837_),
    .X(_1838_));
 sg13g2_a221oi_1 _5687_ (.B2(_1671_),
    .C1(_1677_),
    .B1(_1754_),
    .A1(_1751_),
    .Y(_1839_),
    .A2(_1752_));
 sg13g2_nand3_1 _5688_ (.B(_1753_),
    .C(_1754_),
    .A(_1671_),
    .Y(_1840_));
 sg13g2_nor2_2 _5689_ (.A(_1781_),
    .B(_1839_),
    .Y(_1841_));
 sg13g2_nand2_2 _5690_ (.Y(_1842_),
    .A(_1840_),
    .B(_1841_));
 sg13g2_and2_1 _5691_ (.A(\tt6581_inst.controller_inst.pw_lo_i[18] ),
    .B(net1420),
    .X(_1843_));
 sg13g2_a221oi_1 _5692_ (.B2(\tt6581_inst.controller_inst.pw_lo_i[2] ),
    .C1(_1843_),
    .B1(net1379),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[10] ),
    .Y(_1844_),
    .A2(net1397));
 sg13g2_a21oi_1 _5693_ (.A1(_1840_),
    .A2(_1841_),
    .Y(_1845_),
    .B1(_1844_));
 sg13g2_nand3_1 _5694_ (.B(_1841_),
    .C(_1844_),
    .A(_1840_),
    .Y(_1846_));
 sg13g2_o21ai_1 _5695_ (.B1(_1846_),
    .Y(_1847_),
    .A1(_1838_),
    .A2(_1845_));
 sg13g2_a21o_1 _5696_ (.A2(_1847_),
    .A1(_1826_),
    .B1(_1825_),
    .X(_1848_));
 sg13g2_a21o_1 _5697_ (.A2(_1848_),
    .A1(_1819_),
    .B1(_1820_),
    .X(_1849_));
 sg13g2_a21oi_1 _5698_ (.A1(_1814_),
    .A2(_1849_),
    .Y(_1850_),
    .B1(_1813_));
 sg13g2_a221oi_1 _5699_ (.B2(_1850_),
    .C1(_1807_),
    .B1(_1808_),
    .A1(_1797_),
    .Y(_1851_),
    .A2(_1799_));
 sg13g2_nor3_1 _5700_ (.A(_1795_),
    .B(_1800_),
    .C(_1851_),
    .Y(_1852_));
 sg13g2_nand2_1 _5701_ (.Y(_1853_),
    .A(_1790_),
    .B(_1794_));
 sg13g2_o21ai_1 _5702_ (.B1(_1853_),
    .Y(_1854_),
    .A1(_1785_),
    .A2(_1787_));
 sg13g2_o21ai_1 _5703_ (.B1(_1788_),
    .Y(_1855_),
    .A1(_1852_),
    .A2(_1854_));
 sg13g2_nor2_1 _5704_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][17] ),
    .B(net1365),
    .Y(_1856_));
 sg13g2_nor2_1 _5705_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][17] ),
    .B(net1407),
    .Y(_1857_));
 sg13g2_nor2_1 _5706_ (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][17] ),
    .B(net1386),
    .Y(_1858_));
 sg13g2_nor3_1 _5707_ (.A(_1856_),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_));
 sg13g2_inv_1 _5708_ (.Y(_1860_),
    .A(_1859_));
 sg13g2_nor2_1 _5709_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[0][0] ),
    .B(net1365),
    .Y(_1861_));
 sg13g2_nor2_1 _5710_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[2][0] ),
    .B(net1407),
    .Y(_1862_));
 sg13g2_nor2_1 _5711_ (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[1][0] ),
    .B(net1386),
    .Y(_1863_));
 sg13g2_nor3_1 _5712_ (.A(_1861_),
    .B(_1862_),
    .C(_1863_),
    .Y(_1864_));
 sg13g2_inv_2 _5713_ (.Y(_1865_),
    .A(_1864_));
 sg13g2_o21ai_1 _5714_ (.B1(_1865_),
    .Y(_1866_),
    .A1(_1783_),
    .A2(_1860_));
 sg13g2_nand3b_1 _5715_ (.B(_1859_),
    .C(_1864_),
    .Y(_1867_),
    .A_N(_1783_));
 sg13g2_and3_2 _5716_ (.X(_1868_),
    .A(net1188),
    .B(_1866_),
    .C(_1867_));
 sg13g2_nand3_1 _5717_ (.B(_1866_),
    .C(_1867_),
    .A(net1188),
    .Y(_1869_));
 sg13g2_and2_1 _5718_ (.A(\tt6581_inst.controller_inst.pw_hi_i[3] ),
    .B(net1379),
    .X(_1870_));
 sg13g2_a221oi_1 _5719_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[11] ),
    .C1(_1870_),
    .B1(net1397),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[19] ),
    .Y(_1871_),
    .A2(net1419));
 sg13g2_or2_1 _5720_ (.X(_1872_),
    .B(_1871_),
    .A(_1868_));
 sg13g2_a21oi_1 _5721_ (.A1(_1783_),
    .A2(_1860_),
    .Y(_1873_),
    .B1(_1781_));
 sg13g2_o21ai_1 _5722_ (.B1(_1873_),
    .Y(_1874_),
    .A1(_1783_),
    .A2(_1860_));
 sg13g2_a22oi_1 _5723_ (.Y(_1875_),
    .B1(net1378),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[2] ),
    .A2(net1419),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[18] ));
 sg13g2_o21ai_1 _5724_ (.B1(_1875_),
    .Y(_1876_),
    .A1(_0963_),
    .A2(net1390));
 sg13g2_nor2_1 _5725_ (.A(_1874_),
    .B(_1876_),
    .Y(_1877_));
 sg13g2_xor2_1 _5726_ (.B(_1876_),
    .A(_1874_),
    .X(_1878_));
 sg13g2_and2_1 _5727_ (.A(_1872_),
    .B(_1878_),
    .X(_1879_));
 sg13g2_and2_1 _5728_ (.A(_1868_),
    .B(_1871_),
    .X(_1880_));
 sg13g2_a21o_1 _5729_ (.A2(_1877_),
    .A1(_1872_),
    .B1(_1880_),
    .X(_1881_));
 sg13g2_a21oi_1 _5730_ (.A1(_1855_),
    .A2(_1879_),
    .Y(_1882_),
    .B1(_1881_));
 sg13g2_a21o_1 _5731_ (.A2(_1879_),
    .A1(_1855_),
    .B1(_1881_),
    .X(_1883_));
 sg13g2_nor2_1 _5732_ (.A(net1190),
    .B(net1144),
    .Y(_1884_));
 sg13g2_nor2_1 _5733_ (.A(_1613_),
    .B(_1842_),
    .Y(_1885_));
 sg13g2_a22oi_1 _5734_ (.Y(_1886_),
    .B1(net1379),
    .B2(\tt6581_inst.control_pack[2] ),
    .A2(net1420),
    .A1(\tt6581_inst.control_pack[18] ));
 sg13g2_o21ai_1 _5735_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_0972_),
    .A2(net1391));
 sg13g2_nand2_1 _5736_ (.Y(_1888_),
    .A(_1775_),
    .B(_1887_));
 sg13g2_xnor2_1 _5737_ (.Y(_1889_),
    .A(_1868_),
    .B(_1888_));
 sg13g2_xnor2_1 _5738_ (.Y(_1890_),
    .A(_1828_),
    .B(net1145));
 sg13g2_a21oi_1 _5739_ (.A1(net1215),
    .A2(_1890_),
    .Y(_1891_),
    .B1(_1885_));
 sg13g2_o21ai_1 _5740_ (.B1(_1891_),
    .Y(_1892_),
    .A1(net1190),
    .A2(net1144));
 sg13g2_a22oi_1 _5741_ (.Y(_1893_),
    .B1(\tt6581_inst.svf_inst.reg_band[0] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[0] ),
    .A1(net1535));
 sg13g2_nand2b_1 _5742_ (.Y(_1894_),
    .B(net1490),
    .A_N(_1893_));
 sg13g2_nor3_1 _5743_ (.A(\tt6581_inst.filt_en_mode[0] ),
    .B(_0919_),
    .C(\tt6581_inst.filt_en_mode[2] ),
    .Y(_1895_));
 sg13g2_nor2b_2 _5744_ (.A(\tt6581_inst.filt_en_mode[1] ),
    .B_N(\tt6581_inst.filt_en_mode[2] ),
    .Y(_1896_));
 sg13g2_nor2_2 _5745_ (.A(net1359),
    .B(_1896_),
    .Y(_1897_));
 sg13g2_or2_1 _5746_ (.X(_1898_),
    .B(_1896_),
    .A(net1359));
 sg13g2_nand2_1 _5747_ (.Y(_1899_),
    .A(\tt6581_inst.svf_inst.hp_node[22] ),
    .B(\tt6581_inst.svf_inst.reg_low[22] ));
 sg13g2_xnor2_1 _5748_ (.Y(_1900_),
    .A(\tt6581_inst.svf_inst.hp_node[15] ),
    .B(\tt6581_inst.svf_inst.reg_low[15] ));
 sg13g2_nand2_1 _5749_ (.Y(_1901_),
    .A(\tt6581_inst.svf_inst.hp_node[14] ),
    .B(\tt6581_inst.svf_inst.reg_low[14] ));
 sg13g2_xor2_1 _5750_ (.B(\tt6581_inst.svf_inst.reg_low[14] ),
    .A(\tt6581_inst.svf_inst.hp_node[14] ),
    .X(_1902_));
 sg13g2_nor2b_1 _5751_ (.A(_1900_),
    .B_N(_1902_),
    .Y(_1903_));
 sg13g2_and2_1 _5752_ (.A(\tt6581_inst.svf_inst.hp_node[13] ),
    .B(\tt6581_inst.svf_inst.reg_low[13] ),
    .X(_1904_));
 sg13g2_nor2_1 _5753_ (.A(\tt6581_inst.svf_inst.hp_node[13] ),
    .B(\tt6581_inst.svf_inst.reg_low[13] ),
    .Y(_1905_));
 sg13g2_nor2_1 _5754_ (.A(_1904_),
    .B(_1905_),
    .Y(_1906_));
 sg13g2_and2_1 _5755_ (.A(\tt6581_inst.svf_inst.hp_node[12] ),
    .B(\tt6581_inst.svf_inst.reg_low[12] ),
    .X(_1907_));
 sg13g2_xnor2_1 _5756_ (.Y(_1908_),
    .A(\tt6581_inst.svf_inst.hp_node[12] ),
    .B(\tt6581_inst.svf_inst.reg_low[12] ));
 sg13g2_nor3_1 _5757_ (.A(_1904_),
    .B(_1905_),
    .C(_1908_),
    .Y(_1909_));
 sg13g2_inv_1 _5758_ (.Y(_1910_),
    .A(_1909_));
 sg13g2_nand2_1 _5759_ (.Y(_1911_),
    .A(_1903_),
    .B(_1909_));
 sg13g2_nand2_1 _5760_ (.Y(_1912_),
    .A(\tt6581_inst.svf_inst.hp_node[10] ),
    .B(\tt6581_inst.svf_inst.reg_low[10] ));
 sg13g2_xnor2_1 _5761_ (.Y(_1913_),
    .A(\tt6581_inst.svf_inst.hp_node[10] ),
    .B(\tt6581_inst.svf_inst.reg_low[10] ));
 sg13g2_xor2_1 _5762_ (.B(\tt6581_inst.svf_inst.reg_low[11] ),
    .A(\tt6581_inst.svf_inst.hp_node[11] ),
    .X(_1914_));
 sg13g2_nor2b_1 _5763_ (.A(_1913_),
    .B_N(_1914_),
    .Y(_1915_));
 sg13g2_nand2_1 _5764_ (.Y(_1916_),
    .A(\tt6581_inst.svf_inst.hp_node[9] ),
    .B(net1505));
 sg13g2_nand2_1 _5765_ (.Y(_1917_),
    .A(\tt6581_inst.svf_inst.hp_node[8] ),
    .B(\tt6581_inst.svf_inst.reg_low[8] ));
 sg13g2_nor2_1 _5766_ (.A(\tt6581_inst.svf_inst.hp_node[9] ),
    .B(net1505),
    .Y(_1918_));
 sg13g2_o21ai_1 _5767_ (.B1(_1916_),
    .Y(_1919_),
    .A1(_1917_),
    .A2(_1918_));
 sg13g2_a21oi_1 _5768_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_1920_),
    .B1(_1912_));
 sg13g2_a221oi_1 _5769_ (.B2(_1919_),
    .C1(_1920_),
    .B1(_1915_),
    .A1(\tt6581_inst.svf_inst.hp_node[11] ),
    .Y(_1921_),
    .A2(\tt6581_inst.svf_inst.reg_low[11] ));
 sg13g2_and2_1 _5770_ (.A(\tt6581_inst.svf_inst.hp_node[4] ),
    .B(\tt6581_inst.svf_inst.reg_low[4] ),
    .X(_1922_));
 sg13g2_xnor2_1 _5771_ (.Y(_1923_),
    .A(\tt6581_inst.svf_inst.hp_node[4] ),
    .B(\tt6581_inst.svf_inst.reg_low[4] ));
 sg13g2_nor2_2 _5772_ (.A(\tt6581_inst.svf_inst.hp_node[3] ),
    .B(net1507),
    .Y(_1924_));
 sg13g2_and2_1 _5773_ (.A(\tt6581_inst.svf_inst.hp_node[2] ),
    .B(\tt6581_inst.svf_inst.reg_low[2] ),
    .X(_1925_));
 sg13g2_nand2_1 _5774_ (.Y(_1926_),
    .A(\tt6581_inst.svf_inst.hp_node[1] ),
    .B(net1508));
 sg13g2_nand2_1 _5775_ (.Y(_1927_),
    .A(\tt6581_inst.svf_inst.hp_node[0] ),
    .B(\tt6581_inst.svf_inst.reg_low[0] ));
 sg13g2_nor2_1 _5776_ (.A(\tt6581_inst.svf_inst.hp_node[1] ),
    .B(net1508),
    .Y(_1928_));
 sg13g2_xor2_1 _5777_ (.B(net1508),
    .A(\tt6581_inst.svf_inst.hp_node[1] ),
    .X(_1929_));
 sg13g2_o21ai_1 _5778_ (.B1(_1926_),
    .Y(_1930_),
    .A1(_1927_),
    .A2(_1928_));
 sg13g2_xnor2_1 _5779_ (.Y(_1931_),
    .A(\tt6581_inst.svf_inst.hp_node[2] ),
    .B(\tt6581_inst.svf_inst.reg_low[2] ));
 sg13g2_inv_1 _5780_ (.Y(_1932_),
    .A(_1931_));
 sg13g2_nand2_1 _5781_ (.Y(_1933_),
    .A(_1930_),
    .B(_1932_));
 sg13g2_nand2b_1 _5782_ (.Y(_1934_),
    .B(_1933_),
    .A_N(_1925_));
 sg13g2_a221oi_1 _5783_ (.B2(_1932_),
    .C1(_1925_),
    .B1(_1930_),
    .A1(\tt6581_inst.svf_inst.hp_node[3] ),
    .Y(_1935_),
    .A2(net1507));
 sg13g2_nor3_2 _5784_ (.A(_1923_),
    .B(_1924_),
    .C(_1935_),
    .Y(_1936_));
 sg13g2_nand2_1 _5785_ (.Y(_1937_),
    .A(\tt6581_inst.svf_inst.hp_node[7] ),
    .B(\tt6581_inst.svf_inst.reg_low[7] ));
 sg13g2_nor2_1 _5786_ (.A(\tt6581_inst.svf_inst.hp_node[7] ),
    .B(\tt6581_inst.svf_inst.reg_low[7] ),
    .Y(_1938_));
 sg13g2_xnor2_1 _5787_ (.Y(_1939_),
    .A(\tt6581_inst.svf_inst.hp_node[7] ),
    .B(\tt6581_inst.svf_inst.reg_low[7] ));
 sg13g2_nand2_1 _5788_ (.Y(_1940_),
    .A(\tt6581_inst.svf_inst.hp_node[6] ),
    .B(\tt6581_inst.svf_inst.reg_low[6] ));
 sg13g2_xnor2_1 _5789_ (.Y(_1941_),
    .A(\tt6581_inst.svf_inst.hp_node[6] ),
    .B(\tt6581_inst.svf_inst.reg_low[6] ));
 sg13g2_nor2_1 _5790_ (.A(_1939_),
    .B(_1941_),
    .Y(_1942_));
 sg13g2_nor2_1 _5791_ (.A(\tt6581_inst.svf_inst.hp_node[5] ),
    .B(net1506),
    .Y(_1943_));
 sg13g2_xor2_1 _5792_ (.B(net1506),
    .A(\tt6581_inst.svf_inst.hp_node[5] ),
    .X(_1944_));
 sg13g2_nand2_1 _5793_ (.Y(_1945_),
    .A(_1942_),
    .B(_1944_));
 sg13g2_nor4_2 _5794_ (.A(_1923_),
    .B(_1924_),
    .C(_1935_),
    .Y(_1946_),
    .D(_1945_));
 sg13g2_a21oi_1 _5795_ (.A1(\tt6581_inst.svf_inst.hp_node[5] ),
    .A2(net1506),
    .Y(_1947_),
    .B1(_1922_));
 sg13g2_nor4_1 _5796_ (.A(_1939_),
    .B(_1941_),
    .C(_1943_),
    .D(_1947_),
    .Y(_1948_));
 sg13g2_o21ai_1 _5797_ (.B1(_1937_),
    .Y(_1949_),
    .A1(_1938_),
    .A2(_1940_));
 sg13g2_or2_1 _5798_ (.X(_1950_),
    .B(_1949_),
    .A(_1948_));
 sg13g2_nor2_1 _5799_ (.A(_1946_),
    .B(_1950_),
    .Y(_1951_));
 sg13g2_xnor2_1 _5800_ (.Y(_1952_),
    .A(\tt6581_inst.svf_inst.hp_node[8] ),
    .B(\tt6581_inst.svf_inst.reg_low[8] ));
 sg13g2_xnor2_1 _5801_ (.Y(_1953_),
    .A(\tt6581_inst.svf_inst.hp_node[9] ),
    .B(\tt6581_inst.svf_inst.reg_low[9] ));
 sg13g2_nor2_1 _5802_ (.A(_1952_),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_nand2_1 _5803_ (.Y(_1955_),
    .A(_1915_),
    .B(_1954_));
 sg13g2_inv_1 _5804_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_o21ai_1 _5805_ (.B1(_1956_),
    .Y(_1957_),
    .A1(_1946_),
    .A2(_1950_));
 sg13g2_a21oi_1 _5806_ (.A1(_0929_),
    .A2(_0930_),
    .Y(_1958_),
    .B1(_1901_));
 sg13g2_a21oi_1 _5807_ (.A1(\tt6581_inst.svf_inst.hp_node[15] ),
    .A2(\tt6581_inst.svf_inst.reg_low[15] ),
    .Y(_1959_),
    .B1(_1958_));
 sg13g2_nor2_1 _5808_ (.A(_1904_),
    .B(_1907_),
    .Y(_1960_));
 sg13g2_nor2_1 _5809_ (.A(_1905_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_o21ai_1 _5810_ (.B1(_1959_),
    .Y(_1962_),
    .A1(_1911_),
    .A2(_1921_));
 sg13g2_a21oi_2 _5811_ (.B1(_1962_),
    .Y(_1963_),
    .A2(_1961_),
    .A1(_1903_));
 sg13g2_nor2_1 _5812_ (.A(_1911_),
    .B(_1955_),
    .Y(_1964_));
 sg13g2_o21ai_1 _5813_ (.B1(_1964_),
    .Y(_1965_),
    .A1(_1946_),
    .A2(_1950_));
 sg13g2_nand2_1 _5814_ (.Y(_1966_),
    .A(\tt6581_inst.svf_inst.hp_node[16] ),
    .B(\tt6581_inst.svf_inst.reg_low[16] ));
 sg13g2_xnor2_1 _5815_ (.Y(_1967_),
    .A(\tt6581_inst.svf_inst.hp_node[16] ),
    .B(\tt6581_inst.svf_inst.reg_low[16] ));
 sg13g2_xnor2_1 _5816_ (.Y(_1968_),
    .A(\tt6581_inst.svf_inst.hp_node[17] ),
    .B(\tt6581_inst.svf_inst.reg_low[17] ));
 sg13g2_or2_1 _5817_ (.X(_1969_),
    .B(_1968_),
    .A(_1967_));
 sg13g2_a21o_1 _5818_ (.A2(_1965_),
    .A1(_1963_),
    .B1(_1969_),
    .X(_1970_));
 sg13g2_nor2_1 _5819_ (.A(\tt6581_inst.svf_inst.hp_node[19] ),
    .B(\tt6581_inst.svf_inst.reg_low[19] ),
    .Y(_1971_));
 sg13g2_nand2_1 _5820_ (.Y(_1972_),
    .A(\tt6581_inst.svf_inst.hp_node[18] ),
    .B(\tt6581_inst.svf_inst.reg_low[18] ));
 sg13g2_a22oi_1 _5821_ (.Y(_1973_),
    .B1(\tt6581_inst.svf_inst.hp_node[18] ),
    .B2(\tt6581_inst.svf_inst.reg_low[18] ),
    .A2(\tt6581_inst.svf_inst.reg_low[19] ),
    .A1(\tt6581_inst.svf_inst.hp_node[19] ));
 sg13g2_a21oi_1 _5822_ (.A1(_0926_),
    .A2(_0927_),
    .Y(_1974_),
    .B1(_1966_));
 sg13g2_a21oi_1 _5823_ (.A1(\tt6581_inst.svf_inst.hp_node[17] ),
    .A2(\tt6581_inst.svf_inst.reg_low[17] ),
    .Y(_1975_),
    .B1(_1974_));
 sg13g2_xnor2_1 _5824_ (.Y(_1976_),
    .A(\tt6581_inst.svf_inst.hp_node[19] ),
    .B(\tt6581_inst.svf_inst.reg_low[19] ));
 sg13g2_xnor2_1 _5825_ (.Y(_1977_),
    .A(\tt6581_inst.svf_inst.hp_node[18] ),
    .B(\tt6581_inst.svf_inst.reg_low[18] ));
 sg13g2_nor2_1 _5826_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_nand2b_1 _5827_ (.Y(_1979_),
    .B(_1978_),
    .A_N(_1975_));
 sg13g2_o21ai_1 _5828_ (.B1(_1979_),
    .Y(_1980_),
    .A1(_1971_),
    .A2(_1973_));
 sg13g2_inv_1 _5829_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_nand2b_1 _5830_ (.Y(_1982_),
    .B(_1978_),
    .A_N(_1969_));
 sg13g2_a21oi_1 _5831_ (.A1(_1963_),
    .A2(_1965_),
    .Y(_1983_),
    .B1(_1982_));
 sg13g2_a21o_1 _5832_ (.A2(_1965_),
    .A1(_1963_),
    .B1(_1982_),
    .X(_1984_));
 sg13g2_nand2_1 _5833_ (.Y(_1985_),
    .A(\tt6581_inst.svf_inst.hp_node[20] ),
    .B(\tt6581_inst.svf_inst.reg_low[20] ));
 sg13g2_xor2_1 _5834_ (.B(\tt6581_inst.svf_inst.reg_low[20] ),
    .A(\tt6581_inst.svf_inst.hp_node[20] ),
    .X(_1986_));
 sg13g2_nand2_1 _5835_ (.Y(_1987_),
    .A(\tt6581_inst.svf_inst.hp_node[21] ),
    .B(\tt6581_inst.svf_inst.reg_low[21] ));
 sg13g2_nor2_1 _5836_ (.A(\tt6581_inst.svf_inst.hp_node[21] ),
    .B(\tt6581_inst.svf_inst.reg_low[21] ),
    .Y(_1988_));
 sg13g2_xnor2_1 _5837_ (.Y(_1989_),
    .A(\tt6581_inst.svf_inst.hp_node[21] ),
    .B(\tt6581_inst.svf_inst.reg_low[21] ));
 sg13g2_nand3b_1 _5838_ (.B(_1986_),
    .C(_1987_),
    .Y(_1990_),
    .A_N(_1988_));
 sg13g2_a21oi_1 _5839_ (.A1(_1981_),
    .A2(_1984_),
    .Y(_1991_),
    .B1(_1990_));
 sg13g2_o21ai_1 _5840_ (.B1(_1987_),
    .Y(_1992_),
    .A1(_1985_),
    .A2(_1988_));
 sg13g2_xor2_1 _5841_ (.B(\tt6581_inst.svf_inst.reg_low[22] ),
    .A(\tt6581_inst.svf_inst.hp_node[22] ),
    .X(_1993_));
 sg13g2_o21ai_1 _5842_ (.B1(_1993_),
    .Y(_1994_),
    .A1(_1991_),
    .A2(_1992_));
 sg13g2_xnor2_1 _5843_ (.Y(_1995_),
    .A(\tt6581_inst.svf_inst.reg_low[23] ),
    .B(\tt6581_inst.svf_inst.hp_node[23] ));
 sg13g2_nand3_1 _5844_ (.B(_1994_),
    .C(_1995_),
    .A(_1899_),
    .Y(_1996_));
 sg13g2_a21o_1 _5845_ (.A2(_1994_),
    .A1(_1899_),
    .B1(_1995_),
    .X(_1997_));
 sg13g2_and2_1 _5846_ (.A(\tt6581_inst.filt_en_mode[0] ),
    .B(_1896_),
    .X(_1998_));
 sg13g2_nand3_1 _5847_ (.B(_1997_),
    .C(net1354),
    .A(_1996_),
    .Y(_1999_));
 sg13g2_nor2b_1 _5848_ (.A(\tt6581_inst.filt_en_mode[0] ),
    .B_N(_1896_),
    .Y(_2000_));
 sg13g2_a221oi_1 _5849_ (.B2(\tt6581_inst.svf_inst.hp_node[23] ),
    .C1(net1268),
    .B1(net1351),
    .A1(\tt6581_inst.svf_inst.reg_band[23] ),
    .Y(_2001_),
    .A2(net1359));
 sg13g2_a22oi_1 _5850_ (.Y(_2002_),
    .B1(_1999_),
    .B2(_2001_),
    .A2(net1268),
    .A1(_0918_));
 sg13g2_a21o_1 _5851_ (.A2(_1975_),
    .A1(_1970_),
    .B1(_1977_),
    .X(_2003_));
 sg13g2_a21o_1 _5852_ (.A2(_2003_),
    .A1(_1972_),
    .B1(_1976_),
    .X(_2004_));
 sg13g2_nand3_1 _5853_ (.B(_1976_),
    .C(_2003_),
    .A(_1972_),
    .Y(_2005_));
 sg13g2_nand3_1 _5854_ (.B(_2004_),
    .C(_2005_),
    .A(net1355),
    .Y(_2006_));
 sg13g2_a221oi_1 _5855_ (.B2(\tt6581_inst.svf_inst.hp_node[19] ),
    .C1(net1267),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[19] ),
    .Y(_2007_),
    .A2(net1358));
 sg13g2_a22oi_1 _5856_ (.Y(_2008_),
    .B1(_2006_),
    .B2(_2007_),
    .A2(net1266),
    .A1(_0924_));
 sg13g2_nor2_1 _5857_ (.A(\tt6581_inst.svf_inst.reg_low[17] ),
    .B(_1898_),
    .Y(_2009_));
 sg13g2_a21o_1 _5858_ (.A2(_1965_),
    .A1(_1963_),
    .B1(_1967_),
    .X(_2010_));
 sg13g2_a21oi_1 _5859_ (.A1(_1966_),
    .A2(_2010_),
    .Y(_2011_),
    .B1(_1968_));
 sg13g2_nand3_1 _5860_ (.B(_1968_),
    .C(_2010_),
    .A(_1966_),
    .Y(_2012_));
 sg13g2_nand3b_1 _5861_ (.B(_2012_),
    .C(net1354),
    .Y(_2013_),
    .A_N(_2011_));
 sg13g2_a221oi_1 _5862_ (.B2(\tt6581_inst.svf_inst.hp_node[17] ),
    .C1(net1266),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[17] ),
    .Y(_2014_),
    .A2(net1358));
 sg13g2_a21o_1 _5863_ (.A2(_2014_),
    .A1(_2013_),
    .B1(_2009_),
    .X(_2015_));
 sg13g2_nor2_1 _5864_ (.A(\tt6581_inst.svf_inst.reg_low[18] ),
    .B(_1898_),
    .Y(_2016_));
 sg13g2_nand3_1 _5865_ (.B(_1975_),
    .C(_1977_),
    .A(_1970_),
    .Y(_2017_));
 sg13g2_nand3_1 _5866_ (.B(_2003_),
    .C(_2017_),
    .A(net1354),
    .Y(_2018_));
 sg13g2_a221oi_1 _5867_ (.B2(\tt6581_inst.svf_inst.hp_node[18] ),
    .C1(net1267),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[18] ),
    .Y(_2019_),
    .A2(net1358));
 sg13g2_a21o_1 _5868_ (.A2(_2019_),
    .A1(_2018_),
    .B1(_2016_),
    .X(_2020_));
 sg13g2_a21oi_1 _5869_ (.A1(_1921_),
    .A2(_1957_),
    .Y(_2021_),
    .B1(_1908_));
 sg13g2_a21oi_1 _5870_ (.A1(_1921_),
    .A2(_1957_),
    .Y(_2022_),
    .B1(_1910_));
 sg13g2_or3_1 _5871_ (.A(_1902_),
    .B(_1961_),
    .C(_2022_),
    .X(_2023_));
 sg13g2_o21ai_1 _5872_ (.B1(_1902_),
    .Y(_2024_),
    .A1(_1961_),
    .A2(_2022_));
 sg13g2_nand3_1 _5873_ (.B(_2023_),
    .C(_2024_),
    .A(net1354),
    .Y(_2025_));
 sg13g2_a221oi_1 _5874_ (.B2(\tt6581_inst.svf_inst.hp_node[14] ),
    .C1(net1266),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[14] ),
    .Y(_2026_),
    .A2(net1358));
 sg13g2_a22oi_1 _5875_ (.Y(_2027_),
    .B1(_2025_),
    .B2(_2026_),
    .A2(net1266),
    .A1(_0932_));
 sg13g2_nand3_1 _5876_ (.B(_1965_),
    .C(_1967_),
    .A(_1963_),
    .Y(_2028_));
 sg13g2_nand3_1 _5877_ (.B(_2010_),
    .C(_2028_),
    .A(net1354),
    .Y(_2029_));
 sg13g2_a221oi_1 _5878_ (.B2(\tt6581_inst.svf_inst.hp_node[16] ),
    .C1(net1266),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[16] ),
    .Y(_2030_),
    .A2(net1358));
 sg13g2_a22oi_1 _5879_ (.Y(_2031_),
    .B1(_2029_),
    .B2(_2030_),
    .A2(net1266),
    .A1(_0928_));
 sg13g2_nor2_1 _5880_ (.A(\tt6581_inst.svf_inst.reg_low[13] ),
    .B(_1898_),
    .Y(_2032_));
 sg13g2_or3_1 _5881_ (.A(_1906_),
    .B(_1907_),
    .C(_2021_),
    .X(_2033_));
 sg13g2_o21ai_1 _5882_ (.B1(_1906_),
    .Y(_2034_),
    .A1(_1907_),
    .A2(_2021_));
 sg13g2_nand3_1 _5883_ (.B(_2033_),
    .C(_2034_),
    .A(net1355),
    .Y(_2035_));
 sg13g2_a221oi_1 _5884_ (.B2(\tt6581_inst.svf_inst.hp_node[13] ),
    .C1(net1267),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[13] ),
    .Y(_2036_),
    .A2(net1358));
 sg13g2_a21o_1 _5885_ (.A2(_2036_),
    .A1(_2035_),
    .B1(_2032_),
    .X(_2037_));
 sg13g2_o21ai_1 _5886_ (.B1(_1986_),
    .Y(_2038_),
    .A1(_1980_),
    .A2(_1983_));
 sg13g2_nand3b_1 _5887_ (.B(_1981_),
    .C(_1984_),
    .Y(_2039_),
    .A_N(_1986_));
 sg13g2_nand3_1 _5888_ (.B(_2038_),
    .C(_2039_),
    .A(net1354),
    .Y(_2040_));
 sg13g2_a221oi_1 _5889_ (.B2(\tt6581_inst.svf_inst.hp_node[20] ),
    .C1(net1268),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[20] ),
    .Y(_2041_),
    .A2(net1358));
 sg13g2_a22oi_1 _5890_ (.Y(_2042_),
    .B1(_2040_),
    .B2(_2041_),
    .A2(net1268),
    .A1(_0923_));
 sg13g2_a21o_1 _5891_ (.A2(_2024_),
    .A1(_1901_),
    .B1(_1900_),
    .X(_2043_));
 sg13g2_nand3_1 _5892_ (.B(_1901_),
    .C(_2024_),
    .A(_1900_),
    .Y(_2044_));
 sg13g2_nand3_1 _5893_ (.B(_2043_),
    .C(_2044_),
    .A(net1354),
    .Y(_2045_));
 sg13g2_a221oi_1 _5894_ (.B2(\tt6581_inst.svf_inst.hp_node[15] ),
    .C1(net1266),
    .B1(net1350),
    .A1(\tt6581_inst.svf_inst.reg_band[15] ),
    .Y(_2046_),
    .A2(net1358));
 sg13g2_a22oi_1 _5895_ (.Y(_2047_),
    .B1(_2045_),
    .B2(_2046_),
    .A2(net1266),
    .A1(_0930_));
 sg13g2_a21o_1 _5896_ (.A2(_2038_),
    .A1(_1985_),
    .B1(_1989_),
    .X(_2048_));
 sg13g2_nand3_1 _5897_ (.B(_1989_),
    .C(_2038_),
    .A(_1985_),
    .Y(_2049_));
 sg13g2_nand3_1 _5898_ (.B(_2048_),
    .C(_2049_),
    .A(net1354),
    .Y(_2050_));
 sg13g2_a221oi_1 _5899_ (.B2(\tt6581_inst.svf_inst.hp_node[21] ),
    .C1(net1268),
    .B1(net1351),
    .A1(\tt6581_inst.svf_inst.reg_band[21] ),
    .Y(_2051_),
    .A2(net1359));
 sg13g2_a22oi_1 _5900_ (.Y(_2052_),
    .B1(_2050_),
    .B2(_2051_),
    .A2(net1268),
    .A1(_0922_));
 sg13g2_or3_1 _5901_ (.A(_1991_),
    .B(_1992_),
    .C(_1993_),
    .X(_2053_));
 sg13g2_nand3_1 _5902_ (.B(net1355),
    .C(_2053_),
    .A(_1994_),
    .Y(_2054_));
 sg13g2_a221oi_1 _5903_ (.B2(\tt6581_inst.svf_inst.hp_node[22] ),
    .C1(net1268),
    .B1(net1351),
    .A1(\tt6581_inst.svf_inst.reg_band[22] ),
    .Y(_2055_),
    .A2(net1359));
 sg13g2_a22oi_1 _5904_ (.Y(_2056_),
    .B1(_2054_),
    .B2(_2055_),
    .A2(net1269),
    .A1(_0920_));
 sg13g2_nor3_1 _5905_ (.A(_2015_),
    .B(_2020_),
    .C(_2037_),
    .Y(_2057_));
 sg13g2_nand4_1 _5906_ (.B(_2031_),
    .C(_2042_),
    .A(_2027_),
    .Y(_2058_),
    .D(_2057_));
 sg13g2_nand4_1 _5907_ (.B(_2047_),
    .C(_2052_),
    .A(_2008_),
    .Y(_2059_),
    .D(_2056_));
 sg13g2_o21ai_1 _5908_ (.B1(_2002_),
    .Y(_2060_),
    .A1(_2058_),
    .A2(_2059_));
 sg13g2_inv_1 _5909_ (.Y(_2061_),
    .A(net1154));
 sg13g2_nand3_1 _5910_ (.B(_2020_),
    .C(_2037_),
    .A(_2015_),
    .Y(_2062_));
 sg13g2_nor4_1 _5911_ (.A(_2027_),
    .B(_2031_),
    .C(_2042_),
    .D(_2062_),
    .Y(_2063_));
 sg13g2_nor4_1 _5912_ (.A(_2008_),
    .B(_2047_),
    .C(_2052_),
    .D(_2056_),
    .Y(_2064_));
 sg13g2_a21oi_1 _5913_ (.A1(_2063_),
    .A2(_2064_),
    .Y(_2065_),
    .B1(_2002_));
 sg13g2_nand2_1 _5914_ (.Y(_2066_),
    .A(\tt6581_inst.svf_inst.reg_band[0] ),
    .B(net1360));
 sg13g2_a21oi_1 _5915_ (.A1(\tt6581_inst.svf_inst.hp_node[0] ),
    .A2(_1898_),
    .Y(_2067_),
    .B1(\tt6581_inst.svf_inst.reg_low[0] ));
 sg13g2_a221oi_1 _5916_ (.B2(\tt6581_inst.svf_inst.hp_node[0] ),
    .C1(net1270),
    .B1(net1352),
    .A1(_1927_),
    .Y(_2068_),
    .A2(net1356));
 sg13g2_o21ai_1 _5917_ (.B1(_2066_),
    .Y(_2069_),
    .A1(_2067_),
    .A2(_2068_));
 sg13g2_o21ai_1 _5918_ (.B1(net1153),
    .Y(_2070_),
    .A1(net1151),
    .A2(_2069_));
 sg13g2_nor2_1 _5919_ (.A(_0950_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_a21o_1 _5920_ (.A2(_2070_),
    .A1(_0950_),
    .B1(_0916_),
    .X(_2072_));
 sg13g2_o21ai_1 _5921_ (.B1(_1894_),
    .Y(_2073_),
    .A1(_2071_),
    .A2(_2072_));
 sg13g2_a21o_2 _5922_ (.A2(_1892_),
    .A1(_1619_),
    .B1(_2073_),
    .X(_2074_));
 sg13g2_a22oi_1 _5923_ (.Y(_2075_),
    .B1(_2074_),
    .B2(_1018_),
    .A2(net1224),
    .A1(net817));
 sg13g2_inv_1 _5924_ (.Y(_0299_),
    .A(_2075_));
 sg13g2_xnor2_1 _5925_ (.Y(_2076_),
    .A(_1842_),
    .B(net1145));
 sg13g2_a22oi_1 _5926_ (.Y(_2077_),
    .B1(_2076_),
    .B2(net1215),
    .A2(_1822_),
    .A1(_1612_));
 sg13g2_o21ai_1 _5927_ (.B1(_2077_),
    .Y(_2078_),
    .A1(_1615_),
    .A2(net1144));
 sg13g2_xnor2_1 _5928_ (.Y(_2079_),
    .A(_1927_),
    .B(_1929_));
 sg13g2_nand2_1 _5929_ (.Y(_2080_),
    .A(net1356),
    .B(_2079_));
 sg13g2_a221oi_1 _5930_ (.B2(\tt6581_inst.svf_inst.hp_node[1] ),
    .C1(net1271),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_band[1] ),
    .Y(_2081_),
    .A2(net1360));
 sg13g2_a22oi_1 _5931_ (.Y(_2082_),
    .B1(_2080_),
    .B2(_2081_),
    .A2(net1271),
    .A1(_0943_));
 sg13g2_a21oi_1 _5932_ (.A1(net1153),
    .A2(_2082_),
    .Y(_2083_),
    .B1(net1151));
 sg13g2_nor2_1 _5933_ (.A(_0973_),
    .B(_2083_),
    .Y(_2084_));
 sg13g2_xnor2_1 _5934_ (.Y(_2085_),
    .A(\tt6581_inst.bypass_accum[1] ),
    .B(_2083_));
 sg13g2_a21oi_1 _5935_ (.A1(_2071_),
    .A2(_2085_),
    .Y(_2086_),
    .B1(_0916_));
 sg13g2_o21ai_1 _5936_ (.B1(_2086_),
    .Y(_2087_),
    .A1(_2071_),
    .A2(_2085_));
 sg13g2_a22oi_1 _5937_ (.Y(_2088_),
    .B1(\tt6581_inst.svf_inst.reg_band[1] ),
    .B2(net1430),
    .A2(\tt6581_inst.svf_inst.hp_node[1] ),
    .A1(net1535));
 sg13g2_o21ai_1 _5938_ (.B1(_2087_),
    .Y(_2089_),
    .A1(net1435),
    .A2(_2088_));
 sg13g2_a21o_2 _5939_ (.A2(_2078_),
    .A1(_1619_),
    .B1(_2089_),
    .X(_2090_));
 sg13g2_nand3_1 _5940_ (.B(_1921_),
    .C(_1957_),
    .A(_1908_),
    .Y(_2091_));
 sg13g2_nor2b_1 _5941_ (.A(_2021_),
    .B_N(net1355),
    .Y(_2092_));
 sg13g2_a22oi_1 _5942_ (.Y(_2093_),
    .B1(net1351),
    .B2(\tt6581_inst.svf_inst.hp_node[12] ),
    .A2(net1359),
    .A1(\tt6581_inst.svf_inst.reg_band[12] ));
 sg13g2_nand2_1 _5943_ (.Y(_2094_),
    .A(_1898_),
    .B(_2093_));
 sg13g2_a21oi_1 _5944_ (.A1(_2091_),
    .A2(_2092_),
    .Y(_2095_),
    .B1(_2094_));
 sg13g2_a21oi_1 _5945_ (.A1(_0934_),
    .A2(net1269),
    .Y(_2096_),
    .B1(_2095_));
 sg13g2_a21oi_1 _5946_ (.A1(net1154),
    .A2(_2096_),
    .Y(_2097_),
    .B1(net1152));
 sg13g2_nand2b_1 _5947_ (.Y(_2098_),
    .B(\tt6581_inst.bypass_accum[12] ),
    .A_N(_2097_));
 sg13g2_nand2_1 _5948_ (.Y(_2099_),
    .A(net1507),
    .B(net1270));
 sg13g2_xor2_1 _5949_ (.B(net1507),
    .A(\tt6581_inst.svf_inst.hp_node[3] ),
    .X(_2100_));
 sg13g2_o21ai_1 _5950_ (.B1(net1356),
    .Y(_2101_),
    .A1(_1934_),
    .A2(_2100_));
 sg13g2_a21o_1 _5951_ (.A2(_2100_),
    .A1(_1934_),
    .B1(_2101_),
    .X(_2102_));
 sg13g2_a22oi_1 _5952_ (.Y(_2103_),
    .B1(net1352),
    .B2(\tt6581_inst.svf_inst.hp_node[3] ),
    .A2(net1360),
    .A1(\tt6581_inst.svf_inst.reg_band[3] ));
 sg13g2_nand3_1 _5953_ (.B(_2102_),
    .C(_2103_),
    .A(_2099_),
    .Y(_2104_));
 sg13g2_a21oi_1 _5954_ (.A1(net1153),
    .A2(_2104_),
    .Y(_2105_),
    .B1(net1151));
 sg13g2_nor2b_1 _5955_ (.A(_2105_),
    .B_N(\tt6581_inst.bypass_accum[3] ),
    .Y(_2106_));
 sg13g2_nand2b_1 _5956_ (.Y(_2107_),
    .B(_1931_),
    .A_N(_1930_));
 sg13g2_nand3_1 _5957_ (.B(net1356),
    .C(_2107_),
    .A(_1933_),
    .Y(_2108_));
 sg13g2_a221oi_1 _5958_ (.B2(\tt6581_inst.svf_inst.hp_node[2] ),
    .C1(net1271),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_band[2] ),
    .Y(_2109_),
    .A2(net1360));
 sg13g2_a22oi_1 _5959_ (.Y(_2110_),
    .B1(_2108_),
    .B2(_2109_),
    .A2(net1271),
    .A1(_0942_));
 sg13g2_a21oi_1 _5960_ (.A1(net1153),
    .A2(_2110_),
    .Y(_2111_),
    .B1(net1151));
 sg13g2_nand2b_1 _5961_ (.Y(_2112_),
    .B(\tt6581_inst.bypass_accum[2] ),
    .A_N(_2111_));
 sg13g2_a21oi_1 _5962_ (.A1(_2071_),
    .A2(_2085_),
    .Y(_2113_),
    .B1(_2084_));
 sg13g2_nor2b_1 _5963_ (.A(\tt6581_inst.bypass_accum[2] ),
    .B_N(_2111_),
    .Y(_2114_));
 sg13g2_xnor2_1 _5964_ (.Y(_2115_),
    .A(\tt6581_inst.bypass_accum[2] ),
    .B(_2111_));
 sg13g2_o21ai_1 _5965_ (.B1(_2112_),
    .Y(_2116_),
    .A1(_2113_),
    .A2(_2114_));
 sg13g2_nand2b_1 _5966_ (.Y(_2117_),
    .B(_2105_),
    .A_N(\tt6581_inst.bypass_accum[3] ));
 sg13g2_nand2b_1 _5967_ (.Y(_2118_),
    .B(_2117_),
    .A_N(_2106_));
 sg13g2_a21oi_2 _5968_ (.B1(_2106_),
    .Y(_2119_),
    .A2(_2117_),
    .A1(_2116_));
 sg13g2_nand2_1 _5969_ (.Y(_2120_),
    .A(net1506),
    .B(net1270));
 sg13g2_o21ai_1 _5970_ (.B1(_1944_),
    .Y(_2121_),
    .A1(_1922_),
    .A2(_1936_));
 sg13g2_or3_1 _5971_ (.A(_1922_),
    .B(_1936_),
    .C(_1944_),
    .X(_2122_));
 sg13g2_nand3_1 _5972_ (.B(_2121_),
    .C(_2122_),
    .A(net1357),
    .Y(_2123_));
 sg13g2_a22oi_1 _5973_ (.Y(_2124_),
    .B1(net1353),
    .B2(\tt6581_inst.svf_inst.hp_node[5] ),
    .A2(net1361),
    .A1(\tt6581_inst.svf_inst.reg_band[5] ));
 sg13g2_nand3_1 _5974_ (.B(_2123_),
    .C(_2124_),
    .A(_2120_),
    .Y(_2125_));
 sg13g2_a21oi_1 _5975_ (.A1(net1153),
    .A2(_2125_),
    .Y(_2126_),
    .B1(net1151));
 sg13g2_nand2_1 _5976_ (.Y(_2127_),
    .A(_0977_),
    .B(_2126_));
 sg13g2_nand2b_1 _5977_ (.Y(_2128_),
    .B(\tt6581_inst.bypass_accum[5] ),
    .A_N(_2126_));
 sg13g2_and2_1 _5978_ (.A(_2127_),
    .B(_2128_),
    .X(_2129_));
 sg13g2_o21ai_1 _5979_ (.B1(_1923_),
    .Y(_2130_),
    .A1(_1924_),
    .A2(_1935_));
 sg13g2_nor2b_1 _5980_ (.A(_1936_),
    .B_N(_2130_),
    .Y(_2131_));
 sg13g2_a22oi_1 _5981_ (.Y(_2132_),
    .B1(net1353),
    .B2(\tt6581_inst.svf_inst.hp_node[4] ),
    .A2(net1360),
    .A1(\tt6581_inst.svf_inst.reg_band[4] ));
 sg13g2_nand2_1 _5982_ (.Y(_2133_),
    .A(_1898_),
    .B(_2132_));
 sg13g2_a21oi_1 _5983_ (.A1(net1357),
    .A2(_2131_),
    .Y(_2134_),
    .B1(_2133_));
 sg13g2_a21oi_1 _5984_ (.A1(_0941_),
    .A2(net1270),
    .Y(_2135_),
    .B1(_2134_));
 sg13g2_a21o_1 _5985_ (.A2(_2135_),
    .A1(net1153),
    .B1(net1152),
    .X(_2136_));
 sg13g2_and2_1 _5986_ (.A(\tt6581_inst.bypass_accum[4] ),
    .B(_2136_),
    .X(_2137_));
 sg13g2_xor2_1 _5987_ (.B(_2136_),
    .A(\tt6581_inst.bypass_accum[4] ),
    .X(_2138_));
 sg13g2_nand2_1 _5988_ (.Y(_2139_),
    .A(_2129_),
    .B(_2138_));
 sg13g2_nor2_1 _5989_ (.A(_2119_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_nand2_1 _5990_ (.Y(_2141_),
    .A(_2127_),
    .B(_2137_));
 sg13g2_nand2_1 _5991_ (.Y(_2142_),
    .A(_2128_),
    .B(_2141_));
 sg13g2_nor2b_1 _5992_ (.A(_1936_),
    .B_N(_1947_),
    .Y(_2143_));
 sg13g2_or3_1 _5993_ (.A(_1941_),
    .B(_1943_),
    .C(_2143_),
    .X(_2144_));
 sg13g2_nand3_1 _5994_ (.B(_1940_),
    .C(_2144_),
    .A(_1939_),
    .Y(_2145_));
 sg13g2_a21o_1 _5995_ (.A2(_2144_),
    .A1(_1940_),
    .B1(_1939_),
    .X(_2146_));
 sg13g2_nand3_1 _5996_ (.B(_2145_),
    .C(_2146_),
    .A(net1356),
    .Y(_2147_));
 sg13g2_a221oi_1 _5997_ (.B2(\tt6581_inst.svf_inst.hp_node[7] ),
    .C1(net1270),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_band[7] ),
    .Y(_2148_),
    .A2(net1361));
 sg13g2_a22oi_1 _5998_ (.Y(_2149_),
    .B1(_2147_),
    .B2(_2148_),
    .A2(net1270),
    .A1(_0939_));
 sg13g2_a21oi_1 _5999_ (.A1(net1153),
    .A2(_2149_),
    .Y(_2150_),
    .B1(net1151));
 sg13g2_nand2b_1 _6000_ (.Y(_2151_),
    .B(_2150_),
    .A_N(\tt6581_inst.bypass_accum[7] ));
 sg13g2_nand2b_1 _6001_ (.Y(_2152_),
    .B(\tt6581_inst.bypass_accum[7] ),
    .A_N(_2150_));
 sg13g2_o21ai_1 _6002_ (.B1(_1941_),
    .Y(_2153_),
    .A1(_1943_),
    .A2(_2143_));
 sg13g2_nand3_1 _6003_ (.B(_2144_),
    .C(_2153_),
    .A(net1357),
    .Y(_2154_));
 sg13g2_a221oi_1 _6004_ (.B2(\tt6581_inst.svf_inst.hp_node[6] ),
    .C1(net1270),
    .B1(net1353),
    .A1(\tt6581_inst.svf_inst.reg_band[6] ),
    .Y(_2155_),
    .A2(net1361));
 sg13g2_a22oi_1 _6005_ (.Y(_2156_),
    .B1(_2154_),
    .B2(_2155_),
    .A2(net1270),
    .A1(_0940_));
 sg13g2_a21oi_1 _6006_ (.A1(net1154),
    .A2(_2156_),
    .Y(_2157_),
    .B1(net1151));
 sg13g2_nand2b_1 _6007_ (.Y(_2158_),
    .B(\tt6581_inst.bypass_accum[6] ),
    .A_N(_2157_));
 sg13g2_nand2_1 _6008_ (.Y(_2159_),
    .A(_2152_),
    .B(_2158_));
 sg13g2_a21oi_1 _6009_ (.A1(_2151_),
    .A2(_2159_),
    .Y(_2160_),
    .B1(_2142_));
 sg13g2_o21ai_1 _6010_ (.B1(_2160_),
    .Y(_2161_),
    .A1(_2119_),
    .A2(_2139_));
 sg13g2_nand2b_1 _6011_ (.Y(_2162_),
    .B(_2157_),
    .A_N(\tt6581_inst.bypass_accum[6] ));
 sg13g2_nand2b_1 _6012_ (.Y(_2163_),
    .B(_2152_),
    .A_N(_2162_));
 sg13g2_and2_1 _6013_ (.A(_2151_),
    .B(_2163_),
    .X(_2164_));
 sg13g2_nand2_1 _6014_ (.Y(_2165_),
    .A(_2161_),
    .B(_2164_));
 sg13g2_o21ai_1 _6015_ (.B1(net1356),
    .Y(_2166_),
    .A1(_1951_),
    .A2(_1952_));
 sg13g2_a21o_1 _6016_ (.A2(_1952_),
    .A1(_1951_),
    .B1(_2166_),
    .X(_2167_));
 sg13g2_a221oi_1 _6017_ (.B2(\tt6581_inst.svf_inst.hp_node[8] ),
    .C1(net1272),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_band[8] ),
    .Y(_2168_),
    .A2(net1360));
 sg13g2_a22oi_1 _6018_ (.Y(_2169_),
    .B1(_2167_),
    .B2(_2168_),
    .A2(net1272),
    .A1(_0938_));
 sg13g2_a21oi_1 _6019_ (.A1(net1153),
    .A2(_2169_),
    .Y(_2170_),
    .B1(net1151));
 sg13g2_nand2b_1 _6020_ (.Y(_2171_),
    .B(\tt6581_inst.bypass_accum[8] ),
    .A_N(_2170_));
 sg13g2_xor2_1 _6021_ (.B(_2170_),
    .A(\tt6581_inst.bypass_accum[8] ),
    .X(_2172_));
 sg13g2_o21ai_1 _6022_ (.B1(_1917_),
    .Y(_2173_),
    .A1(_1951_),
    .A2(_1952_));
 sg13g2_xnor2_1 _6023_ (.Y(_2174_),
    .A(_1953_),
    .B(_2173_));
 sg13g2_a22oi_1 _6024_ (.Y(_2175_),
    .B1(net1356),
    .B2(_2174_),
    .A2(net1360),
    .A1(\tt6581_inst.svf_inst.reg_band[9] ));
 sg13g2_a221oi_1 _6025_ (.B2(\tt6581_inst.svf_inst.hp_node[9] ),
    .C1(net1152),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_low[9] ),
    .Y(_2176_),
    .A2(net1272));
 sg13g2_a21oi_2 _6026_ (.B1(_2061_),
    .Y(_2177_),
    .A2(_2176_),
    .A1(_2175_));
 sg13g2_nand2_1 _6027_ (.Y(_2178_),
    .A(\tt6581_inst.bypass_accum[9] ),
    .B(_2177_));
 sg13g2_xnor2_1 _6028_ (.Y(_2179_),
    .A(\tt6581_inst.bypass_accum[9] ),
    .B(_2177_));
 sg13g2_nor2_1 _6029_ (.A(_2172_),
    .B(_2179_),
    .Y(_2180_));
 sg13g2_nand3_1 _6030_ (.B(_2164_),
    .C(_2180_),
    .A(_2161_),
    .Y(_2181_));
 sg13g2_nand2_1 _6031_ (.Y(_2182_),
    .A(_2171_),
    .B(_2178_));
 sg13g2_o21ai_1 _6032_ (.B1(_2182_),
    .Y(_2183_),
    .A1(\tt6581_inst.bypass_accum[9] ),
    .A2(_2177_));
 sg13g2_nand2b_1 _6033_ (.Y(_2184_),
    .B(_2173_),
    .A_N(_1918_));
 sg13g2_a21o_1 _6034_ (.A2(_2184_),
    .A1(_1916_),
    .B1(_1913_),
    .X(_2185_));
 sg13g2_nand3_1 _6035_ (.B(_1916_),
    .C(_2184_),
    .A(_1913_),
    .Y(_2186_));
 sg13g2_nand3_1 _6036_ (.B(_2185_),
    .C(_2186_),
    .A(net1356),
    .Y(_2187_));
 sg13g2_a221oi_1 _6037_ (.B2(\tt6581_inst.svf_inst.hp_node[10] ),
    .C1(net1272),
    .B1(net1352),
    .A1(\tt6581_inst.svf_inst.reg_band[10] ),
    .Y(_2188_),
    .A2(net1360));
 sg13g2_a22oi_1 _6038_ (.Y(_2189_),
    .B1(_2187_),
    .B2(_2188_),
    .A2(net1272),
    .A1(_0937_));
 sg13g2_a21oi_1 _6039_ (.A1(net1154),
    .A2(_2189_),
    .Y(_2190_),
    .B1(net1152));
 sg13g2_nand2b_1 _6040_ (.Y(_2191_),
    .B(\tt6581_inst.bypass_accum[10] ),
    .A_N(_2190_));
 sg13g2_inv_1 _6041_ (.Y(_2192_),
    .A(_2191_));
 sg13g2_xnor2_1 _6042_ (.Y(_2193_),
    .A(\tt6581_inst.bypass_accum[10] ),
    .B(_2190_));
 sg13g2_inv_1 _6043_ (.Y(_2194_),
    .A(_2193_));
 sg13g2_and2_1 _6044_ (.A(_1912_),
    .B(_2185_),
    .X(_2195_));
 sg13g2_xnor2_1 _6045_ (.Y(_2196_),
    .A(_1914_),
    .B(_2195_));
 sg13g2_a22oi_1 _6046_ (.Y(_2197_),
    .B1(net1351),
    .B2(\tt6581_inst.svf_inst.hp_node[11] ),
    .A2(net1359),
    .A1(\tt6581_inst.svf_inst.reg_band[11] ));
 sg13g2_a22oi_1 _6047_ (.Y(_2198_),
    .B1(net1355),
    .B2(_2196_),
    .A2(net1269),
    .A1(\tt6581_inst.svf_inst.reg_low[11] ));
 sg13g2_nand3b_1 _6048_ (.B(_2197_),
    .C(_2198_),
    .Y(_2199_),
    .A_N(net1152));
 sg13g2_and2_1 _6049_ (.A(net1154),
    .B(_2199_),
    .X(_2200_));
 sg13g2_nor2_1 _6050_ (.A(\tt6581_inst.bypass_accum[11] ),
    .B(_2200_),
    .Y(_2201_));
 sg13g2_nand2_1 _6051_ (.Y(_2202_),
    .A(\tt6581_inst.bypass_accum[11] ),
    .B(_2200_));
 sg13g2_nor2b_1 _6052_ (.A(_2201_),
    .B_N(_2202_),
    .Y(_2203_));
 sg13g2_and2_1 _6053_ (.A(_2193_),
    .B(_2203_),
    .X(_2204_));
 sg13g2_inv_1 _6054_ (.Y(_2205_),
    .A(_2204_));
 sg13g2_a21oi_1 _6055_ (.A1(_2181_),
    .A2(_2183_),
    .Y(_2206_),
    .B1(_2205_));
 sg13g2_a21oi_1 _6056_ (.A1(_2191_),
    .A2(_2202_),
    .Y(_2207_),
    .B1(_2201_));
 sg13g2_xnor2_1 _6057_ (.Y(_2208_),
    .A(\tt6581_inst.bypass_accum[12] ),
    .B(_2097_));
 sg13g2_o21ai_1 _6058_ (.B1(_2208_),
    .Y(_2209_),
    .A1(_2206_),
    .A2(_2207_));
 sg13g2_xnor2_1 _6059_ (.Y(_2210_),
    .A(\tt6581_inst.bypass_accum[13] ),
    .B(_2002_));
 sg13g2_nand3_1 _6060_ (.B(_2209_),
    .C(_2210_),
    .A(_2098_),
    .Y(_2211_));
 sg13g2_a21oi_1 _6061_ (.A1(_2098_),
    .A2(_2209_),
    .Y(_2212_),
    .B1(_2210_));
 sg13g2_nand2_1 _6062_ (.Y(_2213_),
    .A(net1492),
    .B(_2211_));
 sg13g2_nor2_1 _6063_ (.A(_2212_),
    .B(_2213_),
    .Y(_2214_));
 sg13g2_nand3b_1 _6064_ (.B(net1492),
    .C(_2211_),
    .Y(_2215_),
    .A_N(_2212_));
 sg13g2_xor2_1 _6065_ (.B(net1145),
    .A(_1874_),
    .X(_2216_));
 sg13g2_nor2_1 _6066_ (.A(_0064_),
    .B(net1368),
    .Y(_2217_));
 sg13g2_nor2_1 _6067_ (.A(_0087_),
    .B(net1388),
    .Y(_2218_));
 sg13g2_nor2_1 _6068_ (.A(_0110_),
    .B(net1410),
    .Y(_2219_));
 sg13g2_nor3_2 _6069_ (.A(_2217_),
    .B(_2218_),
    .C(_2219_),
    .Y(_2220_));
 sg13g2_nand2_1 _6070_ (.Y(_2221_),
    .A(_1610_),
    .B(_2220_));
 sg13g2_o21ai_1 _6071_ (.B1(_2221_),
    .Y(_2222_),
    .A1(_1613_),
    .A2(_1869_));
 sg13g2_a221oi_1 _6072_ (.B2(net1215),
    .C1(_2222_),
    .B1(_2216_),
    .A1(_1616_),
    .Y(_2223_),
    .A2(net1144));
 sg13g2_nor2_1 _6073_ (.A(_1620_),
    .B(_2223_),
    .Y(_2224_));
 sg13g2_nor2_1 _6074_ (.A(_2214_),
    .B(_2224_),
    .Y(_2225_));
 sg13g2_o21ai_1 _6075_ (.B1(_2215_),
    .Y(_2226_),
    .A1(_1620_),
    .A2(_2223_));
 sg13g2_a22oi_1 _6076_ (.Y(_2227_),
    .B1(\tt6581_inst.svf_inst.reg_band[23] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[23] ),
    .A1(net1532));
 sg13g2_nor2_1 _6077_ (.A(net1434),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_nor2_1 _6078_ (.A(net1143),
    .B(_2228_),
    .Y(_2229_));
 sg13g2_or2_1 _6079_ (.X(_2230_),
    .B(_2228_),
    .A(net1143));
 sg13g2_nand2_1 _6080_ (.Y(_2231_),
    .A(_2074_),
    .B(net1140));
 sg13g2_xnor2_1 _6081_ (.Y(_2232_),
    .A(_2090_),
    .B(_2231_));
 sg13g2_nor2_1 _6082_ (.A(net1439),
    .B(net817),
    .Y(_2233_));
 sg13g2_nor2_1 _6083_ (.A(net1224),
    .B(_2233_),
    .Y(_2234_));
 sg13g2_o21ai_1 _6084_ (.B1(_2234_),
    .Y(_2235_),
    .A1(net1538),
    .A2(_2232_));
 sg13g2_o21ai_1 _6085_ (.B1(_2235_),
    .Y(_0300_),
    .A1(_0978_),
    .A2(net1194));
 sg13g2_xor2_1 _6086_ (.B(net1145),
    .A(_1822_),
    .X(_2236_));
 sg13g2_nor2_1 _6087_ (.A(_1613_),
    .B(_1816_),
    .Y(_2237_));
 sg13g2_a22oi_1 _6088_ (.Y(_2238_),
    .B1(net1393),
    .B2(_0836_),
    .A2(net1417),
    .A1(_0833_));
 sg13g2_o21ai_1 _6089_ (.B1(_2238_),
    .Y(_2239_),
    .A1(_0044_),
    .A2(net1367));
 sg13g2_a221oi_1 _6090_ (.B2(_1610_),
    .C1(_2237_),
    .B1(_2239_),
    .A1(net1215),
    .Y(_2240_),
    .A2(_2236_));
 sg13g2_o21ai_1 _6091_ (.B1(_2240_),
    .Y(_2241_),
    .A1(_1615_),
    .A2(net1144));
 sg13g2_xnor2_1 _6092_ (.Y(_2242_),
    .A(_2113_),
    .B(_2115_));
 sg13g2_nand2_1 _6093_ (.Y(_2243_),
    .A(net1492),
    .B(_2242_));
 sg13g2_a22oi_1 _6094_ (.Y(_2244_),
    .B1(\tt6581_inst.svf_inst.reg_band[2] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[2] ),
    .A1(net1534));
 sg13g2_o21ai_1 _6095_ (.B1(_2243_),
    .Y(_2245_),
    .A1(net1435),
    .A2(_2244_));
 sg13g2_a21o_1 _6096_ (.A2(_2241_),
    .A1(_1619_),
    .B1(_2245_),
    .X(_2246_));
 sg13g2_inv_1 _6097_ (.Y(_2247_),
    .A(_2246_));
 sg13g2_nor2_1 _6098_ (.A(_2074_),
    .B(_2090_),
    .Y(_2248_));
 sg13g2_a21oi_1 _6099_ (.A1(_2247_),
    .A2(_2248_),
    .Y(_2249_),
    .B1(net1141));
 sg13g2_o21ai_1 _6100_ (.B1(_2249_),
    .Y(_2250_),
    .A1(_2247_),
    .A2(_2248_));
 sg13g2_a21oi_1 _6101_ (.A1(net1142),
    .A2(_2246_),
    .Y(_2251_),
    .B1(net1538));
 sg13g2_a221oi_1 _6102_ (.B2(_2251_),
    .C1(net1226),
    .B1(_2250_),
    .A1(net1538),
    .Y(_2252_),
    .A2(_0978_));
 sg13g2_a21o_1 _6103_ (.A2(net1226),
    .A1(net541),
    .B1(_2252_),
    .X(_0301_));
 sg13g2_nand2_1 _6104_ (.Y(_2253_),
    .A(net273),
    .B(net1226));
 sg13g2_xnor2_1 _6105_ (.Y(_2254_),
    .A(_1816_),
    .B(net1145));
 sg13g2_a22oi_1 _6106_ (.Y(_2255_),
    .B1(net1393),
    .B2(_0835_),
    .A2(net1417),
    .A1(_0832_));
 sg13g2_o21ai_1 _6107_ (.B1(_2255_),
    .Y(_2256_),
    .A1(_0046_),
    .A2(net1364));
 sg13g2_nor2_1 _6108_ (.A(_1613_),
    .B(_1810_),
    .Y(_2257_));
 sg13g2_a221oi_1 _6109_ (.B2(_1610_),
    .C1(_2257_),
    .B1(_2256_),
    .A1(net1215),
    .Y(_2258_),
    .A2(_2254_));
 sg13g2_o21ai_1 _6110_ (.B1(_2258_),
    .Y(_2259_),
    .A1(_1615_),
    .A2(_1882_));
 sg13g2_xnor2_1 _6111_ (.Y(_2260_),
    .A(_2116_),
    .B(_2118_));
 sg13g2_nand2_1 _6112_ (.Y(_2261_),
    .A(net1492),
    .B(_2260_));
 sg13g2_a22oi_1 _6113_ (.Y(_2262_),
    .B1(\tt6581_inst.svf_inst.reg_band[3] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[3] ),
    .A1(net1534));
 sg13g2_o21ai_1 _6114_ (.B1(_2261_),
    .Y(_2263_),
    .A1(net1435),
    .A2(_2262_));
 sg13g2_a21o_1 _6115_ (.A2(_2259_),
    .A1(_1619_),
    .B1(_2263_),
    .X(_2264_));
 sg13g2_xnor2_1 _6116_ (.Y(_2265_),
    .A(_2249_),
    .B(_2264_));
 sg13g2_nand2_1 _6117_ (.Y(_2266_),
    .A(net1441),
    .B(_2265_));
 sg13g2_o21ai_1 _6118_ (.B1(_2266_),
    .Y(_2267_),
    .A1(net1441),
    .A2(\tt6581_inst.mult_inst.a_reg[2] ));
 sg13g2_o21ai_1 _6119_ (.B1(_2253_),
    .Y(_0302_),
    .A1(net1226),
    .A2(_2267_));
 sg13g2_nand2_1 _6120_ (.Y(_2268_),
    .A(net224),
    .B(net1226));
 sg13g2_xnor2_1 _6121_ (.Y(_2269_),
    .A(_1810_),
    .B(net1145));
 sg13g2_nor2_1 _6122_ (.A(_0049_),
    .B(net1364),
    .Y(_2270_));
 sg13g2_nor2_1 _6123_ (.A(_0072_),
    .B(net1385),
    .Y(_2271_));
 sg13g2_nor2_1 _6124_ (.A(_0095_),
    .B(net1406),
    .Y(_2272_));
 sg13g2_nor3_2 _6125_ (.A(_2270_),
    .B(_2271_),
    .C(_2272_),
    .Y(_2273_));
 sg13g2_nand2b_1 _6126_ (.Y(_2274_),
    .B(_1610_),
    .A_N(_2273_));
 sg13g2_o21ai_1 _6127_ (.B1(_2274_),
    .Y(_2275_),
    .A1(_1613_),
    .A2(_1804_));
 sg13g2_a21oi_1 _6128_ (.A1(net1215),
    .A2(_2269_),
    .Y(_2276_),
    .B1(_2275_));
 sg13g2_o21ai_1 _6129_ (.B1(_2276_),
    .Y(_2277_),
    .A1(net1190),
    .A2(net1144));
 sg13g2_nand2b_1 _6130_ (.Y(_2278_),
    .B(_2119_),
    .A_N(_2138_));
 sg13g2_nor2b_1 _6131_ (.A(_2119_),
    .B_N(_2138_),
    .Y(_2279_));
 sg13g2_nor2_1 _6132_ (.A(_0916_),
    .B(_2279_),
    .Y(_2280_));
 sg13g2_a22oi_1 _6133_ (.Y(_2281_),
    .B1(\tt6581_inst.svf_inst.reg_band[4] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[4] ),
    .A1(net1534));
 sg13g2_nor2_1 _6134_ (.A(net1435),
    .B(_2281_),
    .Y(_2282_));
 sg13g2_a221oi_1 _6135_ (.B2(_2280_),
    .C1(_2282_),
    .B1(_2278_),
    .A1(_1619_),
    .Y(_2283_),
    .A2(_2277_));
 sg13g2_nor4_2 _6136_ (.A(_2074_),
    .B(_2090_),
    .C(_2246_),
    .Y(_2284_),
    .D(_2264_));
 sg13g2_nor2_1 _6137_ (.A(net1142),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_xnor2_1 _6138_ (.Y(_2286_),
    .A(_2283_),
    .B(_2285_));
 sg13g2_nor2_1 _6139_ (.A(net1539),
    .B(_2286_),
    .Y(_2287_));
 sg13g2_o21ai_1 _6140_ (.B1(net1198),
    .Y(_2288_),
    .A1(net1441),
    .A2(\tt6581_inst.mult_inst.a_reg[3] ));
 sg13g2_o21ai_1 _6141_ (.B1(_2268_),
    .Y(_0303_),
    .A1(_2287_),
    .A2(_2288_));
 sg13g2_nand2_1 _6142_ (.Y(_2289_),
    .A(net206),
    .B(net1226));
 sg13g2_xnor2_1 _6143_ (.Y(_2290_),
    .A(_1804_),
    .B(net1145));
 sg13g2_nor2_1 _6144_ (.A(_0053_),
    .B(net1366),
    .Y(_2291_));
 sg13g2_nor2_1 _6145_ (.A(_0076_),
    .B(net1387),
    .Y(_2292_));
 sg13g2_nor2_1 _6146_ (.A(_0099_),
    .B(net1408),
    .Y(_2293_));
 sg13g2_nor3_2 _6147_ (.A(_2291_),
    .B(_2292_),
    .C(_2293_),
    .Y(_2294_));
 sg13g2_nand2b_1 _6148_ (.Y(_2295_),
    .B(_1610_),
    .A_N(_2294_));
 sg13g2_o21ai_1 _6149_ (.B1(_2295_),
    .Y(_2296_),
    .A1(_1613_),
    .A2(_1797_));
 sg13g2_a21o_1 _6150_ (.A2(_2290_),
    .A1(net1215),
    .B1(_2296_),
    .X(_2297_));
 sg13g2_o21ai_1 _6151_ (.B1(_1619_),
    .Y(_2298_),
    .A1(_1884_),
    .A2(_2297_));
 sg13g2_a22oi_1 _6152_ (.Y(_2299_),
    .B1(\tt6581_inst.svf_inst.reg_band[5] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[5] ),
    .A1(net1534));
 sg13g2_nor2_1 _6153_ (.A(net1435),
    .B(_2299_),
    .Y(_2300_));
 sg13g2_nor2_1 _6154_ (.A(_2137_),
    .B(_2279_),
    .Y(_2301_));
 sg13g2_xnor2_1 _6155_ (.Y(_2302_),
    .A(_2129_),
    .B(_2301_));
 sg13g2_a21oi_2 _6156_ (.B1(_2300_),
    .Y(_2303_),
    .A2(_2302_),
    .A1(net1493));
 sg13g2_nand2_1 _6157_ (.Y(_2304_),
    .A(_2298_),
    .B(_2303_));
 sg13g2_a21oi_1 _6158_ (.A1(_2283_),
    .A2(_2284_),
    .Y(_2305_),
    .B1(net1142));
 sg13g2_xor2_1 _6159_ (.B(_2305_),
    .A(_2304_),
    .X(_2306_));
 sg13g2_nor2_1 _6160_ (.A(net1539),
    .B(_2306_),
    .Y(_2307_));
 sg13g2_o21ai_1 _6161_ (.B1(net1198),
    .Y(_2308_),
    .A1(net1441),
    .A2(\tt6581_inst.mult_inst.a_reg[4] ));
 sg13g2_o21ai_1 _6162_ (.B1(_2289_),
    .Y(_0304_),
    .A1(_2307_),
    .A2(_2308_));
 sg13g2_xnor2_1 _6163_ (.Y(_2309_),
    .A(_1797_),
    .B(_1889_));
 sg13g2_nor2_1 _6164_ (.A(_0055_),
    .B(net1366),
    .Y(_2310_));
 sg13g2_nor2_1 _6165_ (.A(_0078_),
    .B(net1387),
    .Y(_2311_));
 sg13g2_nor2_1 _6166_ (.A(_0101_),
    .B(net1408),
    .Y(_2312_));
 sg13g2_nor3_2 _6167_ (.A(_2310_),
    .B(_2311_),
    .C(_2312_),
    .Y(_2313_));
 sg13g2_nor3_1 _6168_ (.A(_1608_),
    .B(_1609_),
    .C(_2313_),
    .Y(_2314_));
 sg13g2_a221oi_1 _6169_ (.B2(_1617_),
    .C1(_2314_),
    .B1(_2309_),
    .A1(_1612_),
    .Y(_2315_),
    .A2(_1793_));
 sg13g2_o21ai_1 _6170_ (.B1(_2315_),
    .Y(_2316_),
    .A1(net1190),
    .A2(net1144));
 sg13g2_and2_1 _6171_ (.A(_2158_),
    .B(_2162_),
    .X(_2317_));
 sg13g2_o21ai_1 _6172_ (.B1(_2317_),
    .Y(_2318_),
    .A1(_2140_),
    .A2(_2142_));
 sg13g2_nor3_1 _6173_ (.A(_2140_),
    .B(_2142_),
    .C(_2317_),
    .Y(_2319_));
 sg13g2_nor2_1 _6174_ (.A(_0916_),
    .B(_2319_),
    .Y(_2320_));
 sg13g2_a22oi_1 _6175_ (.Y(_2321_),
    .B1(\tt6581_inst.svf_inst.reg_band[6] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[6] ),
    .A1(net1534));
 sg13g2_nor2_1 _6176_ (.A(net1435),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_a221oi_1 _6177_ (.B2(_2320_),
    .C1(_2322_),
    .B1(_2318_),
    .A1(_1619_),
    .Y(_2323_),
    .A2(_2316_));
 sg13g2_and3_2 _6178_ (.X(_2324_),
    .A(_2283_),
    .B(_2298_),
    .C(_2303_));
 sg13g2_a21oi_1 _6179_ (.A1(_2284_),
    .A2(_2324_),
    .Y(_2325_),
    .B1(net1142));
 sg13g2_xor2_1 _6180_ (.B(_2325_),
    .A(_2323_),
    .X(_2326_));
 sg13g2_nand3_1 _6181_ (.B(_2323_),
    .C(_2324_),
    .A(_2284_),
    .Y(_2327_));
 sg13g2_nor2_1 _6182_ (.A(net1441),
    .B(net206),
    .Y(_2328_));
 sg13g2_a21oi_1 _6183_ (.A1(net1441),
    .A2(_2326_),
    .Y(_2329_),
    .B1(_2328_));
 sg13g2_mux2_1 _6184_ (.A0(net755),
    .A1(_2329_),
    .S(net1193),
    .X(_0305_));
 sg13g2_nand2_1 _6185_ (.Y(_2330_),
    .A(net271),
    .B(net1227));
 sg13g2_xnor2_1 _6186_ (.Y(_2331_),
    .A(_1794_),
    .B(_1889_));
 sg13g2_nor2_1 _6187_ (.A(_0058_),
    .B(net1364),
    .Y(_2332_));
 sg13g2_nor2_1 _6188_ (.A(_0081_),
    .B(net1385),
    .Y(_2333_));
 sg13g2_nor2_1 _6189_ (.A(_0104_),
    .B(net1406),
    .Y(_2334_));
 sg13g2_nor3_2 _6190_ (.A(_2332_),
    .B(_2333_),
    .C(_2334_),
    .Y(_2335_));
 sg13g2_nor3_1 _6191_ (.A(_1608_),
    .B(_1609_),
    .C(_2335_),
    .Y(_2336_));
 sg13g2_a221oi_1 _6192_ (.B2(_1617_),
    .C1(_2336_),
    .B1(_2331_),
    .A1(_1612_),
    .Y(_2337_),
    .A2(_1785_));
 sg13g2_o21ai_1 _6193_ (.B1(_2337_),
    .Y(_2338_),
    .A1(net1190),
    .A2(net1144));
 sg13g2_nand2_1 _6194_ (.Y(_2339_),
    .A(_2151_),
    .B(_2152_));
 sg13g2_and2_1 _6195_ (.A(_2158_),
    .B(_2318_),
    .X(_2340_));
 sg13g2_o21ai_1 _6196_ (.B1(net1492),
    .Y(_2341_),
    .A1(_2339_),
    .A2(_2340_));
 sg13g2_a21oi_1 _6197_ (.A1(_2339_),
    .A2(_2340_),
    .Y(_2342_),
    .B1(_2341_));
 sg13g2_a22oi_1 _6198_ (.Y(_2343_),
    .B1(\tt6581_inst.svf_inst.reg_band[7] ),
    .B2(net1429),
    .A2(\tt6581_inst.svf_inst.hp_node[7] ),
    .A1(net1534));
 sg13g2_inv_1 _6199_ (.Y(_2344_),
    .A(_2343_));
 sg13g2_a221oi_1 _6200_ (.B2(net1490),
    .C1(_2342_),
    .B1(_2344_),
    .A1(_1619_),
    .Y(_2345_),
    .A2(_2338_));
 sg13g2_and3_1 _6201_ (.X(_2346_),
    .A(net1140),
    .B(_2327_),
    .C(_2345_));
 sg13g2_a21oi_1 _6202_ (.A1(net1140),
    .A2(_2327_),
    .Y(_2347_),
    .B1(_2345_));
 sg13g2_nor3_1 _6203_ (.A(net1539),
    .B(_2346_),
    .C(_2347_),
    .Y(_2348_));
 sg13g2_o21ai_1 _6204_ (.B1(net1193),
    .Y(_2349_),
    .A1(net1440),
    .A2(\tt6581_inst.mult_inst.a_reg[6] ));
 sg13g2_o21ai_1 _6205_ (.B1(_2330_),
    .Y(_0306_),
    .A1(_2348_),
    .A2(_2349_));
 sg13g2_xor2_1 _6206_ (.B(net1145),
    .A(_1785_),
    .X(_2350_));
 sg13g2_a22oi_1 _6207_ (.Y(_2351_),
    .B1(net1395),
    .B2(_0834_),
    .A2(net1417),
    .A1(_0831_));
 sg13g2_o21ai_1 _6208_ (.B1(_2351_),
    .Y(_2352_),
    .A1(_0062_),
    .A2(net1368));
 sg13g2_nand2_1 _6209_ (.Y(_2353_),
    .A(_1610_),
    .B(_2352_));
 sg13g2_o21ai_1 _6210_ (.B1(_2353_),
    .Y(_2354_),
    .A1(_1613_),
    .A2(_1874_));
 sg13g2_a221oi_1 _6211_ (.B2(_1617_),
    .C1(_2354_),
    .B1(_2350_),
    .A1(_1616_),
    .Y(_2355_),
    .A2(_1883_));
 sg13g2_a22oi_1 _6212_ (.Y(_2356_),
    .B1(\tt6581_inst.svf_inst.reg_band[8] ),
    .B2(net1430),
    .A2(\tt6581_inst.svf_inst.hp_node[8] ),
    .A1(net1535));
 sg13g2_inv_1 _6213_ (.Y(_2357_),
    .A(_2356_));
 sg13g2_or2_1 _6214_ (.X(_2358_),
    .B(_2172_),
    .A(_2165_));
 sg13g2_a21oi_1 _6215_ (.A1(_2165_),
    .A2(_2172_),
    .Y(_2359_),
    .B1(_0916_));
 sg13g2_a22oi_1 _6216_ (.Y(_2360_),
    .B1(_2358_),
    .B2(_2359_),
    .A2(_2357_),
    .A1(net1490));
 sg13g2_o21ai_1 _6217_ (.B1(_2360_),
    .Y(_2361_),
    .A1(_1620_),
    .A2(_2355_));
 sg13g2_and2_1 _6218_ (.A(_2323_),
    .B(_2345_),
    .X(_2362_));
 sg13g2_nand3_1 _6219_ (.B(_2324_),
    .C(_2362_),
    .A(_2284_),
    .Y(_2363_));
 sg13g2_o21ai_1 _6220_ (.B1(net1140),
    .Y(_2364_),
    .A1(_2361_),
    .A2(_2363_));
 sg13g2_a21oi_1 _6221_ (.A1(_2361_),
    .A2(_2363_),
    .Y(_2365_),
    .B1(_2364_));
 sg13g2_a21oi_1 _6222_ (.A1(net1142),
    .A2(_2361_),
    .Y(_2366_),
    .B1(_2365_));
 sg13g2_o21ai_1 _6223_ (.B1(net1193),
    .Y(_2367_),
    .A1(net1440),
    .A2(net271));
 sg13g2_a21o_1 _6224_ (.A2(_2366_),
    .A1(net1440),
    .B1(_2367_),
    .X(_2368_));
 sg13g2_o21ai_1 _6225_ (.B1(_2368_),
    .Y(_0307_),
    .A1(_0979_),
    .A2(net1194));
 sg13g2_a22oi_1 _6226_ (.Y(_2369_),
    .B1(\tt6581_inst.svf_inst.reg_band[9] ),
    .B2(net1430),
    .A2(\tt6581_inst.svf_inst.hp_node[9] ),
    .A1(net1535));
 sg13g2_nor2_1 _6227_ (.A(net1435),
    .B(_2369_),
    .Y(_2370_));
 sg13g2_nand3_1 _6228_ (.B(_2179_),
    .C(_2358_),
    .A(_2171_),
    .Y(_2371_));
 sg13g2_a21o_1 _6229_ (.A2(_2358_),
    .A1(_2171_),
    .B1(_2179_),
    .X(_2372_));
 sg13g2_and2_1 _6230_ (.A(net1492),
    .B(_2371_),
    .X(_2373_));
 sg13g2_a21oi_1 _6231_ (.A1(_2372_),
    .A2(_2373_),
    .Y(_2374_),
    .B1(_2370_));
 sg13g2_o21ai_1 _6232_ (.B1(_2374_),
    .Y(_2375_),
    .A1(_1620_),
    .A2(_2223_));
 sg13g2_xnor2_1 _6233_ (.Y(_2376_),
    .A(_2364_),
    .B(_2375_));
 sg13g2_a21oi_1 _6234_ (.A1(net1539),
    .A2(_0979_),
    .Y(_2377_),
    .B1(net1226));
 sg13g2_o21ai_1 _6235_ (.B1(_2377_),
    .Y(_2378_),
    .A1(net1539),
    .A2(_2376_));
 sg13g2_o21ai_1 _6236_ (.B1(_2378_),
    .Y(_0308_),
    .A1(_0980_),
    .A2(net1193));
 sg13g2_a22oi_1 _6237_ (.Y(_2379_),
    .B1(\tt6581_inst.svf_inst.reg_band[10] ),
    .B2(net1430),
    .A2(\tt6581_inst.svf_inst.hp_node[10] ),
    .A1(net1535));
 sg13g2_inv_1 _6238_ (.Y(_2380_),
    .A(_2379_));
 sg13g2_nand3_1 _6239_ (.B(_2183_),
    .C(_2194_),
    .A(_2181_),
    .Y(_2381_));
 sg13g2_a21oi_1 _6240_ (.A1(_2181_),
    .A2(_2183_),
    .Y(_2382_),
    .B1(_2194_));
 sg13g2_nor2_1 _6241_ (.A(_0916_),
    .B(_2382_),
    .Y(_2383_));
 sg13g2_a22oi_1 _6242_ (.Y(_2384_),
    .B1(_2381_),
    .B2(_2383_),
    .A2(_2380_),
    .A1(net1491));
 sg13g2_o21ai_1 _6243_ (.B1(_2384_),
    .Y(_2385_),
    .A1(_1620_),
    .A2(_2223_));
 sg13g2_or3_1 _6244_ (.A(_2361_),
    .B(_2363_),
    .C(_2375_),
    .X(_2386_));
 sg13g2_nand2_1 _6245_ (.Y(_2387_),
    .A(net1140),
    .B(_2386_));
 sg13g2_o21ai_1 _6246_ (.B1(_2230_),
    .Y(_2388_),
    .A1(_2385_),
    .A2(_2386_));
 sg13g2_xnor2_1 _6247_ (.Y(_2389_),
    .A(_2385_),
    .B(_2387_));
 sg13g2_a21oi_1 _6248_ (.A1(net1541),
    .A2(_0980_),
    .Y(_2390_),
    .B1(net1227));
 sg13g2_o21ai_1 _6249_ (.B1(_2390_),
    .Y(_2391_),
    .A1(net1539),
    .A2(_2389_));
 sg13g2_o21ai_1 _6250_ (.B1(_2391_),
    .Y(_0309_),
    .A1(_0981_),
    .A2(net1197));
 sg13g2_nor3_1 _6251_ (.A(_2192_),
    .B(_2203_),
    .C(_2382_),
    .Y(_2392_));
 sg13g2_o21ai_1 _6252_ (.B1(_2203_),
    .Y(_2393_),
    .A1(_2192_),
    .A2(_2382_));
 sg13g2_nor2_1 _6253_ (.A(_0916_),
    .B(_2392_),
    .Y(_2394_));
 sg13g2_a22oi_1 _6254_ (.Y(_2395_),
    .B1(\tt6581_inst.svf_inst.reg_band[11] ),
    .B2(net1428),
    .A2(\tt6581_inst.svf_inst.hp_node[11] ),
    .A1(net1533));
 sg13g2_nor2_1 _6255_ (.A(net1437),
    .B(_2395_),
    .Y(_2396_));
 sg13g2_a21oi_1 _6256_ (.A1(_2393_),
    .A2(_2394_),
    .Y(_2397_),
    .B1(_2396_));
 sg13g2_o21ai_1 _6257_ (.B1(_2397_),
    .Y(_2398_),
    .A1(_1620_),
    .A2(_2223_));
 sg13g2_xor2_1 _6258_ (.B(_2398_),
    .A(_2388_),
    .X(_2399_));
 sg13g2_o21ai_1 _6259_ (.B1(net1197),
    .Y(_2400_),
    .A1(net1440),
    .A2(\tt6581_inst.mult_inst.a_reg[10] ));
 sg13g2_a21oi_1 _6260_ (.A1(net1440),
    .A2(_2399_),
    .Y(_2401_),
    .B1(_2400_));
 sg13g2_a21o_1 _6261_ (.A2(net1227),
    .A1(net529),
    .B1(_2401_),
    .X(_0310_));
 sg13g2_or3_1 _6262_ (.A(_2206_),
    .B(_2207_),
    .C(_2208_),
    .X(_2402_));
 sg13g2_and2_1 _6263_ (.A(net1492),
    .B(_2209_),
    .X(_2403_));
 sg13g2_a22oi_1 _6264_ (.Y(_2404_),
    .B1(\tt6581_inst.svf_inst.reg_band[12] ),
    .B2(net1428),
    .A2(\tt6581_inst.svf_inst.hp_node[12] ),
    .A1(net1533));
 sg13g2_inv_1 _6265_ (.Y(_2405_),
    .A(_2404_));
 sg13g2_a22oi_1 _6266_ (.Y(_2406_),
    .B1(_2405_),
    .B2(net1491),
    .A2(_2403_),
    .A1(_2402_));
 sg13g2_o21ai_1 _6267_ (.B1(_2406_),
    .Y(_2407_),
    .A1(_1620_),
    .A2(_2223_));
 sg13g2_nor4_1 _6268_ (.A(_2361_),
    .B(_2375_),
    .C(_2385_),
    .D(_2398_),
    .Y(_2408_));
 sg13g2_nand4_1 _6269_ (.B(_2324_),
    .C(_2362_),
    .A(_2284_),
    .Y(_2409_),
    .D(_2408_));
 sg13g2_o21ai_1 _6270_ (.B1(net1140),
    .Y(_2410_),
    .A1(_2407_),
    .A2(_2409_));
 sg13g2_a21oi_1 _6271_ (.A1(_2407_),
    .A2(_2409_),
    .Y(_2411_),
    .B1(_2410_));
 sg13g2_a21o_1 _6272_ (.A2(_2407_),
    .A1(net1142),
    .B1(_2411_),
    .X(_2412_));
 sg13g2_a21oi_1 _6273_ (.A1(net1540),
    .A2(_0982_),
    .Y(_2413_),
    .B1(net1227));
 sg13g2_o21ai_1 _6274_ (.B1(_2413_),
    .Y(_2414_),
    .A1(net1540),
    .A2(_2412_));
 sg13g2_o21ai_1 _6275_ (.B1(_2414_),
    .Y(_0311_),
    .A1(_0983_),
    .A2(net1193));
 sg13g2_a22oi_1 _6276_ (.Y(_2415_),
    .B1(\tt6581_inst.svf_inst.reg_band[13] ),
    .B2(net1428),
    .A2(\tt6581_inst.svf_inst.hp_node[13] ),
    .A1(net1533));
 sg13g2_nor2_1 _6277_ (.A(net1437),
    .B(_2415_),
    .Y(_2416_));
 sg13g2_nor2_1 _6278_ (.A(_2226_),
    .B(_2416_),
    .Y(_2417_));
 sg13g2_xnor2_1 _6279_ (.Y(_2418_),
    .A(_2410_),
    .B(_2417_));
 sg13g2_o21ai_1 _6280_ (.B1(net1193),
    .Y(_2419_),
    .A1(net1440),
    .A2(\tt6581_inst.mult_inst.a_reg[12] ));
 sg13g2_a21oi_1 _6281_ (.A1(net1440),
    .A2(_2418_),
    .Y(_2420_),
    .B1(_2419_));
 sg13g2_a21o_1 _6282_ (.A2(net1226),
    .A1(net579),
    .B1(_2420_),
    .X(_0312_));
 sg13g2_a22oi_1 _6283_ (.Y(_2421_),
    .B1(\tt6581_inst.svf_inst.reg_band[14] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[14] ),
    .A1(net1532));
 sg13g2_nor2_1 _6284_ (.A(net1434),
    .B(_2421_),
    .Y(_2422_));
 sg13g2_nor3_2 _6285_ (.A(_2214_),
    .B(_2224_),
    .C(_2422_),
    .Y(_2423_));
 sg13g2_nor3_1 _6286_ (.A(net1143),
    .B(_2407_),
    .C(_2416_),
    .Y(_2424_));
 sg13g2_nor2b_1 _6287_ (.A(_2409_),
    .B_N(_2424_),
    .Y(_2425_));
 sg13g2_nor2_1 _6288_ (.A(net1142),
    .B(_2425_),
    .Y(_2426_));
 sg13g2_a21oi_1 _6289_ (.A1(_2423_),
    .A2(_2425_),
    .Y(_2427_),
    .B1(_2229_));
 sg13g2_xnor2_1 _6290_ (.Y(_2428_),
    .A(_2423_),
    .B(_2426_));
 sg13g2_a21oi_1 _6291_ (.A1(net1540),
    .A2(_0984_),
    .Y(_2429_),
    .B1(net1228));
 sg13g2_o21ai_1 _6292_ (.B1(_2429_),
    .Y(_2430_),
    .A1(net1540),
    .A2(_2428_));
 sg13g2_o21ai_1 _6293_ (.B1(_2430_),
    .Y(_0313_),
    .A1(_0985_),
    .A2(net1193));
 sg13g2_a22oi_1 _6294_ (.Y(_2431_),
    .B1(\tt6581_inst.svf_inst.reg_band[15] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[15] ),
    .A1(net1532));
 sg13g2_inv_1 _6295_ (.Y(_2432_),
    .A(_2431_));
 sg13g2_a21oi_1 _6296_ (.A1(net1491),
    .A2(_2432_),
    .Y(_2433_),
    .B1(_2226_));
 sg13g2_xnor2_1 _6297_ (.Y(_2434_),
    .A(_2427_),
    .B(_2433_));
 sg13g2_a21oi_1 _6298_ (.A1(net1539),
    .A2(_0985_),
    .Y(_2435_),
    .B1(net1228));
 sg13g2_o21ai_1 _6299_ (.B1(_2435_),
    .Y(_2436_),
    .A1(net1539),
    .A2(_2434_));
 sg13g2_o21ai_1 _6300_ (.B1(_2436_),
    .Y(_0314_),
    .A1(_0986_),
    .A2(net1193));
 sg13g2_a22oi_1 _6301_ (.Y(_2437_),
    .B1(\tt6581_inst.svf_inst.reg_band[16] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[16] ),
    .A1(net1532));
 sg13g2_nor2_1 _6302_ (.A(net1434),
    .B(_2437_),
    .Y(_2438_));
 sg13g2_nor2_1 _6303_ (.A(net1143),
    .B(_2438_),
    .Y(_2439_));
 sg13g2_nand4_1 _6304_ (.B(_2423_),
    .C(_2424_),
    .A(_2408_),
    .Y(_2440_),
    .D(_2433_));
 sg13g2_nor2_1 _6305_ (.A(_2363_),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_inv_1 _6306_ (.Y(_2442_),
    .A(_2441_));
 sg13g2_a21oi_1 _6307_ (.A1(_2439_),
    .A2(_2441_),
    .Y(_2443_),
    .B1(net1141));
 sg13g2_o21ai_1 _6308_ (.B1(_2443_),
    .Y(_2444_),
    .A1(_2439_),
    .A2(_2441_));
 sg13g2_a21oi_1 _6309_ (.A1(net1141),
    .A2(_2438_),
    .Y(_2445_),
    .B1(net1537));
 sg13g2_a221oi_1 _6310_ (.B2(_2445_),
    .C1(net1223),
    .B1(_2444_),
    .A1(net1537),
    .Y(_2446_),
    .A2(_0986_));
 sg13g2_a21o_1 _6311_ (.A2(net1223),
    .A1(net1060),
    .B1(_2446_),
    .X(_0315_));
 sg13g2_nand2_1 _6312_ (.Y(_2447_),
    .A(net368),
    .B(net1223));
 sg13g2_a22oi_1 _6313_ (.Y(_2448_),
    .B1(\tt6581_inst.svf_inst.reg_band[17] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[17] ),
    .A1(net1532));
 sg13g2_nor2_1 _6314_ (.A(net1434),
    .B(_2448_),
    .Y(_2449_));
 sg13g2_or2_1 _6315_ (.X(_2450_),
    .B(_2449_),
    .A(net1143));
 sg13g2_xor2_1 _6316_ (.B(_2450_),
    .A(_2443_),
    .X(_2451_));
 sg13g2_nor2_1 _6317_ (.A(net1537),
    .B(_2451_),
    .Y(_2452_));
 sg13g2_o21ai_1 _6318_ (.B1(net1192),
    .Y(_2453_),
    .A1(net1439),
    .A2(\tt6581_inst.mult_inst.a_reg[16] ));
 sg13g2_o21ai_1 _6319_ (.B1(_2447_),
    .Y(_0316_),
    .A1(_2452_),
    .A2(_2453_));
 sg13g2_nand2_1 _6320_ (.Y(_2454_),
    .A(net209),
    .B(net1223));
 sg13g2_a22oi_1 _6321_ (.Y(_2455_),
    .B1(\tt6581_inst.svf_inst.reg_band[18] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[18] ),
    .A1(net1532));
 sg13g2_nor2_1 _6322_ (.A(net1434),
    .B(_2455_),
    .Y(_2456_));
 sg13g2_nor2_1 _6323_ (.A(net1143),
    .B(_2456_),
    .Y(_2457_));
 sg13g2_or2_1 _6324_ (.X(_2458_),
    .B(_2456_),
    .A(net1143));
 sg13g2_nor4_1 _6325_ (.A(_2363_),
    .B(_2438_),
    .C(_2440_),
    .D(_2450_),
    .Y(_2459_));
 sg13g2_a21oi_1 _6326_ (.A1(_2457_),
    .A2(_2459_),
    .Y(_2460_),
    .B1(net1141));
 sg13g2_or2_1 _6327_ (.X(_2461_),
    .B(_2459_),
    .A(_2457_));
 sg13g2_a221oi_1 _6328_ (.B2(_2461_),
    .C1(net1537),
    .B1(_2460_),
    .A1(net1141),
    .Y(_2462_),
    .A2(_2458_));
 sg13g2_o21ai_1 _6329_ (.B1(net1192),
    .Y(_2463_),
    .A1(net1438),
    .A2(\tt6581_inst.mult_inst.a_reg[17] ));
 sg13g2_o21ai_1 _6330_ (.B1(_2454_),
    .Y(_0317_),
    .A1(_2462_),
    .A2(_2463_));
 sg13g2_a22oi_1 _6331_ (.Y(_2464_),
    .B1(\tt6581_inst.svf_inst.reg_band[19] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[19] ),
    .A1(net1532));
 sg13g2_nor2_1 _6332_ (.A(net1434),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nor2_1 _6333_ (.A(net1143),
    .B(_2465_),
    .Y(_2466_));
 sg13g2_xor2_1 _6334_ (.B(_2466_),
    .A(_2460_),
    .X(_2467_));
 sg13g2_o21ai_1 _6335_ (.B1(net1192),
    .Y(_2468_),
    .A1(net1438),
    .A2(net209));
 sg13g2_a21oi_1 _6336_ (.A1(net1438),
    .A2(_2467_),
    .Y(_2469_),
    .B1(_2468_));
 sg13g2_a21o_1 _6337_ (.A2(net1224),
    .A1(net630),
    .B1(_2469_),
    .X(_0318_));
 sg13g2_nand2_1 _6338_ (.Y(_2470_),
    .A(net243),
    .B(net1223));
 sg13g2_a22oi_1 _6339_ (.Y(_2471_),
    .B1(\tt6581_inst.svf_inst.reg_band[20] ),
    .B2(net1427),
    .A2(\tt6581_inst.svf_inst.hp_node[20] ),
    .A1(net1532));
 sg13g2_o21ai_1 _6340_ (.B1(_2225_),
    .Y(_2472_),
    .A1(net1434),
    .A2(_2471_));
 sg13g2_or4_1 _6341_ (.A(_2438_),
    .B(_2450_),
    .C(_2458_),
    .D(_2465_),
    .X(_2473_));
 sg13g2_nor4_1 _6342_ (.A(_2363_),
    .B(_2440_),
    .C(_2472_),
    .D(_2473_),
    .Y(_2474_));
 sg13g2_nor2_1 _6343_ (.A(net1141),
    .B(_2474_),
    .Y(_2475_));
 sg13g2_o21ai_1 _6344_ (.B1(_2472_),
    .Y(_2476_),
    .A1(_2442_),
    .A2(_2473_));
 sg13g2_a221oi_1 _6345_ (.B2(_2476_),
    .C1(net1537),
    .B1(_2475_),
    .A1(net1141),
    .Y(_2477_),
    .A2(_2472_));
 sg13g2_o21ai_1 _6346_ (.B1(net1192),
    .Y(_2478_),
    .A1(net1439),
    .A2(\tt6581_inst.mult_inst.a_reg[19] ));
 sg13g2_o21ai_1 _6347_ (.B1(_2470_),
    .Y(_0319_),
    .A1(_2477_),
    .A2(_2478_));
 sg13g2_a22oi_1 _6348_ (.Y(_2479_),
    .B1(\tt6581_inst.svf_inst.reg_band[21] ),
    .B2(net1428),
    .A2(\tt6581_inst.svf_inst.hp_node[21] ),
    .A1(net1533));
 sg13g2_nand2b_1 _6349_ (.Y(_2480_),
    .B(net1491),
    .A_N(_2479_));
 sg13g2_nand2_1 _6350_ (.Y(_2481_),
    .A(_2225_),
    .B(_2480_));
 sg13g2_xnor2_1 _6351_ (.Y(_2482_),
    .A(_2475_),
    .B(_2481_));
 sg13g2_o21ai_1 _6352_ (.B1(net1192),
    .Y(_2483_),
    .A1(net1438),
    .A2(net243));
 sg13g2_a21oi_1 _6353_ (.A1(net1438),
    .A2(_2482_),
    .Y(_2484_),
    .B1(_2483_));
 sg13g2_a21o_1 _6354_ (.A2(net1223),
    .A1(net550),
    .B1(_2484_),
    .X(_0320_));
 sg13g2_nand2_1 _6355_ (.Y(_2485_),
    .A(net252),
    .B(net1223));
 sg13g2_a22oi_1 _6356_ (.Y(_2486_),
    .B1(\tt6581_inst.svf_inst.reg_band[22] ),
    .B2(net1428),
    .A2(\tt6581_inst.svf_inst.hp_node[22] ),
    .A1(net1533));
 sg13g2_o21ai_1 _6357_ (.B1(_2225_),
    .Y(_2487_),
    .A1(net1434),
    .A2(_2486_));
 sg13g2_nand2_1 _6358_ (.Y(_2488_),
    .A(_2474_),
    .B(_2480_));
 sg13g2_nand2_1 _6359_ (.Y(_2489_),
    .A(net1140),
    .B(_2488_));
 sg13g2_nor2_1 _6360_ (.A(net1141),
    .B(_2487_),
    .Y(_2490_));
 sg13g2_a221oi_1 _6361_ (.B2(_2488_),
    .C1(net1537),
    .B1(_2490_),
    .A1(_2487_),
    .Y(_2491_),
    .A2(_2489_));
 sg13g2_o21ai_1 _6362_ (.B1(net1192),
    .Y(_2492_),
    .A1(net1438),
    .A2(\tt6581_inst.mult_inst.a_reg[21] ));
 sg13g2_o21ai_1 _6363_ (.B1(_2485_),
    .Y(_0321_),
    .A1(_2491_),
    .A2(_2492_));
 sg13g2_nand2_1 _6364_ (.Y(_2493_),
    .A(net776),
    .B(net1224));
 sg13g2_nand3_1 _6365_ (.B(_2480_),
    .C(_2490_),
    .A(_2474_),
    .Y(_2494_));
 sg13g2_nand2_1 _6366_ (.Y(_2495_),
    .A(net1438),
    .B(_2494_));
 sg13g2_o21ai_1 _6367_ (.B1(_2495_),
    .Y(_2496_),
    .A1(net1438),
    .A2(net252));
 sg13g2_o21ai_1 _6368_ (.B1(_2493_),
    .Y(_0322_),
    .A1(net1223),
    .A2(_2496_));
 sg13g2_a22oi_1 _6369_ (.Y(_2497_),
    .B1(net1221),
    .B2(net477),
    .A2(net1287),
    .A1(\tt6581_inst.mult_inst.a_reg[23] ));
 sg13g2_inv_1 _6370_ (.Y(_0323_),
    .A(net478));
 sg13g2_a22oi_1 _6371_ (.Y(_2498_),
    .B1(net1221),
    .B2(net525),
    .A2(net1287),
    .A1(net477));
 sg13g2_inv_1 _6372_ (.Y(_0324_),
    .A(_2498_));
 sg13g2_a22oi_1 _6373_ (.Y(_2499_),
    .B1(net1221),
    .B2(net627),
    .A2(net1287),
    .A1(net525));
 sg13g2_inv_1 _6374_ (.Y(_0325_),
    .A(_2499_));
 sg13g2_a22oi_1 _6375_ (.Y(_2500_),
    .B1(net1221),
    .B2(net583),
    .A2(net1287),
    .A1(\tt6581_inst.mult_inst.a_reg[26] ));
 sg13g2_inv_1 _6376_ (.Y(_0326_),
    .A(net584));
 sg13g2_a22oi_1 _6377_ (.Y(_2501_),
    .B1(net1221),
    .B2(net695),
    .A2(net1287),
    .A1(net583));
 sg13g2_inv_1 _6378_ (.Y(_0327_),
    .A(_2501_));
 sg13g2_a22oi_1 _6379_ (.Y(_2502_),
    .B1(net1221),
    .B2(net519),
    .A2(net1287),
    .A1(\tt6581_inst.mult_inst.a_reg[28] ));
 sg13g2_inv_1 _6380_ (.Y(_0328_),
    .A(net520));
 sg13g2_a22oi_1 _6381_ (.Y(_2503_),
    .B1(net1221),
    .B2(net538),
    .A2(net1287),
    .A1(net519));
 sg13g2_inv_1 _6382_ (.Y(_0329_),
    .A(_2503_));
 sg13g2_a22oi_1 _6383_ (.Y(_2504_),
    .B1(net1221),
    .B2(net816),
    .A2(net1287),
    .A1(net538));
 sg13g2_inv_1 _6384_ (.Y(_0330_),
    .A(_2504_));
 sg13g2_a22oi_1 _6385_ (.Y(_2505_),
    .B1(net1222),
    .B2(net482),
    .A2(net1288),
    .A1(\tt6581_inst.mult_inst.a_reg[31] ));
 sg13g2_inv_1 _6386_ (.Y(_0331_),
    .A(net483));
 sg13g2_a22oi_1 _6387_ (.Y(_2506_),
    .B1(net1222),
    .B2(net511),
    .A2(net1288),
    .A1(net482));
 sg13g2_inv_1 _6388_ (.Y(_0332_),
    .A(_2506_));
 sg13g2_a22oi_1 _6389_ (.Y(_2507_),
    .B1(net1222),
    .B2(net555),
    .A2(net1288),
    .A1(net511));
 sg13g2_inv_1 _6390_ (.Y(_0333_),
    .A(_2507_));
 sg13g2_a22oi_1 _6391_ (.Y(_2508_),
    .B1(net1222),
    .B2(net484),
    .A2(net1289),
    .A1(\tt6581_inst.mult_inst.a_reg[34] ));
 sg13g2_inv_1 _6392_ (.Y(_0334_),
    .A(net485));
 sg13g2_a22oi_1 _6393_ (.Y(_2509_),
    .B1(net1222),
    .B2(net508),
    .A2(net1289),
    .A1(net484));
 sg13g2_inv_1 _6394_ (.Y(_0335_),
    .A(_2509_));
 sg13g2_a22oi_1 _6395_ (.Y(_2510_),
    .B1(net1222),
    .B2(net533),
    .A2(net1289),
    .A1(net508));
 sg13g2_inv_1 _6396_ (.Y(_0336_),
    .A(_2510_));
 sg13g2_a22oi_1 _6397_ (.Y(_2511_),
    .B1(net1225),
    .B2(net259),
    .A2(net1289),
    .A1(\tt6581_inst.mult_inst.a_reg[37] ));
 sg13g2_inv_1 _6398_ (.Y(_0337_),
    .A(net260));
 sg13g2_nor2_1 _6399_ (.A(_1005_),
    .B(net1415),
    .Y(_2512_));
 sg13g2_nor2_1 _6400_ (.A(net132),
    .B(net1346),
    .Y(_2513_));
 sg13g2_nand3b_1 _6401_ (.B(net1544),
    .C(_0037_),
    .Y(_2514_),
    .A_N(net1545));
 sg13g2_o21ai_1 _6402_ (.B1(_2514_),
    .Y(_2515_),
    .A1(_0838_),
    .A2(net1372));
 sg13g2_a21o_2 _6403_ (.A2(net1402),
    .A1(_0040_),
    .B1(_2515_),
    .X(_2516_));
 sg13g2_nand2_1 _6404_ (.Y(_2517_),
    .A(_0041_),
    .B(net1402));
 sg13g2_a22oi_1 _6405_ (.Y(_2518_),
    .B1(net1373),
    .B2(_0043_),
    .A2(net1423),
    .A1(_0038_));
 sg13g2_nand2_2 _6406_ (.Y(_2519_),
    .A(_2517_),
    .B(_2518_));
 sg13g2_or2_1 _6407_ (.X(_2520_),
    .B(_2519_),
    .A(_2516_));
 sg13g2_a22oi_1 _6408_ (.Y(_2521_),
    .B1(net1383),
    .B2(\tt6581_inst.controller_inst.sr_i[4] ),
    .A2(net1401),
    .A1(\tt6581_inst.controller_inst.sr_i[12] ));
 sg13g2_o21ai_1 _6409_ (.B1(_2521_),
    .Y(_2522_),
    .A1(_0875_),
    .A2(net1416));
 sg13g2_nor2_1 _6410_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][16] ),
    .B(net1372),
    .Y(_2523_));
 sg13g2_nor2_1 _6411_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][16] ),
    .B(net1415),
    .Y(_2524_));
 sg13g2_nor2_1 _6412_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][16] ),
    .B(net1392),
    .Y(_2525_));
 sg13g2_nor3_2 _6413_ (.A(_2523_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_));
 sg13g2_or3_1 _6414_ (.A(_2523_),
    .B(_2524_),
    .C(_2525_),
    .X(_2527_));
 sg13g2_nand2_2 _6415_ (.Y(_2528_),
    .A(\tt6581_inst.controller_inst.sr_i[21] ),
    .B(net1423));
 sg13g2_a22oi_1 _6416_ (.Y(_2529_),
    .B1(net1382),
    .B2(\tt6581_inst.controller_inst.sr_i[5] ),
    .A2(net1401),
    .A1(\tt6581_inst.controller_inst.sr_i[13] ));
 sg13g2_nand2_2 _6417_ (.Y(_2530_),
    .A(_2528_),
    .B(_2529_));
 sg13g2_nand2b_1 _6418_ (.Y(_2531_),
    .B(net1403),
    .A_N(\tt6581_inst.envelope_inst.vol_regs[1][17] ));
 sg13g2_a22oi_1 _6419_ (.Y(_2532_),
    .B1(net1373),
    .B2(_0839_),
    .A2(net1423),
    .A1(_0840_));
 sg13g2_and2_1 _6420_ (.A(_2531_),
    .B(_2532_),
    .X(_2533_));
 sg13g2_nand2_2 _6421_ (.Y(_2534_),
    .A(_2531_),
    .B(_2532_));
 sg13g2_nand4_1 _6422_ (.B(_2529_),
    .C(_2531_),
    .A(_2528_),
    .Y(_2535_),
    .D(_2532_));
 sg13g2_nand3_1 _6423_ (.B(_2527_),
    .C(_2535_),
    .A(net1265),
    .Y(_2536_));
 sg13g2_nand2b_2 _6424_ (.Y(_2537_),
    .B(net1423),
    .A_N(\tt6581_inst.envelope_inst.vol_regs[2][23] ));
 sg13g2_a22oi_1 _6425_ (.Y(_2538_),
    .B1(net1373),
    .B2(_0843_),
    .A2(net1402),
    .A1(_0844_));
 sg13g2_nand2_1 _6426_ (.Y(_2539_),
    .A(_2537_),
    .B(_2538_));
 sg13g2_nand2_2 _6427_ (.Y(_2540_),
    .A(\tt6581_inst.controller_inst.sr_i[7] ),
    .B(net1382));
 sg13g2_a22oi_1 _6428_ (.Y(_2541_),
    .B1(net1401),
    .B2(\tt6581_inst.controller_inst.sr_i[15] ),
    .A2(net1425),
    .A1(\tt6581_inst.controller_inst.sr_i[23] ));
 sg13g2_and2_1 _6429_ (.A(_2540_),
    .B(_2541_),
    .X(_2542_));
 sg13g2_nand2_2 _6430_ (.Y(_2543_),
    .A(_2540_),
    .B(_2541_));
 sg13g2_and4_1 _6431_ (.A(_2537_),
    .B(_2538_),
    .C(_2540_),
    .D(_2541_),
    .X(_2544_));
 sg13g2_nand2b_2 _6432_ (.Y(_2545_),
    .B(net1423),
    .A_N(\tt6581_inst.envelope_inst.vol_regs[2][22] ));
 sg13g2_a22oi_1 _6433_ (.Y(_2546_),
    .B1(net1373),
    .B2(_0845_),
    .A2(net1402),
    .A1(_0846_));
 sg13g2_and2_1 _6434_ (.A(_2545_),
    .B(_2546_),
    .X(_2547_));
 sg13g2_nand2_2 _6435_ (.Y(_2548_),
    .A(_2545_),
    .B(_2546_));
 sg13g2_nand2_1 _6436_ (.Y(_2549_),
    .A(\tt6581_inst.controller_inst.sr_i[14] ),
    .B(net1402));
 sg13g2_a22oi_1 _6437_ (.Y(_2550_),
    .B1(net1381),
    .B2(\tt6581_inst.controller_inst.sr_i[6] ),
    .A2(net1422),
    .A1(\tt6581_inst.controller_inst.sr_i[22] ));
 sg13g2_nand2_2 _6438_ (.Y(_2551_),
    .A(_2549_),
    .B(_2550_));
 sg13g2_and4_1 _6439_ (.A(_2545_),
    .B(_2546_),
    .C(_2549_),
    .D(_2550_),
    .X(_2552_));
 sg13g2_a22oi_1 _6440_ (.Y(_2553_),
    .B1(_2540_),
    .B2(_2541_),
    .A2(_2538_),
    .A1(_2537_));
 sg13g2_nand2_1 _6441_ (.Y(_2554_),
    .A(net1263),
    .B(_2543_));
 sg13g2_a22oi_1 _6442_ (.Y(_2555_),
    .B1(_2549_),
    .B2(_2550_),
    .A2(_2546_),
    .A1(_2545_));
 sg13g2_nor4_1 _6443_ (.A(_2544_),
    .B(_2552_),
    .C(_2553_),
    .D(_2555_),
    .Y(_2556_));
 sg13g2_nand2b_1 _6444_ (.Y(_2557_),
    .B(net1423),
    .A_N(\tt6581_inst.envelope_inst.vol_regs[2][21] ));
 sg13g2_a22oi_1 _6445_ (.Y(_2558_),
    .B1(net1373),
    .B2(_0847_),
    .A2(net1403),
    .A1(_0848_));
 sg13g2_nand2_1 _6446_ (.Y(_2559_),
    .A(_2557_),
    .B(_2558_));
 sg13g2_nand2_1 _6447_ (.Y(_2560_),
    .A(_2530_),
    .B(net1261));
 sg13g2_a22oi_1 _6448_ (.Y(_2561_),
    .B1(net1404),
    .B2(_0850_),
    .A2(net1424),
    .A1(_0849_));
 sg13g2_o21ai_1 _6449_ (.B1(_2561_),
    .Y(_2562_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][20] ),
    .A2(net1370));
 sg13g2_nand4_1 _6450_ (.B(_2529_),
    .C(_2557_),
    .A(_2528_),
    .Y(_2563_),
    .D(_2558_));
 sg13g2_xor2_1 _6451_ (.B(net1260),
    .A(net1265),
    .X(_2564_));
 sg13g2_and4_1 _6452_ (.A(_2556_),
    .B(_2560_),
    .C(_2563_),
    .D(_2564_),
    .X(_2565_));
 sg13g2_nand4_1 _6453_ (.B(_2560_),
    .C(_2563_),
    .A(_2556_),
    .Y(_2566_),
    .D(_2564_));
 sg13g2_nor2_1 _6454_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][19] ),
    .B(net1372),
    .Y(_2567_));
 sg13g2_nor2_1 _6455_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][19] ),
    .B(net1415),
    .Y(_2568_));
 sg13g2_nor2_1 _6456_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][19] ),
    .B(net1392),
    .Y(_2569_));
 sg13g2_nor3_2 _6457_ (.A(_2567_),
    .B(_2568_),
    .C(_2569_),
    .Y(_2570_));
 sg13g2_or3_1 _6458_ (.A(_2567_),
    .B(_2568_),
    .C(_2569_),
    .X(_2571_));
 sg13g2_nand2_1 _6459_ (.Y(_2572_),
    .A(_2543_),
    .B(net1258));
 sg13g2_a22oi_1 _6460_ (.Y(_2573_),
    .B1(net1400),
    .B2(_0842_),
    .A2(net1421),
    .A1(_0841_));
 sg13g2_o21ai_1 _6461_ (.B1(_2573_),
    .Y(_2574_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][18] ),
    .A2(net1370));
 sg13g2_inv_2 _6462_ (.Y(_2575_),
    .A(_2574_));
 sg13g2_nor2_1 _6463_ (.A(_2551_),
    .B(net1257),
    .Y(_2576_));
 sg13g2_nor2_1 _6464_ (.A(_2543_),
    .B(net1258),
    .Y(_2577_));
 sg13g2_xor2_1 _6465_ (.B(net1257),
    .A(_2551_),
    .X(_2578_));
 sg13g2_a22oi_1 _6466_ (.Y(_2579_),
    .B1(_2542_),
    .B2(_2570_),
    .A2(_2534_),
    .A1(_2530_));
 sg13g2_and4_1 _6467_ (.A(_2565_),
    .B(_2572_),
    .C(_2578_),
    .D(_2579_),
    .X(_2580_));
 sg13g2_o21ai_1 _6468_ (.B1(_2563_),
    .Y(_2581_),
    .A1(net1265),
    .A2(net1259));
 sg13g2_and2_1 _6469_ (.A(_2560_),
    .B(_2581_),
    .X(_2582_));
 sg13g2_a221oi_1 _6470_ (.B2(_2582_),
    .C1(_2544_),
    .B1(_2556_),
    .A1(_2552_),
    .Y(_2583_),
    .A2(_2554_));
 sg13g2_a21oi_1 _6471_ (.A1(_2572_),
    .A2(_2576_),
    .Y(_2584_),
    .B1(_2577_));
 sg13g2_nand4_1 _6472_ (.B(_2572_),
    .C(_2578_),
    .A(_2536_),
    .Y(_2585_),
    .D(_2579_));
 sg13g2_a21o_1 _6473_ (.A2(_2585_),
    .A1(_2584_),
    .B1(_2566_),
    .X(_2586_));
 sg13g2_xnor2_1 _6474_ (.Y(_2587_),
    .A(net1265),
    .B(_2526_));
 sg13g2_a22oi_1 _6475_ (.Y(_2588_),
    .B1(net1373),
    .B2(_0869_),
    .A2(net1403),
    .A1(_0870_));
 sg13g2_o21ai_1 _6476_ (.B1(_2588_),
    .Y(_2589_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[2][12] ),
    .A2(net1415));
 sg13g2_a22oi_1 _6477_ (.Y(_2590_),
    .B1(net1403),
    .B2(_0874_),
    .A2(net1424),
    .A1(_0873_));
 sg13g2_o21ai_1 _6478_ (.B1(_2590_),
    .Y(_2591_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][14] ),
    .A2(net1372));
 sg13g2_a22oi_1 _6479_ (.Y(_2592_),
    .B1(net1404),
    .B2(_0864_),
    .A2(net1424),
    .A1(_0863_));
 sg13g2_o21ai_1 _6480_ (.B1(_2592_),
    .Y(_2593_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][8] ),
    .A2(net1370));
 sg13g2_a22oi_1 _6481_ (.Y(_2594_),
    .B1(net1404),
    .B2(_0852_),
    .A2(net1424),
    .A1(_0851_));
 sg13g2_o21ai_1 _6482_ (.B1(_2594_),
    .Y(_2595_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][1] ),
    .A2(net1370));
 sg13g2_a22oi_1 _6483_ (.Y(_2596_),
    .B1(net1404),
    .B2(_0854_),
    .A2(net1424),
    .A1(_0853_));
 sg13g2_o21ai_1 _6484_ (.B1(_2596_),
    .Y(_2597_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][5] ),
    .A2(net1371));
 sg13g2_a22oi_1 _6485_ (.Y(_2598_),
    .B1(net1403),
    .B2(_0868_),
    .A2(net1423),
    .A1(_0867_));
 sg13g2_o21ai_1 _6486_ (.B1(_2598_),
    .Y(_2599_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][10] ),
    .A2(net1372));
 sg13g2_a22oi_1 _6487_ (.Y(_2600_),
    .B1(net1405),
    .B2(_0866_),
    .A2(net1425),
    .A1(_0865_));
 sg13g2_o21ai_1 _6488_ (.B1(_2600_),
    .Y(_2601_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][11] ),
    .A2(net1371));
 sg13g2_nor2_1 _6489_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][0] ),
    .B(net1371),
    .Y(_2602_));
 sg13g2_nor2_1 _6490_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][0] ),
    .B(net1415),
    .Y(_2603_));
 sg13g2_nor2_1 _6491_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][0] ),
    .B(net1392),
    .Y(_2604_));
 sg13g2_nor3_1 _6492_ (.A(_2602_),
    .B(_2603_),
    .C(_2604_),
    .Y(_2605_));
 sg13g2_or3_1 _6493_ (.A(_2602_),
    .B(_2603_),
    .C(_2604_),
    .X(_2606_));
 sg13g2_a22oi_1 _6494_ (.Y(_2607_),
    .B1(net1404),
    .B2(_0858_),
    .A2(net1424),
    .A1(_0857_));
 sg13g2_o21ai_1 _6495_ (.B1(_2607_),
    .Y(_2608_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][7] ),
    .A2(net1370));
 sg13g2_a22oi_1 _6496_ (.Y(_2609_),
    .B1(net1403),
    .B2(_0872_),
    .A2(net1424),
    .A1(_0871_));
 sg13g2_o21ai_1 _6497_ (.B1(_2609_),
    .Y(_2610_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][15] ),
    .A2(net1371));
 sg13g2_a22oi_1 _6498_ (.Y(_2611_),
    .B1(_1532_),
    .B2(_0861_),
    .A2(net1404),
    .A1(_0862_));
 sg13g2_o21ai_1 _6499_ (.B1(_2611_),
    .Y(_2612_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[2][9] ),
    .A2(net1415));
 sg13g2_a22oi_1 _6500_ (.Y(_2613_),
    .B1(net1373),
    .B2(_0859_),
    .A2(net1404),
    .A1(_0860_));
 sg13g2_o21ai_1 _6501_ (.B1(_2613_),
    .Y(_2614_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[2][6] ),
    .A2(net1415));
 sg13g2_nor2_1 _6502_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][2] ),
    .B(net1370),
    .Y(_2615_));
 sg13g2_nor2_1 _6503_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][2] ),
    .B(net1415),
    .Y(_2616_));
 sg13g2_nor2_1 _6504_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][2] ),
    .B(net1392),
    .Y(_2617_));
 sg13g2_nor3_2 _6505_ (.A(_2615_),
    .B(_2616_),
    .C(_2617_),
    .Y(_2618_));
 sg13g2_or3_1 _6506_ (.A(_2615_),
    .B(_2616_),
    .C(_2617_),
    .X(_2619_));
 sg13g2_nor2_1 _6507_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][13] ),
    .B(net1371),
    .Y(_2620_));
 sg13g2_nor2_1 _6508_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][13] ),
    .B(net1416),
    .Y(_2621_));
 sg13g2_nor2_1 _6509_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][13] ),
    .B(net1392),
    .Y(_2622_));
 sg13g2_nor3_1 _6510_ (.A(_2620_),
    .B(_2621_),
    .C(_2622_),
    .Y(_2623_));
 sg13g2_or3_1 _6511_ (.A(_2620_),
    .B(_2621_),
    .C(_2622_),
    .X(_2624_));
 sg13g2_nor2_1 _6512_ (.A(\tt6581_inst.envelope_inst.vol_regs[0][3] ),
    .B(net1370),
    .Y(_2625_));
 sg13g2_nor2_1 _6513_ (.A(\tt6581_inst.envelope_inst.vol_regs[2][3] ),
    .B(net1416),
    .Y(_2626_));
 sg13g2_nor2_1 _6514_ (.A(\tt6581_inst.envelope_inst.vol_regs[1][3] ),
    .B(_1043_),
    .Y(_2627_));
 sg13g2_nor3_2 _6515_ (.A(_2625_),
    .B(_2626_),
    .C(_2627_),
    .Y(_2628_));
 sg13g2_a22oi_1 _6516_ (.Y(_2629_),
    .B1(net1404),
    .B2(_0856_),
    .A2(net1425),
    .A1(_0855_));
 sg13g2_o21ai_1 _6517_ (.B1(_2629_),
    .Y(_2630_),
    .A1(\tt6581_inst.envelope_inst.vol_regs[0][4] ),
    .A2(net1370));
 sg13g2_inv_2 _6518_ (.Y(_2631_),
    .A(_2630_));
 sg13g2_and4_1 _6519_ (.A(_2589_),
    .B(_2599_),
    .C(_2614_),
    .D(_2624_),
    .X(_2632_));
 sg13g2_nand4_1 _6520_ (.B(_2608_),
    .C(_2610_),
    .A(_2593_),
    .Y(_2633_),
    .D(_2612_));
 sg13g2_nand3_1 _6521_ (.B(_2601_),
    .C(_2630_),
    .A(_2595_),
    .Y(_2634_));
 sg13g2_nand4_1 _6522_ (.B(_2597_),
    .C(_2606_),
    .A(_2591_),
    .Y(_2635_),
    .D(_2619_));
 sg13g2_nor4_1 _6523_ (.A(_2628_),
    .B(_2633_),
    .C(_2634_),
    .D(_2635_),
    .Y(_2636_));
 sg13g2_and4_1 _6524_ (.A(_2535_),
    .B(_2587_),
    .C(_2632_),
    .D(_2636_),
    .X(_2637_));
 sg13g2_a221oi_1 _6525_ (.B2(_2580_),
    .C1(_2516_),
    .B1(_2637_),
    .A1(_2583_),
    .Y(_2638_),
    .A2(_2586_));
 sg13g2_or4_1 _6526_ (.A(net1263),
    .B(_2548_),
    .C(net1262),
    .D(net1260),
    .X(_2639_));
 sg13g2_or4_1 _6527_ (.A(_2608_),
    .B(_2610_),
    .C(_2612_),
    .D(_2614_),
    .X(_2640_));
 sg13g2_nand4_1 _6528_ (.B(_2623_),
    .C(_2628_),
    .A(_2618_),
    .Y(_2641_),
    .D(_2631_));
 sg13g2_nor4_1 _6529_ (.A(_2527_),
    .B(_2534_),
    .C(net1258),
    .D(net1257),
    .Y(_2642_));
 sg13g2_and2_1 _6530_ (.A(_2516_),
    .B(_2519_),
    .X(_2643_));
 sg13g2_nor4_1 _6531_ (.A(_2589_),
    .B(_2591_),
    .C(_2593_),
    .D(_2595_),
    .Y(_2644_));
 sg13g2_nor4_1 _6532_ (.A(_2597_),
    .B(_2599_),
    .C(_2601_),
    .D(_2606_),
    .Y(_2645_));
 sg13g2_nand4_1 _6533_ (.B(_2643_),
    .C(_2644_),
    .A(_2642_),
    .Y(_2646_),
    .D(_2645_));
 sg13g2_nor4_1 _6534_ (.A(_2639_),
    .B(_2640_),
    .C(_2641_),
    .D(_2646_),
    .Y(_2647_));
 sg13g2_o21ai_1 _6535_ (.B1(_2520_),
    .Y(_2648_),
    .A1(_2638_),
    .A2(_2647_));
 sg13g2_nand2_1 _6536_ (.Y(_2649_),
    .A(\tt6581_inst.control_pack[8] ),
    .B(net1402));
 sg13g2_a22oi_1 _6537_ (.Y(_2650_),
    .B1(net1383),
    .B2(\tt6581_inst.control_pack[0] ),
    .A2(net1421),
    .A1(\tt6581_inst.control_pack[16] ));
 sg13g2_and2_1 _6538_ (.A(_2649_),
    .B(_2650_),
    .X(_2651_));
 sg13g2_nand2_2 _6539_ (.Y(_2652_),
    .A(_2649_),
    .B(_2650_));
 sg13g2_and2_1 _6540_ (.A(_2648_),
    .B(_2652_),
    .X(_2653_));
 sg13g2_nand2_2 _6541_ (.Y(_2654_),
    .A(_2648_),
    .B(_2652_));
 sg13g2_a21oi_1 _6542_ (.A1(net1346),
    .A2(_2654_),
    .Y(_0338_),
    .B1(_2513_));
 sg13g2_xnor2_1 _6543_ (.Y(_2655_),
    .A(_2516_),
    .B(_2519_));
 sg13g2_nor2_1 _6544_ (.A(_2638_),
    .B(_2655_),
    .Y(_2656_));
 sg13g2_nor2_2 _6545_ (.A(_2651_),
    .B(_2656_),
    .Y(_2657_));
 sg13g2_o21ai_1 _6546_ (.B1(_2652_),
    .Y(_2658_),
    .A1(_2638_),
    .A2(_2655_));
 sg13g2_nor2_1 _6547_ (.A(net218),
    .B(net1346),
    .Y(_2659_));
 sg13g2_a21oi_1 _6548_ (.A1(net1346),
    .A2(_2658_),
    .Y(_0339_),
    .B1(_2659_));
 sg13g2_and2_1 _6549_ (.A(net1542),
    .B(net102),
    .X(_2660_));
 sg13g2_or2_1 _6550_ (.X(_2661_),
    .B(\tt6581_inst.svf_inst.cur_state[10] ),
    .A(net1535));
 sg13g2_a22oi_1 _6551_ (.Y(_2662_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[0] ),
    .A2(\tt6581_inst.filt_q_lo[0] ),
    .A1(net1525));
 sg13g2_a22oi_1 _6552_ (.Y(_2663_),
    .B1(_1002_),
    .B2(_2526_),
    .A2(net1493),
    .A1(\tt6581_inst.filt_volume[0] ));
 sg13g2_o21ai_1 _6553_ (.B1(_2663_),
    .Y(_2664_),
    .A1(net1435),
    .A2(_2662_));
 sg13g2_a21oi_1 _6554_ (.A1(net1442),
    .A2(_2664_),
    .Y(_2665_),
    .B1(_2660_));
 sg13g2_nand2_1 _6555_ (.Y(_2666_),
    .A(net229),
    .B(net1231));
 sg13g2_o21ai_1 _6556_ (.B1(_2666_),
    .Y(_0340_),
    .A1(net1231),
    .A2(_2665_));
 sg13g2_nand2_1 _6557_ (.Y(_2667_),
    .A(net102),
    .B(net1229));
 sg13g2_a22oi_1 _6558_ (.Y(_2668_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[1] ),
    .A2(\tt6581_inst.filt_q_lo[1] ),
    .A1(net1524));
 sg13g2_inv_1 _6559_ (.Y(_2669_),
    .A(_2668_));
 sg13g2_a22oi_1 _6560_ (.Y(_2670_),
    .B1(_2669_),
    .B2(net1490),
    .A2(\tt6581_inst.filt_volume[1] ),
    .A1(net1493));
 sg13g2_o21ai_1 _6561_ (.B1(_2670_),
    .Y(_2671_),
    .A1(net1494),
    .A2(_2534_));
 sg13g2_a22oi_1 _6562_ (.Y(_2672_),
    .B1(net1362),
    .B2(\tt6581_inst.filt_f_hi[7] ),
    .A2(\tt6581_inst.filt_q_hi[7] ),
    .A1(net1524));
 sg13g2_nor2_1 _6563_ (.A(net1436),
    .B(_2672_),
    .Y(_2673_));
 sg13g2_nand2b_2 _6564_ (.Y(_2674_),
    .B(net1489),
    .A_N(_2672_));
 sg13g2_nand2_1 _6565_ (.Y(_2675_),
    .A(_2664_),
    .B(net1256));
 sg13g2_xnor2_1 _6566_ (.Y(_2676_),
    .A(_2671_),
    .B(_2675_));
 sg13g2_nor2_1 _6567_ (.A(net1541),
    .B(_2676_),
    .Y(_2677_));
 sg13g2_o21ai_1 _6568_ (.B1(net1196),
    .Y(_2678_),
    .A1(net1442),
    .A2(net86));
 sg13g2_o21ai_1 _6569_ (.B1(_2667_),
    .Y(_0341_),
    .A1(_2677_),
    .A2(_2678_));
 sg13g2_nand2_1 _6570_ (.Y(_2679_),
    .A(net86),
    .B(net1229));
 sg13g2_a22oi_1 _6571_ (.Y(_2680_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[2] ),
    .A2(\tt6581_inst.filt_q_lo[2] ),
    .A1(net1525));
 sg13g2_nand2b_1 _6572_ (.Y(_2681_),
    .B(net1489),
    .A_N(_2680_));
 sg13g2_o21ai_1 _6573_ (.B1(_2681_),
    .Y(_2682_),
    .A1(net1494),
    .A2(_2574_));
 sg13g2_a21oi_1 _6574_ (.A1(net1493),
    .A2(\tt6581_inst.filt_volume[2] ),
    .Y(_2683_),
    .B1(_2682_));
 sg13g2_nor2_1 _6575_ (.A(_2664_),
    .B(_2671_),
    .Y(_2684_));
 sg13g2_nor2_1 _6576_ (.A(_2674_),
    .B(_2684_),
    .Y(_2685_));
 sg13g2_o21ai_1 _6577_ (.B1(net1442),
    .Y(_2686_),
    .A1(_2683_),
    .A2(_2685_));
 sg13g2_a21oi_1 _6578_ (.A1(_2683_),
    .A2(_2685_),
    .Y(_2687_),
    .B1(_2686_));
 sg13g2_o21ai_1 _6579_ (.B1(net1196),
    .Y(_2688_),
    .A1(net1442),
    .A2(\tt6581_inst.mult_inst.b_reg[3] ));
 sg13g2_o21ai_1 _6580_ (.B1(_2679_),
    .Y(_0342_),
    .A1(_2687_),
    .A2(_2688_));
 sg13g2_nand2_1 _6581_ (.Y(_2689_),
    .A(net115),
    .B(net1229));
 sg13g2_a22oi_1 _6582_ (.Y(_2690_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[3] ),
    .A2(\tt6581_inst.filt_q_lo[3] ),
    .A1(net1524));
 sg13g2_inv_1 _6583_ (.Y(_2691_),
    .A(_2690_));
 sg13g2_a22oi_1 _6584_ (.Y(_2692_),
    .B1(_2691_),
    .B2(net1489),
    .A2(\tt6581_inst.filt_volume[3] ),
    .A1(net1493));
 sg13g2_o21ai_1 _6585_ (.B1(_2692_),
    .Y(_2693_),
    .A1(net1494),
    .A2(net1258));
 sg13g2_and2_1 _6586_ (.A(_2683_),
    .B(_2684_),
    .X(_2694_));
 sg13g2_nor2_1 _6587_ (.A(_2674_),
    .B(_2694_),
    .Y(_2695_));
 sg13g2_xor2_1 _6588_ (.B(_2695_),
    .A(_2693_),
    .X(_2696_));
 sg13g2_nor2_1 _6589_ (.A(net1541),
    .B(_2696_),
    .Y(_2697_));
 sg13g2_o21ai_1 _6590_ (.B1(net1196),
    .Y(_2698_),
    .A1(net1443),
    .A2(net100));
 sg13g2_o21ai_1 _6591_ (.B1(_2689_),
    .Y(_0343_),
    .A1(_2697_),
    .A2(_2698_));
 sg13g2_nand2_1 _6592_ (.Y(_2699_),
    .A(net100),
    .B(net1229));
 sg13g2_a22oi_1 _6593_ (.Y(_2700_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[4] ),
    .A2(\tt6581_inst.filt_q_lo[4] ),
    .A1(net1525));
 sg13g2_nand2b_1 _6594_ (.Y(_2701_),
    .B(net1489),
    .A_N(_2700_));
 sg13g2_o21ai_1 _6595_ (.B1(_2701_),
    .Y(_2702_),
    .A1(net1494),
    .A2(_2562_));
 sg13g2_a21oi_1 _6596_ (.A1(net1493),
    .A2(\tt6581_inst.filt_volume[4] ),
    .Y(_2703_),
    .B1(_2702_));
 sg13g2_nor2b_1 _6597_ (.A(_2693_),
    .B_N(_2694_),
    .Y(_2704_));
 sg13g2_nor2_1 _6598_ (.A(_2674_),
    .B(_2704_),
    .Y(_2705_));
 sg13g2_o21ai_1 _6599_ (.B1(net1442),
    .Y(_2706_),
    .A1(_2703_),
    .A2(_2705_));
 sg13g2_a21oi_1 _6600_ (.A1(_2703_),
    .A2(_2705_),
    .Y(_2707_),
    .B1(_2706_));
 sg13g2_o21ai_1 _6601_ (.B1(net1196),
    .Y(_2708_),
    .A1(net1443),
    .A2(net84));
 sg13g2_o21ai_1 _6602_ (.B1(_2699_),
    .Y(_0344_),
    .A1(_2707_),
    .A2(_2708_));
 sg13g2_nand2_1 _6603_ (.Y(_2709_),
    .A(net84),
    .B(net1229));
 sg13g2_a22oi_1 _6604_ (.Y(_2710_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[5] ),
    .A2(\tt6581_inst.filt_q_lo[5] ),
    .A1(net1525));
 sg13g2_nor2_1 _6605_ (.A(net1436),
    .B(_2710_),
    .Y(_2711_));
 sg13g2_a21oi_1 _6606_ (.A1(net1493),
    .A2(\tt6581_inst.filt_volume[5] ),
    .Y(_2712_),
    .B1(_2711_));
 sg13g2_o21ai_1 _6607_ (.B1(_2712_),
    .Y(_2713_),
    .A1(net1494),
    .A2(net1262));
 sg13g2_and2_1 _6608_ (.A(_2703_),
    .B(_2704_),
    .X(_2714_));
 sg13g2_nor2_1 _6609_ (.A(_2674_),
    .B(_2714_),
    .Y(_2715_));
 sg13g2_xor2_1 _6610_ (.B(_2715_),
    .A(_2713_),
    .X(_2716_));
 sg13g2_nor2_1 _6611_ (.A(net1542),
    .B(_2716_),
    .Y(_2717_));
 sg13g2_o21ai_1 _6612_ (.B1(net1196),
    .Y(_2718_),
    .A1(net1442),
    .A2(net75));
 sg13g2_o21ai_1 _6613_ (.B1(_2709_),
    .Y(_0345_),
    .A1(_2717_),
    .A2(_2718_));
 sg13g2_nand2_1 _6614_ (.Y(_2719_),
    .A(net75),
    .B(net1230));
 sg13g2_a22oi_1 _6615_ (.Y(_2720_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[6] ),
    .A2(\tt6581_inst.filt_q_lo[6] ),
    .A1(net1525));
 sg13g2_nand2b_1 _6616_ (.Y(_2721_),
    .B(net1490),
    .A_N(_2720_));
 sg13g2_o21ai_1 _6617_ (.B1(_2721_),
    .Y(_2722_),
    .A1(_0113_),
    .A2(_2548_));
 sg13g2_a21oi_1 _6618_ (.A1(\tt6581_inst.controller_inst.mult_in_mux_o[1] ),
    .A2(\tt6581_inst.filt_volume[6] ),
    .Y(_2723_),
    .B1(_2722_));
 sg13g2_nand2b_1 _6619_ (.Y(_2724_),
    .B(_2714_),
    .A_N(_2713_));
 sg13g2_nand3_1 _6620_ (.B(_2723_),
    .C(_2724_),
    .A(net1256),
    .Y(_2725_));
 sg13g2_a21o_1 _6621_ (.A2(_2724_),
    .A1(net1256),
    .B1(_2723_),
    .X(_2726_));
 sg13g2_nand3_1 _6622_ (.B(_2725_),
    .C(_2726_),
    .A(net1442),
    .Y(_2727_));
 sg13g2_o21ai_1 _6623_ (.B1(_2727_),
    .Y(_2728_),
    .A1(net1442),
    .A2(\tt6581_inst.mult_inst.b_reg[7] ));
 sg13g2_o21ai_1 _6624_ (.B1(_2719_),
    .Y(_0346_),
    .A1(net1229),
    .A2(_2728_));
 sg13g2_nand2_1 _6625_ (.Y(_2729_),
    .A(net96),
    .B(net1229));
 sg13g2_a22oi_1 _6626_ (.Y(_2730_),
    .B1(net1363),
    .B2(\tt6581_inst.filt_f_lo[7] ),
    .A2(\tt6581_inst.filt_q_lo[7] ),
    .A1(net1525));
 sg13g2_nor2_1 _6627_ (.A(net1436),
    .B(_2730_),
    .Y(_2731_));
 sg13g2_a21oi_1 _6628_ (.A1(\tt6581_inst.controller_inst.mult_in_mux_o[1] ),
    .A2(\tt6581_inst.filt_volume[7] ),
    .Y(_2732_),
    .B1(_2731_));
 sg13g2_o21ai_1 _6629_ (.B1(_2732_),
    .Y(_2733_),
    .A1(_0113_),
    .A2(net1264));
 sg13g2_nand3b_1 _6630_ (.B(_2714_),
    .C(_2723_),
    .Y(_2734_),
    .A_N(_2713_));
 sg13g2_nand2_1 _6631_ (.Y(_2735_),
    .A(_2673_),
    .B(_2734_));
 sg13g2_a21oi_1 _6632_ (.A1(_2733_),
    .A2(_2735_),
    .Y(_2736_),
    .B1(net1542));
 sg13g2_o21ai_1 _6633_ (.B1(_2736_),
    .Y(_2737_),
    .A1(_2733_),
    .A2(_2735_));
 sg13g2_o21ai_1 _6634_ (.B1(_2737_),
    .Y(_2738_),
    .A1(net1443),
    .A2(net73));
 sg13g2_o21ai_1 _6635_ (.B1(_2729_),
    .Y(_0347_),
    .A1(net1230),
    .A2(_2738_));
 sg13g2_nand2_1 _6636_ (.Y(_2739_),
    .A(net73),
    .B(net1230));
 sg13g2_nor2_1 _6637_ (.A(_2733_),
    .B(_2734_),
    .Y(_2740_));
 sg13g2_nor2_1 _6638_ (.A(_2674_),
    .B(_2740_),
    .Y(_2741_));
 sg13g2_a22oi_1 _6639_ (.Y(_2742_),
    .B1(net1362),
    .B2(\tt6581_inst.filt_f_hi[0] ),
    .A2(\tt6581_inst.filt_q_hi[0] ),
    .A1(net1524));
 sg13g2_nor2_1 _6640_ (.A(net1436),
    .B(_2742_),
    .Y(_2743_));
 sg13g2_mux2_1 _6641_ (.A0(_2743_),
    .A1(_2742_),
    .S(_2741_),
    .X(_2744_));
 sg13g2_nor2_1 _6642_ (.A(net1542),
    .B(_2744_),
    .Y(_2745_));
 sg13g2_o21ai_1 _6643_ (.B1(net1195),
    .Y(_2746_),
    .A1(net1443),
    .A2(\tt6581_inst.mult_inst.b_reg[9] ));
 sg13g2_o21ai_1 _6644_ (.B1(_2739_),
    .Y(_0348_),
    .A1(_2745_),
    .A2(_2746_));
 sg13g2_nand2_1 _6645_ (.Y(_2747_),
    .A(net110),
    .B(net1230));
 sg13g2_a22oi_1 _6646_ (.Y(_2748_),
    .B1(net1362),
    .B2(\tt6581_inst.filt_f_hi[1] ),
    .A2(\tt6581_inst.filt_q_hi[1] ),
    .A1(net1524));
 sg13g2_nor2_1 _6647_ (.A(net1436),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_a21o_1 _6648_ (.A2(_2742_),
    .A1(_2740_),
    .B1(_2674_),
    .X(_2750_));
 sg13g2_o21ai_1 _6649_ (.B1(net1443),
    .Y(_2751_),
    .A1(_2749_),
    .A2(_2750_));
 sg13g2_a21oi_1 _6650_ (.A1(_2749_),
    .A2(_2750_),
    .Y(_2752_),
    .B1(_2751_));
 sg13g2_o21ai_1 _6651_ (.B1(net1195),
    .Y(_2753_),
    .A1(net1443),
    .A2(\tt6581_inst.mult_inst.b_reg[10] ));
 sg13g2_o21ai_1 _6652_ (.B1(_2747_),
    .Y(_0349_),
    .A1(_2752_),
    .A2(_2753_));
 sg13g2_or4_1 _6653_ (.A(_2733_),
    .B(_2734_),
    .C(_2743_),
    .D(_2749_),
    .X(_2754_));
 sg13g2_nand2_1 _6654_ (.Y(_2755_),
    .A(net1256),
    .B(_2754_));
 sg13g2_and2_1 _6655_ (.A(net1526),
    .B(\tt6581_inst.filt_q_hi[2] ),
    .X(_2756_));
 sg13g2_a21o_1 _6656_ (.A2(net1362),
    .A1(\tt6581_inst.filt_f_hi[2] ),
    .B1(_2756_),
    .X(_2757_));
 sg13g2_nand2_1 _6657_ (.Y(_2758_),
    .A(net1489),
    .B(_2757_));
 sg13g2_mux2_1 _6658_ (.A0(_2757_),
    .A1(_2758_),
    .S(_2755_),
    .X(_2759_));
 sg13g2_o21ai_1 _6659_ (.B1(net1195),
    .Y(_2760_),
    .A1(net1444),
    .A2(net82));
 sg13g2_a21oi_1 _6660_ (.A1(net1444),
    .A2(_2759_),
    .Y(_2761_),
    .B1(_2760_));
 sg13g2_a21o_1 _6661_ (.A2(net1231),
    .A1(net226),
    .B1(_2761_),
    .X(_0350_));
 sg13g2_nand2_1 _6662_ (.Y(_2762_),
    .A(net82),
    .B(net1231));
 sg13g2_o21ai_1 _6663_ (.B1(net1256),
    .Y(_2763_),
    .A1(_2754_),
    .A2(_2757_));
 sg13g2_a22oi_1 _6664_ (.Y(_2764_),
    .B1(net1362),
    .B2(\tt6581_inst.filt_f_hi[3] ),
    .A2(\tt6581_inst.filt_q_hi[3] ),
    .A1(net1524));
 sg13g2_nor2_1 _6665_ (.A(net1436),
    .B(_2764_),
    .Y(_2765_));
 sg13g2_mux2_1 _6666_ (.A0(_2764_),
    .A1(_2765_),
    .S(_2763_),
    .X(_2766_));
 sg13g2_nor2_1 _6667_ (.A(net1541),
    .B(_2766_),
    .Y(_2767_));
 sg13g2_o21ai_1 _6668_ (.B1(net1195),
    .Y(_2768_),
    .A1(net1444),
    .A2(\tt6581_inst.mult_inst.b_reg[12] ));
 sg13g2_o21ai_1 _6669_ (.B1(_2762_),
    .Y(_0351_),
    .A1(_2767_),
    .A2(_2768_));
 sg13g2_nor2_1 _6670_ (.A(_2754_),
    .B(_2765_),
    .Y(_2769_));
 sg13g2_a21o_1 _6671_ (.A2(_2769_),
    .A1(_2758_),
    .B1(_2674_),
    .X(_2770_));
 sg13g2_and2_1 _6672_ (.A(net1524),
    .B(\tt6581_inst.filt_q_hi[4] ),
    .X(_2771_));
 sg13g2_a21o_1 _6673_ (.A2(net1362),
    .A1(\tt6581_inst.filt_f_hi[4] ),
    .B1(_2771_),
    .X(_2772_));
 sg13g2_nand2_1 _6674_ (.Y(_2773_),
    .A(net1489),
    .B(_2772_));
 sg13g2_mux2_1 _6675_ (.A0(_2772_),
    .A1(_2773_),
    .S(_2770_),
    .X(_2774_));
 sg13g2_o21ai_1 _6676_ (.B1(net1195),
    .Y(_2775_),
    .A1(net1444),
    .A2(net79));
 sg13g2_a21oi_1 _6677_ (.A1(net1444),
    .A2(_2774_),
    .Y(_2776_),
    .B1(_2775_));
 sg13g2_a21o_1 _6678_ (.A2(net1231),
    .A1(net251),
    .B1(_2776_),
    .X(_0352_));
 sg13g2_nand2_1 _6679_ (.Y(_2777_),
    .A(net79),
    .B(net1231));
 sg13g2_nand2_1 _6680_ (.Y(_2778_),
    .A(net1256),
    .B(_2772_));
 sg13g2_nand2_1 _6681_ (.Y(_2779_),
    .A(_2770_),
    .B(_2778_));
 sg13g2_a22oi_1 _6682_ (.Y(_2780_),
    .B1(net1362),
    .B2(\tt6581_inst.filt_f_hi[5] ),
    .A2(\tt6581_inst.filt_q_hi[5] ),
    .A1(net1526));
 sg13g2_nand2b_1 _6683_ (.Y(_2781_),
    .B(net1489),
    .A_N(_2780_));
 sg13g2_nand2_1 _6684_ (.Y(_2782_),
    .A(_2779_),
    .B(_2780_));
 sg13g2_o21ai_1 _6685_ (.B1(_2782_),
    .Y(_2783_),
    .A1(_2779_),
    .A2(_2781_));
 sg13g2_nor2_1 _6686_ (.A(net1541),
    .B(_2783_),
    .Y(_2784_));
 sg13g2_o21ai_1 _6687_ (.B1(net1195),
    .Y(_2785_),
    .A1(net1444),
    .A2(\tt6581_inst.mult_inst.b_reg[14] ));
 sg13g2_o21ai_1 _6688_ (.B1(_2777_),
    .Y(_0353_),
    .A1(_2784_),
    .A2(_2785_));
 sg13g2_nand4_1 _6689_ (.B(_2769_),
    .C(_2773_),
    .A(_2758_),
    .Y(_2786_),
    .D(_2781_));
 sg13g2_nand2_1 _6690_ (.Y(_2787_),
    .A(net1256),
    .B(_2786_));
 sg13g2_and2_1 _6691_ (.A(net1524),
    .B(\tt6581_inst.filt_q_hi[6] ),
    .X(_2788_));
 sg13g2_a21o_1 _6692_ (.A2(net1362),
    .A1(\tt6581_inst.filt_f_hi[6] ),
    .B1(_2788_),
    .X(_2789_));
 sg13g2_nand3_1 _6693_ (.B(_2787_),
    .C(_2789_),
    .A(net1489),
    .Y(_2790_));
 sg13g2_nor2_1 _6694_ (.A(_2787_),
    .B(_2789_),
    .Y(_2791_));
 sg13g2_nor2_1 _6695_ (.A(net1541),
    .B(_2791_),
    .Y(_2792_));
 sg13g2_o21ai_1 _6696_ (.B1(net1195),
    .Y(_2793_),
    .A1(net1444),
    .A2(\tt6581_inst.mult_inst.b_reg[15] ));
 sg13g2_a21oi_1 _6697_ (.A1(_2790_),
    .A2(_2792_),
    .Y(_2794_),
    .B1(_2793_));
 sg13g2_a21o_1 _6698_ (.A2(net1227),
    .A1(net237),
    .B1(_2794_),
    .X(_0354_));
 sg13g2_nor4_1 _6699_ (.A(net1541),
    .B(_2674_),
    .C(_2786_),
    .D(_2789_),
    .Y(_2795_));
 sg13g2_a21o_1 _6700_ (.A2(net1231),
    .A1(net239),
    .B1(_2795_),
    .X(_0355_));
 sg13g2_o21ai_1 _6701_ (.B1(net1195),
    .Y(_2796_),
    .A1(net1444),
    .A2(\tt6581_inst.mult_inst.b_reg[0] ));
 sg13g2_o21ai_1 _6702_ (.B1(net435),
    .Y(_2797_),
    .A1(_2233_),
    .A2(net1180));
 sg13g2_nor2_1 _6703_ (.A(net1439),
    .B(net1180),
    .Y(_2798_));
 sg13g2_nand3_1 _6704_ (.B(net229),
    .C(_1009_),
    .A(net1541),
    .Y(_2799_));
 sg13g2_nand2b_1 _6705_ (.Y(_2800_),
    .B(\tt6581_inst.mult_inst.a_reg[0] ),
    .A_N(net435));
 sg13g2_o21ai_1 _6706_ (.B1(net436),
    .Y(_0356_),
    .A1(net1254),
    .A2(_2800_));
 sg13g2_nand2_1 _6707_ (.Y(_2801_),
    .A(net432),
    .B(net1180));
 sg13g2_nand2_1 _6708_ (.Y(_2802_),
    .A(\tt6581_inst.mult_inst.accum[0] ),
    .B(\tt6581_inst.mult_inst.a_reg[0] ));
 sg13g2_nand2_1 _6709_ (.Y(_2803_),
    .A(\tt6581_inst.mult_inst.accum[1] ),
    .B(\tt6581_inst.mult_inst.a_reg[1] ));
 sg13g2_xnor2_1 _6710_ (.Y(_2804_),
    .A(net432),
    .B(\tt6581_inst.mult_inst.a_reg[1] ));
 sg13g2_xnor2_1 _6711_ (.Y(_2805_),
    .A(_2802_),
    .B(_2804_));
 sg13g2_o21ai_1 _6712_ (.B1(_2801_),
    .Y(_0357_),
    .A1(net1254),
    .A2(_2805_));
 sg13g2_nand2_1 _6713_ (.Y(_2806_),
    .A(net307),
    .B(net1180));
 sg13g2_and2_1 _6714_ (.A(net307),
    .B(\tt6581_inst.mult_inst.a_reg[2] ),
    .X(_2807_));
 sg13g2_xor2_1 _6715_ (.B(\tt6581_inst.mult_inst.a_reg[2] ),
    .A(net307),
    .X(_2808_));
 sg13g2_o21ai_1 _6716_ (.B1(_2803_),
    .Y(_2809_),
    .A1(_2802_),
    .A2(_2804_));
 sg13g2_xnor2_1 _6717_ (.Y(_2810_),
    .A(_2808_),
    .B(_2809_));
 sg13g2_o21ai_1 _6718_ (.B1(_2806_),
    .Y(_0358_),
    .A1(net1254),
    .A2(_2810_));
 sg13g2_nand2_1 _6719_ (.Y(_2811_),
    .A(net442),
    .B(net1180));
 sg13g2_nand2_1 _6720_ (.Y(_2812_),
    .A(\tt6581_inst.mult_inst.accum[3] ),
    .B(\tt6581_inst.mult_inst.a_reg[3] ));
 sg13g2_xnor2_1 _6721_ (.Y(_2813_),
    .A(net442),
    .B(net273));
 sg13g2_a21oi_1 _6722_ (.A1(_2808_),
    .A2(_2809_),
    .Y(_2814_),
    .B1(_2807_));
 sg13g2_nor2_1 _6723_ (.A(_2813_),
    .B(_2814_),
    .Y(_2815_));
 sg13g2_a21o_1 _6724_ (.A2(_2814_),
    .A1(_2813_),
    .B1(net1254),
    .X(_2816_));
 sg13g2_o21ai_1 _6725_ (.B1(_2811_),
    .Y(_0359_),
    .A1(_2815_),
    .A2(_2816_));
 sg13g2_nand2_1 _6726_ (.Y(_2817_),
    .A(net275),
    .B(net1180));
 sg13g2_a21oi_1 _6727_ (.A1(\tt6581_inst.mult_inst.accum[3] ),
    .A2(net273),
    .Y(_2818_),
    .B1(_2815_));
 sg13g2_o21ai_1 _6728_ (.B1(_2812_),
    .Y(_2819_),
    .A1(_2813_),
    .A2(_2814_));
 sg13g2_and2_1 _6729_ (.A(\tt6581_inst.mult_inst.accum[4] ),
    .B(\tt6581_inst.mult_inst.a_reg[4] ),
    .X(_2820_));
 sg13g2_or2_1 _6730_ (.X(_2821_),
    .B(\tt6581_inst.mult_inst.a_reg[4] ),
    .A(\tt6581_inst.mult_inst.accum[4] ));
 sg13g2_nand2b_1 _6731_ (.Y(_2822_),
    .B(_2821_),
    .A_N(_2820_));
 sg13g2_nor2_1 _6732_ (.A(_2818_),
    .B(_2822_),
    .Y(_2823_));
 sg13g2_a21o_1 _6733_ (.A2(_2822_),
    .A1(_2818_),
    .B1(net1254),
    .X(_2824_));
 sg13g2_o21ai_1 _6734_ (.B1(_2817_),
    .Y(_0360_),
    .A1(_2823_),
    .A2(_2824_));
 sg13g2_nor2_1 _6735_ (.A(_2820_),
    .B(_2823_),
    .Y(_2825_));
 sg13g2_and2_1 _6736_ (.A(net976),
    .B(net206),
    .X(_2826_));
 sg13g2_nor2_1 _6737_ (.A(net976),
    .B(net206),
    .Y(_2827_));
 sg13g2_o21ai_1 _6738_ (.B1(_2825_),
    .Y(_2828_),
    .A1(_2826_),
    .A2(_2827_));
 sg13g2_nor3_1 _6739_ (.A(_2825_),
    .B(_2826_),
    .C(_2827_),
    .Y(_2829_));
 sg13g2_nor2_1 _6740_ (.A(net1254),
    .B(_2829_),
    .Y(_2830_));
 sg13g2_a22oi_1 _6741_ (.Y(_2831_),
    .B1(_2828_),
    .B2(_2830_),
    .A2(net1179),
    .A1(net976));
 sg13g2_inv_1 _6742_ (.Y(_0361_),
    .A(_2831_));
 sg13g2_nand2_1 _6743_ (.Y(_2832_),
    .A(net255),
    .B(net1179));
 sg13g2_and2_1 _6744_ (.A(\tt6581_inst.mult_inst.accum[6] ),
    .B(\tt6581_inst.mult_inst.a_reg[6] ),
    .X(_2833_));
 sg13g2_xnor2_1 _6745_ (.Y(_2834_),
    .A(net255),
    .B(\tt6581_inst.mult_inst.a_reg[6] ));
 sg13g2_a221oi_1 _6746_ (.B2(_2821_),
    .C1(_2820_),
    .B1(_2819_),
    .A1(\tt6581_inst.mult_inst.accum[5] ),
    .Y(_2835_),
    .A2(\tt6581_inst.mult_inst.a_reg[5] ));
 sg13g2_nor3_1 _6747_ (.A(_2827_),
    .B(_2834_),
    .C(_2835_),
    .Y(_2836_));
 sg13g2_o21ai_1 _6748_ (.B1(_2834_),
    .Y(_2837_),
    .A1(_2827_),
    .A2(_2835_));
 sg13g2_nand2_1 _6749_ (.Y(_2838_),
    .A(net1171),
    .B(_2837_));
 sg13g2_o21ai_1 _6750_ (.B1(_2832_),
    .Y(_0362_),
    .A1(_2836_),
    .A2(_2838_));
 sg13g2_nand2_1 _6751_ (.Y(_2839_),
    .A(net977),
    .B(net271));
 sg13g2_xor2_1 _6752_ (.B(net271),
    .A(net977),
    .X(_2840_));
 sg13g2_o21ai_1 _6753_ (.B1(_2840_),
    .Y(_2841_),
    .A1(_2833_),
    .A2(_2836_));
 sg13g2_nor3_1 _6754_ (.A(_2833_),
    .B(_2836_),
    .C(_2840_),
    .Y(_2842_));
 sg13g2_nor2_1 _6755_ (.A(net1255),
    .B(_2842_),
    .Y(_2843_));
 sg13g2_a22oi_1 _6756_ (.Y(_2844_),
    .B1(_2841_),
    .B2(_2843_),
    .A2(net1179),
    .A1(net977));
 sg13g2_inv_1 _6757_ (.Y(_0363_),
    .A(_2844_));
 sg13g2_xnor2_1 _6758_ (.Y(_2845_),
    .A(net1127),
    .B(net803));
 sg13g2_nand3_1 _6759_ (.B(_2841_),
    .C(_2845_),
    .A(_2839_),
    .Y(_2846_));
 sg13g2_a21oi_1 _6760_ (.A1(_2839_),
    .A2(_2841_),
    .Y(_2847_),
    .B1(_2845_));
 sg13g2_nor2_1 _6761_ (.A(net1255),
    .B(_2847_),
    .Y(_2848_));
 sg13g2_a22oi_1 _6762_ (.Y(_2849_),
    .B1(_2846_),
    .B2(_2848_),
    .A2(net1179),
    .A1(net1127));
 sg13g2_inv_1 _6763_ (.Y(_0364_),
    .A(_2849_));
 sg13g2_xor2_1 _6764_ (.B(\tt6581_inst.mult_inst.a_reg[9] ),
    .A(net556),
    .X(_2850_));
 sg13g2_a21oi_1 _6765_ (.A1(\tt6581_inst.mult_inst.accum[8] ),
    .A2(\tt6581_inst.mult_inst.a_reg[8] ),
    .Y(_2851_),
    .B1(_2850_));
 sg13g2_nand2b_1 _6766_ (.Y(_2852_),
    .B(_2851_),
    .A_N(_2847_));
 sg13g2_nand3_1 _6767_ (.B(\tt6581_inst.mult_inst.a_reg[8] ),
    .C(_2850_),
    .A(\tt6581_inst.mult_inst.accum[8] ),
    .Y(_2853_));
 sg13g2_nand3_1 _6768_ (.B(_2852_),
    .C(_2853_),
    .A(net1171),
    .Y(_2854_));
 sg13g2_a21oi_1 _6769_ (.A1(_2847_),
    .A2(_2850_),
    .Y(_2855_),
    .B1(_2854_));
 sg13g2_a21o_1 _6770_ (.A2(net1179),
    .A1(net556),
    .B1(_2855_),
    .X(_0365_));
 sg13g2_xnor2_1 _6771_ (.Y(_2856_),
    .A(net1536),
    .B(net553));
 sg13g2_inv_1 _6772_ (.Y(_2857_),
    .A(_2856_));
 sg13g2_o21ai_1 _6773_ (.B1(_2853_),
    .Y(_2858_),
    .A1(_0910_),
    .A2(_0980_));
 sg13g2_a21oi_1 _6774_ (.A1(_2847_),
    .A2(_2850_),
    .Y(_2859_),
    .B1(_2858_));
 sg13g2_nand2b_1 _6775_ (.Y(_2860_),
    .B(_2857_),
    .A_N(_2859_));
 sg13g2_a21oi_1 _6776_ (.A1(_2856_),
    .A2(_2859_),
    .Y(_2861_),
    .B1(net1255));
 sg13g2_a22oi_1 _6777_ (.Y(_2862_),
    .B1(_2860_),
    .B2(_2861_),
    .A2(net1178),
    .A1(net1536));
 sg13g2_inv_1 _6778_ (.Y(_0366_),
    .A(_2862_));
 sg13g2_xor2_1 _6779_ (.B(net529),
    .A(\tt6581_inst.mult_inst.accum[11] ),
    .X(_2863_));
 sg13g2_a21oi_1 _6780_ (.A1(net1536),
    .A2(net553),
    .Y(_2864_),
    .B1(_2863_));
 sg13g2_nand3b_1 _6781_ (.B(_2863_),
    .C(_2857_),
    .Y(_2865_),
    .A_N(_2859_));
 sg13g2_nand3_1 _6782_ (.B(net553),
    .C(_2863_),
    .A(net1536),
    .Y(_2866_));
 sg13g2_inv_1 _6783_ (.Y(_2867_),
    .A(_2866_));
 sg13g2_nand3_1 _6784_ (.B(_2865_),
    .C(_2866_),
    .A(net1171),
    .Y(_2868_));
 sg13g2_a21oi_1 _6785_ (.A1(_2860_),
    .A2(_2864_),
    .Y(_2869_),
    .B1(_2868_));
 sg13g2_a21o_1 _6786_ (.A2(net1178),
    .A1(net1074),
    .B1(_2869_),
    .X(_0367_));
 sg13g2_nand2_1 _6787_ (.Y(_2870_),
    .A(net491),
    .B(net1178));
 sg13g2_xnor2_1 _6788_ (.Y(_2871_),
    .A(net491),
    .B(\tt6581_inst.mult_inst.a_reg[12] ));
 sg13g2_a21oi_1 _6789_ (.A1(\tt6581_inst.mult_inst.accum[11] ),
    .A2(\tt6581_inst.mult_inst.a_reg[11] ),
    .Y(_2872_),
    .B1(_2867_));
 sg13g2_nand3_1 _6790_ (.B(_2871_),
    .C(_2872_),
    .A(_2865_),
    .Y(_2873_));
 sg13g2_a21oi_1 _6791_ (.A1(_2865_),
    .A2(_2872_),
    .Y(_2874_),
    .B1(_2871_));
 sg13g2_nand2_1 _6792_ (.Y(_2875_),
    .A(net1171),
    .B(_2873_));
 sg13g2_o21ai_1 _6793_ (.B1(_2870_),
    .Y(_0368_),
    .A1(_2874_),
    .A2(_2875_));
 sg13g2_nand2_1 _6794_ (.Y(_2876_),
    .A(\tt6581_inst.mult_inst.accum[13] ),
    .B(net579));
 sg13g2_xor2_1 _6795_ (.B(net579),
    .A(\tt6581_inst.mult_inst.accum[13] ),
    .X(_2877_));
 sg13g2_a21oi_1 _6796_ (.A1(net491),
    .A2(net674),
    .Y(_2878_),
    .B1(_2877_));
 sg13g2_nand2b_1 _6797_ (.Y(_2879_),
    .B(_2878_),
    .A_N(_2874_));
 sg13g2_nand3_1 _6798_ (.B(net674),
    .C(_2877_),
    .A(net491),
    .Y(_2880_));
 sg13g2_nand3_1 _6799_ (.B(_2879_),
    .C(_2880_),
    .A(net1172),
    .Y(_2881_));
 sg13g2_a21oi_1 _6800_ (.A1(_2874_),
    .A2(_2877_),
    .Y(_2882_),
    .B1(_2881_));
 sg13g2_a21o_1 _6801_ (.A2(net1178),
    .A1(net1110),
    .B1(_2882_),
    .X(_0369_));
 sg13g2_nand2_1 _6802_ (.Y(_2883_),
    .A(net690),
    .B(net1178));
 sg13g2_nor2_1 _6803_ (.A(_0913_),
    .B(_0985_),
    .Y(_2884_));
 sg13g2_xnor2_1 _6804_ (.Y(_2885_),
    .A(net690),
    .B(\tt6581_inst.mult_inst.a_reg[14] ));
 sg13g2_inv_1 _6805_ (.Y(_2886_),
    .A(_2885_));
 sg13g2_nand2_1 _6806_ (.Y(_2887_),
    .A(_2876_),
    .B(_2880_));
 sg13g2_a21oi_1 _6807_ (.A1(_2874_),
    .A2(_2877_),
    .Y(_2888_),
    .B1(_2887_));
 sg13g2_nor2_1 _6808_ (.A(_2885_),
    .B(_2888_),
    .Y(_2889_));
 sg13g2_a21o_1 _6809_ (.A2(_2888_),
    .A1(_2885_),
    .B1(net1255),
    .X(_2890_));
 sg13g2_o21ai_1 _6810_ (.B1(_2883_),
    .Y(_0370_),
    .A1(_2889_),
    .A2(_2890_));
 sg13g2_nand2_1 _6811_ (.Y(_2891_),
    .A(net465),
    .B(net1178));
 sg13g2_xor2_1 _6812_ (.B(\tt6581_inst.mult_inst.a_reg[15] ),
    .A(net465),
    .X(_2892_));
 sg13g2_nand3b_1 _6813_ (.B(_2892_),
    .C(_2886_),
    .Y(_2893_),
    .A_N(_2888_));
 sg13g2_nor3_1 _6814_ (.A(_2884_),
    .B(_2889_),
    .C(_2892_),
    .Y(_2894_));
 sg13g2_nand2_1 _6815_ (.Y(_2895_),
    .A(_2884_),
    .B(_2892_));
 sg13g2_inv_1 _6816_ (.Y(_2896_),
    .A(_2895_));
 sg13g2_nand3_1 _6817_ (.B(_2893_),
    .C(_2895_),
    .A(net1172),
    .Y(_2897_));
 sg13g2_o21ai_1 _6818_ (.B1(_2891_),
    .Y(_0371_),
    .A1(_2894_),
    .A2(_2897_));
 sg13g2_and2_1 _6819_ (.A(net1133),
    .B(net1178),
    .X(_2898_));
 sg13g2_xnor2_1 _6820_ (.Y(_2899_),
    .A(net1133),
    .B(net1060));
 sg13g2_a21oi_1 _6821_ (.A1(net465),
    .A2(net1015),
    .Y(_2900_),
    .B1(_2896_));
 sg13g2_a21oi_1 _6822_ (.A1(_2893_),
    .A2(_2900_),
    .Y(_2901_),
    .B1(_2899_));
 sg13g2_nand3_1 _6823_ (.B(_2899_),
    .C(_2900_),
    .A(_2893_),
    .Y(_2902_));
 sg13g2_nor2_1 _6824_ (.A(net1255),
    .B(_2901_),
    .Y(_2903_));
 sg13g2_a21o_1 _6825_ (.A2(_2903_),
    .A1(_2902_),
    .B1(_2898_),
    .X(_0372_));
 sg13g2_nand2_1 _6826_ (.Y(_2904_),
    .A(\tt6581_inst.mult_inst.accum[17] ),
    .B(\tt6581_inst.mult_inst.a_reg[17] ));
 sg13g2_xor2_1 _6827_ (.B(net368),
    .A(\tt6581_inst.mult_inst.accum[17] ),
    .X(_2905_));
 sg13g2_a21oi_1 _6828_ (.A1(\tt6581_inst.mult_inst.accum[16] ),
    .A2(net1060),
    .Y(_2906_),
    .B1(_2905_));
 sg13g2_nand2b_1 _6829_ (.Y(_2907_),
    .B(_2906_),
    .A_N(_2901_));
 sg13g2_nand3_1 _6830_ (.B(net1060),
    .C(_2905_),
    .A(\tt6581_inst.mult_inst.accum[16] ),
    .Y(_2908_));
 sg13g2_nand3_1 _6831_ (.B(_2907_),
    .C(_2908_),
    .A(net1172),
    .Y(_2909_));
 sg13g2_a21oi_1 _6832_ (.A1(_2901_),
    .A2(_2905_),
    .Y(_2910_),
    .B1(_2909_));
 sg13g2_a21o_1 _6833_ (.A2(net1178),
    .A1(net1099),
    .B1(_2910_),
    .X(_0373_));
 sg13g2_nand2_1 _6834_ (.Y(_2911_),
    .A(_2904_),
    .B(_2908_));
 sg13g2_a21oi_1 _6835_ (.A1(_2901_),
    .A2(_2905_),
    .Y(_2912_),
    .B1(_2911_));
 sg13g2_nand2_1 _6836_ (.Y(_2913_),
    .A(\tt6581_inst.mult_inst.accum[18] ),
    .B(net209));
 sg13g2_xnor2_1 _6837_ (.Y(_2914_),
    .A(net1064),
    .B(net209));
 sg13g2_o21ai_1 _6838_ (.B1(net1171),
    .Y(_2915_),
    .A1(_2912_),
    .A2(_2914_));
 sg13g2_a21oi_1 _6839_ (.A1(_2912_),
    .A2(_2914_),
    .Y(_2916_),
    .B1(_2915_));
 sg13g2_a21o_1 _6840_ (.A2(net1180),
    .A1(net1064),
    .B1(_2916_),
    .X(_0374_));
 sg13g2_o21ai_1 _6841_ (.B1(_2913_),
    .Y(_2917_),
    .A1(_2912_),
    .A2(_2914_));
 sg13g2_and2_1 _6842_ (.A(\tt6581_inst.mult_inst.accum[19] ),
    .B(\tt6581_inst.mult_inst.a_reg[19] ),
    .X(_2918_));
 sg13g2_or2_1 _6843_ (.X(_2919_),
    .B(\tt6581_inst.mult_inst.a_reg[19] ),
    .A(\tt6581_inst.mult_inst.accum[19] ));
 sg13g2_nor2b_1 _6844_ (.A(_2918_),
    .B_N(_2919_),
    .Y(_2920_));
 sg13g2_o21ai_1 _6845_ (.B1(net1171),
    .Y(_2921_),
    .A1(_2917_),
    .A2(_2920_));
 sg13g2_a21oi_1 _6846_ (.A1(_2917_),
    .A2(_2920_),
    .Y(_2922_),
    .B1(_2921_));
 sg13g2_a21o_1 _6847_ (.A2(net1181),
    .A1(net841),
    .B1(_2922_),
    .X(_0375_));
 sg13g2_nand2_1 _6848_ (.Y(_2923_),
    .A(net589),
    .B(net1181));
 sg13g2_and2_1 _6849_ (.A(net589),
    .B(net243),
    .X(_2924_));
 sg13g2_xnor2_1 _6850_ (.Y(_2925_),
    .A(net589),
    .B(net243));
 sg13g2_inv_1 _6851_ (.Y(_2926_),
    .A(_2925_));
 sg13g2_a21oi_1 _6852_ (.A1(_2917_),
    .A2(_2919_),
    .Y(_2927_),
    .B1(_2918_));
 sg13g2_nor2_1 _6853_ (.A(_2925_),
    .B(_2927_),
    .Y(_2928_));
 sg13g2_a21o_1 _6854_ (.A2(_2927_),
    .A1(_2925_),
    .B1(net1254),
    .X(_2929_));
 sg13g2_o21ai_1 _6855_ (.B1(_2923_),
    .Y(_0376_),
    .A1(_2928_),
    .A2(_2929_));
 sg13g2_nand2_1 _6856_ (.Y(_2930_),
    .A(net662),
    .B(net1181));
 sg13g2_nand2_1 _6857_ (.Y(_2931_),
    .A(\tt6581_inst.mult_inst.accum[21] ),
    .B(\tt6581_inst.mult_inst.a_reg[21] ));
 sg13g2_xor2_1 _6858_ (.B(net550),
    .A(net662),
    .X(_2932_));
 sg13g2_nor3_1 _6859_ (.A(_2924_),
    .B(_2928_),
    .C(_2932_),
    .Y(_2933_));
 sg13g2_nand3b_1 _6860_ (.B(_2932_),
    .C(_2926_),
    .Y(_2934_),
    .A_N(_2927_));
 sg13g2_nand2_1 _6861_ (.Y(_2935_),
    .A(_2924_),
    .B(_2932_));
 sg13g2_nand3_1 _6862_ (.B(_2934_),
    .C(_2935_),
    .A(net1171),
    .Y(_2936_));
 sg13g2_o21ai_1 _6863_ (.B1(_2930_),
    .Y(_0377_),
    .A1(_2933_),
    .A2(_2936_));
 sg13g2_nand2_1 _6864_ (.Y(_2937_),
    .A(net495),
    .B(net1181));
 sg13g2_and2_1 _6865_ (.A(_2931_),
    .B(_2935_),
    .X(_2938_));
 sg13g2_nand2_1 _6866_ (.Y(_2939_),
    .A(_2934_),
    .B(_2938_));
 sg13g2_nand2_1 _6867_ (.Y(_2940_),
    .A(net252),
    .B(\tt6581_inst.mult_inst.accum[22] ));
 sg13g2_xor2_1 _6868_ (.B(net495),
    .A(net252),
    .X(_2941_));
 sg13g2_inv_1 _6869_ (.Y(_2942_),
    .A(_2941_));
 sg13g2_a21oi_1 _6870_ (.A1(_2934_),
    .A2(_2938_),
    .Y(_2943_),
    .B1(_2942_));
 sg13g2_a21o_1 _6871_ (.A2(_2938_),
    .A1(_2934_),
    .B1(_2942_),
    .X(_2944_));
 sg13g2_o21ai_1 _6872_ (.B1(net1171),
    .Y(_2945_),
    .A1(_2939_),
    .A2(_2941_));
 sg13g2_o21ai_1 _6873_ (.B1(_2937_),
    .Y(_0378_),
    .A1(_2943_),
    .A2(_2945_));
 sg13g2_and2_1 _6874_ (.A(_2940_),
    .B(_2944_),
    .X(_2946_));
 sg13g2_and2_1 _6875_ (.A(\tt6581_inst.mult_inst.a_reg[23] ),
    .B(\tt6581_inst.mult_inst.accum[23] ),
    .X(_2947_));
 sg13g2_nand2_1 _6876_ (.Y(_2948_),
    .A(net776),
    .B(net1125));
 sg13g2_nor2_1 _6877_ (.A(net776),
    .B(\tt6581_inst.mult_inst.accum[23] ),
    .Y(_2949_));
 sg13g2_a21oi_2 _6878_ (.B1(_2949_),
    .Y(_2950_),
    .A2(_2944_),
    .A1(_2940_));
 sg13g2_o21ai_1 _6879_ (.B1(_2946_),
    .Y(_2951_),
    .A1(_2947_),
    .A2(_2949_));
 sg13g2_a21oi_1 _6880_ (.A1(_2948_),
    .A2(_2950_),
    .Y(_2952_),
    .B1(net1254));
 sg13g2_a22oi_1 _6881_ (.Y(_2953_),
    .B1(_2951_),
    .B2(_2952_),
    .A2(net1181),
    .A1(net1125));
 sg13g2_inv_1 _6882_ (.Y(_0379_),
    .A(net1126));
 sg13g2_nand2_1 _6883_ (.Y(_2954_),
    .A(net477),
    .B(\tt6581_inst.mult_inst.accum[24] ));
 sg13g2_xor2_1 _6884_ (.B(net1122),
    .A(net477),
    .X(_2955_));
 sg13g2_or2_1 _6885_ (.X(_2956_),
    .B(_2950_),
    .A(_2947_));
 sg13g2_nand2_1 _6886_ (.Y(_2957_),
    .A(_2955_),
    .B(_2956_));
 sg13g2_o21ai_1 _6887_ (.B1(net1168),
    .Y(_2958_),
    .A1(_2955_),
    .A2(_2956_));
 sg13g2_inv_1 _6888_ (.Y(_2959_),
    .A(_2958_));
 sg13g2_a22oi_1 _6889_ (.Y(_2960_),
    .B1(_2957_),
    .B2(_2959_),
    .A2(net1175),
    .A1(net1122));
 sg13g2_inv_1 _6890_ (.Y(_0380_),
    .A(_2960_));
 sg13g2_nor2_1 _6891_ (.A(\tt6581_inst.mult_inst.a_reg[25] ),
    .B(\tt6581_inst.mult_inst.accum[25] ),
    .Y(_2961_));
 sg13g2_nand2_1 _6892_ (.Y(_2962_),
    .A(net525),
    .B(net1071));
 sg13g2_nor2b_1 _6893_ (.A(_2961_),
    .B_N(_2962_),
    .Y(_2963_));
 sg13g2_nand2_1 _6894_ (.Y(_2964_),
    .A(_2954_),
    .B(_2957_));
 sg13g2_nand2_1 _6895_ (.Y(_2965_),
    .A(_2963_),
    .B(_2964_));
 sg13g2_o21ai_1 _6896_ (.B1(net1168),
    .Y(_2966_),
    .A1(_2963_),
    .A2(_2964_));
 sg13g2_nor2b_1 _6897_ (.A(_2966_),
    .B_N(_2965_),
    .Y(_2967_));
 sg13g2_a21o_1 _6898_ (.A2(net1175),
    .A1(net1071),
    .B1(_2967_),
    .X(_0381_));
 sg13g2_nand2_1 _6899_ (.Y(_2968_),
    .A(net1098),
    .B(net1175));
 sg13g2_xor2_1 _6900_ (.B(net1098),
    .A(net627),
    .X(_2969_));
 sg13g2_inv_1 _6901_ (.Y(_2970_),
    .A(_2969_));
 sg13g2_nand2_1 _6902_ (.Y(_2971_),
    .A(_2962_),
    .B(_2965_));
 sg13g2_a21oi_1 _6903_ (.A1(_2962_),
    .A2(_2965_),
    .Y(_2972_),
    .B1(_2970_));
 sg13g2_o21ai_1 _6904_ (.B1(net1168),
    .Y(_2973_),
    .A1(_2969_),
    .A2(_2971_));
 sg13g2_o21ai_1 _6905_ (.B1(_2968_),
    .Y(_0382_),
    .A1(_2972_),
    .A2(_2973_));
 sg13g2_or2_1 _6906_ (.X(_2974_),
    .B(\tt6581_inst.mult_inst.accum[27] ),
    .A(\tt6581_inst.mult_inst.a_reg[27] ));
 sg13g2_xnor2_1 _6907_ (.Y(_2975_),
    .A(net583),
    .B(net1090));
 sg13g2_a21oi_1 _6908_ (.A1(net627),
    .A2(\tt6581_inst.mult_inst.accum[26] ),
    .Y(_2976_),
    .B1(_2972_));
 sg13g2_o21ai_1 _6909_ (.B1(net1168),
    .Y(_2977_),
    .A1(_2975_),
    .A2(_2976_));
 sg13g2_a21oi_1 _6910_ (.A1(_2975_),
    .A2(_2976_),
    .Y(_2978_),
    .B1(_2977_));
 sg13g2_a21o_1 _6911_ (.A2(net1175),
    .A1(net1090),
    .B1(_2978_),
    .X(_0383_));
 sg13g2_nand2_1 _6912_ (.Y(_2979_),
    .A(net606),
    .B(net1175));
 sg13g2_nor2_1 _6913_ (.A(_2970_),
    .B(_2975_),
    .Y(_2980_));
 sg13g2_and3_1 _6914_ (.X(_2981_),
    .A(_2955_),
    .B(_2963_),
    .C(_2980_));
 sg13g2_o21ai_1 _6915_ (.B1(_2981_),
    .Y(_2982_),
    .A1(_2947_),
    .A2(_2950_));
 sg13g2_o21ai_1 _6916_ (.B1(_2962_),
    .Y(_2983_),
    .A1(_2954_),
    .A2(_2961_));
 sg13g2_and3_1 _6917_ (.X(_2984_),
    .A(\tt6581_inst.mult_inst.a_reg[26] ),
    .B(\tt6581_inst.mult_inst.accum[26] ),
    .C(_2974_));
 sg13g2_a221oi_1 _6918_ (.B2(_2983_),
    .C1(_2984_),
    .B1(_2980_),
    .A1(\tt6581_inst.mult_inst.a_reg[27] ),
    .Y(_2985_),
    .A2(\tt6581_inst.mult_inst.accum[27] ));
 sg13g2_nand2_1 _6919_ (.Y(_2986_),
    .A(_2982_),
    .B(_2985_));
 sg13g2_xor2_1 _6920_ (.B(net606),
    .A(\tt6581_inst.mult_inst.a_reg[28] ),
    .X(_2987_));
 sg13g2_and2_1 _6921_ (.A(_2986_),
    .B(_2987_),
    .X(_2988_));
 sg13g2_nand2_1 _6922_ (.Y(_2989_),
    .A(_2986_),
    .B(_2987_));
 sg13g2_o21ai_1 _6923_ (.B1(net1168),
    .Y(_2990_),
    .A1(_2986_),
    .A2(_2987_));
 sg13g2_o21ai_1 _6924_ (.B1(_2979_),
    .Y(_0384_),
    .A1(_2988_),
    .A2(_2990_));
 sg13g2_xnor2_1 _6925_ (.Y(_2991_),
    .A(net519),
    .B(net573));
 sg13g2_inv_1 _6926_ (.Y(_2992_),
    .A(_2991_));
 sg13g2_a21oi_1 _6927_ (.A1(\tt6581_inst.mult_inst.a_reg[28] ),
    .A2(\tt6581_inst.mult_inst.accum[28] ),
    .Y(_2993_),
    .B1(_2988_));
 sg13g2_and3_1 _6928_ (.X(_2994_),
    .A(\tt6581_inst.mult_inst.a_reg[28] ),
    .B(\tt6581_inst.mult_inst.accum[28] ),
    .C(_2992_));
 sg13g2_o21ai_1 _6929_ (.B1(net1168),
    .Y(_2995_),
    .A1(_2991_),
    .A2(_2993_));
 sg13g2_a21oi_1 _6930_ (.A1(_2991_),
    .A2(_2993_),
    .Y(_2996_),
    .B1(_2995_));
 sg13g2_a21o_1 _6931_ (.A2(net1175),
    .A1(net573),
    .B1(_2996_),
    .X(_0385_));
 sg13g2_nand2_1 _6932_ (.Y(_2997_),
    .A(net610),
    .B(net1175));
 sg13g2_and2_1 _6933_ (.A(\tt6581_inst.mult_inst.a_reg[30] ),
    .B(\tt6581_inst.mult_inst.accum[30] ),
    .X(_2998_));
 sg13g2_xor2_1 _6934_ (.B(net610),
    .A(net538),
    .X(_2999_));
 sg13g2_inv_1 _6935_ (.Y(_3000_),
    .A(_2999_));
 sg13g2_a21oi_1 _6936_ (.A1(net519),
    .A2(\tt6581_inst.mult_inst.accum[29] ),
    .Y(_3001_),
    .B1(_2994_));
 sg13g2_o21ai_1 _6937_ (.B1(_3001_),
    .Y(_3002_),
    .A1(_2989_),
    .A2(_2991_));
 sg13g2_and2_1 _6938_ (.A(_2999_),
    .B(_3002_),
    .X(_3003_));
 sg13g2_o21ai_1 _6939_ (.B1(net1168),
    .Y(_3004_),
    .A1(_2999_),
    .A2(_3002_));
 sg13g2_o21ai_1 _6940_ (.B1(_2997_),
    .Y(_0386_),
    .A1(_3003_),
    .A2(_3004_));
 sg13g2_xnor2_1 _6941_ (.Y(_3005_),
    .A(net816),
    .B(net1083));
 sg13g2_inv_1 _6942_ (.Y(_3006_),
    .A(_3005_));
 sg13g2_nor2_1 _6943_ (.A(_2998_),
    .B(_3003_),
    .Y(_3007_));
 sg13g2_o21ai_1 _6944_ (.B1(net1168),
    .Y(_3008_),
    .A1(_3005_),
    .A2(_3007_));
 sg13g2_a21oi_1 _6945_ (.A1(_3005_),
    .A2(_3007_),
    .Y(_3009_),
    .B1(_3008_));
 sg13g2_a21o_1 _6946_ (.A2(net1175),
    .A1(net1083),
    .B1(_3009_),
    .X(_0387_));
 sg13g2_nand2_1 _6947_ (.Y(_3010_),
    .A(net482),
    .B(\tt6581_inst.mult_inst.accum[32] ));
 sg13g2_xor2_1 _6948_ (.B(\tt6581_inst.mult_inst.accum[32] ),
    .A(\tt6581_inst.mult_inst.a_reg[32] ),
    .X(_3011_));
 sg13g2_nand4_1 _6949_ (.B(_2992_),
    .C(_2999_),
    .A(_2987_),
    .Y(_3012_),
    .D(_3006_));
 sg13g2_a21oi_1 _6950_ (.A1(_2982_),
    .A2(_2985_),
    .Y(_3013_),
    .B1(_3012_));
 sg13g2_nor3_1 _6951_ (.A(_3000_),
    .B(_3001_),
    .C(_3005_),
    .Y(_3014_));
 sg13g2_o21ai_1 _6952_ (.B1(_2998_),
    .Y(_3015_),
    .A1(\tt6581_inst.mult_inst.a_reg[31] ),
    .A2(\tt6581_inst.mult_inst.accum[31] ));
 sg13g2_a21oi_1 _6953_ (.A1(\tt6581_inst.mult_inst.a_reg[31] ),
    .A2(\tt6581_inst.mult_inst.accum[31] ),
    .Y(_3016_),
    .B1(_3014_));
 sg13g2_and2_1 _6954_ (.A(_3015_),
    .B(_3016_),
    .X(_3017_));
 sg13g2_inv_1 _6955_ (.Y(_3018_),
    .A(_3017_));
 sg13g2_o21ai_1 _6956_ (.B1(_3011_),
    .Y(_3019_),
    .A1(_3013_),
    .A2(_3018_));
 sg13g2_or3_1 _6957_ (.A(_3011_),
    .B(_3013_),
    .C(_3018_),
    .X(_3020_));
 sg13g2_and2_1 _6958_ (.A(net1169),
    .B(_3019_),
    .X(_3021_));
 sg13g2_a22oi_1 _6959_ (.Y(_3022_),
    .B1(_3020_),
    .B2(_3021_),
    .A2(net1176),
    .A1(net1096));
 sg13g2_inv_1 _6960_ (.Y(_0388_),
    .A(net1097));
 sg13g2_nand2_1 _6961_ (.Y(_3023_),
    .A(_3010_),
    .B(_3019_));
 sg13g2_nand2_1 _6962_ (.Y(_3024_),
    .A(net511),
    .B(net997));
 sg13g2_or2_1 _6963_ (.X(_3025_),
    .B(\tt6581_inst.mult_inst.accum[33] ),
    .A(\tt6581_inst.mult_inst.a_reg[33] ));
 sg13g2_and2_1 _6964_ (.A(_3024_),
    .B(_3025_),
    .X(_3026_));
 sg13g2_o21ai_1 _6965_ (.B1(net1169),
    .Y(_3027_),
    .A1(_3023_),
    .A2(_3026_));
 sg13g2_a21oi_1 _6966_ (.A1(_3023_),
    .A2(_3026_),
    .Y(_3028_),
    .B1(_3027_));
 sg13g2_a21o_1 _6967_ (.A2(net1176),
    .A1(net997),
    .B1(_3028_),
    .X(_0389_));
 sg13g2_and2_1 _6968_ (.A(net555),
    .B(\tt6581_inst.mult_inst.accum[34] ),
    .X(_3029_));
 sg13g2_xor2_1 _6969_ (.B(net723),
    .A(net555),
    .X(_3030_));
 sg13g2_nand3_1 _6970_ (.B(_3019_),
    .C(_3024_),
    .A(_3010_),
    .Y(_3031_));
 sg13g2_and2_1 _6971_ (.A(_3025_),
    .B(_3031_),
    .X(_3032_));
 sg13g2_and3_1 _6972_ (.X(_3033_),
    .A(_3025_),
    .B(_3030_),
    .C(_3031_));
 sg13g2_o21ai_1 _6973_ (.B1(net1169),
    .Y(_3034_),
    .A1(_3030_),
    .A2(_3032_));
 sg13g2_nor2_1 _6974_ (.A(_3033_),
    .B(_3034_),
    .Y(_3035_));
 sg13g2_a21oi_1 _6975_ (.A1(net723),
    .A2(net1176),
    .Y(_3036_),
    .B1(_3035_));
 sg13g2_inv_1 _6976_ (.Y(_0390_),
    .A(_3036_));
 sg13g2_nor2_1 _6977_ (.A(_3029_),
    .B(_3033_),
    .Y(_3037_));
 sg13g2_nand2_1 _6978_ (.Y(_3038_),
    .A(net484),
    .B(net706));
 sg13g2_or2_1 _6979_ (.X(_3039_),
    .B(\tt6581_inst.mult_inst.accum[35] ),
    .A(\tt6581_inst.mult_inst.a_reg[35] ));
 sg13g2_nand2_1 _6980_ (.Y(_3040_),
    .A(_3038_),
    .B(_3039_));
 sg13g2_o21ai_1 _6981_ (.B1(net1169),
    .Y(_3041_),
    .A1(_3037_),
    .A2(_3040_));
 sg13g2_a21oi_1 _6982_ (.A1(_3037_),
    .A2(_3040_),
    .Y(_3042_),
    .B1(_3041_));
 sg13g2_a21o_1 _6983_ (.A2(net1176),
    .A1(net706),
    .B1(_3042_),
    .X(_0391_));
 sg13g2_nand2_1 _6984_ (.Y(_3043_),
    .A(net380),
    .B(net1177));
 sg13g2_xnor2_1 _6985_ (.Y(_3044_),
    .A(\tt6581_inst.mult_inst.a_reg[36] ),
    .B(net380));
 sg13g2_o21ai_1 _6986_ (.B1(_3039_),
    .Y(_3045_),
    .A1(_3029_),
    .A2(_3033_));
 sg13g2_a21oi_1 _6987_ (.A1(_3038_),
    .A2(_3045_),
    .Y(_3046_),
    .B1(_3044_));
 sg13g2_nand3_1 _6988_ (.B(_3044_),
    .C(_3045_),
    .A(_3038_),
    .Y(_3047_));
 sg13g2_nand2_1 _6989_ (.Y(_3048_),
    .A(net1170),
    .B(_3047_));
 sg13g2_o21ai_1 _6990_ (.B1(_3043_),
    .Y(_0392_),
    .A1(_3046_),
    .A2(_3048_));
 sg13g2_a21oi_1 _6991_ (.A1(net508),
    .A2(net380),
    .Y(_3049_),
    .B1(_3046_));
 sg13g2_nand2_1 _6992_ (.Y(_3050_),
    .A(\tt6581_inst.mult_inst.a_reg[37] ),
    .B(\tt6581_inst.mult_inst.accum[37] ));
 sg13g2_nor2_1 _6993_ (.A(\tt6581_inst.mult_inst.a_reg[37] ),
    .B(\tt6581_inst.mult_inst.accum[37] ),
    .Y(_3051_));
 sg13g2_xnor2_1 _6994_ (.Y(_3052_),
    .A(net533),
    .B(net1032));
 sg13g2_o21ai_1 _6995_ (.B1(net1170),
    .Y(_3053_),
    .A1(_3049_),
    .A2(_3052_));
 sg13g2_a21oi_1 _6996_ (.A1(_3049_),
    .A2(_3052_),
    .Y(_3054_),
    .B1(_3053_));
 sg13g2_a21o_1 _6997_ (.A2(net1177),
    .A1(net1032),
    .B1(_3054_),
    .X(_0393_));
 sg13g2_nand2_1 _6998_ (.Y(_3055_),
    .A(net211),
    .B(net1177));
 sg13g2_xor2_1 _6999_ (.B(net211),
    .A(\tt6581_inst.mult_inst.a_reg[38] ),
    .X(_3056_));
 sg13g2_a21oi_1 _7000_ (.A1(_3049_),
    .A2(_3050_),
    .Y(_3057_),
    .B1(_3051_));
 sg13g2_and2_1 _7001_ (.A(_3056_),
    .B(_3057_),
    .X(_3058_));
 sg13g2_o21ai_1 _7002_ (.B1(net1170),
    .Y(_3059_),
    .A1(_3056_),
    .A2(_3057_));
 sg13g2_o21ai_1 _7003_ (.B1(_3055_),
    .Y(_0394_),
    .A1(_3058_),
    .A2(_3059_));
 sg13g2_and2_1 _7004_ (.A(net462),
    .B(net138),
    .X(_3060_));
 sg13g2_and2_1 _7005_ (.A(net577),
    .B(_3060_),
    .X(_3061_));
 sg13g2_nand2b_1 _7006_ (.Y(_3062_),
    .B(net35),
    .A_N(net845));
 sg13g2_nor2_2 _7007_ (.A(net826),
    .B(_3062_),
    .Y(_3063_));
 sg13g2_or2_1 _7008_ (.X(_3064_),
    .B(_3062_),
    .A(\tt6581_inst.spi_inst.cs_sync[1] ));
 sg13g2_nand2_2 _7009_ (.Y(_3065_),
    .A(_3061_),
    .B(_3063_));
 sg13g2_nor2_2 _7010_ (.A(net823),
    .B(_3065_),
    .Y(_3066_));
 sg13g2_nand2_1 _7011_ (.Y(_3067_),
    .A(net245),
    .B(_3066_));
 sg13g2_o21ai_1 _7012_ (.B1(net246),
    .Y(_0395_),
    .A1(_0878_),
    .A2(_3066_));
 sg13g2_nand2_1 _7013_ (.Y(_3068_),
    .A(net1521),
    .B(_1110_));
 sg13g2_xnor2_1 _7014_ (.Y(_0396_),
    .A(net383),
    .B(_3068_));
 sg13g2_nor2_1 _7015_ (.A(net1508),
    .B(net1521),
    .Y(_3069_));
 sg13g2_o21ai_1 _7016_ (.B1(net383),
    .Y(_3070_),
    .A1(_1108_),
    .A2(_1109_));
 sg13g2_o21ai_1 _7017_ (.B1(net1508),
    .Y(_3071_),
    .A1(_1122_),
    .A2(_1123_));
 sg13g2_nor3_1 _7018_ (.A(net1508),
    .B(_1122_),
    .C(_1123_),
    .Y(_3072_));
 sg13g2_xnor2_1 _7019_ (.Y(_3073_),
    .A(net1508),
    .B(net1184));
 sg13g2_xnor2_1 _7020_ (.Y(_3074_),
    .A(_3070_),
    .B(_3073_));
 sg13g2_a21oi_1 _7021_ (.A1(net1521),
    .A2(_3074_),
    .Y(_0397_),
    .B1(_3069_));
 sg13g2_and2_1 _7022_ (.A(net991),
    .B(net1182),
    .X(_3075_));
 sg13g2_or2_1 _7023_ (.X(_3076_),
    .B(net1182),
    .A(\tt6581_inst.svf_inst.reg_low[2] ));
 sg13g2_nor2b_1 _7024_ (.A(_3075_),
    .B_N(_3076_),
    .Y(_3077_));
 sg13g2_o21ai_1 _7025_ (.B1(_3071_),
    .Y(_3078_),
    .A1(_3070_),
    .A2(_3072_));
 sg13g2_xnor2_1 _7026_ (.Y(_3079_),
    .A(_3077_),
    .B(_3078_));
 sg13g2_nor2_1 _7027_ (.A(net991),
    .B(net1519),
    .Y(_3080_));
 sg13g2_a21oi_1 _7028_ (.A1(net1520),
    .A2(_3079_),
    .Y(_0398_),
    .B1(_3080_));
 sg13g2_nand2_1 _7029_ (.Y(_3081_),
    .A(net1507),
    .B(net1173));
 sg13g2_xnor2_1 _7030_ (.Y(_3082_),
    .A(net1507),
    .B(net1173));
 sg13g2_a21oi_1 _7031_ (.A1(_3076_),
    .A2(_3078_),
    .Y(_3083_),
    .B1(_3075_));
 sg13g2_xnor2_1 _7032_ (.Y(_3084_),
    .A(_3082_),
    .B(_3083_));
 sg13g2_nor2_1 _7033_ (.A(net1507),
    .B(net1519),
    .Y(_3085_));
 sg13g2_a21oi_1 _7034_ (.A1(net1519),
    .A2(_3084_),
    .Y(_0399_),
    .B1(_3085_));
 sg13g2_and2_1 _7035_ (.A(net971),
    .B(net1166),
    .X(_3086_));
 sg13g2_or2_1 _7036_ (.X(_3087_),
    .B(net1166),
    .A(\tt6581_inst.svf_inst.reg_low[4] ));
 sg13g2_nor2b_1 _7037_ (.A(_3086_),
    .B_N(_3087_),
    .Y(_3088_));
 sg13g2_o21ai_1 _7038_ (.B1(_3081_),
    .Y(_3089_),
    .A1(_3082_),
    .A2(_3083_));
 sg13g2_xnor2_1 _7039_ (.Y(_3090_),
    .A(_3088_),
    .B(_3089_));
 sg13g2_nor2_1 _7040_ (.A(net971),
    .B(net1519),
    .Y(_3091_));
 sg13g2_a21oi_1 _7041_ (.A1(net1519),
    .A2(_3090_),
    .Y(_0400_),
    .B1(_3091_));
 sg13g2_nor2_1 _7042_ (.A(net1506),
    .B(net1519),
    .Y(_3092_));
 sg13g2_a21oi_1 _7043_ (.A1(_3087_),
    .A2(_3089_),
    .Y(_3093_),
    .B1(_3086_));
 sg13g2_nor2_1 _7044_ (.A(net1506),
    .B(net1164),
    .Y(_3094_));
 sg13g2_xnor2_1 _7045_ (.Y(_3095_),
    .A(net1691),
    .B(net1165));
 sg13g2_xnor2_1 _7046_ (.Y(_3096_),
    .A(_3093_),
    .B(_3095_));
 sg13g2_a21oi_1 _7047_ (.A1(net1519),
    .A2(_3096_),
    .Y(_0401_),
    .B1(_3092_));
 sg13g2_nor2_1 _7048_ (.A(_0940_),
    .B(_1188_),
    .Y(_3097_));
 sg13g2_xnor2_1 _7049_ (.Y(_3098_),
    .A(\tt6581_inst.svf_inst.reg_low[6] ),
    .B(_1187_));
 sg13g2_a221oi_1 _7050_ (.B2(_3089_),
    .C1(_3086_),
    .B1(_3087_),
    .A1(\tt6581_inst.svf_inst.reg_low[5] ),
    .Y(_3099_),
    .A2(net1165));
 sg13g2_nor3_1 _7051_ (.A(_3094_),
    .B(_3098_),
    .C(_3099_),
    .Y(_3100_));
 sg13g2_o21ai_1 _7052_ (.B1(_3098_),
    .Y(_3101_),
    .A1(_3094_),
    .A2(_3099_));
 sg13g2_nand2b_1 _7053_ (.Y(_3102_),
    .B(_3101_),
    .A_N(_3100_));
 sg13g2_mux2_1 _7054_ (.A0(_0940_),
    .A1(_3102_),
    .S(net1519),
    .X(_3103_));
 sg13g2_inv_1 _7055_ (.Y(_0402_),
    .A(_3103_));
 sg13g2_nand2_1 _7056_ (.Y(_3104_),
    .A(net1115),
    .B(_1200_));
 sg13g2_xnor2_1 _7057_ (.Y(_3105_),
    .A(\tt6581_inst.svf_inst.reg_low[7] ),
    .B(_1200_));
 sg13g2_inv_1 _7058_ (.Y(_3106_),
    .A(_3105_));
 sg13g2_o21ai_1 _7059_ (.B1(_3106_),
    .Y(_3107_),
    .A1(_3097_),
    .A2(_3100_));
 sg13g2_nor3_1 _7060_ (.A(_3097_),
    .B(_3100_),
    .C(_3106_),
    .Y(_3108_));
 sg13g2_nand3b_1 _7061_ (.B(net1520),
    .C(_3107_),
    .Y(_3109_),
    .A_N(_3108_));
 sg13g2_o21ai_1 _7062_ (.B1(_3109_),
    .Y(_0403_),
    .A1(_0939_),
    .A2(net1520));
 sg13g2_xnor2_1 _7063_ (.Y(_3110_),
    .A(\tt6581_inst.svf_inst.reg_low[8] ),
    .B(_1211_));
 sg13g2_a21oi_1 _7064_ (.A1(_3104_),
    .A2(_3107_),
    .Y(_3111_),
    .B1(_3110_));
 sg13g2_nand3_1 _7065_ (.B(_3107_),
    .C(_3110_),
    .A(_3104_),
    .Y(_3112_));
 sg13g2_nand3b_1 _7066_ (.B(_3112_),
    .C(net1522),
    .Y(_3113_),
    .A_N(_3111_));
 sg13g2_o21ai_1 _7067_ (.B1(_3113_),
    .Y(_0404_),
    .A1(_0938_),
    .A2(net1522));
 sg13g2_a21oi_1 _7068_ (.A1(net1128),
    .A2(_1211_),
    .Y(_3114_),
    .B1(_3111_));
 sg13g2_nor2_1 _7069_ (.A(net1505),
    .B(_1225_),
    .Y(_3115_));
 sg13g2_xor2_1 _7070_ (.B(_1224_),
    .A(net1505),
    .X(_3116_));
 sg13g2_xnor2_1 _7071_ (.Y(_3117_),
    .A(_3114_),
    .B(_3116_));
 sg13g2_nor2_1 _7072_ (.A(net1505),
    .B(net1522),
    .Y(_3118_));
 sg13g2_a21oi_1 _7073_ (.A1(net1522),
    .A2(_3117_),
    .Y(_0405_),
    .B1(net1693));
 sg13g2_and2_1 _7074_ (.A(\tt6581_inst.svf_inst.reg_low[10] ),
    .B(_1239_),
    .X(_3119_));
 sg13g2_xnor2_1 _7075_ (.Y(_3120_),
    .A(net1118),
    .B(_1239_));
 sg13g2_a221oi_1 _7076_ (.B2(net1505),
    .C1(_3111_),
    .B1(_1225_),
    .A1(\tt6581_inst.svf_inst.reg_low[8] ),
    .Y(_3121_),
    .A2(_1211_));
 sg13g2_nor3_1 _7077_ (.A(_3115_),
    .B(_3120_),
    .C(_3121_),
    .Y(_3122_));
 sg13g2_o21ai_1 _7078_ (.B1(_3120_),
    .Y(_3123_),
    .A1(_3115_),
    .A2(_3121_));
 sg13g2_nand3b_1 _7079_ (.B(_3123_),
    .C(net1522),
    .Y(_3124_),
    .A_N(_3122_));
 sg13g2_o21ai_1 _7080_ (.B1(_3124_),
    .Y(_0406_),
    .A1(_0937_),
    .A2(net1522));
 sg13g2_nor2_1 _7081_ (.A(_3119_),
    .B(_3122_),
    .Y(_3125_));
 sg13g2_nand2_1 _7082_ (.Y(_3126_),
    .A(net1076),
    .B(_1253_));
 sg13g2_nand2_1 _7083_ (.Y(_3127_),
    .A(_0936_),
    .B(_1254_));
 sg13g2_nand2_1 _7084_ (.Y(_3128_),
    .A(_3126_),
    .B(_3127_));
 sg13g2_xnor2_1 _7085_ (.Y(_3129_),
    .A(_3125_),
    .B(_3128_));
 sg13g2_nor2_1 _7086_ (.A(net1076),
    .B(net1518),
    .Y(_3130_));
 sg13g2_a21oi_1 _7087_ (.A1(net1518),
    .A2(_3129_),
    .Y(_0407_),
    .B1(net1077));
 sg13g2_and2_1 _7088_ (.A(\tt6581_inst.svf_inst.reg_low[12] ),
    .B(_1267_),
    .X(_3131_));
 sg13g2_xnor2_1 _7089_ (.Y(_3132_),
    .A(net1116),
    .B(_1267_));
 sg13g2_o21ai_1 _7090_ (.B1(_3127_),
    .Y(_3133_),
    .A1(_3119_),
    .A2(_3122_));
 sg13g2_a21oi_1 _7091_ (.A1(_3126_),
    .A2(_3133_),
    .Y(_3134_),
    .B1(_3132_));
 sg13g2_nand3_1 _7092_ (.B(_3132_),
    .C(_3133_),
    .A(_3126_),
    .Y(_3135_));
 sg13g2_nand3b_1 _7093_ (.B(_3135_),
    .C(net1518),
    .Y(_3136_),
    .A_N(_3134_));
 sg13g2_o21ai_1 _7094_ (.B1(_3136_),
    .Y(_0408_),
    .A1(_0934_),
    .A2(net1518));
 sg13g2_nor2_1 _7095_ (.A(_3131_),
    .B(_3134_),
    .Y(_3137_));
 sg13g2_nand2_1 _7096_ (.Y(_3138_),
    .A(net1041),
    .B(_1280_));
 sg13g2_or2_1 _7097_ (.X(_3139_),
    .B(_1280_),
    .A(\tt6581_inst.svf_inst.reg_low[13] ));
 sg13g2_nand2_1 _7098_ (.Y(_3140_),
    .A(_3138_),
    .B(_3139_));
 sg13g2_xnor2_1 _7099_ (.Y(_3141_),
    .A(_3137_),
    .B(_3140_));
 sg13g2_nor2_1 _7100_ (.A(net1041),
    .B(net1523),
    .Y(_3142_));
 sg13g2_a21oi_1 _7101_ (.A1(net1523),
    .A2(_3141_),
    .Y(_0409_),
    .B1(net1042));
 sg13g2_nand2_1 _7102_ (.Y(_3143_),
    .A(\tt6581_inst.svf_inst.reg_low[14] ),
    .B(_1296_));
 sg13g2_xnor2_1 _7103_ (.Y(_3144_),
    .A(net1132),
    .B(_1296_));
 sg13g2_o21ai_1 _7104_ (.B1(_3139_),
    .Y(_3145_),
    .A1(_3131_),
    .A2(_3134_));
 sg13g2_a21o_2 _7105_ (.A2(_3145_),
    .A1(_3138_),
    .B1(_3144_),
    .X(_3146_));
 sg13g2_nand3_1 _7106_ (.B(_3144_),
    .C(_3145_),
    .A(_3138_),
    .Y(_3147_));
 sg13g2_a21oi_1 _7107_ (.A1(_3146_),
    .A2(_3147_),
    .Y(_3148_),
    .B1(_1000_));
 sg13g2_a21oi_1 _7108_ (.A1(_0932_),
    .A2(_1000_),
    .Y(_0410_),
    .B1(_3148_));
 sg13g2_xnor2_1 _7109_ (.Y(_3149_),
    .A(_0930_),
    .B(_1305_));
 sg13g2_nand2_1 _7110_ (.Y(_3150_),
    .A(_3143_),
    .B(_3146_));
 sg13g2_xnor2_1 _7111_ (.Y(_3151_),
    .A(_3149_),
    .B(_3150_));
 sg13g2_nor2_1 _7112_ (.A(net1103),
    .B(net1517),
    .Y(_3152_));
 sg13g2_a21oi_1 _7113_ (.A1(net1517),
    .A2(_3151_),
    .Y(_0411_),
    .B1(_3152_));
 sg13g2_xnor2_1 _7114_ (.Y(_3153_),
    .A(net1065),
    .B(_1320_));
 sg13g2_a22oi_1 _7115_ (.Y(_3154_),
    .B1(_1305_),
    .B2(\tt6581_inst.svf_inst.reg_low[15] ),
    .A2(_1296_),
    .A1(\tt6581_inst.svf_inst.reg_low[14] ));
 sg13g2_a22oi_1 _7116_ (.Y(_3155_),
    .B1(_3146_),
    .B2(_3154_),
    .A2(_1306_),
    .A1(_0930_));
 sg13g2_a221oi_1 _7117_ (.B2(_3154_),
    .C1(_3153_),
    .B1(_3146_),
    .A1(_0930_),
    .Y(_3156_),
    .A2(_1306_));
 sg13g2_xor2_1 _7118_ (.B(_3155_),
    .A(_3153_),
    .X(_3157_));
 sg13g2_nor2_1 _7119_ (.A(net1065),
    .B(net1516),
    .Y(_3158_));
 sg13g2_a21oi_1 _7120_ (.A1(net1516),
    .A2(_3157_),
    .Y(_0412_),
    .B1(_3158_));
 sg13g2_a21oi_1 _7121_ (.A1(\tt6581_inst.svf_inst.reg_low[16] ),
    .A2(_1320_),
    .Y(_3159_),
    .B1(_3156_));
 sg13g2_nor2_1 _7122_ (.A(_0927_),
    .B(_1331_),
    .Y(_3160_));
 sg13g2_inv_1 _7123_ (.Y(_3161_),
    .A(_3160_));
 sg13g2_and2_1 _7124_ (.A(_0927_),
    .B(_1331_),
    .X(_3162_));
 sg13g2_nor2_1 _7125_ (.A(_3160_),
    .B(_3162_),
    .Y(_3163_));
 sg13g2_xor2_1 _7126_ (.B(_3163_),
    .A(_3159_),
    .X(_3164_));
 sg13g2_nor2_1 _7127_ (.A(net1034),
    .B(net1516),
    .Y(_3165_));
 sg13g2_a21oi_1 _7128_ (.A1(net1516),
    .A2(_3164_),
    .Y(_0413_),
    .B1(_3165_));
 sg13g2_xnor2_1 _7129_ (.Y(_3166_),
    .A(_0925_),
    .B(_1343_));
 sg13g2_o21ai_1 _7130_ (.B1(_3161_),
    .Y(_3167_),
    .A1(_3159_),
    .A2(_3162_));
 sg13g2_and2_1 _7131_ (.A(_3166_),
    .B(_3167_),
    .X(_3168_));
 sg13g2_nand2_1 _7132_ (.Y(_3169_),
    .A(net1061),
    .B(_1000_));
 sg13g2_o21ai_1 _7133_ (.B1(net1516),
    .Y(_3170_),
    .A1(_3166_),
    .A2(_3167_));
 sg13g2_o21ai_1 _7134_ (.B1(_3169_),
    .Y(_0414_),
    .A1(_3168_),
    .A2(_3170_));
 sg13g2_nor2_1 _7135_ (.A(net1101),
    .B(_1356_),
    .Y(_3171_));
 sg13g2_xnor2_1 _7136_ (.Y(_3172_),
    .A(_0924_),
    .B(_1355_));
 sg13g2_a21oi_1 _7137_ (.A1(net1061),
    .A2(_1343_),
    .Y(_3173_),
    .B1(_3168_));
 sg13g2_xnor2_1 _7138_ (.Y(_3174_),
    .A(_3172_),
    .B(_3173_));
 sg13g2_nor2_1 _7139_ (.A(net1101),
    .B(net1516),
    .Y(_3175_));
 sg13g2_a21oi_1 _7140_ (.A1(net1516),
    .A2(_3174_),
    .Y(_0415_),
    .B1(_3175_));
 sg13g2_xnor2_1 _7141_ (.Y(_3176_),
    .A(net1113),
    .B(_1372_));
 sg13g2_a221oi_1 _7142_ (.B2(\tt6581_inst.svf_inst.reg_low[19] ),
    .C1(_3168_),
    .B1(_1356_),
    .A1(\tt6581_inst.svf_inst.reg_low[18] ),
    .Y(_3177_),
    .A2(_1343_));
 sg13g2_nor3_1 _7143_ (.A(_3171_),
    .B(_3176_),
    .C(_3177_),
    .Y(_3178_));
 sg13g2_o21ai_1 _7144_ (.B1(_3176_),
    .Y(_3179_),
    .A1(_3171_),
    .A2(_3177_));
 sg13g2_nand3b_1 _7145_ (.B(_3179_),
    .C(net1517),
    .Y(_3180_),
    .A_N(_3178_));
 sg13g2_o21ai_1 _7146_ (.B1(_3180_),
    .Y(_0416_),
    .A1(_0923_),
    .A2(net1517));
 sg13g2_a21oi_1 _7147_ (.A1(\tt6581_inst.svf_inst.reg_low[20] ),
    .A2(_1372_),
    .Y(_3181_),
    .B1(_3178_));
 sg13g2_nand2b_1 _7148_ (.Y(_3182_),
    .B(_1370_),
    .A_N(\tt6581_inst.mult_inst.accum[35] ));
 sg13g2_and2_1 _7149_ (.A(net1500),
    .B(_3182_),
    .X(_3183_));
 sg13g2_xor2_1 _7150_ (.B(_3183_),
    .A(\tt6581_inst.mult_inst.accum[36] ),
    .X(_3184_));
 sg13g2_inv_1 _7151_ (.Y(_3185_),
    .A(_3184_));
 sg13g2_nor2_1 _7152_ (.A(_0922_),
    .B(_3185_),
    .Y(_3186_));
 sg13g2_nor2_1 _7153_ (.A(net1044),
    .B(_3184_),
    .Y(_3187_));
 sg13g2_nor2_1 _7154_ (.A(_3186_),
    .B(_3187_),
    .Y(_3188_));
 sg13g2_xor2_1 _7155_ (.B(_3188_),
    .A(_3181_),
    .X(_3189_));
 sg13g2_nor2_1 _7156_ (.A(net1044),
    .B(net1517),
    .Y(_3190_));
 sg13g2_a21oi_1 _7157_ (.A1(net1518),
    .A2(_3189_),
    .Y(_0417_),
    .B1(_3190_));
 sg13g2_o21ai_1 _7158_ (.B1(net1500),
    .Y(_3191_),
    .A1(\tt6581_inst.mult_inst.accum[36] ),
    .A2(_3182_));
 sg13g2_inv_1 _7159_ (.Y(_3192_),
    .A(_3191_));
 sg13g2_xnor2_1 _7160_ (.Y(_3193_),
    .A(\tt6581_inst.mult_inst.accum[37] ),
    .B(_3191_));
 sg13g2_nand2_1 _7161_ (.Y(_3194_),
    .A(\tt6581_inst.svf_inst.reg_low[22] ),
    .B(_3193_));
 sg13g2_xnor2_1 _7162_ (.Y(_3195_),
    .A(_0920_),
    .B(_3193_));
 sg13g2_nor2_1 _7163_ (.A(_3181_),
    .B(_3187_),
    .Y(_3196_));
 sg13g2_o21ai_1 _7164_ (.B1(_3195_),
    .Y(_3197_),
    .A1(_3186_),
    .A2(_3196_));
 sg13g2_or3_1 _7165_ (.A(_3186_),
    .B(_3195_),
    .C(_3196_),
    .X(_3198_));
 sg13g2_nand3_1 _7166_ (.B(_3197_),
    .C(_3198_),
    .A(net1518),
    .Y(_3199_));
 sg13g2_o21ai_1 _7167_ (.B1(_3199_),
    .Y(_0418_),
    .A1(_0920_),
    .A2(net1518));
 sg13g2_nor2_1 _7168_ (.A(net1024),
    .B(net1517),
    .Y(_3200_));
 sg13g2_nand2_1 _7169_ (.Y(_3201_),
    .A(_3194_),
    .B(_3197_));
 sg13g2_o21ai_1 _7170_ (.B1(net1504),
    .Y(_3202_),
    .A1(\tt6581_inst.mult_inst.accum[37] ),
    .A2(_3192_));
 sg13g2_xor2_1 _7171_ (.B(_3202_),
    .A(\tt6581_inst.mult_inst.accum[38] ),
    .X(_3203_));
 sg13g2_xnor2_1 _7172_ (.Y(_3204_),
    .A(net1024),
    .B(_3203_));
 sg13g2_xnor2_1 _7173_ (.Y(_3205_),
    .A(_3201_),
    .B(_3204_));
 sg13g2_a21oi_1 _7174_ (.A1(net1517),
    .A2(_3205_),
    .Y(_0419_),
    .B1(_3200_));
 sg13g2_nand2_1 _7175_ (.Y(_3206_),
    .A(net1530),
    .B(net1185));
 sg13g2_xnor2_1 _7176_ (.Y(_0420_),
    .A(net123),
    .B(_3206_));
 sg13g2_nor2_1 _7177_ (.A(net827),
    .B(\tt6581_inst.svf_inst.cur_state[5] ),
    .Y(_3207_));
 sg13g2_o21ai_1 _7178_ (.B1(net123),
    .Y(_3208_),
    .A1(_1108_),
    .A2(_1109_));
 sg13g2_o21ai_1 _7179_ (.B1(net1706),
    .Y(_3209_),
    .A1(_1122_),
    .A2(_1123_));
 sg13g2_nor3_1 _7180_ (.A(\tt6581_inst.svf_inst.reg_band[1] ),
    .B(_1122_),
    .C(_1123_),
    .Y(_3210_));
 sg13g2_xnor2_1 _7181_ (.Y(_3211_),
    .A(net827),
    .B(_1124_));
 sg13g2_xnor2_1 _7182_ (.Y(_3212_),
    .A(_3208_),
    .B(_3211_));
 sg13g2_a21oi_1 _7183_ (.A1(net1531),
    .A2(_3212_),
    .Y(_0421_),
    .B1(net828));
 sg13g2_and2_1 _7184_ (.A(net337),
    .B(net1183),
    .X(_3213_));
 sg13g2_or2_1 _7185_ (.X(_3214_),
    .B(net1183),
    .A(\tt6581_inst.svf_inst.reg_band[2] ));
 sg13g2_nand2b_1 _7186_ (.Y(_3215_),
    .B(_3214_),
    .A_N(_3213_));
 sg13g2_o21ai_1 _7187_ (.B1(_3209_),
    .Y(_3216_),
    .A1(_3208_),
    .A2(_3210_));
 sg13g2_nand2b_1 _7188_ (.Y(_3217_),
    .B(_3216_),
    .A_N(_3215_));
 sg13g2_nand2b_1 _7189_ (.Y(_3218_),
    .B(_3215_),
    .A_N(_3216_));
 sg13g2_a21oi_1 _7190_ (.A1(_3217_),
    .A2(_3218_),
    .Y(_3219_),
    .B1(net1431));
 sg13g2_a21oi_1 _7191_ (.A1(_0949_),
    .A2(net1431),
    .Y(_0422_),
    .B1(_3219_));
 sg13g2_nand2_1 _7192_ (.Y(_3220_),
    .A(\tt6581_inst.svf_inst.reg_band[3] ),
    .B(net1173));
 sg13g2_xnor2_1 _7193_ (.Y(_3221_),
    .A(net560),
    .B(net1173));
 sg13g2_a21oi_1 _7194_ (.A1(_3214_),
    .A2(_3216_),
    .Y(_3222_),
    .B1(_3213_));
 sg13g2_xnor2_1 _7195_ (.Y(_3223_),
    .A(_3221_),
    .B(_3222_));
 sg13g2_nor2_1 _7196_ (.A(net560),
    .B(net1530),
    .Y(_3224_));
 sg13g2_a21oi_1 _7197_ (.A1(net1530),
    .A2(_3223_),
    .Y(_0423_),
    .B1(net561));
 sg13g2_and2_1 _7198_ (.A(net371),
    .B(net1167),
    .X(_3225_));
 sg13g2_xor2_1 _7199_ (.B(net1167),
    .A(net371),
    .X(_3226_));
 sg13g2_o21ai_1 _7200_ (.B1(_3220_),
    .Y(_3227_),
    .A1(_3221_),
    .A2(_3222_));
 sg13g2_and2_1 _7201_ (.A(_3226_),
    .B(_3227_),
    .X(_3228_));
 sg13g2_nand2_1 _7202_ (.Y(_3229_),
    .A(net371),
    .B(net1431));
 sg13g2_o21ai_1 _7203_ (.B1(net1530),
    .Y(_3230_),
    .A1(_3226_),
    .A2(_3227_));
 sg13g2_o21ai_1 _7204_ (.B1(_3229_),
    .Y(_0424_),
    .A1(_3228_),
    .A2(_3230_));
 sg13g2_nor2_1 _7205_ (.A(net854),
    .B(net1530),
    .Y(_3231_));
 sg13g2_nor2_1 _7206_ (.A(_3225_),
    .B(_3228_),
    .Y(_3232_));
 sg13g2_nor2_1 _7207_ (.A(\tt6581_inst.svf_inst.reg_band[5] ),
    .B(net1164),
    .Y(_3233_));
 sg13g2_xnor2_1 _7208_ (.Y(_3234_),
    .A(net854),
    .B(net1164));
 sg13g2_xnor2_1 _7209_ (.Y(_3235_),
    .A(_3232_),
    .B(_3234_));
 sg13g2_a21oi_1 _7210_ (.A1(net1530),
    .A2(_3235_),
    .Y(_0425_),
    .B1(net855));
 sg13g2_nand2_1 _7211_ (.Y(_3236_),
    .A(\tt6581_inst.svf_inst.reg_band[6] ),
    .B(_1187_));
 sg13g2_xnor2_1 _7212_ (.Y(_3237_),
    .A(\tt6581_inst.svf_inst.reg_band[6] ),
    .B(_1187_));
 sg13g2_a221oi_1 _7213_ (.B2(_3227_),
    .C1(_3225_),
    .B1(_3226_),
    .A1(\tt6581_inst.svf_inst.reg_band[5] ),
    .Y(_3238_),
    .A2(net1165));
 sg13g2_or3_1 _7214_ (.A(_3233_),
    .B(_3237_),
    .C(_3238_),
    .X(_3239_));
 sg13g2_o21ai_1 _7215_ (.B1(_3237_),
    .Y(_3240_),
    .A1(_3233_),
    .A2(_3238_));
 sg13g2_and2_1 _7216_ (.A(net1530),
    .B(_3240_),
    .X(_3241_));
 sg13g2_a22oi_1 _7217_ (.Y(_3242_),
    .B1(_3239_),
    .B2(_3241_),
    .A2(net1431),
    .A1(net1001));
 sg13g2_inv_1 _7218_ (.Y(_0426_),
    .A(_3242_));
 sg13g2_nand2_1 _7219_ (.Y(_3243_),
    .A(net430),
    .B(_1200_));
 sg13g2_xnor2_1 _7220_ (.Y(_3244_),
    .A(net430),
    .B(_1200_));
 sg13g2_a21o_1 _7221_ (.A2(_3239_),
    .A1(_3236_),
    .B1(_3244_),
    .X(_3245_));
 sg13g2_nand3_1 _7222_ (.B(_3239_),
    .C(_3244_),
    .A(_3236_),
    .Y(_3246_));
 sg13g2_a21oi_1 _7223_ (.A1(_3245_),
    .A2(_3246_),
    .Y(_3247_),
    .B1(net1431));
 sg13g2_a21oi_1 _7224_ (.A1(_0948_),
    .A2(net1431),
    .Y(_0427_),
    .B1(_3247_));
 sg13g2_xnor2_1 _7225_ (.Y(_3248_),
    .A(net880),
    .B(_1211_));
 sg13g2_a21o_2 _7226_ (.A2(_3245_),
    .A1(_3243_),
    .B1(_3248_),
    .X(_3249_));
 sg13g2_nand3_1 _7227_ (.B(_3245_),
    .C(_3248_),
    .A(_3243_),
    .Y(_3250_));
 sg13g2_a21oi_1 _7228_ (.A1(_3249_),
    .A2(_3250_),
    .Y(_3251_),
    .B1(_1001_));
 sg13g2_a21oi_1 _7229_ (.A1(_0947_),
    .A2(_1001_),
    .Y(_0428_),
    .B1(_3251_));
 sg13g2_xnor2_1 _7230_ (.Y(_3252_),
    .A(net818),
    .B(_1224_));
 sg13g2_o21ai_1 _7231_ (.B1(_3249_),
    .Y(_3253_),
    .A1(_0947_),
    .A2(_1212_));
 sg13g2_xnor2_1 _7232_ (.Y(_3254_),
    .A(_3252_),
    .B(_3253_));
 sg13g2_nor2_1 _7233_ (.A(net818),
    .B(net1531),
    .Y(_3255_));
 sg13g2_a21oi_1 _7234_ (.A1(net1531),
    .A2(_3254_),
    .Y(_0429_),
    .B1(net819));
 sg13g2_xnor2_1 _7235_ (.Y(_3256_),
    .A(net912),
    .B(_1239_));
 sg13g2_a22oi_1 _7236_ (.Y(_3257_),
    .B1(_1225_),
    .B2(\tt6581_inst.svf_inst.reg_band[9] ),
    .A2(_1211_),
    .A1(\tt6581_inst.svf_inst.reg_band[8] ));
 sg13g2_a22oi_1 _7237_ (.Y(_3258_),
    .B1(_3249_),
    .B2(_3257_),
    .A2(_1224_),
    .A1(_0946_));
 sg13g2_a221oi_1 _7238_ (.B2(_3257_),
    .C1(_3256_),
    .B1(_3249_),
    .A1(_0946_),
    .Y(_3259_),
    .A2(_1224_));
 sg13g2_xor2_1 _7239_ (.B(_3258_),
    .A(_3256_),
    .X(_3260_));
 sg13g2_nor2_1 _7240_ (.A(net912),
    .B(net1531),
    .Y(_3261_));
 sg13g2_a21oi_1 _7241_ (.A1(net1531),
    .A2(_3260_),
    .Y(_0430_),
    .B1(net913));
 sg13g2_nor2_1 _7242_ (.A(net727),
    .B(net1531),
    .Y(_3262_));
 sg13g2_nand2b_1 _7243_ (.Y(_3263_),
    .B(_1254_),
    .A_N(\tt6581_inst.svf_inst.reg_band[11] ));
 sg13g2_xnor2_1 _7244_ (.Y(_3264_),
    .A(net727),
    .B(_1253_));
 sg13g2_a21oi_1 _7245_ (.A1(\tt6581_inst.svf_inst.reg_band[10] ),
    .A2(_1239_),
    .Y(_3265_),
    .B1(_3259_));
 sg13g2_xnor2_1 _7246_ (.Y(_3266_),
    .A(_3264_),
    .B(_3265_));
 sg13g2_a21oi_1 _7247_ (.A1(net1531),
    .A2(_3266_),
    .Y(_0431_),
    .B1(net728));
 sg13g2_nand2_1 _7248_ (.Y(_3267_),
    .A(\tt6581_inst.svf_inst.reg_band[12] ),
    .B(_1267_));
 sg13g2_xnor2_1 _7249_ (.Y(_3268_),
    .A(net642),
    .B(_1267_));
 sg13g2_a22oi_1 _7250_ (.Y(_3269_),
    .B1(_1253_),
    .B2(\tt6581_inst.svf_inst.reg_band[11] ),
    .A2(_1239_),
    .A1(\tt6581_inst.svf_inst.reg_band[10] ));
 sg13g2_inv_1 _7251_ (.Y(_3270_),
    .A(_3269_));
 sg13g2_o21ai_1 _7252_ (.B1(_3263_),
    .Y(_3271_),
    .A1(_3259_),
    .A2(_3270_));
 sg13g2_xnor2_1 _7253_ (.Y(_3272_),
    .A(_3268_),
    .B(_3271_));
 sg13g2_nor2_1 _7254_ (.A(net642),
    .B(net1529),
    .Y(_3273_));
 sg13g2_a21oi_1 _7255_ (.A1(net1529),
    .A2(_3272_),
    .Y(_0432_),
    .B1(net643));
 sg13g2_o21ai_1 _7256_ (.B1(_3267_),
    .Y(_3274_),
    .A1(_3268_),
    .A2(_3271_));
 sg13g2_nand2_1 _7257_ (.Y(_3275_),
    .A(net937),
    .B(_1280_));
 sg13g2_inv_1 _7258_ (.Y(_3276_),
    .A(_3275_));
 sg13g2_or2_1 _7259_ (.X(_3277_),
    .B(_1280_),
    .A(\tt6581_inst.svf_inst.reg_band[13] ));
 sg13g2_nand2_1 _7260_ (.Y(_3278_),
    .A(_3275_),
    .B(_3277_));
 sg13g2_xnor2_1 _7261_ (.Y(_3279_),
    .A(_3274_),
    .B(_3278_));
 sg13g2_mux2_1 _7262_ (.A0(net937),
    .A1(_3279_),
    .S(net1529),
    .X(_0433_));
 sg13g2_and2_1 _7263_ (.A(net862),
    .B(_1296_),
    .X(_3280_));
 sg13g2_or2_1 _7264_ (.X(_3281_),
    .B(_1296_),
    .A(\tt6581_inst.svf_inst.reg_band[14] ));
 sg13g2_nand2b_1 _7265_ (.Y(_3282_),
    .B(_3281_),
    .A_N(_3280_));
 sg13g2_a21o_1 _7266_ (.A2(_3277_),
    .A1(_3274_),
    .B1(_3276_),
    .X(_3283_));
 sg13g2_xnor2_1 _7267_ (.Y(_3284_),
    .A(_3282_),
    .B(_3283_));
 sg13g2_mux2_1 _7268_ (.A0(net862),
    .A1(_3284_),
    .S(net1529),
    .X(_0434_));
 sg13g2_a21oi_1 _7269_ (.A1(_3281_),
    .A2(_3283_),
    .Y(_3285_),
    .B1(_3280_));
 sg13g2_nand2_1 _7270_ (.Y(_3286_),
    .A(\tt6581_inst.svf_inst.reg_band[15] ),
    .B(_1305_));
 sg13g2_nor2_1 _7271_ (.A(\tt6581_inst.svf_inst.reg_band[15] ),
    .B(_1305_),
    .Y(_3287_));
 sg13g2_xnor2_1 _7272_ (.Y(_3288_),
    .A(net876),
    .B(_1305_));
 sg13g2_xnor2_1 _7273_ (.Y(_3289_),
    .A(_3285_),
    .B(_3288_));
 sg13g2_nor2_1 _7274_ (.A(net876),
    .B(net1527),
    .Y(_3290_));
 sg13g2_a21oi_1 _7275_ (.A1(net1528),
    .A2(_3289_),
    .Y(_0435_),
    .B1(_3290_));
 sg13g2_xnor2_1 _7276_ (.Y(_3291_),
    .A(net789),
    .B(_1320_));
 sg13g2_o21ai_1 _7277_ (.B1(_3286_),
    .Y(_3292_),
    .A1(_3285_),
    .A2(_3287_));
 sg13g2_nor2b_1 _7278_ (.A(_3291_),
    .B_N(_3292_),
    .Y(_3293_));
 sg13g2_xor2_1 _7279_ (.B(_3292_),
    .A(_3291_),
    .X(_3294_));
 sg13g2_nor2_1 _7280_ (.A(net789),
    .B(net1527),
    .Y(_3295_));
 sg13g2_a21oi_1 _7281_ (.A1(net1527),
    .A2(_3294_),
    .Y(_0436_),
    .B1(_3295_));
 sg13g2_a21o_1 _7282_ (.A2(_1320_),
    .A1(\tt6581_inst.svf_inst.reg_band[16] ),
    .B1(_3293_),
    .X(_3296_));
 sg13g2_nand2b_1 _7283_ (.Y(_3297_),
    .B(net536),
    .A_N(_1331_));
 sg13g2_nand2b_1 _7284_ (.Y(_3298_),
    .B(_1331_),
    .A_N(\tt6581_inst.svf_inst.reg_band[17] ));
 sg13g2_nand2_1 _7285_ (.Y(_3299_),
    .A(_3297_),
    .B(_3298_));
 sg13g2_xor2_1 _7286_ (.B(_3299_),
    .A(_3296_),
    .X(_3300_));
 sg13g2_nor2_1 _7287_ (.A(net536),
    .B(net1527),
    .Y(_3301_));
 sg13g2_a21oi_1 _7288_ (.A1(net1527),
    .A2(_3300_),
    .Y(_0437_),
    .B1(_3301_));
 sg13g2_xnor2_1 _7289_ (.Y(_3302_),
    .A(net1021),
    .B(_1343_));
 sg13g2_nand2_1 _7290_ (.Y(_3303_),
    .A(_3296_),
    .B(_3298_));
 sg13g2_a21oi_1 _7291_ (.A1(_3297_),
    .A2(_3303_),
    .Y(_3304_),
    .B1(_3302_));
 sg13g2_and3_1 _7292_ (.X(_3305_),
    .A(_3297_),
    .B(_3302_),
    .C(_3303_));
 sg13g2_nor3_1 _7293_ (.A(net1431),
    .B(_3304_),
    .C(_3305_),
    .Y(_3306_));
 sg13g2_a21o_1 _7294_ (.A2(net1431),
    .A1(net1021),
    .B1(_3306_),
    .X(_0438_));
 sg13g2_a21o_1 _7295_ (.A2(_1343_),
    .A1(net1021),
    .B1(_3304_),
    .X(_3307_));
 sg13g2_nand2_1 _7296_ (.Y(_3308_),
    .A(\tt6581_inst.svf_inst.reg_band[19] ),
    .B(_1356_));
 sg13g2_xnor2_1 _7297_ (.Y(_3309_),
    .A(net1059),
    .B(_1355_));
 sg13g2_xnor2_1 _7298_ (.Y(_3310_),
    .A(_3307_),
    .B(_3309_));
 sg13g2_nor2_1 _7299_ (.A(net1059),
    .B(net1527),
    .Y(_3311_));
 sg13g2_a21oi_1 _7300_ (.A1(net1527),
    .A2(_3310_),
    .Y(_0439_),
    .B1(_3311_));
 sg13g2_nand2_1 _7301_ (.Y(_3312_),
    .A(\tt6581_inst.svf_inst.reg_band[20] ),
    .B(_1372_));
 sg13g2_xnor2_1 _7302_ (.Y(_3313_),
    .A(net1049),
    .B(_1372_));
 sg13g2_o21ai_1 _7303_ (.B1(_3307_),
    .Y(_3314_),
    .A1(\tt6581_inst.svf_inst.reg_band[19] ),
    .A2(_1356_));
 sg13g2_a21o_2 _7304_ (.A2(_3314_),
    .A1(_3308_),
    .B1(_3313_),
    .X(_3315_));
 sg13g2_nand3_1 _7305_ (.B(_3313_),
    .C(_3314_),
    .A(_3308_),
    .Y(_3316_));
 sg13g2_nand3_1 _7306_ (.B(_3315_),
    .C(_3316_),
    .A(net1528),
    .Y(_3317_));
 sg13g2_o21ai_1 _7307_ (.B1(_3317_),
    .Y(_0440_),
    .A1(_0945_),
    .A2(net1528));
 sg13g2_xnor2_1 _7308_ (.Y(_3318_),
    .A(_0944_),
    .B(_3184_));
 sg13g2_nand2_1 _7309_ (.Y(_3319_),
    .A(_3312_),
    .B(_3315_));
 sg13g2_xnor2_1 _7310_ (.Y(_3320_),
    .A(_3318_),
    .B(_3319_));
 sg13g2_nor2_1 _7311_ (.A(net920),
    .B(net1528),
    .Y(_3321_));
 sg13g2_a21oi_1 _7312_ (.A1(net1528),
    .A2(_3320_),
    .Y(_0441_),
    .B1(net921));
 sg13g2_a22oi_1 _7313_ (.Y(_3322_),
    .B1(_3184_),
    .B2(\tt6581_inst.svf_inst.reg_band[21] ),
    .A2(_1372_),
    .A1(\tt6581_inst.svf_inst.reg_band[20] ));
 sg13g2_a22oi_1 _7314_ (.Y(_3323_),
    .B1(_3315_),
    .B2(_3322_),
    .A2(_3185_),
    .A1(_0944_));
 sg13g2_xnor2_1 _7315_ (.Y(_3324_),
    .A(net1089),
    .B(_3193_));
 sg13g2_a221oi_1 _7316_ (.B2(_3322_),
    .C1(_3324_),
    .B1(_3315_),
    .A1(_0944_),
    .Y(_3325_),
    .A2(_3185_));
 sg13g2_xnor2_1 _7317_ (.Y(_3326_),
    .A(_3323_),
    .B(_3324_));
 sg13g2_mux2_1 _7318_ (.A0(net1089),
    .A1(_3326_),
    .S(net1528),
    .X(_0442_));
 sg13g2_a21oi_1 _7319_ (.A1(\tt6581_inst.svf_inst.reg_band[22] ),
    .A2(_3193_),
    .Y(_3327_),
    .B1(_3325_));
 sg13g2_o21ai_1 _7320_ (.B1(net1528),
    .Y(_3328_),
    .A1(_3203_),
    .A2(_3327_));
 sg13g2_a21oi_1 _7321_ (.A1(_3203_),
    .A2(_3327_),
    .Y(_3329_),
    .B1(_3328_));
 sg13g2_xor2_1 _7322_ (.B(_3329_),
    .A(net91),
    .X(_0443_));
 sg13g2_nor2_2 _7323_ (.A(_1005_),
    .B(net1392),
    .Y(_3330_));
 sg13g2_nor2_1 _7324_ (.A(net283),
    .B(net1339),
    .Y(_3331_));
 sg13g2_a21oi_1 _7325_ (.A1(_2654_),
    .A2(net1339),
    .Y(_0444_),
    .B1(_3331_));
 sg13g2_nor2_1 _7326_ (.A(net208),
    .B(net1339),
    .Y(_3332_));
 sg13g2_a21oi_1 _7327_ (.A1(_2658_),
    .A2(net1339),
    .Y(_0445_),
    .B1(_3332_));
 sg13g2_nor2b_2 _7328_ (.A(_1005_),
    .B_N(net1382),
    .Y(_3333_));
 sg13g2_nor2_1 _7329_ (.A(net163),
    .B(net1334),
    .Y(_3334_));
 sg13g2_nor2_1 _7330_ (.A(_2654_),
    .B(_2658_),
    .Y(_3335_));
 sg13g2_nand2b_2 _7331_ (.Y(_3336_),
    .B(_2648_),
    .A_N(_2658_));
 sg13g2_nand2_1 _7332_ (.Y(_3337_),
    .A(\tt6581_inst.ad_pack[15] ),
    .B(net1402));
 sg13g2_a22oi_1 _7333_ (.Y(_3338_),
    .B1(net1380),
    .B2(\tt6581_inst.ad_pack[7] ),
    .A2(net1422),
    .A1(\tt6581_inst.ad_pack[23] ));
 sg13g2_and2_1 _7334_ (.A(_3337_),
    .B(_3338_),
    .X(_3339_));
 sg13g2_nand2_2 _7335_ (.Y(_3340_),
    .A(_3337_),
    .B(_3338_));
 sg13g2_a22oi_1 _7336_ (.Y(_3341_),
    .B1(net1380),
    .B2(\tt6581_inst.ad_pack[4] ),
    .A2(net1401),
    .A1(\tt6581_inst.ad_pack[12] ));
 sg13g2_o21ai_1 _7337_ (.B1(_3341_),
    .Y(_3342_),
    .A1(_0989_),
    .A2(net1416));
 sg13g2_nand2_1 _7338_ (.Y(_3343_),
    .A(\tt6581_inst.ad_pack[14] ),
    .B(net1403));
 sg13g2_a22oi_1 _7339_ (.Y(_3344_),
    .B1(net1380),
    .B2(\tt6581_inst.ad_pack[6] ),
    .A2(net1421),
    .A1(\tt6581_inst.ad_pack[22] ));
 sg13g2_and2_1 _7340_ (.A(_3343_),
    .B(_3344_),
    .X(_3345_));
 sg13g2_nand2_2 _7341_ (.Y(_3346_),
    .A(_3343_),
    .B(_3344_));
 sg13g2_nand2_1 _7342_ (.Y(_3347_),
    .A(\tt6581_inst.ad_pack[5] ),
    .B(net1380));
 sg13g2_a22oi_1 _7343_ (.Y(_3348_),
    .B1(net1400),
    .B2(\tt6581_inst.ad_pack[13] ),
    .A2(net1422),
    .A1(\tt6581_inst.ad_pack[21] ));
 sg13g2_and2_1 _7344_ (.A(_3347_),
    .B(_3348_),
    .X(_3349_));
 sg13g2_nand2_2 _7345_ (.Y(_3350_),
    .A(_3347_),
    .B(_3348_));
 sg13g2_nand2_1 _7346_ (.Y(_3351_),
    .A(_3345_),
    .B(net1251));
 sg13g2_nor2_1 _7347_ (.A(net1158),
    .B(_3351_),
    .Y(_3352_));
 sg13g2_nor3_1 _7348_ (.A(net1158),
    .B(net1252),
    .C(_3351_),
    .Y(_3353_));
 sg13g2_nor2_1 _7349_ (.A(net1252),
    .B(_3346_),
    .Y(_3354_));
 sg13g2_a221oi_1 _7350_ (.B2(_2518_),
    .C1(_2515_),
    .B1(_2517_),
    .A1(_0040_),
    .Y(_3355_),
    .A2(net1402));
 sg13g2_nor2b_1 _7351_ (.A(\tt6581_inst.ad_pack[3] ),
    .B_N(net1247),
    .Y(_3356_));
 sg13g2_o21ai_1 _7352_ (.B1(net1380),
    .Y(_3357_),
    .A1(\tt6581_inst.controller_inst.sr_i[3] ),
    .A2(net1247));
 sg13g2_mux2_1 _7353_ (.A0(\tt6581_inst.controller_inst.sr_i[3] ),
    .A1(\tt6581_inst.ad_pack[3] ),
    .S(net1247),
    .X(_3358_));
 sg13g2_a22oi_1 _7354_ (.Y(_3359_),
    .B1(net1400),
    .B2(\tt6581_inst.ad_pack[11] ),
    .A2(net1422),
    .A1(\tt6581_inst.ad_pack[19] ));
 sg13g2_inv_1 _7355_ (.Y(_3360_),
    .A(_3359_));
 sg13g2_a22oi_1 _7356_ (.Y(_3361_),
    .B1(net1400),
    .B2(\tt6581_inst.controller_inst.sr_i[11] ),
    .A2(net1421),
    .A1(\tt6581_inst.controller_inst.sr_i[19] ));
 sg13g2_nor2_1 _7357_ (.A(net1247),
    .B(_3361_),
    .Y(_3362_));
 sg13g2_mux2_1 _7358_ (.A0(_3361_),
    .A1(_3359_),
    .S(net1247),
    .X(_3363_));
 sg13g2_a221oi_1 _7359_ (.B2(net1247),
    .C1(_3362_),
    .B1(_3360_),
    .A1(net1380),
    .Y(_3364_),
    .A2(_3358_));
 sg13g2_o21ai_1 _7360_ (.B1(_3363_),
    .Y(_3365_),
    .A1(_3356_),
    .A2(_3357_));
 sg13g2_nor2b_1 _7361_ (.A(\tt6581_inst.ad_pack[2] ),
    .B_N(net1248),
    .Y(_3366_));
 sg13g2_o21ai_1 _7362_ (.B1(net1380),
    .Y(_3367_),
    .A1(\tt6581_inst.controller_inst.sr_i[2] ),
    .A2(net1249));
 sg13g2_mux2_1 _7363_ (.A0(\tt6581_inst.controller_inst.sr_i[2] ),
    .A1(\tt6581_inst.ad_pack[2] ),
    .S(net1247),
    .X(_3368_));
 sg13g2_a22oi_1 _7364_ (.Y(_3369_),
    .B1(net1401),
    .B2(\tt6581_inst.ad_pack[10] ),
    .A2(net1422),
    .A1(\tt6581_inst.ad_pack[18] ));
 sg13g2_inv_1 _7365_ (.Y(_3370_),
    .A(_3369_));
 sg13g2_a22oi_1 _7366_ (.Y(_3371_),
    .B1(net1400),
    .B2(\tt6581_inst.controller_inst.sr_i[10] ),
    .A2(net1421),
    .A1(\tt6581_inst.controller_inst.sr_i[18] ));
 sg13g2_nor2_1 _7367_ (.A(net1248),
    .B(_3371_),
    .Y(_3372_));
 sg13g2_mux2_1 _7368_ (.A0(_3371_),
    .A1(_3369_),
    .S(net1247),
    .X(_3373_));
 sg13g2_a221oi_1 _7369_ (.B2(net1249),
    .C1(_3372_),
    .B1(_3370_),
    .A1(net1380),
    .Y(_3374_),
    .A2(_3368_));
 sg13g2_o21ai_1 _7370_ (.B1(_3373_),
    .Y(_3375_),
    .A1(_3366_),
    .A2(_3367_));
 sg13g2_nor2b_1 _7371_ (.A(\tt6581_inst.ad_pack[1] ),
    .B_N(net1250),
    .Y(_3376_));
 sg13g2_o21ai_1 _7372_ (.B1(net1381),
    .Y(_3377_),
    .A1(\tt6581_inst.controller_inst.sr_i[1] ),
    .A2(net1249));
 sg13g2_mux2_1 _7373_ (.A0(\tt6581_inst.controller_inst.sr_i[1] ),
    .A1(\tt6581_inst.ad_pack[1] ),
    .S(net1250),
    .X(_3378_));
 sg13g2_a22oi_1 _7374_ (.Y(_3379_),
    .B1(net1401),
    .B2(\tt6581_inst.ad_pack[9] ),
    .A2(net1422),
    .A1(\tt6581_inst.ad_pack[17] ));
 sg13g2_inv_1 _7375_ (.Y(_3380_),
    .A(_3379_));
 sg13g2_a22oi_1 _7376_ (.Y(_3381_),
    .B1(net1400),
    .B2(\tt6581_inst.controller_inst.sr_i[9] ),
    .A2(net1421),
    .A1(\tt6581_inst.controller_inst.sr_i[17] ));
 sg13g2_nor2_1 _7377_ (.A(net1248),
    .B(_3381_),
    .Y(_3382_));
 sg13g2_mux2_1 _7378_ (.A0(_3381_),
    .A1(_3379_),
    .S(net1248),
    .X(_3383_));
 sg13g2_a221oi_1 _7379_ (.B2(net1249),
    .C1(_3382_),
    .B1(_3380_),
    .A1(net1381),
    .Y(_3384_),
    .A2(_3378_));
 sg13g2_o21ai_1 _7380_ (.B1(_3383_),
    .Y(_3385_),
    .A1(_3376_),
    .A2(_3377_));
 sg13g2_nor2b_1 _7381_ (.A(\tt6581_inst.ad_pack[0] ),
    .B_N(net1250),
    .Y(_3386_));
 sg13g2_o21ai_1 _7382_ (.B1(net1381),
    .Y(_3387_),
    .A1(\tt6581_inst.controller_inst.sr_i[0] ),
    .A2(net1250));
 sg13g2_mux2_1 _7383_ (.A0(\tt6581_inst.controller_inst.sr_i[0] ),
    .A1(\tt6581_inst.ad_pack[0] ),
    .S(net1250),
    .X(_3388_));
 sg13g2_a22oi_1 _7384_ (.Y(_3389_),
    .B1(net1400),
    .B2(\tt6581_inst.ad_pack[8] ),
    .A2(net1421),
    .A1(\tt6581_inst.ad_pack[16] ));
 sg13g2_inv_1 _7385_ (.Y(_3390_),
    .A(_3389_));
 sg13g2_a22oi_1 _7386_ (.Y(_3391_),
    .B1(net1400),
    .B2(\tt6581_inst.controller_inst.sr_i[8] ),
    .A2(net1421),
    .A1(\tt6581_inst.controller_inst.sr_i[16] ));
 sg13g2_nor2_1 _7387_ (.A(net1250),
    .B(_3391_),
    .Y(_3392_));
 sg13g2_mux2_1 _7388_ (.A0(_3391_),
    .A1(_3389_),
    .S(net1250),
    .X(_3393_));
 sg13g2_a221oi_1 _7389_ (.B2(net1250),
    .C1(_3392_),
    .B1(_3390_),
    .A1(net1381),
    .Y(_3394_),
    .A2(_3388_));
 sg13g2_o21ai_1 _7390_ (.B1(_3393_),
    .Y(_3395_),
    .A1(_3386_),
    .A2(_3387_));
 sg13g2_nand2_1 _7391_ (.Y(_3396_),
    .A(net1187),
    .B(_3384_));
 sg13g2_nand4_1 _7392_ (.B(_3374_),
    .C(_3384_),
    .A(net1187),
    .Y(_3397_),
    .D(_3394_));
 sg13g2_nor3_1 _7393_ (.A(net1263),
    .B(net1155),
    .C(_3397_),
    .Y(_3398_));
 sg13g2_a21o_2 _7394_ (.A2(_3353_),
    .A1(_3339_),
    .B1(_3398_),
    .X(_3399_));
 sg13g2_and2_1 _7395_ (.A(_2530_),
    .B(_3399_),
    .X(_3400_));
 sg13g2_xor2_1 _7396_ (.B(_3399_),
    .A(_2530_),
    .X(_3401_));
 sg13g2_and2_1 _7397_ (.A(net1263),
    .B(_2548_),
    .X(_3402_));
 sg13g2_nand2_2 _7398_ (.Y(_3403_),
    .A(net1264),
    .B(_2548_));
 sg13g2_o21ai_1 _7399_ (.B1(net1264),
    .Y(_3404_),
    .A1(_2547_),
    .A2(net1261));
 sg13g2_nor2_1 _7400_ (.A(_3397_),
    .B(net1210),
    .Y(_3405_));
 sg13g2_nand3_1 _7401_ (.B(net1212),
    .C(_3405_),
    .A(net1159),
    .Y(_3406_));
 sg13g2_nor2b_1 _7402_ (.A(_3406_),
    .B_N(net1265),
    .Y(_3407_));
 sg13g2_a21o_1 _7403_ (.A2(_3407_),
    .A1(_3401_),
    .B1(_3400_),
    .X(_3408_));
 sg13g2_nand2_1 _7404_ (.Y(_3409_),
    .A(_2551_),
    .B(_3408_));
 sg13g2_nand3_1 _7405_ (.B(_2551_),
    .C(_3408_),
    .A(_2543_),
    .Y(_3410_));
 sg13g2_nand2b_2 _7406_ (.Y(_3411_),
    .B(_2522_),
    .A_N(_3410_));
 sg13g2_nand2b_1 _7407_ (.Y(_3412_),
    .B(_3410_),
    .A_N(_2522_));
 sg13g2_a21o_1 _7408_ (.A2(_3412_),
    .A1(_3411_),
    .B1(net1259),
    .X(_3413_));
 sg13g2_xnor2_1 _7409_ (.Y(_3414_),
    .A(_2543_),
    .B(_3409_));
 sg13g2_nand2_1 _7410_ (.Y(_3415_),
    .A(net1258),
    .B(_3414_));
 sg13g2_xor2_1 _7411_ (.B(_3408_),
    .A(_2551_),
    .X(_3416_));
 sg13g2_nand2b_1 _7412_ (.Y(_3417_),
    .B(_2575_),
    .A_N(_3416_));
 sg13g2_o21ai_1 _7413_ (.B1(_3417_),
    .Y(_3418_),
    .A1(net1258),
    .A2(_3414_));
 sg13g2_xnor2_1 _7414_ (.Y(_3419_),
    .A(_3401_),
    .B(_3407_));
 sg13g2_xor2_1 _7415_ (.B(_3406_),
    .A(net1265),
    .X(_3420_));
 sg13g2_a22oi_1 _7416_ (.Y(_3421_),
    .B1(_3420_),
    .B2(_2526_),
    .A2(_3419_),
    .A1(_2533_));
 sg13g2_and2_1 _7417_ (.A(_3342_),
    .B(_3345_),
    .X(_3422_));
 sg13g2_xnor2_1 _7418_ (.Y(_3423_),
    .A(net1252),
    .B(_3346_));
 sg13g2_nor2_1 _7419_ (.A(_3345_),
    .B(net1251),
    .Y(_3424_));
 sg13g2_nor3_1 _7420_ (.A(net1253),
    .B(_3423_),
    .C(_3424_),
    .Y(_3425_));
 sg13g2_nor2_1 _7421_ (.A(_3375_),
    .B(_3394_),
    .Y(_3426_));
 sg13g2_nor2b_2 _7422_ (.A(_3396_),
    .B_N(_3426_),
    .Y(_3427_));
 sg13g2_nor2_1 _7423_ (.A(net1262),
    .B(net1212),
    .Y(_3428_));
 sg13g2_nand2_1 _7424_ (.Y(_3429_),
    .A(_3385_),
    .B(_3426_));
 sg13g2_nand4_1 _7425_ (.B(_3374_),
    .C(_3385_),
    .A(net1187),
    .Y(_3430_),
    .D(_3395_));
 sg13g2_nor2_1 _7426_ (.A(net1186),
    .B(_3395_),
    .Y(_3431_));
 sg13g2_nand3_1 _7427_ (.B(_3374_),
    .C(_3431_),
    .A(net1187),
    .Y(_3432_));
 sg13g2_nor2b_1 _7428_ (.A(net1210),
    .B_N(_3432_),
    .Y(_3433_));
 sg13g2_a21oi_1 _7429_ (.A1(net1210),
    .A2(_3430_),
    .Y(_3434_),
    .B1(_3433_));
 sg13g2_a22oi_1 _7430_ (.Y(_3435_),
    .B1(_3434_),
    .B2(net1212),
    .A2(_3428_),
    .A1(_3427_));
 sg13g2_nand2_1 _7431_ (.Y(_3436_),
    .A(net1158),
    .B(_3435_));
 sg13g2_o21ai_1 _7432_ (.B1(_3436_),
    .Y(_3437_),
    .A1(net1158),
    .A2(_3425_));
 sg13g2_inv_1 _7433_ (.Y(_3438_),
    .A(_3437_));
 sg13g2_nand2_1 _7434_ (.Y(_3439_),
    .A(_2624_),
    .B(_3437_));
 sg13g2_nand2_1 _7435_ (.Y(_3440_),
    .A(_2623_),
    .B(_3438_));
 sg13g2_nand2_1 _7436_ (.Y(_3441_),
    .A(_3439_),
    .B(_3440_));
 sg13g2_nand2_1 _7437_ (.Y(_3442_),
    .A(net1210),
    .B(_3432_));
 sg13g2_o21ai_1 _7438_ (.B1(_3442_),
    .Y(_3443_),
    .A1(net1210),
    .A2(_3427_));
 sg13g2_nor2_1 _7439_ (.A(net1209),
    .B(_3430_),
    .Y(_3444_));
 sg13g2_nor2_1 _7440_ (.A(_3396_),
    .B(_3426_),
    .Y(_3445_));
 sg13g2_a21oi_1 _7441_ (.A1(net1210),
    .A2(_3445_),
    .Y(_3446_),
    .B1(_3444_));
 sg13g2_and2_1 _7442_ (.A(net1212),
    .B(_3446_),
    .X(_3447_));
 sg13g2_a21oi_1 _7443_ (.A1(net1213),
    .A2(_3443_),
    .Y(_3448_),
    .B1(_3447_));
 sg13g2_nor2_1 _7444_ (.A(net1253),
    .B(net1251),
    .Y(_3449_));
 sg13g2_nand2_1 _7445_ (.Y(_3450_),
    .A(_3339_),
    .B(_3350_));
 sg13g2_nand2_2 _7446_ (.Y(_3451_),
    .A(_3339_),
    .B(net1252));
 sg13g2_nor2_1 _7447_ (.A(_3345_),
    .B(_3451_),
    .Y(_3452_));
 sg13g2_nor2_1 _7448_ (.A(_3449_),
    .B(_3452_),
    .Y(_3453_));
 sg13g2_nor2_1 _7449_ (.A(net1159),
    .B(_3453_),
    .Y(_3454_));
 sg13g2_a21oi_1 _7450_ (.A1(net1159),
    .A2(_3448_),
    .Y(_3455_),
    .B1(_3454_));
 sg13g2_nor2b_1 _7451_ (.A(_2589_),
    .B_N(_3455_),
    .Y(_3456_));
 sg13g2_nor2_1 _7452_ (.A(_2589_),
    .B(_3455_),
    .Y(_3457_));
 sg13g2_xor2_1 _7453_ (.B(_3455_),
    .A(_2589_),
    .X(_3458_));
 sg13g2_inv_2 _7454_ (.Y(_3459_),
    .A(_3458_));
 sg13g2_a21oi_1 _7455_ (.A1(_3439_),
    .A2(_3440_),
    .Y(_3460_),
    .B1(_3458_));
 sg13g2_o21ai_1 _7456_ (.B1(net1210),
    .Y(_3461_),
    .A1(net1213),
    .A2(_3427_));
 sg13g2_a21oi_1 _7457_ (.A1(net1263),
    .A2(_3397_),
    .Y(_3462_),
    .B1(_3461_));
 sg13g2_a22oi_1 _7458_ (.Y(_3463_),
    .B1(_3462_),
    .B2(net1158),
    .A2(_3352_),
    .A1(_3339_));
 sg13g2_or2_1 _7459_ (.X(_3464_),
    .B(_3463_),
    .A(_2610_));
 sg13g2_nand2_1 _7460_ (.Y(_3465_),
    .A(_2610_),
    .B(_3463_));
 sg13g2_nand2_2 _7461_ (.Y(_3466_),
    .A(_3464_),
    .B(_3465_));
 sg13g2_nor2_1 _7462_ (.A(net1212),
    .B(_3405_),
    .Y(_3467_));
 sg13g2_a21oi_1 _7463_ (.A1(net1212),
    .A2(_3443_),
    .Y(_3468_),
    .B1(_3467_));
 sg13g2_nor4_1 _7464_ (.A(net1158),
    .B(net1252),
    .C(_3346_),
    .D(_3450_),
    .Y(_3469_));
 sg13g2_a21oi_2 _7465_ (.B1(_3469_),
    .Y(_3470_),
    .A2(_3468_),
    .A1(net1158));
 sg13g2_nand2b_1 _7466_ (.Y(_3471_),
    .B(_3470_),
    .A_N(_2591_));
 sg13g2_nor2_1 _7467_ (.A(_2591_),
    .B(_3470_),
    .Y(_3472_));
 sg13g2_inv_1 _7468_ (.Y(_3473_),
    .A(_3472_));
 sg13g2_xnor2_1 _7469_ (.Y(_3474_),
    .A(_2591_),
    .B(_3470_));
 sg13g2_and3_1 _7470_ (.X(_3475_),
    .A(_3460_),
    .B(_3466_),
    .C(_3474_));
 sg13g2_nor2_1 _7471_ (.A(_3374_),
    .B(net1186),
    .Y(_3476_));
 sg13g2_mux2_1 _7472_ (.A0(_3374_),
    .A1(_3395_),
    .S(net1186),
    .X(_3477_));
 sg13g2_o21ai_1 _7473_ (.B1(_3477_),
    .Y(_3478_),
    .A1(_3384_),
    .A2(_3394_));
 sg13g2_a21oi_1 _7474_ (.A1(_3374_),
    .A2(_3394_),
    .Y(_3479_),
    .B1(net1187));
 sg13g2_a21oi_1 _7475_ (.A1(_3365_),
    .A2(_3385_),
    .Y(_3480_),
    .B1(_3479_));
 sg13g2_nand2_1 _7476_ (.Y(_3481_),
    .A(_3478_),
    .B(_3480_));
 sg13g2_nor2_1 _7477_ (.A(net1210),
    .B(_3445_),
    .Y(_3482_));
 sg13g2_a21oi_1 _7478_ (.A1(net1209),
    .A2(_3481_),
    .Y(_3483_),
    .B1(_3482_));
 sg13g2_mux2_1 _7479_ (.A0(_3434_),
    .A1(_3483_),
    .S(net1212),
    .X(_3484_));
 sg13g2_a21oi_2 _7480_ (.B1(_3353_),
    .Y(_3485_),
    .A2(_3484_),
    .A1(net1158));
 sg13g2_nand2b_1 _7481_ (.Y(_3486_),
    .B(_3485_),
    .A_N(_2601_));
 sg13g2_nor2_1 _7482_ (.A(_2601_),
    .B(_3485_),
    .Y(_3487_));
 sg13g2_nand2_1 _7483_ (.Y(_3488_),
    .A(_2601_),
    .B(_3485_));
 sg13g2_nand2b_1 _7484_ (.Y(_3489_),
    .B(_3488_),
    .A_N(_3487_));
 sg13g2_inv_2 _7485_ (.Y(_3490_),
    .A(_3489_));
 sg13g2_nor2_1 _7486_ (.A(_3424_),
    .B(_3451_),
    .Y(_3491_));
 sg13g2_mux2_1 _7487_ (.A0(_3451_),
    .A1(_3491_),
    .S(_3351_),
    .X(_3492_));
 sg13g2_inv_1 _7488_ (.Y(_3493_),
    .A(_3492_));
 sg13g2_a22oi_1 _7489_ (.Y(_3494_),
    .B1(_3478_),
    .B2(net1187),
    .A2(_3426_),
    .A1(net1186));
 sg13g2_a21oi_1 _7490_ (.A1(_3478_),
    .A2(_3480_),
    .Y(_3495_),
    .B1(net1209));
 sg13g2_a21oi_1 _7491_ (.A1(net1209),
    .A2(_3494_),
    .Y(_3496_),
    .B1(_3495_));
 sg13g2_a21oi_1 _7492_ (.A1(net1213),
    .A2(_3446_),
    .Y(_3497_),
    .B1(net1155));
 sg13g2_o21ai_1 _7493_ (.B1(_3497_),
    .Y(_3498_),
    .A1(net1213),
    .A2(_3496_));
 sg13g2_o21ai_1 _7494_ (.B1(_3498_),
    .Y(_3499_),
    .A1(net1161),
    .A2(_3493_));
 sg13g2_or2_1 _7495_ (.X(_3500_),
    .B(_3499_),
    .A(_2599_));
 sg13g2_o21ai_1 _7496_ (.B1(_3486_),
    .Y(_3501_),
    .A1(_3490_),
    .A2(_3500_));
 sg13g2_nand2b_1 _7497_ (.Y(_3502_),
    .B(_3499_),
    .A_N(_2599_));
 sg13g2_nand2b_1 _7498_ (.Y(_3503_),
    .B(_2599_),
    .A_N(_3499_));
 sg13g2_nand2_1 _7499_ (.Y(_3504_),
    .A(_3502_),
    .B(_3503_));
 sg13g2_inv_2 _7500_ (.Y(_3505_),
    .A(_3504_));
 sg13g2_nand2_1 _7501_ (.Y(_3506_),
    .A(_3489_),
    .B(_3504_));
 sg13g2_inv_1 _7502_ (.Y(_3507_),
    .A(_3506_));
 sg13g2_nand2_1 _7503_ (.Y(_3508_),
    .A(_3346_),
    .B(net1251));
 sg13g2_a21oi_1 _7504_ (.A1(_3346_),
    .A2(net1251),
    .Y(_3509_),
    .B1(net1253));
 sg13g2_nand2_1 _7505_ (.Y(_3510_),
    .A(net1253),
    .B(net1251));
 sg13g2_nor2_1 _7506_ (.A(_3339_),
    .B(_3354_),
    .Y(_3511_));
 sg13g2_a221oi_1 _7507_ (.B2(_3509_),
    .C1(_3511_),
    .B1(_3423_),
    .A1(net1253),
    .Y(_3512_),
    .A2(net1251));
 sg13g2_nand3_1 _7508_ (.B(net1186),
    .C(_3394_),
    .A(_3375_),
    .Y(_3513_));
 sg13g2_nor4_1 _7509_ (.A(_3365_),
    .B(_3374_),
    .C(_3385_),
    .D(_3395_),
    .Y(_3514_));
 sg13g2_nor3_1 _7510_ (.A(_3365_),
    .B(net1186),
    .C(_3394_),
    .Y(_3515_));
 sg13g2_nor3_1 _7511_ (.A(_3479_),
    .B(_3514_),
    .C(_3515_),
    .Y(_3516_));
 sg13g2_nand2_1 _7512_ (.Y(_3517_),
    .A(net1208),
    .B(_3516_));
 sg13g2_o21ai_1 _7513_ (.B1(_3517_),
    .Y(_3518_),
    .A1(net1209),
    .A2(_3494_));
 sg13g2_nand2_1 _7514_ (.Y(_3519_),
    .A(net1211),
    .B(_3518_));
 sg13g2_nand2_1 _7515_ (.Y(_3520_),
    .A(net1213),
    .B(_3483_));
 sg13g2_a21oi_1 _7516_ (.A1(_3519_),
    .A2(_3520_),
    .Y(_3521_),
    .B1(net1155));
 sg13g2_a21oi_1 _7517_ (.A1(net1155),
    .A2(_3512_),
    .Y(_3522_),
    .B1(_3521_));
 sg13g2_nand2b_1 _7518_ (.Y(_3523_),
    .B(_3522_),
    .A_N(_2612_));
 sg13g2_and2_1 _7519_ (.A(_2612_),
    .B(_3522_),
    .X(_3524_));
 sg13g2_nor2_1 _7520_ (.A(_2612_),
    .B(_3522_),
    .Y(_3525_));
 sg13g2_nor2_2 _7521_ (.A(_3524_),
    .B(_3525_),
    .Y(_3526_));
 sg13g2_inv_1 _7522_ (.Y(_3527_),
    .A(_3526_));
 sg13g2_xnor2_1 _7523_ (.Y(_3528_),
    .A(_3342_),
    .B(_3349_));
 sg13g2_nor2_1 _7524_ (.A(net1253),
    .B(_3528_),
    .Y(_3529_));
 sg13g2_o21ai_1 _7525_ (.B1(net1253),
    .Y(_3530_),
    .A1(net1252),
    .A2(_3350_));
 sg13g2_nor2_1 _7526_ (.A(_3422_),
    .B(_3530_),
    .Y(_3531_));
 sg13g2_nor2_1 _7527_ (.A(_3529_),
    .B(_3531_),
    .Y(_3532_));
 sg13g2_nand2_1 _7528_ (.Y(_3533_),
    .A(net1213),
    .B(_3496_));
 sg13g2_nand2_1 _7529_ (.Y(_3534_),
    .A(_3365_),
    .B(_3429_));
 sg13g2_nand2_1 _7530_ (.Y(_3535_),
    .A(_3513_),
    .B(_3534_));
 sg13g2_o21ai_1 _7531_ (.B1(_3535_),
    .Y(_3536_),
    .A1(net1187),
    .A2(_3513_));
 sg13g2_mux2_1 _7532_ (.A0(_3516_),
    .A1(_3536_),
    .S(net1208),
    .X(_3537_));
 sg13g2_nand2_1 _7533_ (.Y(_3538_),
    .A(net1211),
    .B(_3537_));
 sg13g2_nand3_1 _7534_ (.B(_3533_),
    .C(_3538_),
    .A(net1161),
    .Y(_3539_));
 sg13g2_o21ai_1 _7535_ (.B1(_3539_),
    .Y(_3540_),
    .A1(net1161),
    .A2(_3532_));
 sg13g2_nand2b_1 _7536_ (.Y(_3541_),
    .B(_3540_),
    .A_N(_2593_));
 sg13g2_nor2_1 _7537_ (.A(_3526_),
    .B(_3541_),
    .Y(_3542_));
 sg13g2_o21ai_1 _7538_ (.B1(_3523_),
    .Y(_3543_),
    .A1(_3526_),
    .A2(_3541_));
 sg13g2_nand3_1 _7539_ (.B(_3451_),
    .C(_3510_),
    .A(_3345_),
    .Y(_3544_));
 sg13g2_nand3_1 _7540_ (.B(net1186),
    .C(_3395_),
    .A(_3375_),
    .Y(_3545_));
 sg13g2_and3_1 _7541_ (.X(_3546_),
    .A(_3429_),
    .B(_3480_),
    .C(_3545_));
 sg13g2_mux2_1 _7542_ (.A0(_3536_),
    .A1(_3546_),
    .S(net1208),
    .X(_3547_));
 sg13g2_nand2_1 _7543_ (.Y(_3548_),
    .A(net1211),
    .B(_3547_));
 sg13g2_a21oi_1 _7544_ (.A1(net1213),
    .A2(_3518_),
    .Y(_3549_),
    .B1(net1155));
 sg13g2_a22oi_1 _7545_ (.Y(_3550_),
    .B1(_3548_),
    .B2(_3549_),
    .A2(_3544_),
    .A1(net1155));
 sg13g2_nand2_1 _7546_ (.Y(_3551_),
    .A(_2608_),
    .B(_3550_));
 sg13g2_or2_1 _7547_ (.X(_3552_),
    .B(_3550_),
    .A(_2608_));
 sg13g2_a21oi_1 _7548_ (.A1(net1252),
    .A2(_3350_),
    .Y(_3553_),
    .B1(_3345_));
 sg13g2_a21oi_1 _7549_ (.A1(_3450_),
    .A2(_3553_),
    .Y(_3554_),
    .B1(_3529_));
 sg13g2_nand3_1 _7550_ (.B(_3385_),
    .C(_3395_),
    .A(_3375_),
    .Y(_3555_));
 sg13g2_nand2_1 _7551_ (.Y(_3556_),
    .A(_3365_),
    .B(_3431_));
 sg13g2_nand3_1 _7552_ (.B(_3555_),
    .C(_3556_),
    .A(_3513_),
    .Y(_3557_));
 sg13g2_nand2_1 _7553_ (.Y(_3558_),
    .A(net1208),
    .B(_3557_));
 sg13g2_o21ai_1 _7554_ (.B1(_3558_),
    .Y(_3559_),
    .A1(net1208),
    .A2(_3546_));
 sg13g2_a21oi_1 _7555_ (.A1(net1211),
    .A2(_3559_),
    .Y(_3560_),
    .B1(net1155));
 sg13g2_o21ai_1 _7556_ (.B1(_3560_),
    .Y(_3561_),
    .A1(_3403_),
    .A2(_3537_));
 sg13g2_o21ai_1 _7557_ (.B1(_3561_),
    .Y(_3562_),
    .A1(net1161),
    .A2(_3554_));
 sg13g2_nor2_1 _7558_ (.A(_2614_),
    .B(_3562_),
    .Y(_3563_));
 sg13g2_a21oi_1 _7559_ (.A1(_3346_),
    .A2(_3449_),
    .Y(_3564_),
    .B1(net1252));
 sg13g2_nor2_1 _7560_ (.A(_3452_),
    .B(_3564_),
    .Y(_3565_));
 sg13g2_nor2_1 _7561_ (.A(net1161),
    .B(_3565_),
    .Y(_3566_));
 sg13g2_a21oi_1 _7562_ (.A1(_3365_),
    .A2(_3476_),
    .Y(_3567_),
    .B1(_3516_));
 sg13g2_mux2_1 _7563_ (.A0(_3557_),
    .A1(_3567_),
    .S(net1209),
    .X(_3568_));
 sg13g2_nor2_1 _7564_ (.A(_3402_),
    .B(_3568_),
    .Y(_3569_));
 sg13g2_a221oi_1 _7565_ (.B2(_3547_),
    .C1(_3569_),
    .B1(_3402_),
    .A1(_2653_),
    .Y(_3570_),
    .A2(_2657_));
 sg13g2_or2_1 _7566_ (.X(_3571_),
    .B(_3570_),
    .A(_3566_));
 sg13g2_nand2b_1 _7567_ (.Y(_3572_),
    .B(_3571_),
    .A_N(_2597_));
 sg13g2_a22oi_1 _7568_ (.Y(_3573_),
    .B1(_3555_),
    .B2(_3479_),
    .A2(_3545_),
    .A1(net1187));
 sg13g2_mux2_1 _7569_ (.A0(_3567_),
    .A1(_3573_),
    .S(net1208),
    .X(_3574_));
 sg13g2_mux2_1 _7570_ (.A0(_3559_),
    .A1(_3574_),
    .S(net1211),
    .X(_3575_));
 sg13g2_nor2_1 _7571_ (.A(_3346_),
    .B(_3528_),
    .Y(_3576_));
 sg13g2_nor2_1 _7572_ (.A(net1253),
    .B(_3576_),
    .Y(_3577_));
 sg13g2_a21oi_1 _7573_ (.A1(_3345_),
    .A2(_3528_),
    .Y(_3578_),
    .B1(_3577_));
 sg13g2_mux2_1 _7574_ (.A0(_3575_),
    .A1(_3578_),
    .S(net1155),
    .X(_3579_));
 sg13g2_nand2_1 _7575_ (.Y(_3580_),
    .A(_2631_),
    .B(_3579_));
 sg13g2_or2_1 _7576_ (.X(_3581_),
    .B(_3579_),
    .A(_2630_));
 sg13g2_xnor2_1 _7577_ (.Y(_3582_),
    .A(_2631_),
    .B(_3579_));
 sg13g2_o21ai_1 _7578_ (.B1(_3430_),
    .Y(_3583_),
    .A1(_3364_),
    .A2(_3477_));
 sg13g2_mux2_1 _7579_ (.A0(_3573_),
    .A1(_3583_),
    .S(net1208),
    .X(_3584_));
 sg13g2_o21ai_1 _7580_ (.B1(_3451_),
    .Y(_3585_),
    .A1(net1251),
    .A2(_3423_));
 sg13g2_nand2b_1 _7581_ (.Y(_3586_),
    .B(_3585_),
    .A_N(net1161));
 sg13g2_nor2_1 _7582_ (.A(_3403_),
    .B(_3568_),
    .Y(_3587_));
 sg13g2_o21ai_1 _7583_ (.B1(net1161),
    .Y(_3588_),
    .A1(_3402_),
    .A2(_3584_));
 sg13g2_o21ai_1 _7584_ (.B1(_3586_),
    .Y(_3589_),
    .A1(_3587_),
    .A2(_3588_));
 sg13g2_or2_1 _7585_ (.X(_3590_),
    .B(_3589_),
    .A(_2628_));
 sg13g2_inv_1 _7586_ (.Y(_3591_),
    .A(_3590_));
 sg13g2_a21o_1 _7587_ (.A2(_3511_),
    .A1(_3508_),
    .B1(_3577_),
    .X(_3592_));
 sg13g2_nand2_1 _7588_ (.Y(_3593_),
    .A(_3365_),
    .B(_3374_));
 sg13g2_nand2_1 _7589_ (.Y(_3594_),
    .A(_3555_),
    .B(_3593_));
 sg13g2_mux4_1 _7590_ (.S0(net1208),
    .A0(_3567_),
    .A1(_3573_),
    .A2(_3583_),
    .A3(_3594_),
    .S1(net1211),
    .X(_3595_));
 sg13g2_mux2_1 _7591_ (.A0(_3592_),
    .A1(_3595_),
    .S(net1162),
    .X(_3596_));
 sg13g2_inv_1 _7592_ (.Y(_3597_),
    .A(_3596_));
 sg13g2_nor2_1 _7593_ (.A(_2619_),
    .B(_3597_),
    .Y(_3598_));
 sg13g2_nand2_1 _7594_ (.Y(_3599_),
    .A(_2619_),
    .B(_3596_));
 sg13g2_inv_1 _7595_ (.Y(_3600_),
    .A(_3599_));
 sg13g2_nand2b_1 _7596_ (.Y(_3601_),
    .B(_2618_),
    .A_N(_3596_));
 sg13g2_and2_1 _7597_ (.A(_3599_),
    .B(_3601_),
    .X(_3602_));
 sg13g2_nand2_1 _7598_ (.Y(_3603_),
    .A(_3599_),
    .B(_3601_));
 sg13g2_and3_1 _7599_ (.X(_3604_),
    .A(net1263),
    .B(_3555_),
    .C(_3593_));
 sg13g2_a22oi_1 _7600_ (.Y(_3605_),
    .B1(_3395_),
    .B2(_3375_),
    .A2(net1186),
    .A1(_3365_));
 sg13g2_and3_1 _7601_ (.X(_3606_),
    .A(net1209),
    .B(_3430_),
    .C(_3605_));
 sg13g2_o21ai_1 _7602_ (.B1(net1211),
    .Y(_3607_),
    .A1(_3604_),
    .A2(_3606_));
 sg13g2_o21ai_1 _7603_ (.B1(_3607_),
    .Y(_3608_),
    .A1(net1211),
    .A2(_3584_));
 sg13g2_a22oi_1 _7604_ (.Y(_3609_),
    .B1(_3423_),
    .B2(_3510_),
    .A2(_3422_),
    .A1(_3340_));
 sg13g2_mux2_1 _7605_ (.A0(_3609_),
    .A1(_3608_),
    .S(net1162),
    .X(_3610_));
 sg13g2_or2_1 _7606_ (.X(_3611_),
    .B(_3610_),
    .A(_2595_));
 sg13g2_o21ai_1 _7607_ (.B1(_3493_),
    .Y(_3612_),
    .A1(_3342_),
    .A2(_3577_));
 sg13g2_nand2b_2 _7608_ (.Y(_3613_),
    .B(_3612_),
    .A_N(net1162));
 sg13g2_and2_1 _7609_ (.A(_2606_),
    .B(_3613_),
    .X(_3614_));
 sg13g2_nor2b_1 _7610_ (.A(_2595_),
    .B_N(_3610_),
    .Y(_3615_));
 sg13g2_xnor2_1 _7611_ (.Y(_3616_),
    .A(_2595_),
    .B(_3610_));
 sg13g2_o21ai_1 _7612_ (.B1(_3611_),
    .Y(_3617_),
    .A1(_3614_),
    .A2(_3616_));
 sg13g2_and2_1 _7613_ (.A(_3603_),
    .B(_3617_),
    .X(_3618_));
 sg13g2_nor2_1 _7614_ (.A(_3598_),
    .B(_3618_),
    .Y(_3619_));
 sg13g2_a221oi_1 _7615_ (.B2(_3617_),
    .C1(_3598_),
    .B1(_3603_),
    .A1(_2628_),
    .Y(_3620_),
    .A2(_3589_));
 sg13g2_or3_1 _7616_ (.A(_3582_),
    .B(_3591_),
    .C(_3620_),
    .X(_3621_));
 sg13g2_nor2_1 _7617_ (.A(_2597_),
    .B(_3571_),
    .Y(_3622_));
 sg13g2_xnor2_1 _7618_ (.Y(_3623_),
    .A(_2597_),
    .B(_3571_));
 sg13g2_xor2_1 _7619_ (.B(_3571_),
    .A(_2597_),
    .X(_3624_));
 sg13g2_a21o_1 _7620_ (.A2(_3621_),
    .A1(_3580_),
    .B1(_3624_),
    .X(_3625_));
 sg13g2_nand2b_1 _7621_ (.Y(_3626_),
    .B(_3562_),
    .A_N(_2614_));
 sg13g2_xnor2_1 _7622_ (.Y(_3627_),
    .A(_2614_),
    .B(_3562_));
 sg13g2_a21oi_1 _7623_ (.A1(_3572_),
    .A2(_3625_),
    .Y(_3628_),
    .B1(_3627_));
 sg13g2_nor2_1 _7624_ (.A(_3563_),
    .B(_3628_),
    .Y(_3629_));
 sg13g2_o21ai_1 _7625_ (.B1(_3551_),
    .Y(_3630_),
    .A1(_3563_),
    .A2(_3628_));
 sg13g2_and2_1 _7626_ (.A(_3552_),
    .B(_3630_),
    .X(_3631_));
 sg13g2_nor2_1 _7627_ (.A(_2593_),
    .B(_3540_),
    .Y(_3632_));
 sg13g2_inv_1 _7628_ (.Y(_3633_),
    .A(_3632_));
 sg13g2_xor2_1 _7629_ (.B(_3540_),
    .A(_2593_),
    .X(_3634_));
 sg13g2_nor2_1 _7630_ (.A(_3631_),
    .B(_3634_),
    .Y(_3635_));
 sg13g2_nor2_1 _7631_ (.A(_3526_),
    .B(_3634_),
    .Y(_3636_));
 sg13g2_nand2_1 _7632_ (.Y(_3637_),
    .A(_3527_),
    .B(_3635_));
 sg13g2_a21oi_1 _7633_ (.A1(_3527_),
    .A2(_3635_),
    .Y(_3638_),
    .B1(_3543_));
 sg13g2_a21oi_1 _7634_ (.A1(_3507_),
    .A2(_3543_),
    .Y(_3639_),
    .B1(_3501_));
 sg13g2_nand2_1 _7635_ (.Y(_3640_),
    .A(_3507_),
    .B(_3636_));
 sg13g2_o21ai_1 _7636_ (.B1(_3639_),
    .Y(_3641_),
    .A1(_3631_),
    .A2(_3640_));
 sg13g2_nor2b_1 _7637_ (.A(_2610_),
    .B_N(_3463_),
    .Y(_3642_));
 sg13g2_nand2_1 _7638_ (.Y(_3643_),
    .A(_3441_),
    .B(_3456_));
 sg13g2_o21ai_1 _7639_ (.B1(_3643_),
    .Y(_3644_),
    .A1(_2624_),
    .A2(_3438_));
 sg13g2_nand2_1 _7640_ (.Y(_3645_),
    .A(_3474_),
    .B(_3644_));
 sg13g2_nand2_1 _7641_ (.Y(_3646_),
    .A(_3471_),
    .B(_3645_));
 sg13g2_a221oi_1 _7642_ (.B2(_3466_),
    .C1(_3642_),
    .B1(_3646_),
    .A1(_3475_),
    .Y(_3647_),
    .A2(_3641_));
 sg13g2_nor2_1 _7643_ (.A(_2526_),
    .B(_3420_),
    .Y(_3648_));
 sg13g2_o21ai_1 _7644_ (.B1(_3421_),
    .Y(_3649_),
    .A1(_3647_),
    .A2(_3648_));
 sg13g2_nand2_1 _7645_ (.Y(_3650_),
    .A(net1257),
    .B(_3416_));
 sg13g2_nand2_1 _7646_ (.Y(_3651_),
    .A(_3415_),
    .B(_3650_));
 sg13g2_nor2_1 _7647_ (.A(_2533_),
    .B(_3419_),
    .Y(_3652_));
 sg13g2_nor2_1 _7648_ (.A(_3651_),
    .B(_3652_),
    .Y(_3653_));
 sg13g2_nor2_1 _7649_ (.A(_3648_),
    .B(_3652_),
    .Y(_3654_));
 sg13g2_a22oi_1 _7650_ (.Y(_3655_),
    .B1(_3649_),
    .B2(_3653_),
    .A2(_3418_),
    .A1(_3415_));
 sg13g2_nand2_1 _7651_ (.Y(_3656_),
    .A(_3421_),
    .B(_3654_));
 sg13g2_nor2b_1 _7652_ (.A(_3589_),
    .B_N(_2628_),
    .Y(_3657_));
 sg13g2_xor2_1 _7653_ (.B(_3589_),
    .A(_2628_),
    .X(_3658_));
 sg13g2_inv_1 _7654_ (.Y(_3659_),
    .A(_3658_));
 sg13g2_nand2_2 _7655_ (.Y(_3660_),
    .A(_3551_),
    .B(_3552_));
 sg13g2_inv_1 _7656_ (.Y(_3661_),
    .A(_3660_));
 sg13g2_and2_1 _7657_ (.A(_2605_),
    .B(_3613_),
    .X(_3662_));
 sg13g2_xnor2_1 _7658_ (.Y(_3663_),
    .A(_2606_),
    .B(_3613_));
 sg13g2_nor4_1 _7659_ (.A(_3616_),
    .B(_3627_),
    .C(_3659_),
    .D(_3663_),
    .Y(_3664_));
 sg13g2_nor4_1 _7660_ (.A(_3582_),
    .B(_3602_),
    .C(_3624_),
    .D(_3660_),
    .Y(_3665_));
 sg13g2_and2_1 _7661_ (.A(_3664_),
    .B(_3665_),
    .X(_3666_));
 sg13g2_nand4_1 _7662_ (.B(_3507_),
    .C(_3636_),
    .A(_3475_),
    .Y(_3667_),
    .D(_3666_));
 sg13g2_nor4_1 _7663_ (.A(_3418_),
    .B(_3651_),
    .C(_3656_),
    .D(_3667_),
    .Y(_3668_));
 sg13g2_o21ai_1 _7664_ (.B1(_3413_),
    .Y(_3669_),
    .A1(_3655_),
    .A2(_3668_));
 sg13g2_nand2b_1 _7665_ (.Y(_3670_),
    .B(_3411_),
    .A_N(_2560_));
 sg13g2_nand3_1 _7666_ (.B(_3411_),
    .C(_3412_),
    .A(net1259),
    .Y(_3671_));
 sg13g2_nand3_1 _7667_ (.B(_3670_),
    .C(_3671_),
    .A(_3669_),
    .Y(_3672_));
 sg13g2_a21oi_1 _7668_ (.A1(_2530_),
    .A2(_3411_),
    .Y(_3673_),
    .B1(net1261));
 sg13g2_a21oi_1 _7669_ (.A1(_2551_),
    .A2(_3411_),
    .Y(_3674_),
    .B1(_2548_));
 sg13g2_nor2_1 _7670_ (.A(_3673_),
    .B(_3674_),
    .Y(_3675_));
 sg13g2_nand2_1 _7671_ (.Y(_3676_),
    .A(_3672_),
    .B(_3675_));
 sg13g2_o21ai_1 _7672_ (.B1(_3411_),
    .Y(_3677_),
    .A1(_2553_),
    .A2(_2555_));
 sg13g2_a21oi_1 _7673_ (.A1(_2543_),
    .A2(_3411_),
    .Y(_3678_),
    .B1(net1263));
 sg13g2_a21o_2 _7674_ (.A2(_3677_),
    .A1(_3676_),
    .B1(_3678_),
    .X(_3679_));
 sg13g2_nor2_2 _7675_ (.A(_2648_),
    .B(_2658_),
    .Y(_3680_));
 sg13g2_nor2_1 _7676_ (.A(_2534_),
    .B(_3399_),
    .Y(_3681_));
 sg13g2_nand2_1 _7677_ (.Y(_3682_),
    .A(_2534_),
    .B(_3399_));
 sg13g2_nand2_1 _7678_ (.Y(_3683_),
    .A(_2526_),
    .B(_3406_));
 sg13g2_nor2_1 _7679_ (.A(_2527_),
    .B(_3406_),
    .Y(_3684_));
 sg13g2_xnor2_1 _7680_ (.Y(_3685_),
    .A(_2526_),
    .B(_3406_));
 sg13g2_inv_2 _7681_ (.Y(_3686_),
    .A(_3685_));
 sg13g2_o21ai_1 _7682_ (.B1(_3683_),
    .Y(_3687_),
    .A1(_3647_),
    .A2(_3685_));
 sg13g2_o21ai_1 _7683_ (.B1(_3682_),
    .Y(_3688_),
    .A1(_3681_),
    .A2(_3687_));
 sg13g2_and2_1 _7684_ (.A(net1257),
    .B(_3688_),
    .X(_3689_));
 sg13g2_and2_1 _7685_ (.A(net1258),
    .B(_3689_),
    .X(_3690_));
 sg13g2_nand2_1 _7686_ (.Y(_3691_),
    .A(_2533_),
    .B(_3399_));
 sg13g2_inv_1 _7687_ (.Y(_3692_),
    .A(_3691_));
 sg13g2_nand2b_2 _7688_ (.Y(_3693_),
    .B(_2534_),
    .A_N(_3399_));
 sg13g2_nand2_2 _7689_ (.Y(_3694_),
    .A(_3691_),
    .B(_3693_));
 sg13g2_nand4_1 _7690_ (.B(net1257),
    .C(_3686_),
    .A(net1258),
    .Y(_3695_),
    .D(_3694_));
 sg13g2_nor2_1 _7691_ (.A(_3667_),
    .B(_3695_),
    .Y(_3696_));
 sg13g2_or2_1 _7692_ (.X(_3697_),
    .B(_3696_),
    .A(_3690_));
 sg13g2_nand4_1 _7693_ (.B(net1259),
    .C(net1213),
    .A(net1261),
    .Y(_3698_),
    .D(_3697_));
 sg13g2_a22oi_1 _7694_ (.Y(_3699_),
    .B1(_3698_),
    .B2(_2651_),
    .A2(_3680_),
    .A1(_3679_));
 sg13g2_inv_2 _7695_ (.Y(_3700_),
    .A(net1138));
 sg13g2_o21ai_1 _7696_ (.B1(net1162),
    .Y(_3701_),
    .A1(_2605_),
    .A2(_3699_));
 sg13g2_a21oi_1 _7697_ (.A1(_3616_),
    .A2(_3662_),
    .Y(_3702_),
    .B1(_3615_));
 sg13g2_a221oi_1 _7698_ (.B2(_3662_),
    .C1(_3615_),
    .B1(_3616_),
    .A1(_2618_),
    .Y(_3703_),
    .A2(_3597_));
 sg13g2_nor3_1 _7699_ (.A(_3600_),
    .B(_3658_),
    .C(_3703_),
    .Y(_3704_));
 sg13g2_o21ai_1 _7700_ (.B1(_3582_),
    .Y(_3705_),
    .A1(_3657_),
    .A2(_3704_));
 sg13g2_a21oi_1 _7701_ (.A1(_3581_),
    .A2(_3705_),
    .Y(_3706_),
    .B1(_3623_));
 sg13g2_o21ai_1 _7702_ (.B1(_3627_),
    .Y(_3707_),
    .A1(_3622_),
    .A2(_3706_));
 sg13g2_a21oi_1 _7703_ (.A1(_3626_),
    .A2(_3707_),
    .Y(_3708_),
    .B1(_3661_));
 sg13g2_nor2b_1 _7704_ (.A(_2608_),
    .B_N(_3550_),
    .Y(_3709_));
 sg13g2_or2_1 _7705_ (.X(_3710_),
    .B(_3709_),
    .A(_3708_));
 sg13g2_o21ai_1 _7706_ (.B1(_3634_),
    .Y(_3711_),
    .A1(_3708_),
    .A2(_3709_));
 sg13g2_nand2_1 _7707_ (.Y(_3712_),
    .A(_3633_),
    .B(_3711_));
 sg13g2_a21oi_1 _7708_ (.A1(_3633_),
    .A2(_3711_),
    .Y(_3713_),
    .B1(_3524_));
 sg13g2_nor2_1 _7709_ (.A(_3525_),
    .B(_3713_),
    .Y(_3714_));
 sg13g2_o21ai_1 _7710_ (.B1(_3502_),
    .Y(_3715_),
    .A1(_3504_),
    .A2(_3714_));
 sg13g2_nor2b_1 _7711_ (.A(_3487_),
    .B_N(_3502_),
    .Y(_3716_));
 sg13g2_o21ai_1 _7712_ (.B1(_3503_),
    .Y(_3717_),
    .A1(_3525_),
    .A2(_3713_));
 sg13g2_a21oi_1 _7713_ (.A1(_3488_),
    .A2(_3715_),
    .Y(_3718_),
    .B1(_3487_));
 sg13g2_a221oi_1 _7714_ (.B2(_3717_),
    .C1(_3459_),
    .B1(_3716_),
    .A1(_2601_),
    .Y(_3719_),
    .A2(_3485_));
 sg13g2_or2_1 _7715_ (.X(_3720_),
    .B(_3719_),
    .A(_3457_));
 sg13g2_o21ai_1 _7716_ (.B1(_3439_),
    .Y(_3721_),
    .A1(_3457_),
    .A2(_3719_));
 sg13g2_and2_1 _7717_ (.A(_3440_),
    .B(_3721_),
    .X(_3722_));
 sg13g2_a21o_1 _7718_ (.A2(_3721_),
    .A1(_3440_),
    .B1(_3474_),
    .X(_3723_));
 sg13g2_and2_1 _7719_ (.A(_3464_),
    .B(_3473_),
    .X(_3724_));
 sg13g2_nand2_1 _7720_ (.Y(_3725_),
    .A(_3723_),
    .B(_3724_));
 sg13g2_nand2_1 _7721_ (.Y(_3726_),
    .A(_3465_),
    .B(_3725_));
 sg13g2_a221oi_1 _7722_ (.B2(_3724_),
    .C1(_3686_),
    .B1(_3723_),
    .A1(_2610_),
    .Y(_3727_),
    .A2(_3463_));
 sg13g2_nor2_1 _7723_ (.A(_3684_),
    .B(_3727_),
    .Y(_3728_));
 sg13g2_or3_1 _7724_ (.A(_3684_),
    .B(_3692_),
    .C(_3727_),
    .X(_3729_));
 sg13g2_nand2_1 _7725_ (.Y(_3730_),
    .A(_3693_),
    .B(_3729_));
 sg13g2_nand4_1 _7726_ (.B(_2575_),
    .C(_3693_),
    .A(_2570_),
    .Y(_3731_),
    .D(_3729_));
 sg13g2_nor3_1 _7727_ (.A(net1261),
    .B(net1259),
    .C(_3731_),
    .Y(_3732_));
 sg13g2_nor2_1 _7728_ (.A(_2639_),
    .B(_3731_),
    .Y(_3733_));
 sg13g2_o21ai_1 _7729_ (.B1(_3701_),
    .Y(_3734_),
    .A1(_3663_),
    .A2(net1136));
 sg13g2_a21oi_1 _7730_ (.A1(net1334),
    .A2(_3734_),
    .Y(_0446_),
    .B1(_3334_));
 sg13g2_xor2_1 _7731_ (.B(_3662_),
    .A(_3616_),
    .X(_3735_));
 sg13g2_o21ai_1 _7732_ (.B1(net1156),
    .Y(_3736_),
    .A1(net1136),
    .A2(_3735_));
 sg13g2_o21ai_1 _7733_ (.B1(net1161),
    .Y(_3737_),
    .A1(_2606_),
    .A2(_3616_));
 sg13g2_a21o_1 _7734_ (.A2(_3616_),
    .A1(_3614_),
    .B1(_3737_),
    .X(_3738_));
 sg13g2_o21ai_1 _7735_ (.B1(_3736_),
    .Y(_3739_),
    .A1(net1138),
    .A2(_3738_));
 sg13g2_mux2_1 _7736_ (.A0(net449),
    .A1(_3739_),
    .S(net1334),
    .X(_0447_));
 sg13g2_xnor2_1 _7737_ (.Y(_3740_),
    .A(_3602_),
    .B(_3702_));
 sg13g2_o21ai_1 _7738_ (.B1(net1157),
    .Y(_3741_),
    .A1(net1136),
    .A2(_3740_));
 sg13g2_nor2_1 _7739_ (.A(_3603_),
    .B(_3617_),
    .Y(_3742_));
 sg13g2_or3_1 _7740_ (.A(net1157),
    .B(_3618_),
    .C(net1138),
    .X(_3743_));
 sg13g2_o21ai_1 _7741_ (.B1(_3741_),
    .Y(_3744_),
    .A1(_3742_),
    .A2(_3743_));
 sg13g2_mux2_1 _7742_ (.A0(net330),
    .A1(_3744_),
    .S(net1336),
    .X(_0448_));
 sg13g2_o21ai_1 _7743_ (.B1(_3658_),
    .Y(_3745_),
    .A1(_3600_),
    .A2(_3703_));
 sg13g2_nor2b_1 _7744_ (.A(_3704_),
    .B_N(_3745_),
    .Y(_3746_));
 sg13g2_o21ai_1 _7745_ (.B1(net1156),
    .Y(_3747_),
    .A1(net1136),
    .A2(_3746_));
 sg13g2_xnor2_1 _7746_ (.Y(_3748_),
    .A(_3619_),
    .B(_3659_));
 sg13g2_o21ai_1 _7747_ (.B1(_3747_),
    .Y(_3749_),
    .A1(net1138),
    .A2(_3748_));
 sg13g2_mux2_1 _7748_ (.A0(net353),
    .A1(_3749_),
    .S(net1334),
    .X(_0449_));
 sg13g2_or3_1 _7749_ (.A(_3582_),
    .B(_3657_),
    .C(_3704_),
    .X(_3750_));
 sg13g2_and2_1 _7750_ (.A(_3705_),
    .B(_3750_),
    .X(_3751_));
 sg13g2_o21ai_1 _7751_ (.B1(net1156),
    .Y(_3752_),
    .A1(net1136),
    .A2(_3751_));
 sg13g2_o21ai_1 _7752_ (.B1(_3582_),
    .Y(_3753_),
    .A1(_3591_),
    .A2(_3620_));
 sg13g2_nand3_1 _7753_ (.B(_3621_),
    .C(_3753_),
    .A(net1163),
    .Y(_3754_));
 sg13g2_o21ai_1 _7754_ (.B1(_3752_),
    .Y(_3755_),
    .A1(net1138),
    .A2(_3754_));
 sg13g2_mux2_1 _7755_ (.A0(net402),
    .A1(_3755_),
    .S(net1336),
    .X(_0450_));
 sg13g2_nand3_1 _7756_ (.B(_3623_),
    .C(_3705_),
    .A(_3581_),
    .Y(_3756_));
 sg13g2_nor2b_1 _7757_ (.A(_3706_),
    .B_N(_3756_),
    .Y(_3757_));
 sg13g2_nor2_1 _7758_ (.A(net1136),
    .B(_3757_),
    .Y(_3758_));
 sg13g2_nand3_1 _7759_ (.B(_3621_),
    .C(_3624_),
    .A(_3580_),
    .Y(_3759_));
 sg13g2_nand4_1 _7760_ (.B(_3625_),
    .C(_3700_),
    .A(net1163),
    .Y(_3760_),
    .D(_3759_));
 sg13g2_o21ai_1 _7761_ (.B1(_3760_),
    .Y(_3761_),
    .A1(net1163),
    .A2(_3758_));
 sg13g2_mux2_1 _7762_ (.A0(net409),
    .A1(_3761_),
    .S(net1334),
    .X(_0451_));
 sg13g2_or3_1 _7763_ (.A(_3622_),
    .B(_3627_),
    .C(_3706_),
    .X(_3762_));
 sg13g2_and2_1 _7764_ (.A(_3707_),
    .B(_3762_),
    .X(_3763_));
 sg13g2_o21ai_1 _7765_ (.B1(net1157),
    .Y(_3764_),
    .A1(net1137),
    .A2(_3763_));
 sg13g2_and3_1 _7766_ (.X(_3765_),
    .A(_3572_),
    .B(_3625_),
    .C(_3627_));
 sg13g2_or3_1 _7767_ (.A(net1156),
    .B(_3628_),
    .C(net1138),
    .X(_3766_));
 sg13g2_o21ai_1 _7768_ (.B1(_3764_),
    .Y(_3767_),
    .A1(_3765_),
    .A2(_3766_));
 sg13g2_nand2_1 _7769_ (.Y(_3768_),
    .A(net1335),
    .B(_3767_));
 sg13g2_o21ai_1 _7770_ (.B1(_3768_),
    .Y(_0452_),
    .A1(_0859_),
    .A2(net1334));
 sg13g2_nand3_1 _7771_ (.B(_3661_),
    .C(_3707_),
    .A(_3626_),
    .Y(_3769_));
 sg13g2_nor2b_1 _7772_ (.A(_3708_),
    .B_N(_3769_),
    .Y(_3770_));
 sg13g2_o21ai_1 _7773_ (.B1(net1156),
    .Y(_3771_),
    .A1(net1136),
    .A2(_3770_));
 sg13g2_xnor2_1 _7774_ (.Y(_3772_),
    .A(_3629_),
    .B(_3660_));
 sg13g2_o21ai_1 _7775_ (.B1(_3771_),
    .Y(_3773_),
    .A1(net1138),
    .A2(_3772_));
 sg13g2_mux2_1 _7776_ (.A0(net422),
    .A1(_3773_),
    .S(net1334),
    .X(_0453_));
 sg13g2_xor2_1 _7777_ (.B(_3710_),
    .A(_3634_),
    .X(_3774_));
 sg13g2_nor2_1 _7778_ (.A(net1136),
    .B(_3774_),
    .Y(_3775_));
 sg13g2_a21oi_1 _7779_ (.A1(_3631_),
    .A2(_3634_),
    .Y(_3776_),
    .B1(net1156));
 sg13g2_nand3b_1 _7780_ (.B(_3700_),
    .C(_3776_),
    .Y(_3777_),
    .A_N(_3635_));
 sg13g2_o21ai_1 _7781_ (.B1(_3777_),
    .Y(_3778_),
    .A1(net1163),
    .A2(_3775_));
 sg13g2_mux2_1 _7782_ (.A0(net299),
    .A1(_3778_),
    .S(net1336),
    .X(_0454_));
 sg13g2_xnor2_1 _7783_ (.Y(_3779_),
    .A(_3527_),
    .B(_3712_));
 sg13g2_nor2_1 _7784_ (.A(net1137),
    .B(_3779_),
    .Y(_3780_));
 sg13g2_nand2_1 _7785_ (.Y(_3781_),
    .A(_3526_),
    .B(_3541_));
 sg13g2_o21ai_1 _7786_ (.B1(_3637_),
    .Y(_3782_),
    .A1(_3635_),
    .A2(_3781_));
 sg13g2_or4_1 _7787_ (.A(net1156),
    .B(_3542_),
    .C(net1138),
    .D(_3782_),
    .X(_3783_));
 sg13g2_o21ai_1 _7788_ (.B1(_3783_),
    .Y(_3784_),
    .A1(net1163),
    .A2(_3780_));
 sg13g2_nand2_1 _7789_ (.Y(_3785_),
    .A(net1335),
    .B(_3784_));
 sg13g2_o21ai_1 _7790_ (.B1(_3785_),
    .Y(_0455_),
    .A1(_0861_),
    .A2(net1334));
 sg13g2_nor2_1 _7791_ (.A(net214),
    .B(net1331),
    .Y(_3786_));
 sg13g2_xnor2_1 _7792_ (.Y(_3787_),
    .A(_3505_),
    .B(_3714_));
 sg13g2_nor2_2 _7793_ (.A(net1160),
    .B(net1137),
    .Y(_3788_));
 sg13g2_inv_2 _7794_ (.Y(_3789_),
    .A(net1135));
 sg13g2_xnor2_1 _7795_ (.Y(_3790_),
    .A(_3505_),
    .B(_3638_));
 sg13g2_o21ai_1 _7796_ (.B1(net1160),
    .Y(_3791_),
    .A1(net1139),
    .A2(_3790_));
 sg13g2_o21ai_1 _7797_ (.B1(_3791_),
    .Y(_3792_),
    .A1(_3787_),
    .A2(_3789_));
 sg13g2_a21oi_1 _7798_ (.A1(net1331),
    .A2(_3792_),
    .Y(_0456_),
    .B1(_3786_));
 sg13g2_o21ai_1 _7799_ (.B1(_3500_),
    .Y(_3793_),
    .A1(_3505_),
    .A2(_3638_));
 sg13g2_xnor2_1 _7800_ (.Y(_3794_),
    .A(_3490_),
    .B(_3793_));
 sg13g2_nand2_1 _7801_ (.Y(_3795_),
    .A(_3700_),
    .B(_3794_));
 sg13g2_xnor2_1 _7802_ (.Y(_3796_),
    .A(_3490_),
    .B(_3715_));
 sg13g2_a22oi_1 _7803_ (.Y(_3797_),
    .B1(_3796_),
    .B2(net1135),
    .A2(_3795_),
    .A1(net1163));
 sg13g2_mux2_1 _7804_ (.A0(net325),
    .A1(_3797_),
    .S(net1335),
    .X(_0457_));
 sg13g2_xnor2_1 _7805_ (.Y(_3798_),
    .A(_3458_),
    .B(_3718_));
 sg13g2_o21ai_1 _7806_ (.B1(net1156),
    .Y(_3799_),
    .A1(net1137),
    .A2(_3798_));
 sg13g2_xnor2_1 _7807_ (.Y(_3800_),
    .A(_3459_),
    .B(_3641_));
 sg13g2_o21ai_1 _7808_ (.B1(_3799_),
    .Y(_3801_),
    .A1(net1139),
    .A2(_3800_));
 sg13g2_nand2_1 _7809_ (.Y(_3802_),
    .A(net1332),
    .B(_3801_));
 sg13g2_o21ai_1 _7810_ (.B1(_3802_),
    .Y(_0458_),
    .A1(_0869_),
    .A2(net1332));
 sg13g2_xnor2_1 _7811_ (.Y(_3803_),
    .A(_3441_),
    .B(_3720_));
 sg13g2_nor2_1 _7812_ (.A(net1137),
    .B(_3803_),
    .Y(_3804_));
 sg13g2_or2_1 _7813_ (.X(_3805_),
    .B(_3456_),
    .A(_3441_));
 sg13g2_a21oi_1 _7814_ (.A1(_3459_),
    .A2(_3641_),
    .Y(_3806_),
    .B1(_3805_));
 sg13g2_and2_1 _7815_ (.A(_3460_),
    .B(_3641_),
    .X(_3807_));
 sg13g2_nand2_1 _7816_ (.Y(_3808_),
    .A(net1160),
    .B(_3643_));
 sg13g2_or4_1 _7817_ (.A(net1139),
    .B(_3806_),
    .C(_3807_),
    .D(_3808_),
    .X(_3809_));
 sg13g2_o21ai_1 _7818_ (.B1(_3809_),
    .Y(_3810_),
    .A1(net1160),
    .A2(_3804_));
 sg13g2_mux2_1 _7819_ (.A0(net427),
    .A1(_3810_),
    .S(net1335),
    .X(_0459_));
 sg13g2_nor2_1 _7820_ (.A(net221),
    .B(net1331),
    .Y(_3811_));
 sg13g2_xor2_1 _7821_ (.B(_3722_),
    .A(_3474_),
    .X(_3812_));
 sg13g2_or3_1 _7822_ (.A(_3474_),
    .B(_3644_),
    .C(_3807_),
    .X(_3813_));
 sg13g2_o21ai_1 _7823_ (.B1(_3474_),
    .Y(_3814_),
    .A1(_3644_),
    .A2(_3807_));
 sg13g2_nand2_1 _7824_ (.Y(_3815_),
    .A(_3813_),
    .B(_3814_));
 sg13g2_o21ai_1 _7825_ (.B1(net1160),
    .Y(_3816_),
    .A1(net1139),
    .A2(_3815_));
 sg13g2_o21ai_1 _7826_ (.B1(_3816_),
    .Y(_3817_),
    .A1(_3789_),
    .A2(_3812_));
 sg13g2_a21oi_1 _7827_ (.A1(net1331),
    .A2(_3817_),
    .Y(_0460_),
    .B1(_3811_));
 sg13g2_nand2_1 _7828_ (.Y(_3818_),
    .A(_3471_),
    .B(_3814_));
 sg13g2_xor2_1 _7829_ (.B(_3818_),
    .A(_3466_),
    .X(_3819_));
 sg13g2_nand2_1 _7830_ (.Y(_3820_),
    .A(_3700_),
    .B(_3819_));
 sg13g2_nand2_1 _7831_ (.Y(_3821_),
    .A(_3473_),
    .B(_3723_));
 sg13g2_xor2_1 _7832_ (.B(_3821_),
    .A(_3466_),
    .X(_3822_));
 sg13g2_a22oi_1 _7833_ (.Y(_3823_),
    .B1(_3822_),
    .B2(net1135),
    .A2(_3820_),
    .A1(net1160));
 sg13g2_mux2_1 _7834_ (.A0(net332),
    .A1(_3823_),
    .S(net1332),
    .X(_0461_));
 sg13g2_nor2_1 _7835_ (.A(net257),
    .B(net1331),
    .Y(_3824_));
 sg13g2_xnor2_1 _7836_ (.Y(_3825_),
    .A(_3686_),
    .B(_3726_));
 sg13g2_nand2_1 _7837_ (.Y(_3826_),
    .A(net1265),
    .B(_3680_));
 sg13g2_o21ai_1 _7838_ (.B1(_2653_),
    .Y(_3827_),
    .A1(net1265),
    .A2(_2657_));
 sg13g2_o21ai_1 _7839_ (.B1(_3827_),
    .Y(_3828_),
    .A1(_3679_),
    .A2(_3826_));
 sg13g2_nand2_1 _7840_ (.Y(_3829_),
    .A(net1139),
    .B(_3826_));
 sg13g2_xnor2_1 _7841_ (.Y(_3830_),
    .A(_3647_),
    .B(_3686_));
 sg13g2_a21oi_1 _7842_ (.A1(_3829_),
    .A2(_3830_),
    .Y(_3831_),
    .B1(_3828_));
 sg13g2_a21o_2 _7843_ (.A2(_3825_),
    .A1(net1135),
    .B1(_3831_),
    .X(_3832_));
 sg13g2_a21oi_1 _7844_ (.A1(net1332),
    .A2(_3832_),
    .Y(_0462_),
    .B1(_3824_));
 sg13g2_nand2_1 _7845_ (.Y(_3833_),
    .A(_2530_),
    .B(_3680_));
 sg13g2_nor2_1 _7846_ (.A(_3679_),
    .B(_3833_),
    .Y(_3834_));
 sg13g2_o21ai_1 _7847_ (.B1(_2653_),
    .Y(_3835_),
    .A1(_2530_),
    .A2(_2657_));
 sg13g2_nor2b_1 _7848_ (.A(_3834_),
    .B_N(_3835_),
    .Y(_3836_));
 sg13g2_nand2_1 _7849_ (.Y(_3837_),
    .A(net1139),
    .B(_3833_));
 sg13g2_xor2_1 _7850_ (.B(_3694_),
    .A(_3687_),
    .X(_3838_));
 sg13g2_nand2_1 _7851_ (.Y(_3839_),
    .A(_3837_),
    .B(_3838_));
 sg13g2_xnor2_1 _7852_ (.Y(_3840_),
    .A(_3694_),
    .B(_3728_));
 sg13g2_a22oi_1 _7853_ (.Y(_3841_),
    .B1(_3840_),
    .B2(net1135),
    .A2(_3839_),
    .A1(_3836_));
 sg13g2_mux2_1 _7854_ (.A0(net428),
    .A1(_3841_),
    .S(net1331),
    .X(_0463_));
 sg13g2_xnor2_1 _7855_ (.Y(_3842_),
    .A(net1257),
    .B(_3730_));
 sg13g2_o21ai_1 _7856_ (.B1(_2653_),
    .Y(_3843_),
    .A1(_2551_),
    .A2(_2657_));
 sg13g2_nand2_1 _7857_ (.Y(_3844_),
    .A(_2551_),
    .B(_3680_));
 sg13g2_and2_1 _7858_ (.A(net1139),
    .B(_3844_),
    .X(_3845_));
 sg13g2_xnor2_1 _7859_ (.Y(_3846_),
    .A(_2575_),
    .B(_3688_));
 sg13g2_o21ai_1 _7860_ (.B1(_3846_),
    .Y(_3847_),
    .A1(_3679_),
    .A2(_3844_));
 sg13g2_nand2b_1 _7861_ (.Y(_3848_),
    .B(_3847_),
    .A_N(_3845_));
 sg13g2_a22oi_1 _7862_ (.Y(_3849_),
    .B1(_3843_),
    .B2(_3848_),
    .A2(_3842_),
    .A1(net1135));
 sg13g2_mux2_1 _7863_ (.A0(net365),
    .A1(_3849_),
    .S(net1336),
    .X(_0464_));
 sg13g2_o21ai_1 _7864_ (.B1(_2571_),
    .Y(_3850_),
    .A1(net1257),
    .A2(_3730_));
 sg13g2_nand2_1 _7865_ (.Y(_3851_),
    .A(_3731_),
    .B(_3850_));
 sg13g2_o21ai_1 _7866_ (.B1(_2653_),
    .Y(_3852_),
    .A1(_2543_),
    .A2(_2657_));
 sg13g2_nand2_1 _7867_ (.Y(_3853_),
    .A(_2543_),
    .B(_3680_));
 sg13g2_nand2_1 _7868_ (.Y(_3854_),
    .A(net1139),
    .B(_3853_));
 sg13g2_nor2b_1 _7869_ (.A(_3854_),
    .B_N(_3852_),
    .Y(_3855_));
 sg13g2_o21ai_1 _7870_ (.B1(_3852_),
    .Y(_3856_),
    .A1(_3679_),
    .A2(_3853_));
 sg13g2_inv_1 _7871_ (.Y(_3857_),
    .A(_3856_));
 sg13g2_xnor2_1 _7872_ (.Y(_3858_),
    .A(_2570_),
    .B(_3689_));
 sg13g2_a221oi_1 _7873_ (.B2(_3858_),
    .C1(_3855_),
    .B1(_3857_),
    .A1(net1135),
    .Y(_3859_),
    .A2(_3851_));
 sg13g2_mux2_1 _7874_ (.A0(net459),
    .A1(_3859_),
    .S(net1331),
    .X(_0465_));
 sg13g2_xnor2_1 _7875_ (.Y(_3860_),
    .A(net1260),
    .B(_3731_));
 sg13g2_xnor2_1 _7876_ (.Y(_3861_),
    .A(net1260),
    .B(_3690_));
 sg13g2_a21oi_1 _7877_ (.A1(_3829_),
    .A2(_3861_),
    .Y(_3862_),
    .B1(_3828_));
 sg13g2_a21oi_2 _7878_ (.B1(_3862_),
    .Y(_3863_),
    .A2(_3860_),
    .A1(_3788_));
 sg13g2_mux2_1 _7879_ (.A0(net328),
    .A1(_3863_),
    .S(net1336),
    .X(_0466_));
 sg13g2_o21ai_1 _7880_ (.B1(net1261),
    .Y(_3864_),
    .A1(net1259),
    .A2(_3731_));
 sg13g2_nand2b_1 _7881_ (.Y(_3865_),
    .B(_3864_),
    .A_N(_3732_));
 sg13g2_and3_2 _7882_ (.X(_3866_),
    .A(net1261),
    .B(net1259),
    .C(_3690_));
 sg13g2_a21oi_1 _7883_ (.A1(net1259),
    .A2(_3690_),
    .Y(_3867_),
    .B1(net1261));
 sg13g2_o21ai_1 _7884_ (.B1(_3837_),
    .Y(_3868_),
    .A1(_3866_),
    .A2(_3867_));
 sg13g2_a22oi_1 _7885_ (.Y(_3869_),
    .B1(_3868_),
    .B2(_3836_),
    .A2(_3865_),
    .A1(net1135));
 sg13g2_mux2_1 _7886_ (.A0(net423),
    .A1(_3869_),
    .S(net1331),
    .X(_0467_));
 sg13g2_nor2_1 _7887_ (.A(net194),
    .B(net1333),
    .Y(_3870_));
 sg13g2_xnor2_1 _7888_ (.Y(_3871_),
    .A(_2548_),
    .B(_3732_));
 sg13g2_and2_1 _7889_ (.A(_2548_),
    .B(_3866_),
    .X(_3872_));
 sg13g2_xnor2_1 _7890_ (.Y(_3873_),
    .A(_2547_),
    .B(_3866_));
 sg13g2_o21ai_1 _7891_ (.B1(_3843_),
    .Y(_3874_),
    .A1(_3845_),
    .A2(_3873_));
 sg13g2_o21ai_1 _7892_ (.B1(_3874_),
    .Y(_3875_),
    .A1(_3789_),
    .A2(_3871_));
 sg13g2_a21oi_1 _7893_ (.A1(net1333),
    .A2(_3875_),
    .Y(_0468_),
    .B1(_3870_));
 sg13g2_nor2_1 _7894_ (.A(net185),
    .B(net1333),
    .Y(_3876_));
 sg13g2_xnor2_1 _7895_ (.Y(_3877_),
    .A(net1263),
    .B(_3872_));
 sg13g2_a21oi_1 _7896_ (.A1(_3854_),
    .A2(_3877_),
    .Y(_3878_),
    .B1(_3856_));
 sg13g2_a221oi_1 _7897_ (.B2(_3732_),
    .C1(net1160),
    .B1(_2547_),
    .A1(_2537_),
    .Y(_3879_),
    .A2(_2538_));
 sg13g2_or2_1 _7898_ (.X(_3880_),
    .B(_3879_),
    .A(_3878_));
 sg13g2_a21oi_1 _7899_ (.A1(net1333),
    .A2(_3880_),
    .Y(_0469_),
    .B1(_3876_));
 sg13g2_nor2_1 _7900_ (.A(net143),
    .B(net1333),
    .Y(_3881_));
 sg13g2_a21oi_1 _7901_ (.A1(_2654_),
    .A2(net1333),
    .Y(_0470_),
    .B1(_3881_));
 sg13g2_nor2_1 _7902_ (.A(net176),
    .B(net1333),
    .Y(_3882_));
 sg13g2_a21oi_1 _7903_ (.A1(_2658_),
    .A2(net1333),
    .Y(_0471_),
    .B1(_3882_));
 sg13g2_nor2_1 _7904_ (.A(net153),
    .B(net1341),
    .Y(_3883_));
 sg13g2_a21oi_1 _7905_ (.A1(net1341),
    .A2(_3734_),
    .Y(_0472_),
    .B1(_3883_));
 sg13g2_mux2_1 _7906_ (.A0(net343),
    .A1(_3739_),
    .S(net1340),
    .X(_0473_));
 sg13g2_mux2_1 _7907_ (.A0(net417),
    .A1(_3744_),
    .S(net1342),
    .X(_0474_));
 sg13g2_mux2_1 _7908_ (.A0(net438),
    .A1(_3749_),
    .S(net1341),
    .X(_0475_));
 sg13g2_nand2_1 _7909_ (.Y(_3884_),
    .A(net1342),
    .B(_3755_));
 sg13g2_o21ai_1 _7910_ (.B1(_3884_),
    .Y(_0476_),
    .A1(_0856_),
    .A2(net1342));
 sg13g2_mux2_1 _7911_ (.A0(net356),
    .A1(_3761_),
    .S(net1341),
    .X(_0477_));
 sg13g2_nand2_1 _7912_ (.Y(_3885_),
    .A(net1340),
    .B(_3767_));
 sg13g2_o21ai_1 _7913_ (.B1(_3885_),
    .Y(_0478_),
    .A1(_0860_),
    .A2(net1340));
 sg13g2_mux2_1 _7914_ (.A0(net390),
    .A1(_3773_),
    .S(net1340),
    .X(_0479_));
 sg13g2_mux2_1 _7915_ (.A0(net268),
    .A1(_3778_),
    .S(net1342),
    .X(_0480_));
 sg13g2_nand2_1 _7916_ (.Y(_3886_),
    .A(net1340),
    .B(_3784_));
 sg13g2_o21ai_1 _7917_ (.B1(_3886_),
    .Y(_0481_),
    .A1(_0862_),
    .A2(net1340));
 sg13g2_nor2_1 _7918_ (.A(net131),
    .B(net1337),
    .Y(_3887_));
 sg13g2_a21oi_1 _7919_ (.A1(net1337),
    .A2(_3792_),
    .Y(_0482_),
    .B1(_3887_));
 sg13g2_mux2_1 _7920_ (.A0(net411),
    .A1(_3797_),
    .S(net1340),
    .X(_0483_));
 sg13g2_nand2_1 _7921_ (.Y(_3888_),
    .A(net1338),
    .B(_3801_));
 sg13g2_o21ai_1 _7922_ (.B1(_3888_),
    .Y(_0484_),
    .A1(_0870_),
    .A2(net1338));
 sg13g2_mux2_1 _7923_ (.A0(net388),
    .A1(_3810_),
    .S(net1340),
    .X(_0485_));
 sg13g2_nor2_1 _7924_ (.A(net121),
    .B(net1337),
    .Y(_3889_));
 sg13g2_a21oi_1 _7925_ (.A1(net1337),
    .A2(_3817_),
    .Y(_0486_),
    .B1(_3889_));
 sg13g2_mux2_1 _7926_ (.A0(net370),
    .A1(_3823_),
    .S(net1338),
    .X(_0487_));
 sg13g2_nor2_1 _7927_ (.A(net222),
    .B(net1338),
    .Y(_3890_));
 sg13g2_a21oi_1 _7928_ (.A1(net1337),
    .A2(_3832_),
    .Y(_0488_),
    .B1(_3890_));
 sg13g2_mux2_1 _7929_ (.A0(net265),
    .A1(_3841_),
    .S(net1337),
    .X(_0489_));
 sg13g2_mux2_1 _7930_ (.A0(net301),
    .A1(_3849_),
    .S(net1342),
    .X(_0490_));
 sg13g2_mux2_1 _7931_ (.A0(net309),
    .A1(_3859_),
    .S(net1337),
    .X(_0491_));
 sg13g2_mux2_1 _7932_ (.A0(net286),
    .A1(_3863_),
    .S(net1342),
    .X(_0492_));
 sg13g2_mux2_1 _7933_ (.A0(net410),
    .A1(_3869_),
    .S(net1337),
    .X(_0493_));
 sg13g2_nor2_1 _7934_ (.A(net165),
    .B(net1339),
    .Y(_3891_));
 sg13g2_a21oi_1 _7935_ (.A1(net1339),
    .A2(_3875_),
    .Y(_0494_),
    .B1(_3891_));
 sg13g2_nor2_1 _7936_ (.A(net215),
    .B(net1339),
    .Y(_3892_));
 sg13g2_a21oi_1 _7937_ (.A1(net1339),
    .A2(_3880_),
    .Y(_0495_),
    .B1(_3892_));
 sg13g2_nor2_1 _7938_ (.A(net186),
    .B(net1347),
    .Y(_3893_));
 sg13g2_a21oi_1 _7939_ (.A1(net1349),
    .A2(_3734_),
    .Y(_0496_),
    .B1(_3893_));
 sg13g2_mux2_1 _7940_ (.A0(net287),
    .A1(_3739_),
    .S(net1347),
    .X(_0497_));
 sg13g2_mux2_1 _7941_ (.A0(net429),
    .A1(_3744_),
    .S(net1348),
    .X(_0498_));
 sg13g2_mux2_1 _7942_ (.A0(net351),
    .A1(_3749_),
    .S(net1348),
    .X(_0499_));
 sg13g2_nand2_1 _7943_ (.Y(_3894_),
    .A(net1348),
    .B(_3755_));
 sg13g2_o21ai_1 _7944_ (.B1(_3894_),
    .Y(_0500_),
    .A1(_0855_),
    .A2(net1348));
 sg13g2_mux2_1 _7945_ (.A0(net339),
    .A1(_3761_),
    .S(net1347),
    .X(_0501_));
 sg13g2_mux2_1 _7946_ (.A0(net395),
    .A1(_3767_),
    .S(net1347),
    .X(_0502_));
 sg13g2_mux2_1 _7947_ (.A0(net324),
    .A1(_3773_),
    .S(net1347),
    .X(_0503_));
 sg13g2_mux2_1 _7948_ (.A0(net331),
    .A1(_3778_),
    .S(net1348),
    .X(_0504_));
 sg13g2_mux2_1 _7949_ (.A0(net378),
    .A1(_3784_),
    .S(net1347),
    .X(_0505_));
 sg13g2_nor2_1 _7950_ (.A(net122),
    .B(net1344),
    .Y(_3895_));
 sg13g2_a21oi_1 _7951_ (.A1(net1344),
    .A2(_3792_),
    .Y(_0506_),
    .B1(_3895_));
 sg13g2_mux2_1 _7952_ (.A0(net403),
    .A1(_3797_),
    .S(net1347),
    .X(_0507_));
 sg13g2_mux2_1 _7953_ (.A0(net379),
    .A1(_3801_),
    .S(net1345),
    .X(_0508_));
 sg13g2_mux2_1 _7954_ (.A0(net304),
    .A1(_3810_),
    .S(net1347),
    .X(_0509_));
 sg13g2_nor2_1 _7955_ (.A(net160),
    .B(net1344),
    .Y(_3896_));
 sg13g2_a21oi_1 _7956_ (.A1(net1344),
    .A2(_3817_),
    .Y(_0510_),
    .B1(_3896_));
 sg13g2_mux2_1 _7957_ (.A0(net346),
    .A1(_3823_),
    .S(net1345),
    .X(_0511_));
 sg13g2_nor2_1 _7958_ (.A(net333),
    .B(net1345),
    .Y(_3897_));
 sg13g2_a21oi_1 _7959_ (.A1(net1344),
    .A2(_3832_),
    .Y(_0512_),
    .B1(_3897_));
 sg13g2_mux2_1 _7960_ (.A0(net377),
    .A1(_3841_),
    .S(net1344),
    .X(_0513_));
 sg13g2_mux2_1 _7961_ (.A0(net393),
    .A1(_3849_),
    .S(net1348),
    .X(_0514_));
 sg13g2_mux2_1 _7962_ (.A0(net440),
    .A1(_3859_),
    .S(net1344),
    .X(_0515_));
 sg13g2_mux2_1 _7963_ (.A0(net282),
    .A1(_3863_),
    .S(net1348),
    .X(_0516_));
 sg13g2_mux2_1 _7964_ (.A0(net316),
    .A1(_3869_),
    .S(net1344),
    .X(_0517_));
 sg13g2_nor2_1 _7965_ (.A(net219),
    .B(net1346),
    .Y(_3898_));
 sg13g2_a21oi_1 _7966_ (.A1(net1346),
    .A2(_3875_),
    .Y(_0518_),
    .B1(_3898_));
 sg13g2_nor2_1 _7967_ (.A(net126),
    .B(net1346),
    .Y(_3899_));
 sg13g2_a21oi_1 _7968_ (.A1(net1346),
    .A2(_3880_),
    .Y(_0519_),
    .B1(_3899_));
 sg13g2_nor2_1 _7969_ (.A(net1502),
    .B(_1018_),
    .Y(_3900_));
 sg13g2_xnor2_1 _7970_ (.Y(_3901_),
    .A(net1140),
    .B(net1256));
 sg13g2_a21oi_1 _7971_ (.A1(_1018_),
    .A2(_3901_),
    .Y(_0520_),
    .B1(_3900_));
 sg13g2_nor2b_1 _7972_ (.A(_1017_),
    .B_N(net1377),
    .Y(_3902_));
 sg13g2_or2_1 _7973_ (.X(_3903_),
    .B(_1728_),
    .A(_1724_));
 sg13g2_and3_1 _7974_ (.X(_3904_),
    .A(_1729_),
    .B(net1189),
    .C(_3903_));
 sg13g2_mux2_1 _7975_ (.A0(net298),
    .A1(_3904_),
    .S(net1330),
    .X(_0521_));
 sg13g2_xor2_1 _7976_ (.B(_1730_),
    .A(_1729_),
    .X(_3905_));
 sg13g2_and2_1 _7977_ (.A(net1189),
    .B(_3905_),
    .X(_3906_));
 sg13g2_mux2_1 _7978_ (.A0(net397),
    .A1(_3906_),
    .S(net1330),
    .X(_0522_));
 sg13g2_nor2_1 _7979_ (.A(net192),
    .B(net1328),
    .Y(_3907_));
 sg13g2_xor2_1 _7980_ (.B(_1733_),
    .A(_1731_),
    .X(_3908_));
 sg13g2_nand2b_1 _7981_ (.Y(_3909_),
    .B(_1782_),
    .A_N(_3908_));
 sg13g2_a21oi_1 _7982_ (.A1(net1328),
    .A2(_3909_),
    .Y(_0523_),
    .B1(_3907_));
 sg13g2_nand2b_1 _7983_ (.Y(_3910_),
    .B(_1734_),
    .A_N(_1736_));
 sg13g2_nand3_1 _7984_ (.B(net1189),
    .C(_3910_),
    .A(_1737_),
    .Y(_3911_));
 sg13g2_nor2_1 _7985_ (.A(net189),
    .B(net1327),
    .Y(_3912_));
 sg13g2_a21oi_1 _7986_ (.A1(net1327),
    .A2(_3911_),
    .Y(_0524_),
    .B1(_3912_));
 sg13g2_nor2_1 _7987_ (.A(net170),
    .B(net1327),
    .Y(_3913_));
 sg13g2_xnor2_1 _7988_ (.Y(_3914_),
    .A(_1738_),
    .B(_1740_));
 sg13g2_nand2_1 _7989_ (.Y(_3915_),
    .A(net1189),
    .B(_3914_));
 sg13g2_a21oi_1 _7990_ (.A1(net1327),
    .A2(_3915_),
    .Y(_0525_),
    .B1(_3913_));
 sg13g2_nand2b_1 _7991_ (.Y(_3916_),
    .B(_1741_),
    .A_N(_1743_));
 sg13g2_nand3_1 _7992_ (.B(net1189),
    .C(_3916_),
    .A(_1744_),
    .Y(_3917_));
 sg13g2_nor2_1 _7993_ (.A(net202),
    .B(net1327),
    .Y(_3918_));
 sg13g2_a21oi_1 _7994_ (.A1(net1327),
    .A2(_3917_),
    .Y(_0526_),
    .B1(_3918_));
 sg13g2_xnor2_1 _7995_ (.Y(_3919_),
    .A(_1745_),
    .B(_1746_));
 sg13g2_nand2_1 _7996_ (.Y(_3920_),
    .A(net1189),
    .B(_3919_));
 sg13g2_nor2_1 _7997_ (.A(net151),
    .B(net1328),
    .Y(_3921_));
 sg13g2_a21oi_1 _7998_ (.A1(net1328),
    .A2(_3920_),
    .Y(_0527_),
    .B1(_3921_));
 sg13g2_nor2_1 _7999_ (.A(net191),
    .B(net1329),
    .Y(_3922_));
 sg13g2_a21oi_1 _8000_ (.A1(_1833_),
    .A2(net1329),
    .Y(_0528_),
    .B1(_3922_));
 sg13g2_nor2_1 _8001_ (.A(net156),
    .B(net1322),
    .Y(_3923_));
 sg13g2_a21oi_1 _8002_ (.A1(_1828_),
    .A2(net1322),
    .Y(_0529_),
    .B1(_3923_));
 sg13g2_nor2_1 _8003_ (.A(net228),
    .B(net1322),
    .Y(_3924_));
 sg13g2_a21oi_1 _8004_ (.A1(_1842_),
    .A2(net1322),
    .Y(_0530_),
    .B1(_3924_));
 sg13g2_mux2_1 _8005_ (.A0(net445),
    .A1(_1822_),
    .S(net1323),
    .X(_0531_));
 sg13g2_nor2_1 _8006_ (.A(net171),
    .B(net1325),
    .Y(_3925_));
 sg13g2_a21oi_1 _8007_ (.A1(_1816_),
    .A2(net1325),
    .Y(_0532_),
    .B1(_3925_));
 sg13g2_nor2_1 _8008_ (.A(net127),
    .B(net1320),
    .Y(_3926_));
 sg13g2_a21oi_1 _8009_ (.A1(_1810_),
    .A2(net1320),
    .Y(_0533_),
    .B1(_3926_));
 sg13g2_nor2_1 _8010_ (.A(net327),
    .B(net1324),
    .Y(_3927_));
 sg13g2_a21oi_1 _8011_ (.A1(_1804_),
    .A2(net1324),
    .Y(_0534_),
    .B1(_3927_));
 sg13g2_nor2_1 _8012_ (.A(net261),
    .B(net1325),
    .Y(_3928_));
 sg13g2_a21oi_1 _8013_ (.A1(_1797_),
    .A2(net1325),
    .Y(_0535_),
    .B1(_3928_));
 sg13g2_nor2_1 _8014_ (.A(net128),
    .B(net1324),
    .Y(_3929_));
 sg13g2_a21oi_1 _8015_ (.A1(_1794_),
    .A2(net1324),
    .Y(_0536_),
    .B1(_3929_));
 sg13g2_mux2_1 _8016_ (.A0(net297),
    .A1(_1785_),
    .S(net1324),
    .X(_0537_));
 sg13g2_nor2_1 _8017_ (.A(net164),
    .B(net1322),
    .Y(_3930_));
 sg13g2_a21oi_1 _8018_ (.A1(_1874_),
    .A2(net1322),
    .Y(_0538_),
    .B1(_3930_));
 sg13g2_nor2_2 _8019_ (.A(_1017_),
    .B(net1390),
    .Y(_3931_));
 sg13g2_mux2_1 _8020_ (.A0(net457),
    .A1(_3904_),
    .S(net1319),
    .X(_0539_));
 sg13g2_nand2_1 _8021_ (.Y(_3932_),
    .A(_3906_),
    .B(net1319));
 sg13g2_o21ai_1 _8022_ (.B1(_3932_),
    .Y(_0540_),
    .A1(_0906_),
    .A2(net1319));
 sg13g2_nor2_1 _8023_ (.A(net149),
    .B(net1317),
    .Y(_3933_));
 sg13g2_a21oi_1 _8024_ (.A1(_3909_),
    .A2(net1317),
    .Y(_0541_),
    .B1(_3933_));
 sg13g2_nor2_1 _8025_ (.A(net159),
    .B(net1316),
    .Y(_3934_));
 sg13g2_a21oi_1 _8026_ (.A1(_3911_),
    .A2(net1316),
    .Y(_0542_),
    .B1(_3934_));
 sg13g2_nor2_1 _8027_ (.A(net248),
    .B(net1316),
    .Y(_3935_));
 sg13g2_a21oi_1 _8028_ (.A1(_3915_),
    .A2(net1316),
    .Y(_0543_),
    .B1(_3935_));
 sg13g2_nor2_1 _8029_ (.A(net204),
    .B(net1316),
    .Y(_3936_));
 sg13g2_a21oi_1 _8030_ (.A1(_3917_),
    .A2(net1316),
    .Y(_0544_),
    .B1(_3936_));
 sg13g2_nor2_1 _8031_ (.A(net183),
    .B(net1317),
    .Y(_3937_));
 sg13g2_a21oi_1 _8032_ (.A1(_3920_),
    .A2(net1317),
    .Y(_0545_),
    .B1(_3937_));
 sg13g2_nor2_1 _8033_ (.A(net190),
    .B(net1318),
    .Y(_3938_));
 sg13g2_a21oi_1 _8034_ (.A1(_1833_),
    .A2(net1315),
    .Y(_0546_),
    .B1(_3938_));
 sg13g2_nor2_1 _8035_ (.A(net155),
    .B(net1310),
    .Y(_3939_));
 sg13g2_a21oi_1 _8036_ (.A1(_1828_),
    .A2(net1311),
    .Y(_0547_),
    .B1(_3939_));
 sg13g2_nor2_1 _8037_ (.A(net196),
    .B(net1310),
    .Y(_3940_));
 sg13g2_a21oi_1 _8038_ (.A1(_1842_),
    .A2(net1310),
    .Y(_0548_),
    .B1(_3940_));
 sg13g2_nand2_1 _8039_ (.Y(_3941_),
    .A(_1822_),
    .B(net1311));
 sg13g2_o21ai_1 _8040_ (.B1(_3941_),
    .Y(_0549_),
    .A1(_0962_),
    .A2(net1311));
 sg13g2_nor2_1 _8041_ (.A(net145),
    .B(net1314),
    .Y(_3942_));
 sg13g2_a21oi_1 _8042_ (.A1(_1816_),
    .A2(net1314),
    .Y(_0550_),
    .B1(_3942_));
 sg13g2_nor2_1 _8043_ (.A(net158),
    .B(net1308),
    .Y(_3943_));
 sg13g2_a21oi_1 _8044_ (.A1(_1810_),
    .A2(net1308),
    .Y(_0551_),
    .B1(_3943_));
 sg13g2_nor2_1 _8045_ (.A(net135),
    .B(net1313),
    .Y(_3944_));
 sg13g2_a21oi_1 _8046_ (.A1(_1804_),
    .A2(net1313),
    .Y(_0552_),
    .B1(_3944_));
 sg13g2_nor2_1 _8047_ (.A(net162),
    .B(net1314),
    .Y(_3945_));
 sg13g2_a21oi_1 _8048_ (.A1(_1797_),
    .A2(net1314),
    .Y(_0553_),
    .B1(_3945_));
 sg13g2_nor2_1 _8049_ (.A(net173),
    .B(net1313),
    .Y(_3946_));
 sg13g2_a21oi_1 _8050_ (.A1(_1794_),
    .A2(net1313),
    .Y(_0554_),
    .B1(_3946_));
 sg13g2_mux2_1 _8051_ (.A0(net419),
    .A1(_1785_),
    .S(net1313),
    .X(_0555_));
 sg13g2_nor2_1 _8052_ (.A(net180),
    .B(net1310),
    .Y(_3947_));
 sg13g2_a21oi_1 _8053_ (.A1(_1874_),
    .A2(net1310),
    .Y(_0556_),
    .B1(_3947_));
 sg13g2_nor2_1 _8054_ (.A(net1413),
    .B(_1017_),
    .Y(_3948_));
 sg13g2_mux2_1 _8055_ (.A0(net340),
    .A1(_3904_),
    .S(net1307),
    .X(_0557_));
 sg13g2_nand2_1 _8056_ (.Y(_3949_),
    .A(_3906_),
    .B(net1307));
 sg13g2_o21ai_1 _8057_ (.B1(_3949_),
    .Y(_0558_),
    .A1(_0905_),
    .A2(net1304));
 sg13g2_nor2_1 _8058_ (.A(net199),
    .B(net1304),
    .Y(_3950_));
 sg13g2_a21oi_1 _8059_ (.A1(_3909_),
    .A2(net1305),
    .Y(_0559_),
    .B1(_3950_));
 sg13g2_nor2_1 _8060_ (.A(net152),
    .B(net1304),
    .Y(_3951_));
 sg13g2_a21oi_1 _8061_ (.A1(_3911_),
    .A2(net1304),
    .Y(_0560_),
    .B1(_3951_));
 sg13g2_nor2_1 _8062_ (.A(net157),
    .B(net1305),
    .Y(_3952_));
 sg13g2_a21oi_1 _8063_ (.A1(_3915_),
    .A2(net1305),
    .Y(_0561_),
    .B1(_3952_));
 sg13g2_nor2_1 _8064_ (.A(net134),
    .B(net1305),
    .Y(_3953_));
 sg13g2_a21oi_1 _8065_ (.A1(_3917_),
    .A2(net1305),
    .Y(_0562_),
    .B1(_3953_));
 sg13g2_nor2_1 _8066_ (.A(net236),
    .B(net1304),
    .Y(_3954_));
 sg13g2_a21oi_1 _8067_ (.A1(_3920_),
    .A2(net1304),
    .Y(_0563_),
    .B1(_3954_));
 sg13g2_nor2_1 _8068_ (.A(net197),
    .B(net1303),
    .Y(_3955_));
 sg13g2_a21oi_1 _8069_ (.A1(_1833_),
    .A2(net1303),
    .Y(_0564_),
    .B1(_3955_));
 sg13g2_nor2_1 _8070_ (.A(net168),
    .B(net1297),
    .Y(_3956_));
 sg13g2_a21oi_1 _8071_ (.A1(_1828_),
    .A2(net1297),
    .Y(_0565_),
    .B1(_3956_));
 sg13g2_nor2_1 _8072_ (.A(net250),
    .B(net1297),
    .Y(_3957_));
 sg13g2_a21oi_1 _8073_ (.A1(_1842_),
    .A2(net1297),
    .Y(_0566_),
    .B1(_3957_));
 sg13g2_nand2_1 _8074_ (.Y(_3958_),
    .A(_1822_),
    .B(net1298));
 sg13g2_o21ai_1 _8075_ (.B1(_3958_),
    .Y(_0567_),
    .A1(_0961_),
    .A2(net1298));
 sg13g2_nor2_1 _8076_ (.A(net146),
    .B(net1302),
    .Y(_3959_));
 sg13g2_a21oi_1 _8077_ (.A1(_1816_),
    .A2(net1302),
    .Y(_0568_),
    .B1(_3959_));
 sg13g2_nor2_1 _8078_ (.A(net227),
    .B(net1300),
    .Y(_3960_));
 sg13g2_a21oi_1 _8079_ (.A1(_1810_),
    .A2(net1300),
    .Y(_0569_),
    .B1(_3960_));
 sg13g2_nor2_1 _8080_ (.A(net232),
    .B(net1300),
    .Y(_3961_));
 sg13g2_a21oi_1 _8081_ (.A1(_1804_),
    .A2(net1300),
    .Y(_0570_),
    .B1(_3961_));
 sg13g2_nor2_1 _8082_ (.A(net140),
    .B(net1301),
    .Y(_3962_));
 sg13g2_a21oi_1 _8083_ (.A1(_1797_),
    .A2(net1301),
    .Y(_0571_),
    .B1(_3962_));
 sg13g2_nor2_1 _8084_ (.A(net174),
    .B(net1300),
    .Y(_3963_));
 sg13g2_a21oi_1 _8085_ (.A1(_1794_),
    .A2(net1301),
    .Y(_0572_),
    .B1(_3963_));
 sg13g2_mux2_1 _8086_ (.A0(net303),
    .A1(_1785_),
    .S(net1301),
    .X(_0573_));
 sg13g2_nor2_1 _8087_ (.A(net150),
    .B(net1297),
    .Y(_3964_));
 sg13g2_a21oi_1 _8088_ (.A1(_1874_),
    .A2(net1297),
    .Y(_0574_),
    .B1(_3964_));
 sg13g2_nand3_1 _8089_ (.B(_1840_),
    .C(_1841_),
    .A(_1669_),
    .Y(_3965_));
 sg13g2_and2_1 _8090_ (.A(_0089_),
    .B(net1395),
    .X(_3966_));
 sg13g2_a221oi_1 _8091_ (.B2(_0066_),
    .C1(_3966_),
    .B1(net1374),
    .A1(_0112_),
    .Y(_3967_),
    .A2(net1417));
 sg13g2_a22oi_1 _8092_ (.Y(_3968_),
    .B1(net1395),
    .B2(_0084_),
    .A2(net1418),
    .A1(_0107_));
 sg13g2_o21ai_1 _8093_ (.B1(_3968_),
    .Y(_3969_),
    .A1(_0837_),
    .A2(net1367));
 sg13g2_xor2_1 _8094_ (.B(_3969_),
    .A(_3967_),
    .X(_3970_));
 sg13g2_nor2_1 _8095_ (.A(net1149),
    .B(_3970_),
    .Y(_3971_));
 sg13g2_a21oi_1 _8096_ (.A1(_2239_),
    .A2(net1150),
    .Y(_3972_),
    .B1(_3971_));
 sg13g2_mux2_1 _8097_ (.A0(net420),
    .A1(_3972_),
    .S(net1326),
    .X(_0575_));
 sg13g2_nor2_1 _8098_ (.A(_0045_),
    .B(net1365),
    .Y(_3973_));
 sg13g2_nor2_1 _8099_ (.A(_0068_),
    .B(net1386),
    .Y(_3974_));
 sg13g2_nor2_1 _8100_ (.A(_0091_),
    .B(net1407),
    .Y(_3975_));
 sg13g2_nor3_1 _8101_ (.A(_3973_),
    .B(_3974_),
    .C(_3975_),
    .Y(_3976_));
 sg13g2_nand2_1 _8102_ (.Y(_3977_),
    .A(net1147),
    .B(_3976_));
 sg13g2_o21ai_1 _8103_ (.B1(_3977_),
    .Y(_3978_),
    .A1(_2239_),
    .A2(net1147));
 sg13g2_mux2_1 _8104_ (.A0(net415),
    .A1(_3978_),
    .S(net1322),
    .X(_0576_));
 sg13g2_nor2_1 _8105_ (.A(net1147),
    .B(_3976_),
    .Y(_3979_));
 sg13g2_a21oi_1 _8106_ (.A1(_2256_),
    .A2(net1147),
    .Y(_3980_),
    .B1(_3979_));
 sg13g2_mux2_1 _8107_ (.A0(net382),
    .A1(_3980_),
    .S(net1320),
    .X(_0577_));
 sg13g2_nor2_1 _8108_ (.A(_0047_),
    .B(net1364),
    .Y(_3981_));
 sg13g2_nor2_1 _8109_ (.A(_0070_),
    .B(net1385),
    .Y(_3982_));
 sg13g2_nor2_1 _8110_ (.A(_0093_),
    .B(net1406),
    .Y(_3983_));
 sg13g2_nor3_1 _8111_ (.A(_3981_),
    .B(_3982_),
    .C(_3983_),
    .Y(_3984_));
 sg13g2_nand2_1 _8112_ (.Y(_3985_),
    .A(net1146),
    .B(_3984_));
 sg13g2_o21ai_1 _8113_ (.B1(_3985_),
    .Y(_3986_),
    .A1(_2256_),
    .A2(net1146));
 sg13g2_mux2_1 _8114_ (.A0(net373),
    .A1(_3986_),
    .S(net1320),
    .X(_0578_));
 sg13g2_nor2_1 _8115_ (.A(_0048_),
    .B(net1364),
    .Y(_3987_));
 sg13g2_nor2_1 _8116_ (.A(_0071_),
    .B(net1385),
    .Y(_3988_));
 sg13g2_nor2_1 _8117_ (.A(_0094_),
    .B(net1406),
    .Y(_3989_));
 sg13g2_nor3_1 _8118_ (.A(_3987_),
    .B(_3988_),
    .C(_3989_),
    .Y(_3990_));
 sg13g2_mux2_1 _8119_ (.A0(_3984_),
    .A1(_3990_),
    .S(net1146),
    .X(_3991_));
 sg13g2_mux2_1 _8120_ (.A0(net294),
    .A1(_3991_),
    .S(net1320),
    .X(_0579_));
 sg13g2_mux2_1 _8121_ (.A0(_3990_),
    .A1(_2273_),
    .S(net1146),
    .X(_3992_));
 sg13g2_mux2_1 _8122_ (.A0(net450),
    .A1(_3992_),
    .S(net1320),
    .X(_0580_));
 sg13g2_nor2_1 _8123_ (.A(_0050_),
    .B(net1364),
    .Y(_3993_));
 sg13g2_nor2_1 _8124_ (.A(_0073_),
    .B(net1385),
    .Y(_3994_));
 sg13g2_nor2_1 _8125_ (.A(_0096_),
    .B(net1406),
    .Y(_3995_));
 sg13g2_nor3_1 _8126_ (.A(_3993_),
    .B(_3994_),
    .C(_3995_),
    .Y(_3996_));
 sg13g2_mux2_1 _8127_ (.A0(_2273_),
    .A1(_3996_),
    .S(net1146),
    .X(_3997_));
 sg13g2_mux2_1 _8128_ (.A0(net434),
    .A1(_3997_),
    .S(net1321),
    .X(_0581_));
 sg13g2_nor2_1 _8129_ (.A(_0051_),
    .B(net1364),
    .Y(_3998_));
 sg13g2_nor2_1 _8130_ (.A(_0074_),
    .B(net1385),
    .Y(_3999_));
 sg13g2_nor2_1 _8131_ (.A(_0097_),
    .B(net1406),
    .Y(_4000_));
 sg13g2_nor3_1 _8132_ (.A(_3998_),
    .B(_3999_),
    .C(_4000_),
    .Y(_4001_));
 sg13g2_mux2_1 _8133_ (.A0(_3996_),
    .A1(_4001_),
    .S(net1147),
    .X(_4002_));
 sg13g2_mux2_1 _8134_ (.A0(net345),
    .A1(_4002_),
    .S(net1321),
    .X(_0582_));
 sg13g2_nor2_1 _8135_ (.A(_0052_),
    .B(net1366),
    .Y(_4003_));
 sg13g2_nor2_1 _8136_ (.A(_0075_),
    .B(net1387),
    .Y(_4004_));
 sg13g2_nor2_1 _8137_ (.A(_0098_),
    .B(net1408),
    .Y(_4005_));
 sg13g2_nor3_1 _8138_ (.A(_4003_),
    .B(_4004_),
    .C(_4005_),
    .Y(_4006_));
 sg13g2_mux2_1 _8139_ (.A0(_4001_),
    .A1(_4006_),
    .S(net1148),
    .X(_4007_));
 sg13g2_mux2_1 _8140_ (.A0(net349),
    .A1(_4007_),
    .S(net1321),
    .X(_0583_));
 sg13g2_mux2_1 _8141_ (.A0(_4006_),
    .A1(_2294_),
    .S(net1148),
    .X(_4008_));
 sg13g2_mux2_1 _8142_ (.A0(net341),
    .A1(_4008_),
    .S(net1324),
    .X(_0584_));
 sg13g2_nor2_1 _8143_ (.A(_0054_),
    .B(net1366),
    .Y(_4009_));
 sg13g2_nor2_1 _8144_ (.A(_0077_),
    .B(net1387),
    .Y(_4010_));
 sg13g2_nor2_1 _8145_ (.A(_0100_),
    .B(net1408),
    .Y(_4011_));
 sg13g2_nor3_1 _8146_ (.A(_4009_),
    .B(_4010_),
    .C(_4011_),
    .Y(_4012_));
 sg13g2_mux2_1 _8147_ (.A0(_2294_),
    .A1(_4012_),
    .S(net1148),
    .X(_4013_));
 sg13g2_mux2_1 _8148_ (.A0(net336),
    .A1(_4013_),
    .S(net1324),
    .X(_0585_));
 sg13g2_mux2_1 _8149_ (.A0(_4012_),
    .A1(_2313_),
    .S(net1148),
    .X(_4014_));
 sg13g2_mux2_1 _8150_ (.A0(net326),
    .A1(_4014_),
    .S(net1324),
    .X(_0586_));
 sg13g2_nor2_1 _8151_ (.A(_0056_),
    .B(net1364),
    .Y(_4015_));
 sg13g2_nor2_1 _8152_ (.A(_0079_),
    .B(net1385),
    .Y(_4016_));
 sg13g2_nor2_1 _8153_ (.A(_0102_),
    .B(net1406),
    .Y(_4017_));
 sg13g2_nor3_1 _8154_ (.A(_4015_),
    .B(_4016_),
    .C(_4017_),
    .Y(_4018_));
 sg13g2_mux2_1 _8155_ (.A0(_2313_),
    .A1(_4018_),
    .S(net1146),
    .X(_4019_));
 sg13g2_mux2_1 _8156_ (.A0(net404),
    .A1(_4019_),
    .S(net1320),
    .X(_0587_));
 sg13g2_nor2_1 _8157_ (.A(_0057_),
    .B(net1365),
    .Y(_4020_));
 sg13g2_nor2_1 _8158_ (.A(_0080_),
    .B(net1385),
    .Y(_4021_));
 sg13g2_nor2_1 _8159_ (.A(_0103_),
    .B(net1406),
    .Y(_4022_));
 sg13g2_nor3_1 _8160_ (.A(_4020_),
    .B(_4021_),
    .C(_4022_),
    .Y(_4023_));
 sg13g2_mux2_1 _8161_ (.A0(_4018_),
    .A1(_4023_),
    .S(net1146),
    .X(_4024_));
 sg13g2_mux2_1 _8162_ (.A0(net401),
    .A1(_4024_),
    .S(net1321),
    .X(_0588_));
 sg13g2_mux2_1 _8163_ (.A0(_4023_),
    .A1(_2335_),
    .S(net1146),
    .X(_4025_));
 sg13g2_mux2_1 _8164_ (.A0(net317),
    .A1(_4025_),
    .S(net1320),
    .X(_0589_));
 sg13g2_nor2_1 _8165_ (.A(_0059_),
    .B(net1365),
    .Y(_4026_));
 sg13g2_nor2_1 _8166_ (.A(_0082_),
    .B(net1386),
    .Y(_4027_));
 sg13g2_nor2_1 _8167_ (.A(_0105_),
    .B(net1407),
    .Y(_4028_));
 sg13g2_nor3_1 _8168_ (.A(_4026_),
    .B(_4027_),
    .C(_4028_),
    .Y(_4029_));
 sg13g2_mux2_1 _8169_ (.A0(_2335_),
    .A1(_4029_),
    .S(net1150),
    .X(_4030_));
 sg13g2_mux2_1 _8170_ (.A0(net473),
    .A1(_4030_),
    .S(net1322),
    .X(_0590_));
 sg13g2_nor2_1 _8171_ (.A(_0060_),
    .B(net1367),
    .Y(_4031_));
 sg13g2_nor2_1 _8172_ (.A(_0083_),
    .B(net1388),
    .Y(_4032_));
 sg13g2_nor2_1 _8173_ (.A(_0106_),
    .B(net1410),
    .Y(_4033_));
 sg13g2_nor3_1 _8174_ (.A(_4031_),
    .B(_4032_),
    .C(_4033_),
    .Y(_4034_));
 sg13g2_mux2_1 _8175_ (.A0(_4029_),
    .A1(_4034_),
    .S(net1150),
    .X(_4035_));
 sg13g2_mux2_1 _8176_ (.A0(net344),
    .A1(_4035_),
    .S(net1326),
    .X(_0591_));
 sg13g2_mux2_1 _8177_ (.A0(_4034_),
    .A1(_3969_),
    .S(net1149),
    .X(_4036_));
 sg13g2_nand2_1 _8178_ (.Y(_4037_),
    .A(net1326),
    .B(_4036_));
 sg13g2_o21ai_1 _8179_ (.B1(_4037_),
    .Y(_0592_),
    .A1(_0837_),
    .A2(net1326));
 sg13g2_nor2_1 _8180_ (.A(net1149),
    .B(_3969_),
    .Y(_4038_));
 sg13g2_a21oi_1 _8181_ (.A1(_2352_),
    .A2(net1150),
    .Y(_4039_),
    .B1(_4038_));
 sg13g2_mux2_1 _8182_ (.A0(net342),
    .A1(_4039_),
    .S(net1328),
    .X(_0593_));
 sg13g2_nor2_1 _8183_ (.A(_0063_),
    .B(net1368),
    .Y(_4040_));
 sg13g2_nor2_1 _8184_ (.A(_0086_),
    .B(net1388),
    .Y(_4041_));
 sg13g2_nor2_1 _8185_ (.A(_0109_),
    .B(net1411),
    .Y(_4042_));
 sg13g2_nor3_1 _8186_ (.A(_4040_),
    .B(_4041_),
    .C(_4042_),
    .Y(_4043_));
 sg13g2_nand2_1 _8187_ (.Y(_4044_),
    .A(net1149),
    .B(_4043_));
 sg13g2_o21ai_1 _8188_ (.B1(_4044_),
    .Y(_4045_),
    .A1(_2352_),
    .A2(net1149));
 sg13g2_mux2_1 _8189_ (.A0(net414),
    .A1(_4045_),
    .S(net1327),
    .X(_0594_));
 sg13g2_mux2_1 _8190_ (.A0(_4043_),
    .A1(_2220_),
    .S(net1149),
    .X(_4046_));
 sg13g2_mux2_1 _8191_ (.A0(net387),
    .A1(_4046_),
    .S(net1327),
    .X(_0595_));
 sg13g2_nor2_1 _8192_ (.A(_0065_),
    .B(net1367),
    .Y(_4047_));
 sg13g2_nor2_1 _8193_ (.A(_0088_),
    .B(net1388),
    .Y(_4048_));
 sg13g2_nor2_1 _8194_ (.A(net1707),
    .B(net1410),
    .Y(_4049_));
 sg13g2_nor3_1 _8195_ (.A(_4047_),
    .B(_4048_),
    .C(_4049_),
    .Y(_4050_));
 sg13g2_mux2_1 _8196_ (.A0(_2220_),
    .A1(_4050_),
    .S(net1149),
    .X(_4051_));
 sg13g2_mux2_1 _8197_ (.A0(net329),
    .A1(_4051_),
    .S(net1326),
    .X(_0596_));
 sg13g2_nor2_1 _8198_ (.A(net1150),
    .B(_4050_),
    .Y(_4052_));
 sg13g2_a21oi_1 _8199_ (.A1(net1149),
    .A2(_3967_),
    .Y(_4053_),
    .B1(_4052_));
 sg13g2_mux2_1 _8200_ (.A0(net306),
    .A1(_4053_),
    .S(net1326),
    .X(_0597_));
 sg13g2_nand2_1 _8201_ (.Y(_4054_),
    .A(net1315),
    .B(_3972_));
 sg13g2_o21ai_1 _8202_ (.B1(_4054_),
    .Y(_0598_),
    .A1(_0836_),
    .A2(net1315));
 sg13g2_mux2_1 _8203_ (.A0(net292),
    .A1(_3978_),
    .S(net1310),
    .X(_0599_));
 sg13g2_nand2_1 _8204_ (.Y(_4055_),
    .A(net1308),
    .B(_3980_));
 sg13g2_o21ai_1 _8205_ (.B1(_4055_),
    .Y(_0600_),
    .A1(_0835_),
    .A2(net1310));
 sg13g2_mux2_1 _8206_ (.A0(net334),
    .A1(_3986_),
    .S(net1308),
    .X(_0601_));
 sg13g2_mux2_1 _8207_ (.A0(net348),
    .A1(_3991_),
    .S(net1308),
    .X(_0602_));
 sg13g2_mux2_1 _8208_ (.A0(net396),
    .A1(_3992_),
    .S(net1308),
    .X(_0603_));
 sg13g2_mux2_1 _8209_ (.A0(net312),
    .A1(_3997_),
    .S(net1309),
    .X(_0604_));
 sg13g2_mux2_1 _8210_ (.A0(net385),
    .A1(_4002_),
    .S(net1309),
    .X(_0605_));
 sg13g2_mux2_1 _8211_ (.A0(net456),
    .A1(_4007_),
    .S(net1309),
    .X(_0606_));
 sg13g2_mux2_1 _8212_ (.A0(net412),
    .A1(_4008_),
    .S(net1313),
    .X(_0607_));
 sg13g2_mux2_1 _8213_ (.A0(net408),
    .A1(_4013_),
    .S(net1313),
    .X(_0608_));
 sg13g2_mux2_1 _8214_ (.A0(net350),
    .A1(_4014_),
    .S(net1313),
    .X(_0609_));
 sg13g2_mux2_1 _8215_ (.A0(net293),
    .A1(_4019_),
    .S(net1308),
    .X(_0610_));
 sg13g2_mux2_1 _8216_ (.A0(net413),
    .A1(_4024_),
    .S(net1309),
    .X(_0611_));
 sg13g2_mux2_1 _8217_ (.A0(net364),
    .A1(_4025_),
    .S(net1308),
    .X(_0612_));
 sg13g2_mux2_1 _8218_ (.A0(net302),
    .A1(_4030_),
    .S(net1310),
    .X(_0613_));
 sg13g2_mux2_1 _8219_ (.A0(net355),
    .A1(_4035_),
    .S(net1315),
    .X(_0614_));
 sg13g2_mux2_1 _8220_ (.A0(net444),
    .A1(_4036_),
    .S(net1315),
    .X(_0615_));
 sg13g2_nand2_1 _8221_ (.Y(_4056_),
    .A(net1317),
    .B(_4039_));
 sg13g2_o21ai_1 _8222_ (.B1(_4056_),
    .Y(_0616_),
    .A1(_0834_),
    .A2(net1317));
 sg13g2_mux2_1 _8223_ (.A0(net416),
    .A1(_4045_),
    .S(net1316),
    .X(_0617_));
 sg13g2_mux2_1 _8224_ (.A0(net305),
    .A1(_4046_),
    .S(net1316),
    .X(_0618_));
 sg13g2_mux2_1 _8225_ (.A0(net398),
    .A1(_4051_),
    .S(net1315),
    .X(_0619_));
 sg13g2_mux2_1 _8226_ (.A0(net281),
    .A1(_4053_),
    .S(net1315),
    .X(_0620_));
 sg13g2_nand2_1 _8227_ (.Y(_4057_),
    .A(net1303),
    .B(_3972_));
 sg13g2_o21ai_1 _8228_ (.B1(_4057_),
    .Y(_0621_),
    .A1(_0833_),
    .A2(net1303));
 sg13g2_mux2_1 _8229_ (.A0(net321),
    .A1(_3978_),
    .S(net1297),
    .X(_0622_));
 sg13g2_nand2_1 _8230_ (.Y(_4058_),
    .A(net1296),
    .B(_3980_));
 sg13g2_o21ai_1 _8231_ (.B1(_4058_),
    .Y(_0623_),
    .A1(_0832_),
    .A2(net1296));
 sg13g2_mux2_1 _8232_ (.A0(net376),
    .A1(_3986_),
    .S(net1296),
    .X(_0624_));
 sg13g2_mux2_1 _8233_ (.A0(net426),
    .A1(_3991_),
    .S(net1296),
    .X(_0625_));
 sg13g2_mux2_1 _8234_ (.A0(net311),
    .A1(_3992_),
    .S(net1296),
    .X(_0626_));
 sg13g2_mux2_1 _8235_ (.A0(net421),
    .A1(_3997_),
    .S(net1299),
    .X(_0627_));
 sg13g2_mux2_1 _8236_ (.A0(net352),
    .A1(_4002_),
    .S(net1299),
    .X(_0628_));
 sg13g2_mux2_1 _8237_ (.A0(net295),
    .A1(_4007_),
    .S(net1299),
    .X(_0629_));
 sg13g2_mux2_1 _8238_ (.A0(net418),
    .A1(_4008_),
    .S(net1300),
    .X(_0630_));
 sg13g2_mux2_1 _8239_ (.A0(net315),
    .A1(_4013_),
    .S(net1300),
    .X(_0631_));
 sg13g2_mux2_1 _8240_ (.A0(net296),
    .A1(_4014_),
    .S(net1300),
    .X(_0632_));
 sg13g2_mux2_1 _8241_ (.A0(net405),
    .A1(_4019_),
    .S(net1296),
    .X(_0633_));
 sg13g2_mux2_1 _8242_ (.A0(net363),
    .A1(_4024_),
    .S(net1296),
    .X(_0634_));
 sg13g2_mux2_1 _8243_ (.A0(net323),
    .A1(_4025_),
    .S(net1296),
    .X(_0635_));
 sg13g2_mux2_1 _8244_ (.A0(net338),
    .A1(_4030_),
    .S(net1297),
    .X(_0636_));
 sg13g2_mux2_1 _8245_ (.A0(net384),
    .A1(_4035_),
    .S(net1303),
    .X(_0637_));
 sg13g2_mux2_1 _8246_ (.A0(net362),
    .A1(_4036_),
    .S(net1303),
    .X(_0638_));
 sg13g2_nand2_1 _8247_ (.Y(_4059_),
    .A(net1304),
    .B(_4039_));
 sg13g2_o21ai_1 _8248_ (.B1(_4059_),
    .Y(_0639_),
    .A1(_0831_),
    .A2(net1304));
 sg13g2_mux2_1 _8249_ (.A0(net300),
    .A1(_4045_),
    .S(net1305),
    .X(_0640_));
 sg13g2_mux2_1 _8250_ (.A0(net441),
    .A1(_4046_),
    .S(net1305),
    .X(_0641_));
 sg13g2_mux2_1 _8251_ (.A0(net354),
    .A1(_4051_),
    .S(net1303),
    .X(_0642_));
 sg13g2_mux2_1 _8252_ (.A0(net347),
    .A1(_4053_),
    .S(net1303),
    .X(_0643_));
 sg13g2_nor2_1 _8253_ (.A(net507),
    .B(net1323),
    .Y(_4060_));
 sg13g2_a21oi_1 _8254_ (.A1(_1869_),
    .A2(net1323),
    .Y(_0644_),
    .B1(_4060_));
 sg13g2_nor2_1 _8255_ (.A(net147),
    .B(net1326),
    .Y(_4061_));
 sg13g2_a21oi_1 _8256_ (.A1(_1865_),
    .A2(net1326),
    .Y(_0645_),
    .B1(_4061_));
 sg13g2_nor2_1 _8257_ (.A(net310),
    .B(net1311),
    .Y(_4062_));
 sg13g2_a21oi_1 _8258_ (.A1(_1869_),
    .A2(net1311),
    .Y(_0646_),
    .B1(_4062_));
 sg13g2_nor2_1 _8259_ (.A(net136),
    .B(net1318),
    .Y(_4063_));
 sg13g2_a21oi_1 _8260_ (.A1(_1865_),
    .A2(net1315),
    .Y(_0647_),
    .B1(_4063_));
 sg13g2_nand2_1 _8261_ (.Y(_4064_),
    .A(\tt6581_inst.accum_en ),
    .B(\tt6581_inst.accum_in_mux ));
 sg13g2_nand2_1 _8262_ (.Y(_4065_),
    .A(net1502),
    .B(_1075_));
 sg13g2_xnor2_1 _8263_ (.Y(_4066_),
    .A(\tt6581_inst.mult_inst.accum[8] ),
    .B(_4065_));
 sg13g2_nand2_1 _8264_ (.Y(_4067_),
    .A(\tt6581_inst.filter_accum[0] ),
    .B(_4066_));
 sg13g2_nor2_1 _8265_ (.A(_4064_),
    .B(_4067_),
    .Y(_4068_));
 sg13g2_a21oi_2 _8266_ (.B1(net124),
    .Y(_4069_),
    .A2(\tt6581_inst.accum_in_mux ),
    .A1(\tt6581_inst.accum_en ));
 sg13g2_inv_4 _8267_ (.A(_4069_),
    .Y(_4070_));
 sg13g2_a21oi_1 _8268_ (.A1(_4066_),
    .A2(_4070_),
    .Y(_4071_),
    .B1(\tt6581_inst.filter_accum[0] ));
 sg13g2_nor3_1 _8269_ (.A(net124),
    .B(_4068_),
    .C(_4071_),
    .Y(_0648_));
 sg13g2_o21ai_1 _8270_ (.B1(net1502),
    .Y(_4072_),
    .A1(\tt6581_inst.mult_inst.accum[8] ),
    .A2(_1075_));
 sg13g2_xnor2_1 _8271_ (.Y(_4073_),
    .A(_0910_),
    .B(_4072_));
 sg13g2_nor2_1 _8272_ (.A(_0990_),
    .B(_4073_),
    .Y(_4074_));
 sg13g2_xnor2_1 _8273_ (.Y(_4075_),
    .A(net955),
    .B(_4073_));
 sg13g2_nor2b_1 _8274_ (.A(_4067_),
    .B_N(_4075_),
    .Y(_4076_));
 sg13g2_a21oi_1 _8275_ (.A1(\tt6581_inst.filter_accum[0] ),
    .A2(_4066_),
    .Y(_4077_),
    .B1(_4075_));
 sg13g2_or2_1 _8276_ (.X(_4078_),
    .B(_4064_),
    .A(\tt6581_inst.accum_rst ));
 sg13g2_or3_1 _8277_ (.A(_4076_),
    .B(_4077_),
    .C(net1295),
    .X(_4079_));
 sg13g2_o21ai_1 _8278_ (.B1(_4079_),
    .Y(_0649_),
    .A1(_0990_),
    .A2(_4070_));
 sg13g2_or2_1 _8279_ (.X(_4080_),
    .B(_4076_),
    .A(_4074_));
 sg13g2_nand2_1 _8280_ (.Y(_4081_),
    .A(net1501),
    .B(_1076_));
 sg13g2_xnor2_1 _8281_ (.Y(_4082_),
    .A(_0911_),
    .B(_4081_));
 sg13g2_xnor2_1 _8282_ (.Y(_4083_),
    .A(net1536),
    .B(_4081_));
 sg13g2_xnor2_1 _8283_ (.Y(_4084_),
    .A(net1011),
    .B(_4082_));
 sg13g2_and2_1 _8284_ (.A(_4080_),
    .B(_4084_),
    .X(_4085_));
 sg13g2_nor2_1 _8285_ (.A(_4080_),
    .B(_4084_),
    .Y(_4086_));
 sg13g2_nor3_1 _8286_ (.A(net1295),
    .B(_4085_),
    .C(_4086_),
    .Y(_4087_));
 sg13g2_a21o_1 _8287_ (.A2(_4069_),
    .A1(net1011),
    .B1(_4087_),
    .X(_0650_));
 sg13g2_o21ai_1 _8288_ (.B1(net1502),
    .Y(_4088_),
    .A1(\tt6581_inst.mult_inst.accum[10] ),
    .A2(_1076_));
 sg13g2_xnor2_1 _8289_ (.Y(_4089_),
    .A(\tt6581_inst.mult_inst.accum[11] ),
    .B(_4088_));
 sg13g2_nand2_1 _8290_ (.Y(_4090_),
    .A(net1038),
    .B(_4089_));
 sg13g2_xnor2_1 _8291_ (.Y(_4091_),
    .A(net1038),
    .B(_4089_));
 sg13g2_a21oi_1 _8292_ (.A1(net1011),
    .A2(_4083_),
    .Y(_4092_),
    .B1(_4085_));
 sg13g2_or2_1 _8293_ (.X(_4093_),
    .B(_4092_),
    .A(_4091_));
 sg13g2_a21oi_1 _8294_ (.A1(_4091_),
    .A2(_4092_),
    .Y(_4094_),
    .B1(net1295));
 sg13g2_a22oi_1 _8295_ (.Y(_4095_),
    .B1(_4093_),
    .B2(_4094_),
    .A2(_4069_),
    .A1(net1038));
 sg13g2_inv_1 _8296_ (.Y(_0651_),
    .A(net1039));
 sg13g2_xnor2_1 _8297_ (.Y(_4096_),
    .A(net1087),
    .B(_1080_));
 sg13g2_a21oi_1 _8298_ (.A1(_4090_),
    .A2(_4093_),
    .Y(_4097_),
    .B1(_4096_));
 sg13g2_nand3_1 _8299_ (.B(_4093_),
    .C(_4096_),
    .A(_4090_),
    .Y(_4098_));
 sg13g2_nor2_1 _8300_ (.A(net1294),
    .B(_4097_),
    .Y(_4099_));
 sg13g2_a22oi_1 _8301_ (.Y(_4100_),
    .B1(_4098_),
    .B2(_4099_),
    .A2(_4069_),
    .A1(net1087));
 sg13g2_inv_1 _8302_ (.Y(_0652_),
    .A(net1088));
 sg13g2_a21oi_1 _8303_ (.A1(\tt6581_inst.filter_accum[4] ),
    .A2(_1080_),
    .Y(_4101_),
    .B1(_4097_));
 sg13g2_nand2_1 _8304_ (.Y(_4102_),
    .A(\tt6581_inst.filter_accum[5] ),
    .B(net1191));
 sg13g2_xnor2_1 _8305_ (.Y(_4103_),
    .A(net1054),
    .B(_1090_));
 sg13g2_a21oi_1 _8306_ (.A1(_4101_),
    .A2(_4103_),
    .Y(_4104_),
    .B1(net1295));
 sg13g2_o21ai_1 _8307_ (.B1(_4104_),
    .Y(_4105_),
    .A1(_4101_),
    .A2(_4103_));
 sg13g2_o21ai_1 _8308_ (.B1(_4105_),
    .Y(_0653_),
    .A1(_0991_),
    .A2(_4070_));
 sg13g2_nand2_1 _8309_ (.Y(_4106_),
    .A(net474),
    .B(_4069_));
 sg13g2_xnor2_1 _8310_ (.Y(_4107_),
    .A(net474),
    .B(_1097_));
 sg13g2_nand2_1 _8311_ (.Y(_4108_),
    .A(_4101_),
    .B(_4102_));
 sg13g2_o21ai_1 _8312_ (.B1(_4108_),
    .Y(_4109_),
    .A1(\tt6581_inst.filter_accum[5] ),
    .A2(_1090_));
 sg13g2_nor2_1 _8313_ (.A(_4107_),
    .B(_4109_),
    .Y(_4110_));
 sg13g2_a21o_1 _8314_ (.A2(_4109_),
    .A1(_4107_),
    .B1(net1295),
    .X(_4111_));
 sg13g2_o21ai_1 _8315_ (.B1(net475),
    .Y(_0654_),
    .A1(_4110_),
    .A2(_4111_));
 sg13g2_nand2_1 _8316_ (.Y(_4112_),
    .A(net543),
    .B(_4069_));
 sg13g2_xnor2_1 _8317_ (.Y(_4113_),
    .A(net543),
    .B(net1185));
 sg13g2_a21oi_1 _8318_ (.A1(net474),
    .A2(_1097_),
    .Y(_4114_),
    .B1(_4110_));
 sg13g2_nor2_1 _8319_ (.A(_4113_),
    .B(_4114_),
    .Y(_4115_));
 sg13g2_a21o_1 _8320_ (.A2(_4114_),
    .A1(_4113_),
    .B1(net1294),
    .X(_4116_));
 sg13g2_o21ai_1 _8321_ (.B1(net544),
    .Y(_0655_),
    .A1(_4115_),
    .A2(_4116_));
 sg13g2_nand2_1 _8322_ (.Y(_4117_),
    .A(net608),
    .B(_4069_));
 sg13g2_xnor2_1 _8323_ (.Y(_4118_),
    .A(net608),
    .B(net1184));
 sg13g2_a21oi_1 _8324_ (.A1(net543),
    .A2(net1185),
    .Y(_4119_),
    .B1(_4115_));
 sg13g2_nor2_1 _8325_ (.A(_4118_),
    .B(_4119_),
    .Y(_4120_));
 sg13g2_a21o_1 _8326_ (.A2(_4119_),
    .A1(_4118_),
    .B1(net1294),
    .X(_4121_));
 sg13g2_o21ai_1 _8327_ (.B1(net609),
    .Y(_0656_),
    .A1(_4120_),
    .A2(_4121_));
 sg13g2_a21o_1 _8328_ (.A2(net1184),
    .A1(net608),
    .B1(_4120_),
    .X(_4122_));
 sg13g2_xnor2_1 _8329_ (.Y(_4123_),
    .A(_0992_),
    .B(net1182));
 sg13g2_a21oi_1 _8330_ (.A1(_4122_),
    .A2(_4123_),
    .Y(_4124_),
    .B1(net1294));
 sg13g2_o21ai_1 _8331_ (.B1(_4124_),
    .Y(_4125_),
    .A1(_4122_),
    .A2(_4123_));
 sg13g2_o21ai_1 _8332_ (.B1(_4125_),
    .Y(_0657_),
    .A1(_0992_),
    .A2(_4070_));
 sg13g2_nand2_1 _8333_ (.Y(_4126_),
    .A(net645),
    .B(_4069_));
 sg13g2_xnor2_1 _8334_ (.Y(_4127_),
    .A(net645),
    .B(net1173));
 sg13g2_a21o_1 _8335_ (.A2(net1182),
    .A1(\tt6581_inst.filter_accum[9] ),
    .B1(_4122_),
    .X(_4128_));
 sg13g2_o21ai_1 _8336_ (.B1(_4128_),
    .Y(_4129_),
    .A1(\tt6581_inst.filter_accum[9] ),
    .A2(net1182));
 sg13g2_nor2_1 _8337_ (.A(_4127_),
    .B(_4129_),
    .Y(_4130_));
 sg13g2_a21o_1 _8338_ (.A2(_4129_),
    .A1(_4127_),
    .B1(net1294),
    .X(_4131_));
 sg13g2_o21ai_1 _8339_ (.B1(net646),
    .Y(_0658_),
    .A1(_4130_),
    .A2(_4131_));
 sg13g2_a21o_1 _8340_ (.A2(net1173),
    .A1(net645),
    .B1(_4130_),
    .X(_4132_));
 sg13g2_xnor2_1 _8341_ (.Y(_4133_),
    .A(_0993_),
    .B(net1167));
 sg13g2_a21oi_1 _8342_ (.A1(_4132_),
    .A2(_4133_),
    .Y(_4134_),
    .B1(net1294));
 sg13g2_o21ai_1 _8343_ (.B1(_4134_),
    .Y(_4135_),
    .A1(_4132_),
    .A2(_4133_));
 sg13g2_o21ai_1 _8344_ (.B1(_4135_),
    .Y(_0659_),
    .A1(_0993_),
    .A2(_4070_));
 sg13g2_xnor2_1 _8345_ (.Y(_4136_),
    .A(net1019),
    .B(net1165));
 sg13g2_a21o_1 _8346_ (.A2(net1167),
    .A1(\tt6581_inst.filter_accum[11] ),
    .B1(_4132_),
    .X(_4137_));
 sg13g2_o21ai_1 _8347_ (.B1(_4137_),
    .Y(_4138_),
    .A1(\tt6581_inst.filter_accum[11] ),
    .A2(net1167));
 sg13g2_nor2_1 _8348_ (.A(_4136_),
    .B(_4138_),
    .Y(_4139_));
 sg13g2_a21oi_1 _8349_ (.A1(_4136_),
    .A2(_4138_),
    .Y(_4140_),
    .B1(net1294));
 sg13g2_nand2b_1 _8350_ (.Y(_4141_),
    .B(_4140_),
    .A_N(_4139_));
 sg13g2_o21ai_1 _8351_ (.B1(_4141_),
    .Y(_0660_),
    .A1(_0994_),
    .A2(_4070_));
 sg13g2_a21oi_1 _8352_ (.A1(net1019),
    .A2(net1165),
    .Y(_4142_),
    .B1(_4139_));
 sg13g2_xnor2_1 _8353_ (.Y(_4143_),
    .A(net1130),
    .B(_1187_));
 sg13g2_a21oi_1 _8354_ (.A1(_4142_),
    .A2(_4143_),
    .Y(_4144_),
    .B1(net1294));
 sg13g2_o21ai_1 _8355_ (.B1(_4144_),
    .Y(_4145_),
    .A1(_4142_),
    .A2(_4143_));
 sg13g2_o21ai_1 _8356_ (.B1(_4145_),
    .Y(_0661_),
    .A1(_0995_),
    .A2(_4070_));
 sg13g2_nand2_2 _8357_ (.Y(_4146_),
    .A(\tt6581_inst.reg_addr[4] ),
    .B(_1048_));
 sg13g2_nand3_1 _8358_ (.B(_1048_),
    .C(_1050_),
    .A(\tt6581_inst.reg_addr[4] ),
    .Y(_4147_));
 sg13g2_nor2_1 _8359_ (.A(_1047_),
    .B(_4147_),
    .Y(_4148_));
 sg13g2_and2_1 _8360_ (.A(net1445),
    .B(net1246),
    .X(_4149_));
 sg13g2_mux2_1 _8361_ (.A0(net1123),
    .A1(net1485),
    .S(net1207),
    .X(_0662_));
 sg13g2_nand2_1 _8362_ (.Y(_4150_),
    .A(net1483),
    .B(net1207));
 sg13g2_o21ai_1 _8363_ (.B1(_4150_),
    .Y(_0663_),
    .A1(_0919_),
    .A2(net1207));
 sg13g2_mux2_1 _8364_ (.A0(net965),
    .A1(net1476),
    .S(net1207),
    .X(_0664_));
 sg13g2_mux2_1 _8365_ (.A0(net593),
    .A1(net1471),
    .S(net1207),
    .X(_0665_));
 sg13g2_mux2_1 _8366_ (.A0(net873),
    .A1(net1468),
    .S(net1207),
    .X(_0666_));
 sg13g2_mux2_1 _8367_ (.A0(net764),
    .A1(net1464),
    .S(net1207),
    .X(_0667_));
 sg13g2_mux2_1 _8368_ (.A0(net322),
    .A1(net1457),
    .S(net1207),
    .X(_0668_));
 sg13g2_mux2_1 _8369_ (.A0(net357),
    .A1(net1454),
    .S(_4149_),
    .X(_0669_));
 sg13g2_nor2_1 _8370_ (.A(net389),
    .B(net1298),
    .Y(_4151_));
 sg13g2_a21oi_1 _8371_ (.A1(_1869_),
    .A2(net1298),
    .Y(_0670_),
    .B1(_4151_));
 sg13g2_nor2_1 _8372_ (.A(net141),
    .B(net1306),
    .Y(_4152_));
 sg13g2_a21oi_1 _8373_ (.A1(_1865_),
    .A2(net1306),
    .Y(_0671_),
    .B1(_4152_));
 sg13g2_nor3_2 _8374_ (.A(_1047_),
    .B(_1067_),
    .C(_4146_),
    .Y(_4153_));
 sg13g2_and2_1 _8375_ (.A(net1447),
    .B(net1245),
    .X(_4154_));
 sg13g2_mux2_1 _8376_ (.A0(net890),
    .A1(net1488),
    .S(_4154_),
    .X(_0672_));
 sg13g2_mux2_1 _8377_ (.A0(net772),
    .A1(net1483),
    .S(_4154_),
    .X(_0673_));
 sg13g2_mux2_1 _8378_ (.A0(net924),
    .A1(net1477),
    .S(_4154_),
    .X(_0674_));
 sg13g2_mux2_1 _8379_ (.A0(net795),
    .A1(net1471),
    .S(_4154_),
    .X(_0675_));
 sg13g2_mux2_1 _8380_ (.A0(net704),
    .A1(net1468),
    .S(_4154_),
    .X(_0676_));
 sg13g2_mux2_1 _8381_ (.A0(net810),
    .A1(net1465),
    .S(_4154_),
    .X(_0677_));
 sg13g2_mux2_1 _8382_ (.A0(net635),
    .A1(net1459),
    .S(_4154_),
    .X(_0678_));
 sg13g2_mux2_1 _8383_ (.A0(net969),
    .A1(net1455),
    .S(_4154_),
    .X(_0679_));
 sg13g2_nor2_1 _8384_ (.A(_1057_),
    .B(_1379_),
    .Y(_4155_));
 sg13g2_nand2_1 _8385_ (.Y(_4156_),
    .A(net1446),
    .B(net1244));
 sg13g2_mux2_1 _8386_ (.A0(net1486),
    .A1(net886),
    .S(net1206),
    .X(_0680_));
 sg13g2_nor2_1 _8387_ (.A(net1482),
    .B(net1205),
    .Y(_4157_));
 sg13g2_a21oi_1 _8388_ (.A1(_0904_),
    .A2(net1205),
    .Y(_0681_),
    .B1(_4157_));
 sg13g2_nor2_1 _8389_ (.A(net1479),
    .B(net1206),
    .Y(_4158_));
 sg13g2_a21oi_1 _8390_ (.A1(_0903_),
    .A2(net1206),
    .Y(_0682_),
    .B1(_4158_));
 sg13g2_nor2_1 _8391_ (.A(net1474),
    .B(net1206),
    .Y(_4159_));
 sg13g2_a21oi_1 _8392_ (.A1(_0902_),
    .A2(net1206),
    .Y(_0683_),
    .B1(_4159_));
 sg13g2_nor2_1 _8393_ (.A(net1466),
    .B(net1205),
    .Y(_4160_));
 sg13g2_a21oi_1 _8394_ (.A1(_0901_),
    .A2(net1205),
    .Y(_0684_),
    .B1(_4160_));
 sg13g2_nor2_1 _8395_ (.A(net1462),
    .B(net1205),
    .Y(_4161_));
 sg13g2_a21oi_1 _8396_ (.A1(_0900_),
    .A2(net1205),
    .Y(_0685_),
    .B1(_4161_));
 sg13g2_nor2_1 _8397_ (.A(net1458),
    .B(net1206),
    .Y(_4162_));
 sg13g2_a21oi_1 _8398_ (.A1(_0897_),
    .A2(net1206),
    .Y(_0686_),
    .B1(_4162_));
 sg13g2_nor2_1 _8399_ (.A(net1454),
    .B(net1205),
    .Y(_4163_));
 sg13g2_a21oi_1 _8400_ (.A1(_0896_),
    .A2(net1205),
    .Y(_0687_),
    .B1(_4163_));
 sg13g2_nor2_2 _8401_ (.A(_1066_),
    .B(_1379_),
    .Y(_4164_));
 sg13g2_nand2_1 _8402_ (.Y(_4165_),
    .A(net1445),
    .B(net1243));
 sg13g2_nor2_1 _8403_ (.A(net1485),
    .B(net1203),
    .Y(_4166_));
 sg13g2_a21oi_1 _8404_ (.A1(_0893_),
    .A2(net1203),
    .Y(_0688_),
    .B1(_4166_));
 sg13g2_nor2_1 _8405_ (.A(net1481),
    .B(net1203),
    .Y(_4167_));
 sg13g2_a21oi_1 _8406_ (.A1(_0890_),
    .A2(net1203),
    .Y(_0689_),
    .B1(_4167_));
 sg13g2_nor2_1 _8407_ (.A(net1476),
    .B(net1204),
    .Y(_4168_));
 sg13g2_a21oi_1 _8408_ (.A1(_0960_),
    .A2(net1204),
    .Y(_0690_),
    .B1(_4168_));
 sg13g2_nor2_1 _8409_ (.A(net1471),
    .B(net1204),
    .Y(_4169_));
 sg13g2_a21oi_1 _8410_ (.A1(_0957_),
    .A2(net1204),
    .Y(_0691_),
    .B1(_4169_));
 sg13g2_mux2_1 _8411_ (.A0(net1468),
    .A1(net1022),
    .S(net1203),
    .X(_0692_));
 sg13g2_mux2_1 _8412_ (.A0(net1463),
    .A1(net992),
    .S(net1203),
    .X(_0693_));
 sg13g2_mux2_1 _8413_ (.A0(net1458),
    .A1(net894),
    .S(net1203),
    .X(_0694_));
 sg13g2_mux2_1 _8414_ (.A0(net1453),
    .A1(net837),
    .S(net1203),
    .X(_0695_));
 sg13g2_nor3_1 _8415_ (.A(net1451),
    .B(net1449),
    .C(_4147_),
    .Y(_4170_));
 sg13g2_nand2_2 _8416_ (.Y(_4171_),
    .A(net1447),
    .B(net1242));
 sg13g2_mux2_1 _8417_ (.A0(net1488),
    .A1(net604),
    .S(_4171_),
    .X(_0696_));
 sg13g2_mux2_1 _8418_ (.A0(net1483),
    .A1(net742),
    .S(_4171_),
    .X(_0697_));
 sg13g2_mux2_1 _8419_ (.A0(net1476),
    .A1(net843),
    .S(_4171_),
    .X(_0698_));
 sg13g2_mux2_1 _8420_ (.A0(net1472),
    .A1(net623),
    .S(_4171_),
    .X(_0699_));
 sg13g2_mux2_1 _8421_ (.A0(net1469),
    .A1(net782),
    .S(_4171_),
    .X(_0700_));
 sg13g2_mux2_1 _8422_ (.A0(net1464),
    .A1(net726),
    .S(_4171_),
    .X(_0701_));
 sg13g2_mux2_1 _8423_ (.A0(net1459),
    .A1(net632),
    .S(_4171_),
    .X(_0702_));
 sg13g2_mux2_1 _8424_ (.A0(net1455),
    .A1(net683),
    .S(_4171_),
    .X(_0703_));
 sg13g2_nor4_1 _8425_ (.A(net1451),
    .B(net1449),
    .C(_1056_),
    .D(_4146_),
    .Y(_4172_));
 sg13g2_nand2_2 _8426_ (.Y(_4173_),
    .A(net1445),
    .B(net1241));
 sg13g2_nor2_1 _8427_ (.A(net1486),
    .B(net1202),
    .Y(_4174_));
 sg13g2_a21oi_1 _8428_ (.A1(_0969_),
    .A2(net1202),
    .Y(_0704_),
    .B1(_4174_));
 sg13g2_mux2_1 _8429_ (.A0(net1481),
    .A1(net1031),
    .S(net1202),
    .X(_0705_));
 sg13g2_mux2_1 _8430_ (.A0(net1478),
    .A1(net650),
    .S(_4173_),
    .X(_0706_));
 sg13g2_mux2_1 _8431_ (.A0(net1473),
    .A1(net655),
    .S(net1202),
    .X(_0707_));
 sg13g2_nor2_1 _8432_ (.A(net1466),
    .B(net1202),
    .Y(_4175_));
 sg13g2_a21oi_1 _8433_ (.A1(_0968_),
    .A2(net1202),
    .Y(_0708_),
    .B1(_4175_));
 sg13g2_mux2_1 _8434_ (.A0(net1462),
    .A1(net653),
    .S(net1202),
    .X(_0709_));
 sg13g2_nor2_1 _8435_ (.A(net1457),
    .B(_4173_),
    .Y(_4176_));
 sg13g2_a21oi_1 _8436_ (.A1(_0966_),
    .A2(_4173_),
    .Y(_0710_),
    .B1(_4176_));
 sg13g2_mux2_1 _8437_ (.A0(net1454),
    .A1(net681),
    .S(net1202),
    .X(_0711_));
 sg13g2_nor3_1 _8438_ (.A(_1047_),
    .B(_1056_),
    .C(_4146_),
    .Y(_4177_));
 sg13g2_and2_1 _8439_ (.A(net1447),
    .B(_4177_),
    .X(_4178_));
 sg13g2_mux2_1 _8440_ (.A0(net896),
    .A1(net1485),
    .S(_4178_),
    .X(_0712_));
 sg13g2_mux2_1 _8441_ (.A0(net885),
    .A1(net1481),
    .S(_4178_),
    .X(_0713_));
 sg13g2_mux2_1 _8442_ (.A0(net888),
    .A1(net1476),
    .S(_4178_),
    .X(_0714_));
 sg13g2_mux2_1 _8443_ (.A0(net587),
    .A1(net1471),
    .S(_4178_),
    .X(_0715_));
 sg13g2_mux2_1 _8444_ (.A0(net497),
    .A1(net1468),
    .S(_4178_),
    .X(_0716_));
 sg13g2_mux2_1 _8445_ (.A0(net361),
    .A1(net1464),
    .S(_4178_),
    .X(_0717_));
 sg13g2_mux2_1 _8446_ (.A0(net318),
    .A1(net1459),
    .S(_4178_),
    .X(_0718_));
 sg13g2_mux2_1 _8447_ (.A0(net319),
    .A1(net1455),
    .S(_4178_),
    .X(_0719_));
 sg13g2_nor3_1 _8448_ (.A(_1056_),
    .B(_1057_),
    .C(_4146_),
    .Y(_4179_));
 sg13g2_nand2_2 _8449_ (.Y(_4180_),
    .A(net1446),
    .B(net1239));
 sg13g2_mux2_1 _8450_ (.A0(net1487),
    .A1(net565),
    .S(_4180_),
    .X(_0720_));
 sg13g2_mux2_1 _8451_ (.A0(net1482),
    .A1(net905),
    .S(_4180_),
    .X(_0721_));
 sg13g2_mux2_1 _8452_ (.A0(net1478),
    .A1(net590),
    .S(_4180_),
    .X(_0722_));
 sg13g2_mux2_1 _8453_ (.A0(net1473),
    .A1(net467),
    .S(_4180_),
    .X(_0723_));
 sg13g2_mux2_1 _8454_ (.A0(net1467),
    .A1(net616),
    .S(_4180_),
    .X(_0724_));
 sg13g2_mux2_1 _8455_ (.A0(net1463),
    .A1(net981),
    .S(_4180_),
    .X(_0725_));
 sg13g2_mux2_1 _8456_ (.A0(net1461),
    .A1(net612),
    .S(_4180_),
    .X(_0726_));
 sg13g2_mux2_1 _8457_ (.A0(net1453),
    .A1(net750),
    .S(_4180_),
    .X(_0727_));
 sg13g2_nor3_1 _8458_ (.A(_1066_),
    .B(_1067_),
    .C(_4146_),
    .Y(_4181_));
 sg13g2_nand2_2 _8459_ (.Y(_4182_),
    .A(net1447),
    .B(net1238));
 sg13g2_mux2_1 _8460_ (.A0(net1487),
    .A1(net663),
    .S(_4182_),
    .X(_0728_));
 sg13g2_mux2_1 _8461_ (.A0(net1483),
    .A1(net769),
    .S(_4182_),
    .X(_0729_));
 sg13g2_mux2_1 _8462_ (.A0(net1480),
    .A1(net1003),
    .S(_4182_),
    .X(_0730_));
 sg13g2_mux2_1 _8463_ (.A0(net1472),
    .A1(net833),
    .S(_4182_),
    .X(_0731_));
 sg13g2_mux2_1 _8464_ (.A0(net1469),
    .A1(net859),
    .S(_4182_),
    .X(_0732_));
 sg13g2_mux2_1 _8465_ (.A0(net1464),
    .A1(net1000),
    .S(_4182_),
    .X(_0733_));
 sg13g2_mux2_1 _8466_ (.A0(net1459),
    .A1(net804),
    .S(_4182_),
    .X(_0734_));
 sg13g2_mux2_1 _8467_ (.A0(net1455),
    .A1(net730),
    .S(_4182_),
    .X(_0735_));
 sg13g2_nor3_1 _8468_ (.A(_1056_),
    .B(_1066_),
    .C(_4146_),
    .Y(_4183_));
 sg13g2_nand2_2 _8469_ (.Y(_4184_),
    .A(net1448),
    .B(net1237));
 sg13g2_mux2_1 _8470_ (.A0(net1488),
    .A1(net857),
    .S(net1201),
    .X(_0736_));
 sg13g2_mux2_1 _8471_ (.A0(net1484),
    .A1(net980),
    .S(net1201),
    .X(_0737_));
 sg13g2_mux2_1 _8472_ (.A0(net1479),
    .A1(net985),
    .S(net1201),
    .X(_0738_));
 sg13g2_mux2_1 _8473_ (.A0(net1474),
    .A1(net1062),
    .S(net1201),
    .X(_0739_));
 sg13g2_nor2_1 _8474_ (.A(net1470),
    .B(net1201),
    .Y(_4185_));
 sg13g2_a21oi_1 _8475_ (.A1(_0989_),
    .A2(net1201),
    .Y(_0740_),
    .B1(_4185_));
 sg13g2_mux2_1 _8476_ (.A0(net1465),
    .A1(net660),
    .S(_4184_),
    .X(_0741_));
 sg13g2_mux2_1 _8477_ (.A0(net1459),
    .A1(net784),
    .S(net1201),
    .X(_0742_));
 sg13g2_mux2_1 _8478_ (.A0(net1456),
    .A1(net898),
    .S(net1201),
    .X(_0743_));
 sg13g2_nor3_1 _8479_ (.A(_1057_),
    .B(_1067_),
    .C(_4146_),
    .Y(_4186_));
 sg13g2_nand2_2 _8480_ (.Y(_4187_),
    .A(net1447),
    .B(net1236));
 sg13g2_mux2_1 _8481_ (.A0(net1488),
    .A1(net915),
    .S(_4187_),
    .X(_0744_));
 sg13g2_mux2_1 _8482_ (.A0(net1483),
    .A1(net902),
    .S(_4187_),
    .X(_0745_));
 sg13g2_mux2_1 _8483_ (.A0(net1476),
    .A1(net978),
    .S(_4187_),
    .X(_0746_));
 sg13g2_mux2_1 _8484_ (.A0(net1472),
    .A1(net918),
    .S(_4187_),
    .X(_0747_));
 sg13g2_mux2_1 _8485_ (.A0(net1469),
    .A1(net699),
    .S(_4187_),
    .X(_0748_));
 sg13g2_mux2_1 _8486_ (.A0(net1464),
    .A1(net923),
    .S(_4187_),
    .X(_0749_));
 sg13g2_mux2_1 _8487_ (.A0(net1457),
    .A1(net736),
    .S(_4187_),
    .X(_0750_));
 sg13g2_mux2_1 _8488_ (.A0(net1455),
    .A1(net793),
    .S(_4187_),
    .X(_0751_));
 sg13g2_nor4_2 _8489_ (.A(net1451),
    .B(net1449),
    .C(_1067_),
    .Y(_4188_),
    .D(_4146_));
 sg13g2_nand2_2 _8490_ (.Y(_4189_),
    .A(net1448),
    .B(_4188_));
 sg13g2_mux2_1 _8491_ (.A0(net1487),
    .A1(net599),
    .S(net1200),
    .X(_0752_));
 sg13g2_mux2_1 _8492_ (.A0(net1484),
    .A1(net658),
    .S(net1200),
    .X(_0753_));
 sg13g2_mux2_1 _8493_ (.A0(net1480),
    .A1(net883),
    .S(net1200),
    .X(_0754_));
 sg13g2_mux2_1 _8494_ (.A0(net1474),
    .A1(net702),
    .S(net1200),
    .X(_0755_));
 sg13g2_nor2_1 _8495_ (.A(net1470),
    .B(net1200),
    .Y(_4190_));
 sg13g2_a21oi_1 _8496_ (.A1(_0875_),
    .A2(net1200),
    .Y(_0756_),
    .B1(_4190_));
 sg13g2_mux2_1 _8497_ (.A0(net1465),
    .A1(net1111),
    .S(net1200),
    .X(_0757_));
 sg13g2_mux2_1 _8498_ (.A0(net1460),
    .A1(net983),
    .S(net1200),
    .X(_0758_));
 sg13g2_mux2_1 _8499_ (.A0(net1455),
    .A1(net943),
    .S(_4189_),
    .X(_0759_));
 sg13g2_nor2_2 _8500_ (.A(_1057_),
    .B(_4147_),
    .Y(_4191_));
 sg13g2_nand2_2 _8501_ (.Y(_4192_),
    .A(net1447),
    .B(net1234));
 sg13g2_mux2_1 _8502_ (.A0(net1488),
    .A1(net651),
    .S(_4192_),
    .X(_0760_));
 sg13g2_mux2_1 _8503_ (.A0(net1483),
    .A1(net846),
    .S(_4192_),
    .X(_0761_));
 sg13g2_mux2_1 _8504_ (.A0(net1477),
    .A1(net839),
    .S(_4192_),
    .X(_0762_));
 sg13g2_mux2_1 _8505_ (.A0(net1472),
    .A1(net713),
    .S(_4192_),
    .X(_0763_));
 sg13g2_mux2_1 _8506_ (.A0(net1469),
    .A1(net984),
    .S(_4192_),
    .X(_0764_));
 sg13g2_mux2_1 _8507_ (.A0(net1465),
    .A1(net779),
    .S(_4192_),
    .X(_0765_));
 sg13g2_mux2_1 _8508_ (.A0(net1460),
    .A1(net732),
    .S(_4192_),
    .X(_0766_));
 sg13g2_mux2_1 _8509_ (.A0(net1456),
    .A1(net908),
    .S(_4192_),
    .X(_0767_));
 sg13g2_nor3_2 _8510_ (.A(_0877_),
    .B(_0878_),
    .C(_3065_),
    .Y(_4193_));
 sg13g2_mux2_1 _8511_ (.A0(net1485),
    .A1(net806),
    .S(net1199),
    .X(_0768_));
 sg13g2_mux2_1 _8512_ (.A0(net1484),
    .A1(net783),
    .S(net1199),
    .X(_0769_));
 sg13g2_mux2_1 _8513_ (.A0(net1479),
    .A1(net724),
    .S(_4193_),
    .X(_0770_));
 sg13g2_mux2_1 _8514_ (.A0(net1473),
    .A1(net771),
    .S(net1199),
    .X(_0771_));
 sg13g2_mux2_1 _8515_ (.A0(net1467),
    .A1(net277),
    .S(net1199),
    .X(_0772_));
 sg13g2_mux2_1 _8516_ (.A0(net1462),
    .A1(net974),
    .S(net1199),
    .X(_0773_));
 sg13g2_mux2_1 _8517_ (.A0(net1458),
    .A1(net648),
    .S(net1199),
    .X(_0774_));
 sg13g2_mux2_1 _8518_ (.A0(net1454),
    .A1(net245),
    .S(net1199),
    .X(_0775_));
 sg13g2_mux2_1 _8519_ (.A0(net1452),
    .A1(net806),
    .S(net1214),
    .X(_0776_));
 sg13g2_mux2_1 _8520_ (.A0(net1450),
    .A1(net783),
    .S(net1214),
    .X(_0777_));
 sg13g2_mux2_1 _8521_ (.A0(net765),
    .A1(net724),
    .S(net1214),
    .X(_0778_));
 sg13g2_mux2_1 _8522_ (.A0(net812),
    .A1(net771),
    .S(net1214),
    .X(_0779_));
 sg13g2_nand2_1 _8523_ (.Y(_4194_),
    .A(net277),
    .B(net1214));
 sg13g2_o21ai_1 _8524_ (.B1(net278),
    .Y(_0780_),
    .A1(_0879_),
    .A2(net1214));
 sg13g2_mux2_1 _8525_ (.A0(net531),
    .A1(\tt6581_inst.spi_inst.shift_reg[4] ),
    .S(net1214),
    .X(_0781_));
 sg13g2_mux2_1 _8526_ (.A0(net509),
    .A1(\tt6581_inst.spi_inst.shift_reg[5] ),
    .S(net1214),
    .X(_0782_));
 sg13g2_nor2b_2 _8527_ (.A(net35),
    .B_N(\tt6581_inst.spi_inst.sclk_sync[2] ),
    .Y(_4195_));
 sg13g2_nor2b_2 _8528_ (.A(\tt6581_inst.spi_inst.cs_sync[1] ),
    .B_N(_4195_),
    .Y(_4196_));
 sg13g2_nand2b_2 _8529_ (.Y(_4197_),
    .B(_4195_),
    .A_N(\tt6581_inst.spi_inst.cs_sync[1] ));
 sg13g2_nand2_1 _8530_ (.Y(_4198_),
    .A(net177),
    .B(_4197_));
 sg13g2_a22oi_1 _8531_ (.Y(_4199_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[0] ),
    .A2(net1246),
    .A1(\tt6581_inst.filt_en_mode[0] ));
 sg13g2_nand2_1 _8532_ (.Y(_4200_),
    .A(\tt6581_inst.controller_inst.pw_hi_i[8] ),
    .B(net1274));
 sg13g2_a22oi_1 _8533_ (.Y(_4201_),
    .B1(net1239),
    .B2(\tt6581_inst.control_pack[16] ),
    .A2(net1275),
    .A1(\tt6581_inst.control_pack[0] ));
 sg13g2_a22oi_1 _8534_ (.Y(_4202_),
    .B1(net1237),
    .B2(\tt6581_inst.ad_pack[16] ),
    .A2(net1280),
    .A1(\tt6581_inst.controller_inst.sr_i[0] ));
 sg13g2_a22oi_1 _8535_ (.Y(_4203_),
    .B1(net1235),
    .B2(\tt6581_inst.controller_inst.sr_i[16] ),
    .A2(net1238),
    .A1(\tt6581_inst.filt_q_lo[0] ));
 sg13g2_a22oi_1 _8536_ (.Y(_4204_),
    .B1(net1236),
    .B2(\tt6581_inst.filt_f_hi[0] ),
    .A2(net1241),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[16] ));
 sg13g2_a22oi_1 _8537_ (.Y(_4205_),
    .B1(net1281),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[0] ),
    .A2(net1282),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[8] ));
 sg13g2_nand3_1 _8538_ (.B(_4204_),
    .C(_4205_),
    .A(_4203_),
    .Y(_4206_));
 sg13g2_a221oi_1 _8539_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[0] ),
    .C1(_4206_),
    .B1(_1397_),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[0] ),
    .Y(_4207_),
    .A2(net1285));
 sg13g2_a22oi_1 _8540_ (.Y(_4208_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[0] ),
    .A2(net1243),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[16] ));
 sg13g2_a22oi_1 _8541_ (.Y(_4209_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[0] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[0] ));
 sg13g2_a22oi_1 _8542_ (.Y(_4210_),
    .B1(net1279),
    .B2(\tt6581_inst.controller_inst.sr_i[8] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[8] ));
 sg13g2_nand4_1 _8543_ (.B(_4208_),
    .C(_4209_),
    .A(_4200_),
    .Y(_4211_),
    .D(_4210_));
 sg13g2_a22oi_1 _8544_ (.Y(_4212_),
    .B1(net1276),
    .B2(\tt6581_inst.control_pack[8] ),
    .A2(net1278),
    .A1(\tt6581_inst.ad_pack[8] ));
 sg13g2_a22oi_1 _8545_ (.Y(_4213_),
    .B1(net1244),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[16] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[8] ));
 sg13g2_nand3_1 _8546_ (.B(_4212_),
    .C(_4213_),
    .A(_4199_),
    .Y(_4214_));
 sg13g2_a221oi_1 _8547_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[16] ),
    .C1(_4214_),
    .B1(net1240),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[0] ),
    .Y(_4215_),
    .A2(net1283));
 sg13g2_nand4_1 _8548_ (.B(_4202_),
    .C(_4207_),
    .A(_4201_),
    .Y(_4216_),
    .D(_4215_));
 sg13g2_nor2_1 _8549_ (.A(net462),
    .B(net138),
    .Y(_4217_));
 sg13g2_nand2_1 _8550_ (.Y(_4218_),
    .A(_4195_),
    .B(_4217_));
 sg13g2_nor4_2 _8551_ (.A(\tt6581_inst.spi_inst.bit_cnt[2] ),
    .B(_0877_),
    .C(\tt6581_inst.spi_inst.is_write_cmd ),
    .Y(_4219_),
    .D(_4218_));
 sg13g2_o21ai_1 _8552_ (.B1(net1232),
    .Y(_4220_),
    .A1(_4211_),
    .A2(_4216_));
 sg13g2_o21ai_1 _8553_ (.B1(net178),
    .Y(_0783_),
    .A1(\tt6581_inst.spi_inst.cs_sync[1] ),
    .A2(_4220_));
 sg13g2_nand2_1 _8554_ (.Y(_4221_),
    .A(net117),
    .B(_4197_));
 sg13g2_nand2_1 _8555_ (.Y(_4222_),
    .A(\tt6581_inst.controller_inst.freq_lo_i[9] ),
    .B(_1068_));
 sg13g2_a22oi_1 _8556_ (.Y(_4223_),
    .B1(net1235),
    .B2(\tt6581_inst.controller_inst.sr_i[17] ),
    .A2(net1281),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[1] ));
 sg13g2_a22oi_1 _8557_ (.Y(_4224_),
    .B1(net1236),
    .B2(\tt6581_inst.filt_f_hi[1] ),
    .A2(net1280),
    .A1(\tt6581_inst.controller_inst.sr_i[1] ));
 sg13g2_a22oi_1 _8558_ (.Y(_4225_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[1] ),
    .A2(net1241),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[17] ));
 sg13g2_a22oi_1 _8559_ (.Y(_4226_),
    .B1(net1273),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[1] ),
    .A2(net1275),
    .A1(\tt6581_inst.control_pack[1] ));
 sg13g2_nand3_1 _8560_ (.B(_4225_),
    .C(_4226_),
    .A(_4224_),
    .Y(_4227_));
 sg13g2_a221oi_1 _8561_ (.B2(\tt6581_inst.ad_pack[17] ),
    .C1(_4227_),
    .B1(net1237),
    .A1(\tt6581_inst.control_pack[17] ),
    .Y(_4228_),
    .A2(net1239));
 sg13g2_a22oi_1 _8562_ (.Y(_4229_),
    .B1(net1283),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[1] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[9] ));
 sg13g2_a22oi_1 _8563_ (.Y(_4230_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[1] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[1] ));
 sg13g2_a22oi_1 _8564_ (.Y(_4231_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[1] ),
    .A2(net1278),
    .A1(\tt6581_inst.ad_pack[9] ));
 sg13g2_a22oi_1 _8565_ (.Y(_4232_),
    .B1(net1243),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[17] ),
    .A2(net1244),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[17] ));
 sg13g2_a22oi_1 _8566_ (.Y(_4233_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[1] ),
    .A2(_1380_),
    .A1(\tt6581_inst.controller_inst.sr_i[9] ));
 sg13g2_nand4_1 _8567_ (.B(_4231_),
    .C(_4232_),
    .A(_4230_),
    .Y(_4234_),
    .D(_4233_));
 sg13g2_a22oi_1 _8568_ (.Y(_4235_),
    .B1(net1274),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[9] ),
    .A2(net1285),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[1] ));
 sg13g2_a22oi_1 _8569_ (.Y(_4236_),
    .B1(net1276),
    .B2(\tt6581_inst.control_pack[9] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[9] ));
 sg13g2_nand4_1 _8570_ (.B(_4229_),
    .C(_4235_),
    .A(net1232),
    .Y(_4237_),
    .D(_4236_));
 sg13g2_a221oi_1 _8571_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[17] ),
    .C1(_4237_),
    .B1(net1240),
    .A1(\tt6581_inst.filt_en_mode[1] ),
    .Y(_4238_),
    .A2(net1246));
 sg13g2_nand4_1 _8572_ (.B(_4223_),
    .C(_4228_),
    .A(_4222_),
    .Y(_4239_),
    .D(_4238_));
 sg13g2_nor2_1 _8573_ (.A(_4234_),
    .B(_4239_),
    .Y(_4240_));
 sg13g2_o21ai_1 _8574_ (.B1(_4196_),
    .Y(_4241_),
    .A1(\tt6581_inst.spi_inst.data_out_reg[0] ),
    .A2(net1233));
 sg13g2_o21ai_1 _8575_ (.B1(net118),
    .Y(_0784_),
    .A1(_4240_),
    .A2(_4241_));
 sg13g2_nand2_1 _8576_ (.Y(_4242_),
    .A(net107),
    .B(_4197_));
 sg13g2_o21ai_1 _8577_ (.B1(_4196_),
    .Y(_4243_),
    .A1(\tt6581_inst.spi_inst.data_out_reg[1] ),
    .A2(net1233));
 sg13g2_a22oi_1 _8578_ (.Y(_4244_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[2] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[2] ));
 sg13g2_nand2_1 _8579_ (.Y(_4245_),
    .A(\tt6581_inst.controller_inst.sr_i[2] ),
    .B(net1280));
 sg13g2_a22oi_1 _8580_ (.Y(_4246_),
    .B1(net1279),
    .B2(\tt6581_inst.controller_inst.sr_i[10] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[10] ));
 sg13g2_a22oi_1 _8581_ (.Y(_4247_),
    .B1(net1237),
    .B2(\tt6581_inst.ad_pack[18] ),
    .A2(net1275),
    .A1(\tt6581_inst.control_pack[2] ));
 sg13g2_a22oi_1 _8582_ (.Y(_4248_),
    .B1(net1235),
    .B2(\tt6581_inst.controller_inst.sr_i[18] ),
    .A2(net1282),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[10] ));
 sg13g2_a22oi_1 _8583_ (.Y(_4249_),
    .B1(_4179_),
    .B2(\tt6581_inst.control_pack[18] ),
    .A2(_1071_),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[2] ));
 sg13g2_a22oi_1 _8584_ (.Y(_4250_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[2] ),
    .A2(net1241),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[18] ));
 sg13g2_nand3_1 _8585_ (.B(_4249_),
    .C(_4250_),
    .A(_4248_),
    .Y(_4251_));
 sg13g2_a221oi_1 _8586_ (.B2(\tt6581_inst.filt_f_hi[2] ),
    .C1(_4251_),
    .B1(net1236),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[2] ),
    .Y(_4252_),
    .A2(net1285));
 sg13g2_a22oi_1 _8587_ (.Y(_4253_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[2] ),
    .A2(_4164_),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[18] ));
 sg13g2_a22oi_1 _8588_ (.Y(_4254_),
    .B1(net1274),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[10] ),
    .A2(net1283),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[2] ));
 sg13g2_a22oi_1 _8589_ (.Y(_4255_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[18] ),
    .A2(_1060_),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[10] ));
 sg13g2_nand4_1 _8590_ (.B(_4253_),
    .C(_4254_),
    .A(_4246_),
    .Y(_4256_),
    .D(_4255_));
 sg13g2_a22oi_1 _8591_ (.Y(_4257_),
    .B1(net1273),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[2] ),
    .A2(net1278),
    .A1(\tt6581_inst.ad_pack[10] ));
 sg13g2_a22oi_1 _8592_ (.Y(_4258_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[2] ),
    .A2(net1246),
    .A1(\tt6581_inst.filt_en_mode[2] ));
 sg13g2_nand4_1 _8593_ (.B(_4244_),
    .C(_4257_),
    .A(net1232),
    .Y(_4259_),
    .D(_4258_));
 sg13g2_a221oi_1 _8594_ (.B2(\tt6581_inst.controller_inst.freq_lo_i[18] ),
    .C1(_4259_),
    .B1(_4155_),
    .A1(\tt6581_inst.control_pack[10] ),
    .Y(_4260_),
    .A2(_1386_));
 sg13g2_nand4_1 _8595_ (.B(_4247_),
    .C(_4252_),
    .A(_4245_),
    .Y(_4261_),
    .D(_4260_));
 sg13g2_nor2_1 _8596_ (.A(_4256_),
    .B(_4261_),
    .Y(_4262_));
 sg13g2_o21ai_1 _8597_ (.B1(net108),
    .Y(_0785_),
    .A1(_4243_),
    .A2(_4262_));
 sg13g2_nand2_1 _8598_ (.Y(_4263_),
    .A(net93),
    .B(_4197_));
 sg13g2_a22oi_1 _8599_ (.Y(_4264_),
    .B1(_1391_),
    .B2(\tt6581_inst.control_pack[3] ),
    .A2(net1285),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[3] ));
 sg13g2_nand2_1 _8600_ (.Y(_4265_),
    .A(\tt6581_inst.controller_inst.freq_lo_i[11] ),
    .B(net1282));
 sg13g2_a22oi_1 _8601_ (.Y(_4266_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[3] ),
    .A2(_1384_),
    .A1(\tt6581_inst.ad_pack[3] ));
 sg13g2_a22oi_1 _8602_ (.Y(_4267_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[19] ),
    .A2(net1283),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[3] ));
 sg13g2_a22oi_1 _8603_ (.Y(_4268_),
    .B1(net1279),
    .B2(\tt6581_inst.controller_inst.sr_i[11] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[11] ));
 sg13g2_a22oi_1 _8604_ (.Y(_4269_),
    .B1(_4181_),
    .B2(\tt6581_inst.filt_q_lo[3] ),
    .A2(net1241),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[19] ));
 sg13g2_a22oi_1 _8605_ (.Y(_4270_),
    .B1(net1280),
    .B2(\tt6581_inst.controller_inst.sr_i[3] ),
    .A2(net1281),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[3] ));
 sg13g2_a22oi_1 _8606_ (.Y(_4271_),
    .B1(net1235),
    .B2(\tt6581_inst.controller_inst.sr_i[19] ),
    .A2(net1273),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[3] ));
 sg13g2_nand3_1 _8607_ (.B(_4270_),
    .C(_4271_),
    .A(_4264_),
    .Y(_4272_));
 sg13g2_a221oi_1 _8608_ (.B2(\tt6581_inst.filt_f_hi[3] ),
    .C1(_4272_),
    .B1(net1236),
    .A1(\tt6581_inst.control_pack[19] ),
    .Y(_4273_),
    .A2(net1239));
 sg13g2_a22oi_1 _8609_ (.Y(_4274_),
    .B1(net1244),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[19] ),
    .A2(net1246),
    .A1(\tt6581_inst.controller_inst.filt_en_i[0] ));
 sg13g2_a22oi_1 _8610_ (.Y(_4275_),
    .B1(net1276),
    .B2(\tt6581_inst.control_pack[11] ),
    .A2(net1278),
    .A1(\tt6581_inst.ad_pack[11] ));
 sg13g2_a22oi_1 _8611_ (.Y(_4276_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[3] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[11] ));
 sg13g2_nand4_1 _8612_ (.B(_4274_),
    .C(_4275_),
    .A(_4266_),
    .Y(_4277_),
    .D(_4276_));
 sg13g2_a22oi_1 _8613_ (.Y(_4278_),
    .B1(net1237),
    .B2(\tt6581_inst.ad_pack[19] ),
    .A2(net1274),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[11] ));
 sg13g2_nand4_1 _8614_ (.B(_4267_),
    .C(_4268_),
    .A(net1232),
    .Y(_4279_),
    .D(_4278_));
 sg13g2_a221oi_1 _8615_ (.B2(\tt6581_inst.filt_volume[3] ),
    .C1(_4279_),
    .B1(net1234),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[19] ),
    .Y(_4280_),
    .A2(net1243));
 sg13g2_nand4_1 _8616_ (.B(_4269_),
    .C(_4273_),
    .A(_4265_),
    .Y(_4281_),
    .D(_4280_));
 sg13g2_nor2_1 _8617_ (.A(_4277_),
    .B(_4281_),
    .Y(_4282_));
 sg13g2_o21ai_1 _8618_ (.B1(_4196_),
    .Y(_4283_),
    .A1(\tt6581_inst.spi_inst.data_out_reg[2] ),
    .A2(net1233));
 sg13g2_o21ai_1 _8619_ (.B1(net94),
    .Y(_0786_),
    .A1(_4282_),
    .A2(_4283_));
 sg13g2_nand2_1 _8620_ (.Y(_4284_),
    .A(net97),
    .B(_4197_));
 sg13g2_nand2_1 _8621_ (.Y(_4285_),
    .A(\tt6581_inst.controller_inst.freq_lo_i[12] ),
    .B(net1282));
 sg13g2_a22oi_1 _8622_ (.Y(_4286_),
    .B1(net1246),
    .B2(\tt6581_inst.controller_inst.filt_en_i[1] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[4] ));
 sg13g2_a22oi_1 _8623_ (.Y(_4287_),
    .B1(net1244),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[20] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[12] ));
 sg13g2_a22oi_1 _8624_ (.Y(_4288_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[4] ),
    .A2(net1241),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[20] ));
 sg13g2_a22oi_1 _8625_ (.Y(_4289_),
    .B1(net1273),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[4] ),
    .A2(net1275),
    .A1(\tt6581_inst.control_pack[4] ));
 sg13g2_a22oi_1 _8626_ (.Y(_4290_),
    .B1(net1236),
    .B2(\tt6581_inst.filt_f_hi[4] ),
    .A2(net1237),
    .A1(\tt6581_inst.ad_pack[20] ));
 sg13g2_a22oi_1 _8627_ (.Y(_4291_),
    .B1(net1280),
    .B2(\tt6581_inst.controller_inst.sr_i[4] ),
    .A2(_1058_),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[4] ));
 sg13g2_nand3_1 _8628_ (.B(_4290_),
    .C(_4291_),
    .A(_4289_),
    .Y(_4292_));
 sg13g2_a221oi_1 _8629_ (.B2(\tt6581_inst.controller_inst.sr_i[20] ),
    .C1(_4292_),
    .B1(net1235),
    .A1(\tt6581_inst.control_pack[20] ),
    .Y(_4293_),
    .A2(net1239));
 sg13g2_nand3_1 _8630_ (.B(_4288_),
    .C(_4293_),
    .A(_4285_),
    .Y(_4294_));
 sg13g2_a22oi_1 _8631_ (.Y(_4295_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[4] ),
    .A2(net1274),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[12] ));
 sg13g2_a22oi_1 _8632_ (.Y(_4296_),
    .B1(net1278),
    .B2(\tt6581_inst.ad_pack[12] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[12] ));
 sg13g2_a22oi_1 _8633_ (.Y(_4297_),
    .B1(net1243),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[20] ),
    .A2(net1279),
    .A1(\tt6581_inst.controller_inst.sr_i[12] ));
 sg13g2_a22oi_1 _8634_ (.Y(_4298_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[20] ),
    .A2(_1064_),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[4] ));
 sg13g2_nand4_1 _8635_ (.B(_4296_),
    .C(_4297_),
    .A(_4295_),
    .Y(_4299_),
    .D(_4298_));
 sg13g2_a22oi_1 _8636_ (.Y(_4300_),
    .B1(net1276),
    .B2(\tt6581_inst.control_pack[12] ),
    .A2(net1281),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[4] ));
 sg13g2_nand2_1 _8637_ (.Y(_4301_),
    .A(net1232),
    .B(_4300_));
 sg13g2_a22oi_1 _8638_ (.Y(_4302_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[4] ),
    .A2(_4153_),
    .A1(\tt6581_inst.filt_f_lo[4] ));
 sg13g2_nand3_1 _8639_ (.B(_4287_),
    .C(_4302_),
    .A(_4286_),
    .Y(_4303_));
 sg13g2_nor4_1 _8640_ (.A(_4294_),
    .B(_4299_),
    .C(_4301_),
    .D(_4303_),
    .Y(_4304_));
 sg13g2_o21ai_1 _8641_ (.B1(_4196_),
    .Y(_4305_),
    .A1(net93),
    .A2(net1233));
 sg13g2_o21ai_1 _8642_ (.B1(net98),
    .Y(_0787_),
    .A1(_4304_),
    .A2(_4305_));
 sg13g2_nand2_1 _8643_ (.Y(_4306_),
    .A(net88),
    .B(_4197_));
 sg13g2_nand2_1 _8644_ (.Y(_4307_),
    .A(\tt6581_inst.controller_inst.freq_lo_i[13] ),
    .B(net1282));
 sg13g2_a22oi_1 _8645_ (.Y(_4308_),
    .B1(net1246),
    .B2(\tt6581_inst.controller_inst.filt_en_i[2] ),
    .A2(net1283),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[5] ));
 sg13g2_a22oi_1 _8646_ (.Y(_4309_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[5] ),
    .A2(_1382_),
    .A1(\tt6581_inst.ad_pack[13] ));
 sg13g2_a22oi_1 _8647_ (.Y(_4310_),
    .B1(net1236),
    .B2(\tt6581_inst.filt_f_hi[5] ),
    .A2(net1280),
    .A1(\tt6581_inst.controller_inst.sr_i[5] ));
 sg13g2_a22oi_1 _8648_ (.Y(_4311_),
    .B1(net1281),
    .B2(\tt6581_inst.controller_inst.freq_lo_i[5] ),
    .A2(net1285),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[5] ));
 sg13g2_a22oi_1 _8649_ (.Y(_4312_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[5] ),
    .A2(net1239),
    .A1(\tt6581_inst.control_pack[21] ));
 sg13g2_a22oi_1 _8650_ (.Y(_4313_),
    .B1(net1241),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[21] ),
    .A2(net1273),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[5] ));
 sg13g2_nand3_1 _8651_ (.B(_4312_),
    .C(_4313_),
    .A(_4311_),
    .Y(_4314_));
 sg13g2_a221oi_1 _8652_ (.B2(\tt6581_inst.controller_inst.sr_i[21] ),
    .C1(_4314_),
    .B1(net1235),
    .A1(\tt6581_inst.ad_pack[21] ),
    .Y(_4315_),
    .A2(net1237));
 sg13g2_a22oi_1 _8653_ (.Y(_4316_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[21] ),
    .A2(net1276),
    .A1(\tt6581_inst.control_pack[13] ));
 sg13g2_a22oi_1 _8654_ (.Y(_4317_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[5] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[5] ));
 sg13g2_a22oi_1 _8655_ (.Y(_4318_),
    .B1(net1243),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[21] ),
    .A2(net1279),
    .A1(\tt6581_inst.controller_inst.sr_i[13] ));
 sg13g2_a22oi_1 _8656_ (.Y(_4319_),
    .B1(net1242),
    .B2(\tt6581_inst.filt_q_hi[5] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[13] ));
 sg13g2_nand4_1 _8657_ (.B(_4317_),
    .C(_4318_),
    .A(_4316_),
    .Y(_4320_),
    .D(_4319_));
 sg13g2_a22oi_1 _8658_ (.Y(_4321_),
    .B1(net1275),
    .B2(\tt6581_inst.control_pack[5] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[13] ));
 sg13g2_nand4_1 _8659_ (.B(_4308_),
    .C(_4309_),
    .A(net1232),
    .Y(_4322_),
    .D(_4321_));
 sg13g2_a221oi_1 _8660_ (.B2(\tt6581_inst.controller_inst.freq_lo_i[21] ),
    .C1(_4322_),
    .B1(net1244),
    .A1(\tt6581_inst.controller_inst.pw_hi_i[13] ),
    .Y(_4323_),
    .A2(_1393_));
 sg13g2_nand4_1 _8661_ (.B(_4310_),
    .C(_4315_),
    .A(_4307_),
    .Y(_4324_),
    .D(_4323_));
 sg13g2_nor2_1 _8662_ (.A(_4320_),
    .B(_4324_),
    .Y(_4325_));
 sg13g2_o21ai_1 _8663_ (.B1(_4196_),
    .Y(_4326_),
    .A1(\tt6581_inst.spi_inst.data_out_reg[4] ),
    .A2(net1233));
 sg13g2_o21ai_1 _8664_ (.B1(net89),
    .Y(_0788_),
    .A1(_4325_),
    .A2(_4326_));
 sg13g2_nand2_1 _8665_ (.Y(_4327_),
    .A(net104),
    .B(_4197_));
 sg13g2_o21ai_1 _8666_ (.B1(_4196_),
    .Y(_4328_),
    .A1(net88),
    .A2(net1233));
 sg13g2_nand2_1 _8667_ (.Y(_4329_),
    .A(\tt6581_inst.controller_inst.freq_lo_i[14] ),
    .B(net1282));
 sg13g2_a22oi_1 _8668_ (.Y(_4330_),
    .B1(net1273),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[6] ),
    .A2(net1281),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[6] ));
 sg13g2_a22oi_1 _8669_ (.Y(_4331_),
    .B1(net1239),
    .B2(\tt6581_inst.control_pack[22] ),
    .A2(net1275),
    .A1(\tt6581_inst.control_pack[6] ));
 sg13g2_a22oi_1 _8670_ (.Y(_4332_),
    .B1(net1236),
    .B2(\tt6581_inst.filt_f_hi[6] ),
    .A2(net1285),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[6] ));
 sg13g2_a22oi_1 _8671_ (.Y(_4333_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[6] ),
    .A2(_4172_),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[22] ));
 sg13g2_nand3_1 _8672_ (.B(_4332_),
    .C(_4333_),
    .A(_4331_),
    .Y(_4334_));
 sg13g2_a221oi_1 _8673_ (.B2(\tt6581_inst.controller_inst.sr_i[22] ),
    .C1(_4334_),
    .B1(net1235),
    .A1(\tt6581_inst.controller_inst.sr_i[6] ),
    .Y(_4335_),
    .A2(net1280));
 sg13g2_a22oi_1 _8674_ (.Y(_4336_),
    .B1(net1245),
    .B2(\tt6581_inst.filt_f_lo[6] ),
    .A2(net1283),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[6] ));
 sg13g2_a22oi_1 _8675_ (.Y(_4337_),
    .B1(net1246),
    .B2(\tt6581_inst.filt_en_mode[6] ),
    .A2(_1052_),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[14] ));
 sg13g2_a22oi_1 _8676_ (.Y(_4338_),
    .B1(net1276),
    .B2(\tt6581_inst.control_pack[14] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[14] ));
 sg13g2_a22oi_1 _8677_ (.Y(_4339_),
    .B1(net1243),
    .B2(\tt6581_inst.controller_inst.freq_hi_i[22] ),
    .A2(net1278),
    .A1(\tt6581_inst.ad_pack[14] ));
 sg13g2_a22oi_1 _8678_ (.Y(_4340_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[22] ),
    .A2(net1242),
    .A1(\tt6581_inst.filt_q_hi[6] ));
 sg13g2_a22oi_1 _8679_ (.Y(_4341_),
    .B1(_4191_),
    .B2(\tt6581_inst.filt_volume[6] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[6] ));
 sg13g2_nand4_1 _8680_ (.B(_4339_),
    .C(_4340_),
    .A(_4338_),
    .Y(_4342_),
    .D(_4341_));
 sg13g2_a22oi_1 _8681_ (.Y(_4343_),
    .B1(net1237),
    .B2(\tt6581_inst.ad_pack[22] ),
    .A2(net1244),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[22] ));
 sg13g2_nand4_1 _8682_ (.B(_4336_),
    .C(_4337_),
    .A(net1232),
    .Y(_4344_),
    .D(_4343_));
 sg13g2_a221oi_1 _8683_ (.B2(\tt6581_inst.controller_inst.pw_hi_i[14] ),
    .C1(_4344_),
    .B1(net1274),
    .A1(\tt6581_inst.controller_inst.sr_i[14] ),
    .Y(_4345_),
    .A2(net1279));
 sg13g2_nand4_1 _8684_ (.B(_4330_),
    .C(_4335_),
    .A(_4329_),
    .Y(_4346_),
    .D(_4345_));
 sg13g2_nor2_1 _8685_ (.A(_4342_),
    .B(_4346_),
    .Y(_4347_));
 sg13g2_o21ai_1 _8686_ (.B1(net105),
    .Y(_0789_),
    .A1(_4328_),
    .A2(_4347_));
 sg13g2_nand2_1 _8687_ (.Y(_4348_),
    .A(net69),
    .B(_4197_));
 sg13g2_nand2_1 _8688_ (.Y(_4349_),
    .A(\tt6581_inst.controller_inst.pw_lo_i[7] ),
    .B(net1285));
 sg13g2_a22oi_1 _8689_ (.Y(_4350_),
    .B1(net1240),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[23] ),
    .A2(net1245),
    .A1(\tt6581_inst.filt_f_lo[7] ));
 sg13g2_a22oi_1 _8690_ (.Y(_4351_),
    .B1(_4170_),
    .B2(\tt6581_inst.filt_q_hi[7] ),
    .A2(net1277),
    .A1(\tt6581_inst.ad_pack[7] ));
 sg13g2_a22oi_1 _8691_ (.Y(_4352_),
    .B1(net1274),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[15] ),
    .A2(net1279),
    .A1(\tt6581_inst.controller_inst.sr_i[15] ));
 sg13g2_a22oi_1 _8692_ (.Y(_4353_),
    .B1(net1273),
    .B2(\tt6581_inst.controller_inst.pw_hi_i[7] ),
    .A2(net1282),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[15] ));
 sg13g2_a22oi_1 _8693_ (.Y(_4354_),
    .B1(_4186_),
    .B2(\tt6581_inst.filt_f_hi[7] ),
    .A2(net1281),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[7] ));
 sg13g2_a22oi_1 _8694_ (.Y(_4355_),
    .B1(net1235),
    .B2(\tt6581_inst.controller_inst.sr_i[23] ),
    .A2(_4183_),
    .A1(\tt6581_inst.ad_pack[23] ));
 sg13g2_a22oi_1 _8695_ (.Y(_4356_),
    .B1(net1238),
    .B2(\tt6581_inst.filt_q_lo[7] ),
    .A2(_1377_),
    .A1(\tt6581_inst.controller_inst.sr_i[7] ));
 sg13g2_nand3_1 _8696_ (.B(_4355_),
    .C(_4356_),
    .A(_4354_),
    .Y(_4357_));
 sg13g2_a221oi_1 _8697_ (.B2(\tt6581_inst.control_pack[23] ),
    .C1(_4357_),
    .B1(net1239),
    .A1(\tt6581_inst.control_pack[7] ),
    .Y(_4358_),
    .A2(net1275));
 sg13g2_a22oi_1 _8698_ (.Y(_4359_),
    .B1(net1234),
    .B2(\tt6581_inst.filt_volume[7] ),
    .A2(net1244),
    .A1(\tt6581_inst.controller_inst.freq_lo_i[23] ));
 sg13g2_a22oi_1 _8699_ (.Y(_4360_),
    .B1(_4148_),
    .B2(\tt6581_inst.filt_en_mode[7] ),
    .A2(net1286),
    .A1(\tt6581_inst.controller_inst.pw_lo_i[15] ));
 sg13g2_a22oi_1 _8700_ (.Y(_4361_),
    .B1(net1278),
    .B2(\tt6581_inst.ad_pack[15] ),
    .A2(net1284),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[15] ));
 sg13g2_nand4_1 _8701_ (.B(_4359_),
    .C(_4360_),
    .A(_4350_),
    .Y(_4362_),
    .D(_4361_));
 sg13g2_a22oi_1 _8702_ (.Y(_4363_),
    .B1(net1241),
    .B2(\tt6581_inst.controller_inst.pw_lo_i[23] ),
    .A2(net1276),
    .A1(\tt6581_inst.control_pack[15] ));
 sg13g2_nand4_1 _8703_ (.B(_4351_),
    .C(_4352_),
    .A(net1232),
    .Y(_4364_),
    .D(_4363_));
 sg13g2_a221oi_1 _8704_ (.B2(\tt6581_inst.controller_inst.freq_hi_i[23] ),
    .C1(_4364_),
    .B1(net1243),
    .A1(\tt6581_inst.controller_inst.freq_hi_i[7] ),
    .Y(_4365_),
    .A2(net1283));
 sg13g2_nand4_1 _8705_ (.B(_4353_),
    .C(_4358_),
    .A(_4349_),
    .Y(_4366_),
    .D(_4365_));
 sg13g2_nor2_1 _8706_ (.A(_4362_),
    .B(_4366_),
    .Y(_4367_));
 sg13g2_o21ai_1 _8707_ (.B1(_4196_),
    .Y(_4368_),
    .A1(\tt6581_inst.spi_inst.data_out_reg[6] ),
    .A2(net1233));
 sg13g2_o21ai_1 _8708_ (.B1(net70),
    .Y(_0790_),
    .A1(_4367_),
    .A2(_4368_));
 sg13g2_a21o_1 _8709_ (.A2(_3063_),
    .A1(net1446),
    .B1(net1199),
    .X(_0791_));
 sg13g2_a21oi_1 _8710_ (.A1(\tt6581_inst.spi_inst.bit_cnt[3] ),
    .A2(_3061_),
    .Y(_4369_),
    .B1(_3062_));
 sg13g2_nor2_1 _8711_ (.A(\tt6581_inst.spi_inst.cs_sync[1] ),
    .B(_4369_),
    .Y(_4370_));
 sg13g2_nand2_1 _8712_ (.Y(_4371_),
    .A(net138),
    .B(_4370_));
 sg13g2_o21ai_1 _8713_ (.B1(_4371_),
    .Y(_0792_),
    .A1(net138),
    .A2(net1343));
 sg13g2_nor3_1 _8714_ (.A(_3060_),
    .B(net1343),
    .C(_4217_),
    .Y(_4372_));
 sg13g2_a21o_1 _8715_ (.A2(_4370_),
    .A1(net462),
    .B1(_4372_),
    .X(_0793_));
 sg13g2_nor2_1 _8716_ (.A(net577),
    .B(_3060_),
    .Y(_4373_));
 sg13g2_nor3_1 _8717_ (.A(_3061_),
    .B(_3064_),
    .C(_4373_),
    .Y(_4374_));
 sg13g2_a21o_1 _8718_ (.A2(_4370_),
    .A1(net577),
    .B1(_4374_),
    .X(_0794_));
 sg13g2_o21ai_1 _8719_ (.B1(_3065_),
    .Y(_0795_),
    .A1(\tt6581_inst.spi_inst.cs_sync[1] ),
    .A2(_0877_));
 sg13g2_mux2_1 _8720_ (.A0(net806),
    .A1(net783),
    .S(net1343),
    .X(_0796_));
 sg13g2_mux2_1 _8721_ (.A0(net783),
    .A1(net724),
    .S(net1343),
    .X(_0797_));
 sg13g2_mux2_1 _8722_ (.A0(net724),
    .A1(net771),
    .S(net1343),
    .X(_0798_));
 sg13g2_mux2_1 _8723_ (.A0(net771),
    .A1(net277),
    .S(net1343),
    .X(_0799_));
 sg13g2_mux2_1 _8724_ (.A0(net277),
    .A1(net974),
    .S(net1343),
    .X(_0800_));
 sg13g2_mux2_1 _8725_ (.A0(\tt6581_inst.spi_inst.shift_reg[4] ),
    .A1(net648),
    .S(net1343),
    .X(_0801_));
 sg13g2_mux2_1 _8726_ (.A0(net245),
    .A1(net648),
    .S(_3063_),
    .X(_0802_));
 sg13g2_mux2_1 _8727_ (.A0(net964),
    .A1(_4066_),
    .S(net1498),
    .X(_0803_));
 sg13g2_nor2_1 _8728_ (.A(net458),
    .B(net1498),
    .Y(_4375_));
 sg13g2_a21oi_1 _8729_ (.A1(net1498),
    .A2(_4073_),
    .Y(_0804_),
    .B1(_4375_));
 sg13g2_nor2_1 _8730_ (.A(net446),
    .B(net1498),
    .Y(_4376_));
 sg13g2_a21oi_1 _8731_ (.A1(net1498),
    .A2(_4082_),
    .Y(_0805_),
    .B1(_4376_));
 sg13g2_mux2_1 _8732_ (.A0(net666),
    .A1(_4089_),
    .S(net1498),
    .X(_0806_));
 sg13g2_mux2_1 _8733_ (.A0(net685),
    .A1(_1080_),
    .S(net1498),
    .X(_0807_));
 sg13g2_mux2_1 _8734_ (.A0(net815),
    .A1(net1191),
    .S(net1498),
    .X(_0808_));
 sg13g2_mux2_1 _8735_ (.A0(net928),
    .A1(_1097_),
    .S(net1499),
    .X(_0809_));
 sg13g2_mux2_1 _8736_ (.A0(net832),
    .A1(net1185),
    .S(net1499),
    .X(_0810_));
 sg13g2_mux2_1 _8737_ (.A0(net942),
    .A1(net1184),
    .S(net1499),
    .X(_0811_));
 sg13g2_mux2_1 _8738_ (.A0(net1030),
    .A1(net1182),
    .S(net1499),
    .X(_0812_));
 sg13g2_mux2_1 _8739_ (.A0(net767),
    .A1(net1174),
    .S(net1499),
    .X(_0813_));
 sg13g2_mux2_1 _8740_ (.A0(net917),
    .A1(net1166),
    .S(net1499),
    .X(_0814_));
 sg13g2_mux2_1 _8741_ (.A0(net850),
    .A1(net1164),
    .S(net1499),
    .X(_0815_));
 sg13g2_nor2_1 _8742_ (.A(\tt6581_inst.delta_sigma_inst.audio[17] ),
    .B(net62),
    .Y(_4377_));
 sg13g2_a21oi_1 _8743_ (.A1(net62),
    .A2(_1188_),
    .Y(_0816_),
    .B1(_4377_));
 sg13g2_nand2b_2 _8744_ (.Y(_4378_),
    .B(\tt6581_inst.accum_en ),
    .A_N(\tt6581_inst.accum_in_mux ));
 sg13g2_nand2_1 _8745_ (.Y(_4379_),
    .A(net129),
    .B(_4066_));
 sg13g2_nor2_1 _8746_ (.A(_4378_),
    .B(_4379_),
    .Y(_4380_));
 sg13g2_nor2b_2 _8747_ (.A(net124),
    .B_N(_4378_),
    .Y(_4381_));
 sg13g2_inv_4 _8748_ (.A(net1293),
    .Y(_4382_));
 sg13g2_a21oi_1 _8749_ (.A1(_4066_),
    .A2(_4382_),
    .Y(_4383_),
    .B1(net129));
 sg13g2_nor3_1 _8750_ (.A(net124),
    .B(_4380_),
    .C(_4383_),
    .Y(_0817_));
 sg13g2_nand2b_1 _8751_ (.Y(_4384_),
    .B(net631),
    .A_N(_4073_));
 sg13g2_xnor2_1 _8752_ (.Y(_4385_),
    .A(_0973_),
    .B(_4073_));
 sg13g2_or2_1 _8753_ (.X(_4386_),
    .B(_4378_),
    .A(\tt6581_inst.accum_rst ));
 sg13g2_a21oi_1 _8754_ (.A1(_4379_),
    .A2(_4385_),
    .Y(_4387_),
    .B1(net1292));
 sg13g2_o21ai_1 _8755_ (.B1(_4387_),
    .Y(_4388_),
    .A1(_4379_),
    .A2(_4385_));
 sg13g2_o21ai_1 _8756_ (.B1(_4388_),
    .Y(_0818_),
    .A1(_0973_),
    .A2(_4382_));
 sg13g2_o21ai_1 _8757_ (.B1(_4384_),
    .Y(_4389_),
    .A1(_4379_),
    .A2(_4385_));
 sg13g2_xnor2_1 _8758_ (.Y(_4390_),
    .A(net1079),
    .B(_4082_));
 sg13g2_and2_1 _8759_ (.A(_4389_),
    .B(_4390_),
    .X(_4391_));
 sg13g2_nor2_1 _8760_ (.A(_4389_),
    .B(_4390_),
    .Y(_4392_));
 sg13g2_nor3_1 _8761_ (.A(net1291),
    .B(_4391_),
    .C(_4392_),
    .Y(_4393_));
 sg13g2_a21o_1 _8762_ (.A2(net1293),
    .A1(net1079),
    .B1(_4393_),
    .X(_0819_));
 sg13g2_nand2_1 _8763_ (.Y(_4394_),
    .A(net1005),
    .B(_4089_));
 sg13g2_xnor2_1 _8764_ (.Y(_4395_),
    .A(net1005),
    .B(_4089_));
 sg13g2_a21oi_1 _8765_ (.A1(\tt6581_inst.bypass_accum[2] ),
    .A2(_4083_),
    .Y(_4396_),
    .B1(_4391_));
 sg13g2_or2_1 _8766_ (.X(_4397_),
    .B(_4396_),
    .A(_4395_));
 sg13g2_a21oi_1 _8767_ (.A1(_4395_),
    .A2(_4396_),
    .Y(_4398_),
    .B1(net1291));
 sg13g2_a22oi_1 _8768_ (.Y(_4399_),
    .B1(_4397_),
    .B2(_4398_),
    .A2(net1293),
    .A1(net1005));
 sg13g2_inv_1 _8769_ (.Y(_0820_),
    .A(net1006));
 sg13g2_xnor2_1 _8770_ (.Y(_4400_),
    .A(net1048),
    .B(_1080_));
 sg13g2_a21oi_1 _8771_ (.A1(_4394_),
    .A2(_4397_),
    .Y(_4401_),
    .B1(_4400_));
 sg13g2_nand3_1 _8772_ (.B(_4397_),
    .C(_4400_),
    .A(_4394_),
    .Y(_4402_));
 sg13g2_nor2_1 _8773_ (.A(net1292),
    .B(_4401_),
    .Y(_4403_));
 sg13g2_a22oi_1 _8774_ (.Y(_4404_),
    .B1(_4402_),
    .B2(_4403_),
    .A2(net1293),
    .A1(net1048));
 sg13g2_inv_1 _8775_ (.Y(_0821_),
    .A(_4404_));
 sg13g2_a21oi_1 _8776_ (.A1(\tt6581_inst.bypass_accum[4] ),
    .A2(_1080_),
    .Y(_4405_),
    .B1(_4401_));
 sg13g2_nand2_1 _8777_ (.Y(_4406_),
    .A(\tt6581_inst.bypass_accum[5] ),
    .B(net1191));
 sg13g2_xnor2_1 _8778_ (.Y(_4407_),
    .A(net1026),
    .B(net1191));
 sg13g2_a21oi_1 _8779_ (.A1(_4405_),
    .A2(_4407_),
    .Y(_4408_),
    .B1(net1292));
 sg13g2_o21ai_1 _8780_ (.B1(_4408_),
    .Y(_4409_),
    .A1(_4405_),
    .A2(_4407_));
 sg13g2_o21ai_1 _8781_ (.B1(_4409_),
    .Y(_0822_),
    .A1(_0977_),
    .A2(_4382_));
 sg13g2_nand2_1 _8782_ (.Y(_4410_),
    .A(net359),
    .B(net1293));
 sg13g2_xnor2_1 _8783_ (.Y(_4411_),
    .A(net359),
    .B(_1097_));
 sg13g2_nand2_1 _8784_ (.Y(_4412_),
    .A(_4405_),
    .B(_4406_));
 sg13g2_o21ai_1 _8785_ (.B1(_4412_),
    .Y(_4413_),
    .A1(\tt6581_inst.bypass_accum[5] ),
    .A2(net1191));
 sg13g2_nor2_1 _8786_ (.A(_4411_),
    .B(_4413_),
    .Y(_4414_));
 sg13g2_a21o_1 _8787_ (.A2(_4413_),
    .A1(_4411_),
    .B1(net1292),
    .X(_4415_));
 sg13g2_o21ai_1 _8788_ (.B1(_4410_),
    .Y(_0823_),
    .A1(_4414_),
    .A2(_4415_));
 sg13g2_nand2_1 _8789_ (.Y(_4416_),
    .A(net399),
    .B(_4381_));
 sg13g2_xnor2_1 _8790_ (.Y(_4417_),
    .A(net399),
    .B(net1185));
 sg13g2_a21oi_1 _8791_ (.A1(net359),
    .A2(_1097_),
    .Y(_4418_),
    .B1(_4414_));
 sg13g2_nor2_1 _8792_ (.A(_4417_),
    .B(_4418_),
    .Y(_4419_));
 sg13g2_a21o_1 _8793_ (.A2(_4418_),
    .A1(_4417_),
    .B1(net1292),
    .X(_4420_));
 sg13g2_o21ai_1 _8794_ (.B1(net400),
    .Y(_0824_),
    .A1(_4419_),
    .A2(_4420_));
 sg13g2_nand2_1 _8795_ (.Y(_4421_),
    .A(net480),
    .B(net1293));
 sg13g2_xnor2_1 _8796_ (.Y(_4422_),
    .A(net480),
    .B(net1184));
 sg13g2_a21oi_1 _8797_ (.A1(net399),
    .A2(net1185),
    .Y(_4423_),
    .B1(_4419_));
 sg13g2_nor2_1 _8798_ (.A(_4422_),
    .B(_4423_),
    .Y(_4424_));
 sg13g2_a21o_1 _8799_ (.A2(_4423_),
    .A1(_4422_),
    .B1(net1291),
    .X(_4425_));
 sg13g2_o21ai_1 _8800_ (.B1(_4421_),
    .Y(_0825_),
    .A1(_4424_),
    .A2(_4425_));
 sg13g2_a21oi_1 _8801_ (.A1(net480),
    .A2(net1184),
    .Y(_4426_),
    .B1(_4424_));
 sg13g2_nand2_1 _8802_ (.Y(_4427_),
    .A(\tt6581_inst.bypass_accum[9] ),
    .B(net1183));
 sg13g2_xnor2_1 _8803_ (.Y(_4428_),
    .A(net1068),
    .B(net1183));
 sg13g2_a21oi_1 _8804_ (.A1(_4426_),
    .A2(_4428_),
    .Y(_4429_),
    .B1(net1291));
 sg13g2_o21ai_1 _8805_ (.B1(_4429_),
    .Y(_4430_),
    .A1(_4426_),
    .A2(_4428_));
 sg13g2_o21ai_1 _8806_ (.B1(_4430_),
    .Y(_0826_),
    .A1(_0976_),
    .A2(_4382_));
 sg13g2_nand2_1 _8807_ (.Y(_4431_),
    .A(net517),
    .B(net1293));
 sg13g2_xnor2_1 _8808_ (.Y(_4432_),
    .A(net517),
    .B(net1174));
 sg13g2_nand2_1 _8809_ (.Y(_4433_),
    .A(_4426_),
    .B(_4427_));
 sg13g2_o21ai_1 _8810_ (.B1(_4433_),
    .Y(_4434_),
    .A1(\tt6581_inst.bypass_accum[9] ),
    .A2(net1183));
 sg13g2_nor2_1 _8811_ (.A(_4432_),
    .B(_4434_),
    .Y(_4435_));
 sg13g2_a21o_1 _8812_ (.A2(_4434_),
    .A1(_4432_),
    .B1(net1291),
    .X(_4436_));
 sg13g2_o21ai_1 _8813_ (.B1(_4431_),
    .Y(_0827_),
    .A1(_4435_),
    .A2(_4436_));
 sg13g2_a21o_1 _8814_ (.A2(net1174),
    .A1(net517),
    .B1(_4435_),
    .X(_4437_));
 sg13g2_xnor2_1 _8815_ (.Y(_4438_),
    .A(_0975_),
    .B(net1166));
 sg13g2_a21oi_1 _8816_ (.A1(_4437_),
    .A2(_4438_),
    .Y(_4439_),
    .B1(net1291));
 sg13g2_o21ai_1 _8817_ (.B1(_4439_),
    .Y(_4440_),
    .A1(_4437_),
    .A2(_4438_));
 sg13g2_o21ai_1 _8818_ (.B1(_4440_),
    .Y(_0828_),
    .A1(_0975_),
    .A2(_4382_));
 sg13g2_nand2_1 _8819_ (.Y(_4441_),
    .A(net486),
    .B(net1293));
 sg13g2_xnor2_1 _8820_ (.Y(_4442_),
    .A(net486),
    .B(net1164));
 sg13g2_a21o_1 _8821_ (.A2(net1166),
    .A1(\tt6581_inst.bypass_accum[11] ),
    .B1(_4437_),
    .X(_4443_));
 sg13g2_o21ai_1 _8822_ (.B1(_4443_),
    .Y(_4444_),
    .A1(\tt6581_inst.bypass_accum[11] ),
    .A2(net1166));
 sg13g2_nor2_1 _8823_ (.A(_4442_),
    .B(_4444_),
    .Y(_4445_));
 sg13g2_a21o_1 _8824_ (.A2(_4444_),
    .A1(_4442_),
    .B1(net1291),
    .X(_4446_));
 sg13g2_o21ai_1 _8825_ (.B1(_4441_),
    .Y(_0829_),
    .A1(_4445_),
    .A2(_4446_));
 sg13g2_a21oi_1 _8826_ (.A1(net486),
    .A2(net1164),
    .Y(_4447_),
    .B1(_4445_));
 sg13g2_xnor2_1 _8827_ (.Y(_4448_),
    .A(net571),
    .B(_1187_));
 sg13g2_a21oi_1 _8828_ (.A1(_4447_),
    .A2(_4448_),
    .Y(_4449_),
    .B1(net1291));
 sg13g2_o21ai_1 _8829_ (.B1(_4449_),
    .Y(_4450_),
    .A1(_4447_),
    .A2(_4448_));
 sg13g2_o21ai_1 _8830_ (.B1(_4450_),
    .Y(_0830_),
    .A1(_0974_),
    .A2(_4382_));
 sg13g2_dfrbpq_2 _8831_ (.RESET_B(net1592),
    .D(net1047),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8832_ (.RESET_B(net1591),
    .D(net745),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[9] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8833_ (.RESET_B(net1609),
    .D(_0119_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[10] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _8834_ (.RESET_B(net1609),
    .D(net596),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[11] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8835_ (.RESET_B(net1591),
    .D(net701),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _8836_ (.RESET_B(net1591),
    .D(net513),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8837_ (.RESET_B(net1609),
    .D(_0123_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[14] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8838_ (.RESET_B(net1603),
    .D(net601),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[15] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _8839_ (.RESET_B(net1599),
    .D(net1029),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _8840_ (.RESET_B(net1592),
    .D(_0126_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _8841_ (.RESET_B(net1609),
    .D(_0127_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8842_ (.RESET_B(net1616),
    .D(_0128_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _8843_ (.RESET_B(net1591),
    .D(net995),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _8844_ (.RESET_B(net1599),
    .D(net953),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _8845_ (.RESET_B(net1604),
    .D(_0131_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8846_ (.RESET_B(net1604),
    .D(net524),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8847_ (.RESET_B(net1603),
    .D(net786),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[8] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8848_ (.RESET_B(net1602),
    .D(net740),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[9] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _8849_ (.RESET_B(net1606),
    .D(_0135_),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8850_ (.RESET_B(net1607),
    .D(net582),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8851_ (.RESET_B(net1606),
    .D(net988),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8852_ (.RESET_B(net1605),
    .D(net620),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8853_ (.RESET_B(net1602),
    .D(_0139_),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8854_ (.RESET_B(net1605),
    .D(net540),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[15] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8855_ (.RESET_B(net1603),
    .D(net709),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8856_ (.RESET_B(net1603),
    .D(net622),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8857_ (.RESET_B(net1605),
    .D(_0143_),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8858_ (.RESET_B(net1607),
    .D(net629),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _8859_ (.RESET_B(net1606),
    .D(net836),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8860_ (.RESET_B(net1606),
    .D(net927),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _8861_ (.RESET_B(net1606),
    .D(net552),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _8862_ (.RESET_B(net1602),
    .D(net576),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8863_ (.RESET_B(net1613),
    .D(net263),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8864_ (.RESET_B(net1616),
    .D(_0150_),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _8865_ (.RESET_B(net1616),
    .D(net809),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[10] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8866_ (.RESET_B(net1616),
    .D(_0152_),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[11] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _8867_ (.RESET_B(net1611),
    .D(net930),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[12] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8868_ (.RESET_B(net1611),
    .D(net735),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[13] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _8869_ (.RESET_B(net1612),
    .D(net698),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[14] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _8870_ (.RESET_B(net1611),
    .D(net754),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[15] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _8871_ (.RESET_B(net1613),
    .D(net800),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _8872_ (.RESET_B(net1617),
    .D(net757),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _8873_ (.RESET_B(net1616),
    .D(_0159_),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8874_ (.RESET_B(net1617),
    .D(_0160_),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _8875_ (.RESET_B(net1598),
    .D(net634),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8876_ (.RESET_B(net1598),
    .D(net798),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _8877_ (.RESET_B(net1612),
    .D(net677),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _8878_ (.RESET_B(net1598),
    .D(_0164_),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _8879_ (.RESET_B(net1648),
    .D(net641),
    .Q(\tt6581_inst.svf_inst.hp_node[0] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8880_ (.RESET_B(net1648),
    .D(_0166_),
    .Q(\tt6581_inst.svf_inst.hp_node[1] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8881_ (.RESET_B(net1647),
    .D(net598),
    .Q(\tt6581_inst.svf_inst.hp_node[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8882_ (.RESET_B(net1642),
    .D(_0168_),
    .Q(\tt6581_inst.svf_inst.hp_node[3] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _8883_ (.RESET_B(net1641),
    .D(net749),
    .Q(\tt6581_inst.svf_inst.hp_node[4] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _8884_ (.RESET_B(net1640),
    .D(_0170_),
    .Q(\tt6581_inst.svf_inst.hp_node[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _8885_ (.RESET_B(net1626),
    .D(net717),
    .Q(\tt6581_inst.svf_inst.hp_node[6] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8886_ (.RESET_B(net1626),
    .D(net849),
    .Q(\tt6581_inst.svf_inst.hp_node[7] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8887_ (.RESET_B(net1624),
    .D(net866),
    .Q(\tt6581_inst.svf_inst.hp_node[8] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8888_ (.RESET_B(net1624),
    .D(net1010),
    .Q(\tt6581_inst.svf_inst.hp_node[9] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _8889_ (.RESET_B(net1624),
    .D(net959),
    .Q(\tt6581_inst.svf_inst.hp_node[10] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _8890_ (.RESET_B(net1574),
    .D(_0176_),
    .Q(\tt6581_inst.svf_inst.hp_node[11] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _8891_ (.RESET_B(net1574),
    .D(net722),
    .Q(\tt6581_inst.svf_inst.hp_node[12] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _8892_ (.RESET_B(net1574),
    .D(net893),
    .Q(\tt6581_inst.svf_inst.hp_node[13] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _8893_ (.RESET_B(net1572),
    .D(_0179_),
    .Q(\tt6581_inst.svf_inst.hp_node[14] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _8894_ (.RESET_B(net1572),
    .D(net1095),
    .Q(\tt6581_inst.svf_inst.hp_node[15] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _8895_ (.RESET_B(net1572),
    .D(_0181_),
    .Q(\tt6581_inst.svf_inst.hp_node[16] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _8896_ (.RESET_B(net1558),
    .D(_0182_),
    .Q(\tt6581_inst.svf_inst.hp_node[17] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _8897_ (.RESET_B(net1558),
    .D(_0183_),
    .Q(\tt6581_inst.svf_inst.hp_node[18] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _8898_ (.RESET_B(net1558),
    .D(_0184_),
    .Q(\tt6581_inst.svf_inst.hp_node[19] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _8899_ (.RESET_B(net1559),
    .D(_0185_),
    .Q(\tt6581_inst.svf_inst.hp_node[20] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _8900_ (.RESET_B(net1573),
    .D(_0186_),
    .Q(\tt6581_inst.svf_inst.hp_node[21] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _8901_ (.RESET_B(net1566),
    .D(net501),
    .Q(\tt6581_inst.svf_inst.hp_node[22] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _8902_ (.RESET_B(net1577),
    .D(_0188_),
    .Q(\tt6581_inst.svf_inst.hp_node[23] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _8903_ (.RESET_B(net1672),
    .D(_0189_),
    .Q(\tt6581_inst.controller_inst.sr_i[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8904_ (.RESET_B(net1672),
    .D(_0190_),
    .Q(\tt6581_inst.controller_inst.sr_i[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8905_ (.RESET_B(net1673),
    .D(net1067),
    .Q(\tt6581_inst.controller_inst.sr_i[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8906_ (.RESET_B(net1671),
    .D(net1093),
    .Q(\tt6581_inst.controller_inst.sr_i[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8907_ (.RESET_B(net1671),
    .D(_0193_),
    .Q(\tt6581_inst.controller_inst.sr_i[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _8908_ (.RESET_B(net1665),
    .D(net861),
    .Q(\tt6581_inst.controller_inst.sr_i[5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8909_ (.RESET_B(net1672),
    .D(_0195_),
    .Q(\tt6581_inst.controller_inst.sr_i[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8910_ (.RESET_B(net1668),
    .D(net949),
    .Q(\tt6581_inst.controller_inst.sr_i[7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8911_ (.RESET_B(net1669),
    .D(_0197_),
    .Q(\tt6581_inst.controller_inst.sr_i[8] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _8912_ (.RESET_B(net1670),
    .D(_0198_),
    .Q(\tt6581_inst.controller_inst.sr_i[9] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8913_ (.RESET_B(net1669),
    .D(net1014),
    .Q(\tt6581_inst.controller_inst.sr_i[10] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8914_ (.RESET_B(net1669),
    .D(net907),
    .Q(\tt6581_inst.controller_inst.sr_i[11] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _8915_ (.RESET_B(net1663),
    .D(net679),
    .Q(\tt6581_inst.controller_inst.sr_i[12] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _8916_ (.RESET_B(net1667),
    .D(_0202_),
    .Q(\tt6581_inst.controller_inst.sr_i[13] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _8917_ (.RESET_B(net1665),
    .D(_0203_),
    .Q(\tt6581_inst.controller_inst.sr_i[14] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _8918_ (.RESET_B(net1665),
    .D(net941),
    .Q(\tt6581_inst.controller_inst.sr_i[15] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8919_ (.RESET_B(net1648),
    .D(net37),
    .Q(_0036_),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8920_ (.RESET_B(net1636),
    .D(_0000_),
    .Q(\tt6581_inst.controller_inst.cur_state[1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _8921_ (.RESET_B(net1650),
    .D(net56),
    .Q(\tt6581_inst.controller_inst.cur_state[2] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8922_ (.RESET_B(net1651),
    .D(net58),
    .Q(\tt6581_inst.controller_inst.cur_state[3] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8923_ (.RESET_B(net1648),
    .D(net61),
    .Q(\tt6581_inst.controller_inst.cur_state[4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8924_ (.RESET_B(net1636),
    .D(_0002_),
    .Q(\tt6581_inst.controller_inst.cur_state[5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _8925_ (.RESET_B(net1651),
    .D(_0012_),
    .Q(\tt6581_inst.controller_inst.cur_state[6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8926_ (.RESET_B(net1637),
    .D(_0013_),
    .Q(\tt6581_inst.controller_inst.cur_state[7] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _8927_ (.RESET_B(net1650),
    .D(net78),
    .Q(\tt6581_inst.controller_inst.cur_state[8] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8928_ (.RESET_B(net1650),
    .D(_0004_),
    .Q(\tt6581_inst.controller_inst.cur_state[9] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _8929_ (.RESET_B(net1636),
    .D(_0009_),
    .Q(\tt6581_inst.controller_inst.cur_state[10] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _8930_ (.RESET_B(net1670),
    .D(_0205_),
    .Q(\tt6581_inst.ad_pack[8] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _8931_ (.RESET_B(net1672),
    .D(_0206_),
    .Q(\tt6581_inst.ad_pack[9] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _8932_ (.RESET_B(net1672),
    .D(net932),
    .Q(\tt6581_inst.ad_pack[10] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _8933_ (.RESET_B(net1670),
    .D(net761),
    .Q(\tt6581_inst.ad_pack[11] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _8934_ (.RESET_B(net1662),
    .D(net752),
    .Q(\tt6581_inst.ad_pack[12] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8935_ (.RESET_B(net1666),
    .D(net951),
    .Q(\tt6581_inst.ad_pack[13] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _8936_ (.RESET_B(net1665),
    .D(_0211_),
    .Q(\tt6581_inst.ad_pack[14] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _8937_ (.RESET_B(net1665),
    .D(_0212_),
    .Q(\tt6581_inst.ad_pack[15] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8938_ (.RESET_B(net1668),
    .D(_0213_),
    .Q(\tt6581_inst.ad_pack[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8939_ (.RESET_B(net1666),
    .D(_0214_),
    .Q(\tt6581_inst.ad_pack[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _8940_ (.RESET_B(net1672),
    .D(net1057),
    .Q(\tt6581_inst.ad_pack[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8941_ (.RESET_B(net1672),
    .D(net1052),
    .Q(\tt6581_inst.ad_pack[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _8942_ (.RESET_B(net1666),
    .D(net665),
    .Q(\tt6581_inst.ad_pack[4] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8943_ (.RESET_B(net1665),
    .D(net693),
    .Q(\tt6581_inst.ad_pack[5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _8944_ (.RESET_B(net1666),
    .D(_0219_),
    .Q(\tt6581_inst.ad_pack[6] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _8945_ (.RESET_B(net1666),
    .D(net638),
    .Q(\tt6581_inst.ad_pack[7] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _8946_ (.RESET_B(net1662),
    .D(net775),
    .Q(\tt6581_inst.control_pack[8] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _8947_ (.RESET_B(net1591),
    .D(net788),
    .Q(\tt6581_inst.control_pack[9] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8948_ (.RESET_B(net1616),
    .D(net461),
    .Q(\tt6581_inst.control_pack[10] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8949_ (.RESET_B(net1669),
    .D(net407),
    .Q(\tt6581_inst.control_pack[11] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _8950_ (.RESET_B(net1598),
    .D(net868),
    .Q(\tt6581_inst.control_pack[12] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _8951_ (.RESET_B(net1602),
    .D(net935),
    .Q(\tt6581_inst.control_pack[13] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _8952_ (.RESET_B(net1602),
    .D(_0227_),
    .Q(\tt6581_inst.control_pack[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _8953_ (.RESET_B(net1591),
    .D(net231),
    .Q(\tt6581_inst.control_pack[15] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8954_ (.RESET_B(net1617),
    .D(net853),
    .Q(\tt6581_inst.control_pack[0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8955_ (.RESET_B(net1598),
    .D(net738),
    .Q(\tt6581_inst.control_pack[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8956_ (.RESET_B(net1617),
    .D(_0231_),
    .Q(\tt6581_inst.control_pack[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8957_ (.RESET_B(net1616),
    .D(_0232_),
    .Q(\tt6581_inst.control_pack[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _8958_ (.RESET_B(net1611),
    .D(net689),
    .Q(\tt6581_inst.control_pack[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _8959_ (.RESET_B(net1604),
    .D(net592),
    .Q(\tt6581_inst.control_pack[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8960_ (.RESET_B(net1604),
    .D(net586),
    .Q(\tt6581_inst.control_pack[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _8961_ (.RESET_B(net1603),
    .D(net626),
    .Q(\tt6581_inst.control_pack[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _8962_ (.RESET_B(net1604),
    .D(net270),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8963_ (.RESET_B(net1603),
    .D(net568),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8964_ (.RESET_B(net1602),
    .D(net235),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _8965_ (.RESET_B(net1609),
    .D(net904),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[11] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8966_ (.RESET_B(net1608),
    .D(net375),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[12] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _8967_ (.RESET_B(net1610),
    .D(_0242_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[13] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8968_ (.RESET_B(net1610),
    .D(_0243_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[14] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _8969_ (.RESET_B(net1610),
    .D(net314),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[15] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _8970_ (.RESET_B(net1612),
    .D(net879),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8971_ (.RESET_B(net1611),
    .D(net505),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _8972_ (.RESET_B(net1612),
    .D(_0247_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8973_ (.RESET_B(net1612),
    .D(_0248_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _8974_ (.RESET_B(net1611),
    .D(net490),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _8975_ (.RESET_B(net1611),
    .D(net452),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _8976_ (.RESET_B(net1612),
    .D(net289),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _8977_ (.RESET_B(net1611),
    .D(net392),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _8978_ (.RESET_B(net1643),
    .D(net113),
    .Q(\tt6581_inst.delta_sigma_inst.en ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _8979_ (.RESET_B(net1655),
    .D(_0253_),
    .Q(pdm),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _8980_ (.RESET_B(net1650),
    .D(net570),
    .Q(\tt6581_inst.controller_inst.cur_voice[0] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _8981_ (.RESET_B(net1651),
    .D(_0255_),
    .Q(\tt6581_inst.controller_inst.cur_voice[1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _8982_ (.RESET_B(net1643),
    .D(net217),
    .Q(\tt6581_inst.delta_sigma_inst.e1[0] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _8983_ (.RESET_B(net1643),
    .D(net472),
    .Q(\tt6581_inst.delta_sigma_inst.e1[1] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _8984_ (.RESET_B(net1645),
    .D(_0258_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[2] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8985_ (.RESET_B(net1643),
    .D(net763),
    .Q(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _8986_ (.RESET_B(net1644),
    .D(_0260_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[4] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _8987_ (.RESET_B(net1645),
    .D(_0261_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[5] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8988_ (.RESET_B(net1645),
    .D(_0262_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8989_ (.RESET_B(net1645),
    .D(_0263_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _8990_ (.RESET_B(net1654),
    .D(_0264_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8991_ (.RESET_B(net1654),
    .D(_0265_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[9] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8992_ (.RESET_B(net1654),
    .D(_0266_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[10] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _8993_ (.RESET_B(net1654),
    .D(_0267_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[11] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _8994_ (.RESET_B(net1656),
    .D(_0268_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _8995_ (.RESET_B(net1653),
    .D(_0269_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[13] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8996_ (.RESET_B(net1653),
    .D(_0270_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[14] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _8997_ (.RESET_B(net1655),
    .D(_0271_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[15] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _8998_ (.RESET_B(net1655),
    .D(_0272_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[16] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _8999_ (.RESET_B(net1655),
    .D(_0273_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[17] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _9000_ (.RESET_B(net1655),
    .D(_0274_),
    .Q(\tt6581_inst.delta_sigma_inst.e1[18] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _9001_ (.RESET_B(net1643),
    .D(net45),
    .Q(\tt6581_inst.delta_sigma_inst.cnt[0] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _9002_ (.RESET_B(net1643),
    .D(_0021_),
    .Q(\tt6581_inst.delta_sigma_inst.cnt[1] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _9003_ (.RESET_B(net1643),
    .D(_0022_),
    .Q(\tt6581_inst.delta_sigma_inst.cnt[2] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9004_ (.RESET_B(net1646),
    .D(_0275_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[0] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _9005_ (.RESET_B(net1646),
    .D(_0276_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[1] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _9006_ (.RESET_B(net1646),
    .D(_0277_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[2] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _9007_ (.RESET_B(net1643),
    .D(net712),
    .Q(\tt6581_inst.delta_sigma_inst.e2[3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _9008_ (.RESET_B(net1644),
    .D(_0279_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _9009_ (.RESET_B(net1644),
    .D(_0280_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[5] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9010_ (.RESET_B(net1645),
    .D(net668),
    .Q(\tt6581_inst.delta_sigma_inst.e2[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _9011_ (.RESET_B(net1645),
    .D(_0282_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _9012_ (.RESET_B(net1645),
    .D(net687),
    .Q(\tt6581_inst.delta_sigma_inst.e2[8] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _9013_ (.RESET_B(net1654),
    .D(_0284_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[9] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _9014_ (.RESET_B(net1654),
    .D(_0285_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[10] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _9015_ (.RESET_B(net1654),
    .D(_0286_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[11] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _9016_ (.RESET_B(net1656),
    .D(net673),
    .Q(\tt6581_inst.delta_sigma_inst.e2[12] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _9017_ (.RESET_B(net1656),
    .D(_0288_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[13] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _9018_ (.RESET_B(net1653),
    .D(_0289_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[14] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _9019_ (.RESET_B(net1655),
    .D(_0290_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[15] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _9020_ (.RESET_B(net1655),
    .D(_0291_),
    .Q(\tt6581_inst.delta_sigma_inst.e2[16] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _9021_ (.RESET_B(net1655),
    .D(net425),
    .Q(\tt6581_inst.delta_sigma_inst.e2[17] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _9022_ (.RESET_B(net1656),
    .D(net188),
    .Q(\tt6581_inst.delta_sigma_inst.e2[18] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _9023_ (.RESET_B(net1577),
    .D(net1192),
    .Q(\tt6581_inst.mult_inst.cur_state ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _9024_ (.RESET_B(net1577),
    .D(_0294_),
    .Q(\tt6581_inst.mult_inst.iter[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _9025_ (.RESET_B(net1577),
    .D(_0295_),
    .Q(\tt6581_inst.mult_inst.iter[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _9026_ (.RESET_B(net1577),
    .D(_0296_),
    .Q(\tt6581_inst.mult_inst.iter[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _9027_ (.RESET_B(net1577),
    .D(_0297_),
    .Q(\tt6581_inst.mult_inst.iter[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _9028_ (.RESET_B(net1577),
    .D(net66),
    .Q(\tt6581_inst.mult_inst.iter[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _9029_ (.RESET_B(net1577),
    .D(_0299_),
    .Q(\tt6581_inst.mult_inst.a_reg[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _9030_ (.RESET_B(net1578),
    .D(net973),
    .Q(\tt6581_inst.mult_inst.a_reg[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _9031_ (.RESET_B(net1583),
    .D(net542),
    .Q(\tt6581_inst.mult_inst.a_reg[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _9032_ (.RESET_B(net1581),
    .D(net274),
    .Q(\tt6581_inst.mult_inst.a_reg[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _9033_ (.RESET_B(net1581),
    .D(net225),
    .Q(\tt6581_inst.mult_inst.a_reg[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9034_ (.RESET_B(net1583),
    .D(net207),
    .Q(\tt6581_inst.mult_inst.a_reg[5] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _9035_ (.RESET_B(net1583),
    .D(_0305_),
    .Q(\tt6581_inst.mult_inst.a_reg[6] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _9036_ (.RESET_B(net1583),
    .D(net272),
    .Q(\tt6581_inst.mult_inst.a_reg[7] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _9037_ (.RESET_B(net1629),
    .D(_0307_),
    .Q(\tt6581_inst.mult_inst.a_reg[8] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _9038_ (.RESET_B(net1629),
    .D(net872),
    .Q(\tt6581_inst.mult_inst.a_reg[9] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _9039_ (.RESET_B(net1629),
    .D(net554),
    .Q(\tt6581_inst.mult_inst.a_reg[10] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _9040_ (.RESET_B(net1629),
    .D(net530),
    .Q(\tt6581_inst.mult_inst.a_reg[11] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9041_ (.RESET_B(net1629),
    .D(_0311_),
    .Q(\tt6581_inst.mult_inst.a_reg[12] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _9042_ (.RESET_B(net1629),
    .D(net580),
    .Q(\tt6581_inst.mult_inst.a_reg[13] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _9043_ (.RESET_B(net1583),
    .D(_0313_),
    .Q(\tt6581_inst.mult_inst.a_reg[14] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _9044_ (.RESET_B(net1583),
    .D(net1016),
    .Q(\tt6581_inst.mult_inst.a_reg[15] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _9045_ (.RESET_B(net1578),
    .D(_0315_),
    .Q(\tt6581_inst.mult_inst.a_reg[16] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _9046_ (.RESET_B(net1575),
    .D(net369),
    .Q(\tt6581_inst.mult_inst.a_reg[17] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _9047_ (.RESET_B(net1575),
    .D(net210),
    .Q(\tt6581_inst.mult_inst.a_reg[18] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _9048_ (.RESET_B(net1578),
    .D(_0318_),
    .Q(\tt6581_inst.mult_inst.a_reg[19] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _9049_ (.RESET_B(net1573),
    .D(net244),
    .Q(\tt6581_inst.mult_inst.a_reg[20] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _9050_ (.RESET_B(net1573),
    .D(_0320_),
    .Q(\tt6581_inst.mult_inst.a_reg[21] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _9051_ (.RESET_B(net1573),
    .D(net253),
    .Q(\tt6581_inst.mult_inst.a_reg[22] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _9052_ (.RESET_B(net1573),
    .D(_0322_),
    .Q(\tt6581_inst.mult_inst.a_reg[23] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _9053_ (.RESET_B(net1553),
    .D(_0323_),
    .Q(\tt6581_inst.mult_inst.a_reg[24] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _9054_ (.RESET_B(net1553),
    .D(_0324_),
    .Q(\tt6581_inst.mult_inst.a_reg[25] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _9055_ (.RESET_B(net1553),
    .D(_0325_),
    .Q(\tt6581_inst.mult_inst.a_reg[26] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _9056_ (.RESET_B(net1553),
    .D(_0326_),
    .Q(\tt6581_inst.mult_inst.a_reg[27] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _9057_ (.RESET_B(net1553),
    .D(_0327_),
    .Q(\tt6581_inst.mult_inst.a_reg[28] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9058_ (.RESET_B(net1553),
    .D(_0328_),
    .Q(\tt6581_inst.mult_inst.a_reg[29] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9059_ (.RESET_B(net1553),
    .D(_0329_),
    .Q(\tt6581_inst.mult_inst.a_reg[30] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9060_ (.RESET_B(net1555),
    .D(_0330_),
    .Q(\tt6581_inst.mult_inst.a_reg[31] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9061_ (.RESET_B(net1555),
    .D(_0331_),
    .Q(\tt6581_inst.mult_inst.a_reg[32] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _9062_ (.RESET_B(net1555),
    .D(_0332_),
    .Q(\tt6581_inst.mult_inst.a_reg[33] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _9063_ (.RESET_B(net1555),
    .D(_0333_),
    .Q(\tt6581_inst.mult_inst.a_reg[34] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _9064_ (.RESET_B(net1555),
    .D(_0334_),
    .Q(\tt6581_inst.mult_inst.a_reg[35] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _9065_ (.RESET_B(net1555),
    .D(_0335_),
    .Q(\tt6581_inst.mult_inst.a_reg[36] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _9066_ (.RESET_B(net1560),
    .D(_0336_),
    .Q(\tt6581_inst.mult_inst.a_reg[37] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _9067_ (.RESET_B(net1562),
    .D(_0337_),
    .Q(\tt6581_inst.mult_inst.a_reg[38] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _9068_ (.RESET_B(net1675),
    .D(net133),
    .Q(_0037_),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9069_ (.RESET_B(net1675),
    .D(_0339_),
    .Q(_0038_),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9070_ (.RESET_B(net1632),
    .D(_0340_),
    .Q(\tt6581_inst.mult_inst.b_reg[0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9071_ (.RESET_B(net1637),
    .D(net103),
    .Q(\tt6581_inst.mult_inst.b_reg[1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9072_ (.RESET_B(net1637),
    .D(net87),
    .Q(\tt6581_inst.mult_inst.b_reg[2] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9073_ (.RESET_B(net1637),
    .D(net116),
    .Q(\tt6581_inst.mult_inst.b_reg[3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9074_ (.RESET_B(net1637),
    .D(net101),
    .Q(\tt6581_inst.mult_inst.b_reg[4] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9075_ (.RESET_B(net1638),
    .D(net85),
    .Q(\tt6581_inst.mult_inst.b_reg[5] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9076_ (.RESET_B(net1638),
    .D(net76),
    .Q(\tt6581_inst.mult_inst.b_reg[6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9077_ (.RESET_B(net1636),
    .D(_0347_),
    .Q(\tt6581_inst.mult_inst.b_reg[7] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9078_ (.RESET_B(net1638),
    .D(net74),
    .Q(\tt6581_inst.mult_inst.b_reg[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9079_ (.RESET_B(net1636),
    .D(net111),
    .Q(\tt6581_inst.mult_inst.b_reg[9] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9080_ (.RESET_B(net1632),
    .D(_0350_),
    .Q(\tt6581_inst.mult_inst.b_reg[10] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9081_ (.RESET_B(net1632),
    .D(net83),
    .Q(\tt6581_inst.mult_inst.b_reg[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _9082_ (.RESET_B(net1632),
    .D(_0352_),
    .Q(\tt6581_inst.mult_inst.b_reg[12] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _9083_ (.RESET_B(net1631),
    .D(net80),
    .Q(\tt6581_inst.mult_inst.b_reg[13] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _9084_ (.RESET_B(net1631),
    .D(net238),
    .Q(\tt6581_inst.mult_inst.b_reg[14] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _9085_ (.RESET_B(net1631),
    .D(net240),
    .Q(\tt6581_inst.mult_inst.b_reg[15] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _9086_ (.RESET_B(net1578),
    .D(net437),
    .Q(\tt6581_inst.mult_inst.accum[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _9087_ (.RESET_B(net1580),
    .D(net433),
    .Q(\tt6581_inst.mult_inst.accum[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _9088_ (.RESET_B(net1581),
    .D(net308),
    .Q(\tt6581_inst.mult_inst.accum[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _9089_ (.RESET_B(net1581),
    .D(net443),
    .Q(\tt6581_inst.mult_inst.accum[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9090_ (.RESET_B(net1582),
    .D(net276),
    .Q(\tt6581_inst.mult_inst.accum[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9091_ (.RESET_B(net1582),
    .D(_0361_),
    .Q(\tt6581_inst.mult_inst.accum[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9092_ (.RESET_B(net1582),
    .D(net256),
    .Q(\tt6581_inst.mult_inst.accum[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9093_ (.RESET_B(net1631),
    .D(_0363_),
    .Q(\tt6581_inst.mult_inst.accum[7] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _9094_ (.RESET_B(net1631),
    .D(_0364_),
    .Q(\tt6581_inst.mult_inst.accum[8] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _9095_ (.RESET_B(net1631),
    .D(net557),
    .Q(\tt6581_inst.mult_inst.accum[9] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _9096_ (.RESET_B(net1629),
    .D(_0366_),
    .Q(\tt6581_inst.mult_inst.accum[10] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _9097_ (.RESET_B(net1630),
    .D(net1075),
    .Q(\tt6581_inst.mult_inst.accum[11] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _9098_ (.RESET_B(net1630),
    .D(net492),
    .Q(\tt6581_inst.mult_inst.accum[12] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9099_ (.RESET_B(net1630),
    .D(_0369_),
    .Q(\tt6581_inst.mult_inst.accum[13] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9100_ (.RESET_B(net1630),
    .D(net691),
    .Q(\tt6581_inst.mult_inst.accum[14] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9101_ (.RESET_B(net1630),
    .D(net466),
    .Q(\tt6581_inst.mult_inst.accum[15] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9102_ (.RESET_B(net1628),
    .D(_0372_),
    .Q(\tt6581_inst.mult_inst.accum[16] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9103_ (.RESET_B(net1625),
    .D(net1100),
    .Q(\tt6581_inst.mult_inst.accum[17] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _9104_ (.RESET_B(net1576),
    .D(_0374_),
    .Q(\tt6581_inst.mult_inst.accum[18] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9105_ (.RESET_B(net1575),
    .D(net842),
    .Q(\tt6581_inst.mult_inst.accum[19] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9106_ (.RESET_B(net1575),
    .D(_0376_),
    .Q(\tt6581_inst.mult_inst.accum[20] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9107_ (.RESET_B(net1575),
    .D(_0377_),
    .Q(\tt6581_inst.mult_inst.accum[21] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9108_ (.RESET_B(net1575),
    .D(net496),
    .Q(\tt6581_inst.mult_inst.accum[22] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9109_ (.RESET_B(net1574),
    .D(_0379_),
    .Q(\tt6581_inst.mult_inst.accum[23] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9110_ (.RESET_B(net1554),
    .D(_0380_),
    .Q(\tt6581_inst.mult_inst.accum[24] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9111_ (.RESET_B(net1554),
    .D(_0381_),
    .Q(\tt6581_inst.mult_inst.accum[25] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9112_ (.RESET_B(net1554),
    .D(_0382_),
    .Q(\tt6581_inst.mult_inst.accum[26] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9113_ (.RESET_B(net1554),
    .D(net1091),
    .Q(\tt6581_inst.mult_inst.accum[27] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9114_ (.RESET_B(net1554),
    .D(net607),
    .Q(\tt6581_inst.mult_inst.accum[28] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9115_ (.RESET_B(net1554),
    .D(net574),
    .Q(\tt6581_inst.mult_inst.accum[29] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9116_ (.RESET_B(net1554),
    .D(net611),
    .Q(\tt6581_inst.mult_inst.accum[30] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9117_ (.RESET_B(net1553),
    .D(net1084),
    .Q(\tt6581_inst.mult_inst.accum[31] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9118_ (.RESET_B(net1555),
    .D(_0388_),
    .Q(\tt6581_inst.mult_inst.accum[32] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _9119_ (.RESET_B(net1556),
    .D(net998),
    .Q(\tt6581_inst.mult_inst.accum[33] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9120_ (.RESET_B(net1556),
    .D(_0390_),
    .Q(\tt6581_inst.mult_inst.accum[34] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9121_ (.RESET_B(net1556),
    .D(net707),
    .Q(\tt6581_inst.mult_inst.accum[35] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9122_ (.RESET_B(net1556),
    .D(net381),
    .Q(\tt6581_inst.mult_inst.accum[36] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9123_ (.RESET_B(net1562),
    .D(_0393_),
    .Q(\tt6581_inst.mult_inst.accum[37] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9124_ (.RESET_B(net1562),
    .D(net212),
    .Q(\tt6581_inst.mult_inst.accum[38] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _9125_ (.RESET_B(net1636),
    .D(net43),
    .Q(_0039_),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _9126_ (.RESET_B(net1634),
    .D(_0016_),
    .Q(\tt6581_inst.svf_inst.cur_state[1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _9127_ (.RESET_B(net1566),
    .D(net1510),
    .Q(\tt6581_inst.svf_inst.cur_state[2] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _9128_ (.RESET_B(net1634),
    .D(_0017_),
    .Q(\tt6581_inst.svf_inst.cur_state[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _9129_ (.RESET_B(net1635),
    .D(net1521),
    .Q(\tt6581_inst.controller_inst.filt_ready_i ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _9130_ (.RESET_B(net1634),
    .D(net52),
    .Q(\tt6581_inst.svf_inst.cur_state[5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _9131_ (.RESET_B(net1637),
    .D(net39),
    .Q(\tt6581_inst.svf_inst.cur_state[6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9132_ (.RESET_B(net1648),
    .D(net54),
    .Q(\tt6581_inst.svf_inst.cur_state[7] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _9133_ (.RESET_B(net1634),
    .D(_0018_),
    .Q(\tt6581_inst.svf_inst.cur_state[8] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _9134_ (.RESET_B(net1648),
    .D(net50),
    .Q(\tt6581_inst.svf_inst.cur_state[9] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _9135_ (.RESET_B(net1635),
    .D(net1530),
    .Q(\tt6581_inst.svf_inst.cur_state[10] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _9136_ (.RESET_B(net1620),
    .D(net247),
    .Q(\tt6581_inst.spi_inst.is_write_cmd ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _9137_ (.RESET_B(net1648),
    .D(_0396_),
    .Q(\tt6581_inst.svf_inst.reg_low[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9138_ (.RESET_B(net1647),
    .D(net1697),
    .Q(\tt6581_inst.svf_inst.reg_low[1] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _9139_ (.RESET_B(net1642),
    .D(_0398_),
    .Q(\tt6581_inst.svf_inst.reg_low[2] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _9140_ (.RESET_B(net1642),
    .D(_0399_),
    .Q(\tt6581_inst.svf_inst.reg_low[3] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _9141_ (.RESET_B(net1640),
    .D(_0400_),
    .Q(\tt6581_inst.svf_inst.reg_low[4] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _9142_ (.RESET_B(net1640),
    .D(_0401_),
    .Q(\tt6581_inst.svf_inst.reg_low[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _9143_ (.RESET_B(net1626),
    .D(_0402_),
    .Q(\tt6581_inst.svf_inst.reg_low[6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9144_ (.RESET_B(net1626),
    .D(_0403_),
    .Q(\tt6581_inst.svf_inst.reg_low[7] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9145_ (.RESET_B(net1625),
    .D(net1129),
    .Q(\tt6581_inst.svf_inst.reg_low[8] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _9146_ (.RESET_B(net1624),
    .D(net1694),
    .Q(\tt6581_inst.svf_inst.reg_low[9] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _9147_ (.RESET_B(net1624),
    .D(net1119),
    .Q(\tt6581_inst.svf_inst.reg_low[10] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _9148_ (.RESET_B(net1574),
    .D(net1078),
    .Q(\tt6581_inst.svf_inst.reg_low[11] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _9149_ (.RESET_B(net1574),
    .D(net1117),
    .Q(\tt6581_inst.svf_inst.reg_low[12] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _9150_ (.RESET_B(net1572),
    .D(net1043),
    .Q(\tt6581_inst.svf_inst.reg_low[13] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _9151_ (.RESET_B(net1572),
    .D(_0410_),
    .Q(\tt6581_inst.svf_inst.reg_low[14] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _9152_ (.RESET_B(net1572),
    .D(net1104),
    .Q(\tt6581_inst.svf_inst.reg_low[15] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _9153_ (.RESET_B(net1558),
    .D(_0412_),
    .Q(\tt6581_inst.svf_inst.reg_low[16] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9154_ (.RESET_B(net1558),
    .D(net1035),
    .Q(\tt6581_inst.svf_inst.reg_low[17] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _9155_ (.RESET_B(net1558),
    .D(_0414_),
    .Q(\tt6581_inst.svf_inst.reg_low[18] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _9156_ (.RESET_B(net1559),
    .D(net1102),
    .Q(\tt6581_inst.svf_inst.reg_low[19] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _9157_ (.RESET_B(net1559),
    .D(net1114),
    .Q(\tt6581_inst.svf_inst.reg_low[20] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _9158_ (.RESET_B(net1559),
    .D(net1045),
    .Q(\tt6581_inst.svf_inst.reg_low[21] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _9159_ (.RESET_B(net1566),
    .D(net1082),
    .Q(\tt6581_inst.svf_inst.reg_low[22] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _9160_ (.RESET_B(net1566),
    .D(net1025),
    .Q(\tt6581_inst.svf_inst.reg_low[23] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _9161_ (.RESET_B(net1634),
    .D(_0420_),
    .Q(\tt6581_inst.svf_inst.reg_band[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _9162_ (.RESET_B(net1634),
    .D(net829),
    .Q(\tt6581_inst.svf_inst.reg_band[1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _9163_ (.RESET_B(net1627),
    .D(_0422_),
    .Q(\tt6581_inst.svf_inst.reg_band[2] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9164_ (.RESET_B(net1627),
    .D(net562),
    .Q(\tt6581_inst.svf_inst.reg_band[3] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9165_ (.RESET_B(net1626),
    .D(net372),
    .Q(\tt6581_inst.svf_inst.reg_band[4] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9166_ (.RESET_B(net1626),
    .D(net856),
    .Q(\tt6581_inst.svf_inst.reg_band[5] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _9167_ (.RESET_B(net1626),
    .D(_0426_),
    .Q(\tt6581_inst.svf_inst.reg_band[6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9168_ (.RESET_B(net1624),
    .D(net431),
    .Q(\tt6581_inst.svf_inst.reg_band[7] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _9169_ (.RESET_B(net1624),
    .D(_0428_),
    .Q(\tt6581_inst.svf_inst.reg_band[8] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _9170_ (.RESET_B(net1624),
    .D(net820),
    .Q(\tt6581_inst.svf_inst.reg_band[9] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _9171_ (.RESET_B(net1574),
    .D(net914),
    .Q(\tt6581_inst.svf_inst.reg_band[10] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _9172_ (.RESET_B(net1576),
    .D(net729),
    .Q(\tt6581_inst.svf_inst.reg_band[11] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _9173_ (.RESET_B(net1574),
    .D(net644),
    .Q(\tt6581_inst.svf_inst.reg_band[12] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _9174_ (.RESET_B(net1572),
    .D(net938),
    .Q(\tt6581_inst.svf_inst.reg_band[13] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _9175_ (.RESET_B(net1573),
    .D(net863),
    .Q(\tt6581_inst.svf_inst.reg_band[14] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _9176_ (.RESET_B(net1572),
    .D(net877),
    .Q(\tt6581_inst.svf_inst.reg_band[15] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _9177_ (.RESET_B(net1573),
    .D(net790),
    .Q(\tt6581_inst.svf_inst.reg_band[16] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _9178_ (.RESET_B(net1558),
    .D(net537),
    .Q(\tt6581_inst.svf_inst.reg_band[17] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _9179_ (.RESET_B(net1558),
    .D(_0438_),
    .Q(\tt6581_inst.svf_inst.reg_band[18] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _9180_ (.RESET_B(net1559),
    .D(_0439_),
    .Q(\tt6581_inst.svf_inst.reg_band[19] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _9181_ (.RESET_B(net1559),
    .D(net1050),
    .Q(\tt6581_inst.svf_inst.reg_band[20] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _9182_ (.RESET_B(net1567),
    .D(net922),
    .Q(\tt6581_inst.svf_inst.reg_band[21] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _9183_ (.RESET_B(net1567),
    .D(_0442_),
    .Q(\tt6581_inst.svf_inst.reg_band[22] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _9184_ (.RESET_B(net1566),
    .D(net92),
    .Q(\tt6581_inst.svf_inst.reg_band[23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _9185_ (.RESET_B(net1650),
    .D(\tt6581_inst.envelope_inst.nxt_state[0] ),
    .Q(\tt6581_inst.envelope_inst.cur_state[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9186_ (.RESET_B(net1650),
    .D(\tt6581_inst.envelope_inst.nxt_state[1] ),
    .Q(\tt6581_inst.envelope_inst.cur_state[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _9187_ (.RESET_B(net1675),
    .D(net284),
    .Q(_0040_),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9188_ (.RESET_B(net1675),
    .D(_0445_),
    .Q(_0041_),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9189_ (.RESET_B(net1683),
    .D(_0446_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9190_ (.RESET_B(net1685),
    .D(_0447_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9191_ (.RESET_B(net1682),
    .D(_0448_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9192_ (.RESET_B(net1685),
    .D(_0449_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9193_ (.RESET_B(net1682),
    .D(_0450_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9194_ (.RESET_B(net1686),
    .D(_0451_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9195_ (.RESET_B(net1686),
    .D(_0452_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9196_ (.RESET_B(net1687),
    .D(_0453_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9197_ (.RESET_B(net1684),
    .D(_0454_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][8] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9198_ (.RESET_B(net1687),
    .D(_0455_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9199_ (.RESET_B(net1678),
    .D(_0456_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][10] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9200_ (.RESET_B(net1687),
    .D(_0457_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][11] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9201_ (.RESET_B(net1680),
    .D(_0458_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][12] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9202_ (.RESET_B(net1680),
    .D(_0459_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _9203_ (.RESET_B(net1678),
    .D(_0460_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][14] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9204_ (.RESET_B(net1680),
    .D(_0461_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][15] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _9205_ (.RESET_B(net1678),
    .D(_0462_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][16] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9206_ (.RESET_B(net1677),
    .D(_0463_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][17] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9207_ (.RESET_B(net1673),
    .D(_0464_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _9208_ (.RESET_B(net1677),
    .D(_0465_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9209_ (.RESET_B(net1682),
    .D(_0466_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][20] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9210_ (.RESET_B(net1677),
    .D(_0467_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][21] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9211_ (.RESET_B(net1675),
    .D(_0468_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][22] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _9212_ (.RESET_B(net1676),
    .D(_0469_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[0][23] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9213_ (.RESET_B(net1675),
    .D(net144),
    .Q(_0042_),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9214_ (.RESET_B(net1675),
    .D(_0471_),
    .Q(_0043_),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9215_ (.RESET_B(net1683),
    .D(_0472_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9216_ (.RESET_B(net1685),
    .D(_0473_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9217_ (.RESET_B(net1682),
    .D(_0474_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][2] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9218_ (.RESET_B(net1685),
    .D(_0475_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9219_ (.RESET_B(net1682),
    .D(_0476_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9220_ (.RESET_B(net1686),
    .D(_0477_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9221_ (.RESET_B(net1686),
    .D(_0478_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9222_ (.RESET_B(net1685),
    .D(_0479_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9223_ (.RESET_B(net1684),
    .D(_0480_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][8] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9224_ (.RESET_B(net1687),
    .D(_0481_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9225_ (.RESET_B(net1678),
    .D(_0482_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][10] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9226_ (.RESET_B(net1687),
    .D(_0483_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][11] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9227_ (.RESET_B(net1680),
    .D(_0484_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][12] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9228_ (.RESET_B(net1687),
    .D(_0485_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][13] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9229_ (.RESET_B(net1678),
    .D(_0486_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9230_ (.RESET_B(net1680),
    .D(_0487_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][15] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9231_ (.RESET_B(net1679),
    .D(_0488_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][16] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9232_ (.RESET_B(net1679),
    .D(_0489_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][17] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9233_ (.RESET_B(net1673),
    .D(_0490_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _9234_ (.RESET_B(net1677),
    .D(_0491_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9235_ (.RESET_B(net1682),
    .D(_0492_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][20] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9236_ (.RESET_B(net1677),
    .D(_0493_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][21] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9237_ (.RESET_B(net1676),
    .D(_0494_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][22] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9238_ (.RESET_B(net1676),
    .D(_0495_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[1][23] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9239_ (.RESET_B(net1683),
    .D(_0496_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9240_ (.RESET_B(net1685),
    .D(_0497_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9241_ (.RESET_B(net1682),
    .D(_0498_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][2] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9242_ (.RESET_B(net1685),
    .D(_0499_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9243_ (.RESET_B(net1683),
    .D(_0500_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _9244_ (.RESET_B(net1686),
    .D(_0501_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _9245_ (.RESET_B(net1686),
    .D(_0502_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9246_ (.RESET_B(net1685),
    .D(_0503_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _9247_ (.RESET_B(net1684),
    .D(_0504_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][8] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9248_ (.RESET_B(net1687),
    .D(_0505_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9249_ (.RESET_B(net1678),
    .D(_0506_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][10] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9250_ (.RESET_B(net1687),
    .D(_0507_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][11] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _9251_ (.RESET_B(net1680),
    .D(_0508_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][12] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9252_ (.RESET_B(net1681),
    .D(_0509_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _9253_ (.RESET_B(net1678),
    .D(_0510_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9254_ (.RESET_B(net1680),
    .D(_0511_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][15] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _9255_ (.RESET_B(net1678),
    .D(_0512_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][16] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _9256_ (.RESET_B(net1677),
    .D(_0513_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][17] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9257_ (.RESET_B(net1673),
    .D(_0514_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _9258_ (.RESET_B(net1677),
    .D(_0515_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9259_ (.RESET_B(net1682),
    .D(_0516_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][20] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _9260_ (.RESET_B(net1677),
    .D(_0517_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][21] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9261_ (.RESET_B(net1675),
    .D(_0518_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][22] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _9262_ (.RESET_B(net1676),
    .D(_0519_),
    .Q(\tt6581_inst.envelope_inst.vol_regs[2][23] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _9263_ (.RESET_B(net1652),
    .D(net41),
    .Q(\tt6581_inst.multi_voice_inst.cur_state[0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _9264_ (.RESET_B(net1652),
    .D(net48),
    .Q(\tt6581_inst.multi_voice_inst.cur_state[1] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _9265_ (.RESET_B(net1651),
    .D(_0024_),
    .Q(\tt6581_inst.controller_inst.voice_ready_i ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _9266_ (.RESET_B(net1629),
    .D(_0520_),
    .Q(\tt6581_inst.mult_inst.neg_result ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _9267_ (.RESET_B(net1600),
    .D(_0521_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _9268_ (.RESET_B(net1600),
    .D(_0522_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9269_ (.RESET_B(net1600),
    .D(_0523_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9270_ (.RESET_B(net1597),
    .D(_0524_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9271_ (.RESET_B(net1597),
    .D(_0525_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _9272_ (.RESET_B(net1594),
    .D(_0526_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9273_ (.RESET_B(net1595),
    .D(_0527_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _9274_ (.RESET_B(net1589),
    .D(_0528_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _9275_ (.RESET_B(net1589),
    .D(_0529_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][8] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9276_ (.RESET_B(net1588),
    .D(_0530_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9277_ (.RESET_B(net1587),
    .D(_0531_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9278_ (.RESET_B(net1593),
    .D(_0532_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9279_ (.RESET_B(net1568),
    .D(_0533_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9280_ (.RESET_B(net1568),
    .D(_0534_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][13] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9281_ (.RESET_B(net1579),
    .D(_0535_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9282_ (.RESET_B(net1579),
    .D(_0536_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9283_ (.RESET_B(net1579),
    .D(_0537_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _9284_ (.RESET_B(net1585),
    .D(_0538_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[0][17] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9285_ (.RESET_B(net1600),
    .D(_0539_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9286_ (.RESET_B(net1600),
    .D(_0540_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9287_ (.RESET_B(net1600),
    .D(_0541_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9288_ (.RESET_B(net1597),
    .D(_0542_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9289_ (.RESET_B(net1597),
    .D(_0543_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _9290_ (.RESET_B(net1597),
    .D(_0544_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9291_ (.RESET_B(net1595),
    .D(_0545_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _9292_ (.RESET_B(net1595),
    .D(_0546_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9293_ (.RESET_B(net1590),
    .D(_0547_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][8] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9294_ (.RESET_B(net1585),
    .D(_0548_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][9] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9295_ (.RESET_B(net1587),
    .D(_0549_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9296_ (.RESET_B(net1593),
    .D(_0550_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9297_ (.RESET_B(net1568),
    .D(_0551_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9298_ (.RESET_B(net1568),
    .D(_0552_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][13] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9299_ (.RESET_B(net1579),
    .D(_0553_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9300_ (.RESET_B(net1580),
    .D(_0554_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][15] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _9301_ (.RESET_B(net1579),
    .D(_0555_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _9302_ (.RESET_B(net1585),
    .D(_0556_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[1][17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9303_ (.RESET_B(net1601),
    .D(_0557_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9304_ (.RESET_B(net1600),
    .D(_0558_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9305_ (.RESET_B(net1600),
    .D(_0559_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9306_ (.RESET_B(net1597),
    .D(_0560_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9307_ (.RESET_B(net1597),
    .D(_0561_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _9308_ (.RESET_B(net1601),
    .D(_0562_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9309_ (.RESET_B(net1599),
    .D(_0563_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _9310_ (.RESET_B(net1589),
    .D(_0564_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _9311_ (.RESET_B(net1587),
    .D(_0565_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][8] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _9312_ (.RESET_B(net1587),
    .D(_0566_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9313_ (.RESET_B(net1587),
    .D(_0567_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9314_ (.RESET_B(net1593),
    .D(_0568_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][11] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _9315_ (.RESET_B(net1568),
    .D(_0569_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9316_ (.RESET_B(net1568),
    .D(_0570_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9317_ (.RESET_B(net1579),
    .D(_0571_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9318_ (.RESET_B(net1579),
    .D(_0572_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _9319_ (.RESET_B(net1579),
    .D(_0573_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _9320_ (.RESET_B(net1585),
    .D(_0574_),
    .Q(\tt6581_inst.multi_voice_inst.phase_regs[2][17] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9321_ (.RESET_B(net1588),
    .D(_0575_),
    .Q(_0044_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9322_ (.RESET_B(net1586),
    .D(_0576_),
    .Q(_0045_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9323_ (.RESET_B(net1563),
    .D(_0577_),
    .Q(_0046_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9324_ (.RESET_B(net1563),
    .D(_0578_),
    .Q(_0047_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9325_ (.RESET_B(net1560),
    .D(_0579_),
    .Q(_0048_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9326_ (.RESET_B(net1563),
    .D(_0580_),
    .Q(_0049_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9327_ (.RESET_B(net1564),
    .D(_0581_),
    .Q(_0050_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9328_ (.RESET_B(net1561),
    .D(_0582_),
    .Q(_0051_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9329_ (.RESET_B(net1568),
    .D(_0583_),
    .Q(_0052_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9330_ (.RESET_B(net1569),
    .D(_0584_),
    .Q(_0053_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9331_ (.RESET_B(net1566),
    .D(_0585_),
    .Q(_0054_),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _9332_ (.RESET_B(net1568),
    .D(_0586_),
    .Q(_0055_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9333_ (.RESET_B(net1564),
    .D(_0587_),
    .Q(_0056_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9334_ (.RESET_B(net1564),
    .D(_0588_),
    .Q(_0057_),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9335_ (.RESET_B(net1563),
    .D(_0589_),
    .Q(_0058_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9336_ (.RESET_B(net1586),
    .D(_0590_),
    .Q(_0059_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9337_ (.RESET_B(net1588),
    .D(_0591_),
    .Q(_0060_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9338_ (.RESET_B(net1588),
    .D(_0592_),
    .Q(_0061_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9339_ (.RESET_B(net1595),
    .D(_0593_),
    .Q(_0062_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9340_ (.RESET_B(net1594),
    .D(_0594_),
    .Q(_0063_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9341_ (.RESET_B(net1594),
    .D(_0595_),
    .Q(_0064_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9342_ (.RESET_B(net1594),
    .D(_0596_),
    .Q(_0065_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9343_ (.RESET_B(net1595),
    .D(_0597_),
    .Q(_0066_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9344_ (.RESET_B(net1588),
    .D(_0598_),
    .Q(_0067_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9345_ (.RESET_B(net1585),
    .D(_0599_),
    .Q(_0068_),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9346_ (.RESET_B(net1585),
    .D(net201),
    .Q(_0069_),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9347_ (.RESET_B(net1563),
    .D(_0601_),
    .Q(_0070_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9348_ (.RESET_B(net1561),
    .D(_0602_),
    .Q(_0071_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9349_ (.RESET_B(net1563),
    .D(_0603_),
    .Q(_0072_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9350_ (.RESET_B(net1564),
    .D(_0604_),
    .Q(_0073_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9351_ (.RESET_B(net1561),
    .D(_0605_),
    .Q(_0074_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9352_ (.RESET_B(net1567),
    .D(_0606_),
    .Q(_0075_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9353_ (.RESET_B(net1569),
    .D(_0607_),
    .Q(_0076_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9354_ (.RESET_B(net1566),
    .D(_0608_),
    .Q(_0077_),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _9355_ (.RESET_B(net1566),
    .D(_0609_),
    .Q(_0078_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9356_ (.RESET_B(net1564),
    .D(_0610_),
    .Q(_0079_),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9357_ (.RESET_B(net1564),
    .D(_0611_),
    .Q(_0080_),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _9358_ (.RESET_B(net1565),
    .D(_0612_),
    .Q(_0081_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9359_ (.RESET_B(net1586),
    .D(_0613_),
    .Q(_0082_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9360_ (.RESET_B(net1589),
    .D(_0614_),
    .Q(_0083_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9361_ (.RESET_B(net1588),
    .D(_0615_),
    .Q(_0084_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9362_ (.RESET_B(net1596),
    .D(_0616_),
    .Q(_0085_),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _9363_ (.RESET_B(net1594),
    .D(_0617_),
    .Q(_0086_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9364_ (.RESET_B(net1596),
    .D(_0618_),
    .Q(_0087_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9365_ (.RESET_B(net1594),
    .D(_0619_),
    .Q(_0088_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9366_ (.RESET_B(net1595),
    .D(_0620_),
    .Q(_0089_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9367_ (.RESET_B(net1588),
    .D(_0621_),
    .Q(_0090_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9368_ (.RESET_B(net1585),
    .D(_0622_),
    .Q(_0091_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9369_ (.RESET_B(net1585),
    .D(net182),
    .Q(_0092_),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9370_ (.RESET_B(net1563),
    .D(_0624_),
    .Q(_0093_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9371_ (.RESET_B(net1561),
    .D(_0625_),
    .Q(_0094_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9372_ (.RESET_B(net1563),
    .D(_0626_),
    .Q(_0095_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _9373_ (.RESET_B(net1564),
    .D(_0627_),
    .Q(_0096_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9374_ (.RESET_B(net1561),
    .D(_0628_),
    .Q(_0097_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9375_ (.RESET_B(net1567),
    .D(_0629_),
    .Q(_0098_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9376_ (.RESET_B(net1569),
    .D(_0630_),
    .Q(_0099_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9377_ (.RESET_B(net1567),
    .D(_0631_),
    .Q(_0100_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _9378_ (.RESET_B(net1569),
    .D(_0632_),
    .Q(_0101_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _9379_ (.RESET_B(net1564),
    .D(_0633_),
    .Q(_0102_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9380_ (.RESET_B(net1565),
    .D(_0634_),
    .Q(_0103_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9381_ (.RESET_B(net1565),
    .D(_0635_),
    .Q(_0104_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _9382_ (.RESET_B(net1586),
    .D(_0636_),
    .Q(_0105_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _9383_ (.RESET_B(net1589),
    .D(_0637_),
    .Q(_0106_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9384_ (.RESET_B(net1588),
    .D(_0638_),
    .Q(_0107_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9385_ (.RESET_B(net1595),
    .D(_0639_),
    .Q(_0108_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9386_ (.RESET_B(net1596),
    .D(_0640_),
    .Q(_0109_),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _9387_ (.RESET_B(net1594),
    .D(_0641_),
    .Q(_0110_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9388_ (.RESET_B(net1594),
    .D(_0642_),
    .Q(_0111_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _9389_ (.RESET_B(net1595),
    .D(_0643_),
    .Q(_0112_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _9390_ (.RESET_B(net1587),
    .D(_0644_),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[0][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _9391_ (.RESET_B(net1589),
    .D(net148),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[0][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9392_ (.RESET_B(net1590),
    .D(_0646_),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[1][0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9393_ (.RESET_B(net1592),
    .D(net137),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[1][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _9394_ (.RESET_B(net1648),
    .D(\tt6581_inst.controller_inst.cur_state[0] ),
    .Q(\tt6581_inst.accum_rst ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9395_ (.RESET_B(net1649),
    .D(net31),
    .Q(\tt6581_inst.audio_valid ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9396_ (.RESET_B(net1650),
    .D(net34),
    .Q(\tt6581_inst.accum_en ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _9397_ (.RESET_B(net1636),
    .D(net32),
    .Q(\tt6581_inst.controller_inst.filt_start_o ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _9398_ (.RESET_B(net1650),
    .D(_0019_),
    .Q(\tt6581_inst.accum_in_mux ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _9399_ (.RESET_B(net1649),
    .D(net125),
    .Q(\tt6581_inst.filter_accum[0] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _9400_ (.RESET_B(net1649),
    .D(net956),
    .Q(\tt6581_inst.filter_accum[1] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _9401_ (.RESET_B(net1642),
    .D(net1012),
    .Q(\tt6581_inst.filter_accum[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _9402_ (.RESET_B(net1642),
    .D(_0651_),
    .Q(\tt6581_inst.filter_accum[3] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _9403_ (.RESET_B(net1642),
    .D(_0652_),
    .Q(\tt6581_inst.filter_accum[4] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9404_ (.RESET_B(net1640),
    .D(net1055),
    .Q(\tt6581_inst.filter_accum[5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9405_ (.RESET_B(net1641),
    .D(net476),
    .Q(\tt6581_inst.filter_accum[6] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9406_ (.RESET_B(net1641),
    .D(_0655_),
    .Q(\tt6581_inst.filter_accum[7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9407_ (.RESET_B(net1641),
    .D(_0656_),
    .Q(\tt6581_inst.filter_accum[8] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9408_ (.RESET_B(net1641),
    .D(net1121),
    .Q(\tt6581_inst.filter_accum[9] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _9409_ (.RESET_B(net1640),
    .D(net647),
    .Q(\tt6581_inst.filter_accum[10] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _9410_ (.RESET_B(net1640),
    .D(net1109),
    .Q(\tt6581_inst.filter_accum[11] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _9411_ (.RESET_B(net1640),
    .D(net1020),
    .Q(\tt6581_inst.filter_accum[12] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _9412_ (.RESET_B(net1640),
    .D(net1131),
    .Q(\tt6581_inst.filter_accum[13] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _9413_ (.RESET_B(net1637),
    .D(_0116_),
    .Q(_0113_),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _9414_ (.RESET_B(net1637),
    .D(_0014_),
    .Q(\tt6581_inst.controller_inst.mult_in_mux_o[1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _9415_ (.RESET_B(net1636),
    .D(_0015_),
    .Q(\tt6581_inst.controller_inst.mult_in_mux_o[2] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _9416_ (.RESET_B(net1651),
    .D(net29),
    .Q(\tt6581_inst.controller_inst.voice_start_o ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _9417_ (.RESET_B(net1651),
    .D(net30),
    .Q(\tt6581_inst.controller_inst.env_start_o ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _9418_ (.RESET_B(net1635),
    .D(net33),
    .Q(\tt6581_inst.controller_inst.mult_start_o ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _9419_ (.RESET_B(net1581),
    .D(net1124),
    .Q(\tt6581_inst.filt_en_mode[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _9420_ (.RESET_B(net1581),
    .D(_0663_),
    .Q(\tt6581_inst.filt_en_mode[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9421_ (.RESET_B(net1582),
    .D(_0664_),
    .Q(\tt6581_inst.filt_en_mode[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9422_ (.RESET_B(net1608),
    .D(net594),
    .Q(\tt6581_inst.controller_inst.filt_en_i[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _9423_ (.RESET_B(net1581),
    .D(net874),
    .Q(\tt6581_inst.controller_inst.filt_en_i[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _9424_ (.RESET_B(net1581),
    .D(_0667_),
    .Q(\tt6581_inst.controller_inst.filt_en_i[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _9425_ (.RESET_B(net1609),
    .D(_0668_),
    .Q(\tt6581_inst.filt_en_mode[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _9426_ (.RESET_B(net1610),
    .D(net358),
    .Q(\tt6581_inst.filt_en_mode[7] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _9427_ (.RESET_B(net1590),
    .D(_0670_),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[2][0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _9428_ (.RESET_B(net1589),
    .D(net142),
    .Q(\tt6581_inst.multi_voice_inst.phase_last_msb[2][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _9429_ (.RESET_B(net1660),
    .D(net891),
    .Q(\tt6581_inst.filt_f_lo[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _9430_ (.RESET_B(net1662),
    .D(net773),
    .Q(\tt6581_inst.filt_f_lo[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _9431_ (.RESET_B(net1666),
    .D(net925),
    .Q(\tt6581_inst.filt_f_lo[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _9432_ (.RESET_B(net1663),
    .D(net796),
    .Q(\tt6581_inst.filt_f_lo[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _9433_ (.RESET_B(net1667),
    .D(net705),
    .Q(\tt6581_inst.filt_f_lo[4] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _9434_ (.RESET_B(net1666),
    .D(net811),
    .Q(\tt6581_inst.filt_f_lo[5] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _9435_ (.RESET_B(net1659),
    .D(_0678_),
    .Q(\tt6581_inst.filt_f_lo[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _9436_ (.RESET_B(net1659),
    .D(_0679_),
    .Q(\tt6581_inst.filt_f_lo[7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _9437_ (.RESET_B(net1598),
    .D(net887),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[16] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _9438_ (.RESET_B(net1599),
    .D(net564),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[17] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _9439_ (.RESET_B(net1617),
    .D(net547),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[18] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _9440_ (.RESET_B(net1617),
    .D(net1018),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[19] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _9441_ (.RESET_B(net1599),
    .D(net528),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[20] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _9442_ (.RESET_B(net1599),
    .D(net670),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _9443_ (.RESET_B(net1612),
    .D(net522),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[22] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _9444_ (.RESET_B(net1598),
    .D(net719),
    .Q(\tt6581_inst.controller_inst.freq_lo_i[23] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _9445_ (.RESET_B(net1602),
    .D(net494),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[16] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _9446_ (.RESET_B(net1593),
    .D(net455),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[17] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _9447_ (.RESET_B(net1606),
    .D(_0690_),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[18] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _9448_ (.RESET_B(net1607),
    .D(net448),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[19] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _9449_ (.RESET_B(net1608),
    .D(net1023),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[20] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _9450_ (.RESET_B(net1602),
    .D(net993),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[21] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _9451_ (.RESET_B(net1608),
    .D(net895),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[22] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _9452_ (.RESET_B(net1593),
    .D(_0695_),
    .Q(\tt6581_inst.controller_inst.freq_hi_i[23] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _9453_ (.RESET_B(net1659),
    .D(net605),
    .Q(\tt6581_inst.filt_q_hi[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _9454_ (.RESET_B(net1661),
    .D(net743),
    .Q(\tt6581_inst.filt_q_hi[1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _9455_ (.RESET_B(net1608),
    .D(_0698_),
    .Q(\tt6581_inst.filt_q_hi[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9456_ (.RESET_B(net1661),
    .D(net624),
    .Q(\tt6581_inst.filt_q_hi[3] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _9457_ (.RESET_B(net1661),
    .D(_0700_),
    .Q(\tt6581_inst.filt_q_hi[4] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9458_ (.RESET_B(net1659),
    .D(_0701_),
    .Q(\tt6581_inst.filt_q_hi[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _9459_ (.RESET_B(net1659),
    .D(_0702_),
    .Q(\tt6581_inst.filt_q_hi[6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _9460_ (.RESET_B(net1661),
    .D(net684),
    .Q(\tt6581_inst.filt_q_hi[7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _9461_ (.RESET_B(net1592),
    .D(net615),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[16] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _9462_ (.RESET_B(net1592),
    .D(_0705_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[17] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _9463_ (.RESET_B(net1609),
    .D(_0706_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[18] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _9464_ (.RESET_B(net1610),
    .D(_0707_),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[19] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _9465_ (.RESET_B(net1592),
    .D(net549),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[20] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _9466_ (.RESET_B(net1591),
    .D(net654),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _9467_ (.RESET_B(net1604),
    .D(net367),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[22] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _9468_ (.RESET_B(net1591),
    .D(net682),
    .Q(\tt6581_inst.controller_inst.pw_lo_i[23] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _9469_ (.RESET_B(net1609),
    .D(net897),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[16] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _9470_ (.RESET_B(net1605),
    .D(_0713_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[17] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _9471_ (.RESET_B(net1607),
    .D(_0714_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[18] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _9472_ (.RESET_B(net1606),
    .D(net588),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[19] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _9473_ (.RESET_B(net1606),
    .D(net498),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[20] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _9474_ (.RESET_B(net1608),
    .D(_0717_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[21] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _9475_ (.RESET_B(net1660),
    .D(_0718_),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[22] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _9476_ (.RESET_B(net1660),
    .D(net320),
    .Q(\tt6581_inst.controller_inst.pw_hi_i[23] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _9477_ (.RESET_B(net1669),
    .D(_0720_),
    .Q(\tt6581_inst.control_pack[16] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _9478_ (.RESET_B(net1598),
    .D(_0721_),
    .Q(\tt6581_inst.control_pack[17] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _9479_ (.RESET_B(net1616),
    .D(_0722_),
    .Q(\tt6581_inst.control_pack[18] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _9480_ (.RESET_B(net1617),
    .D(_0723_),
    .Q(\tt6581_inst.control_pack[19] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _9481_ (.RESET_B(net1612),
    .D(net617),
    .Q(\tt6581_inst.control_pack[20] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _9482_ (.RESET_B(net1604),
    .D(net982),
    .Q(\tt6581_inst.control_pack[21] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _9483_ (.RESET_B(net1603),
    .D(net613),
    .Q(\tt6581_inst.control_pack[22] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _9484_ (.RESET_B(net1603),
    .D(_0727_),
    .Q(\tt6581_inst.control_pack[23] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _9485_ (.RESET_B(net1663),
    .D(_0728_),
    .Q(\tt6581_inst.filt_q_lo[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _9486_ (.RESET_B(net1662),
    .D(net770),
    .Q(\tt6581_inst.filt_q_lo[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _9487_ (.RESET_B(net1664),
    .D(net1004),
    .Q(\tt6581_inst.filt_q_lo[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _9488_ (.RESET_B(net1663),
    .D(net834),
    .Q(\tt6581_inst.filt_q_lo[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _9489_ (.RESET_B(net1662),
    .D(_0732_),
    .Q(\tt6581_inst.filt_q_lo[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _9490_ (.RESET_B(net1662),
    .D(_0733_),
    .Q(\tt6581_inst.filt_q_lo[5] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _9491_ (.RESET_B(net1663),
    .D(_0734_),
    .Q(\tt6581_inst.filt_q_lo[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _9492_ (.RESET_B(net1663),
    .D(net731),
    .Q(\tt6581_inst.filt_q_lo[7] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _9493_ (.RESET_B(net1670),
    .D(net858),
    .Q(\tt6581_inst.ad_pack[16] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _9494_ (.RESET_B(net1670),
    .D(_0737_),
    .Q(\tt6581_inst.ad_pack[17] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _9495_ (.RESET_B(net1673),
    .D(net986),
    .Q(\tt6581_inst.ad_pack[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _9496_ (.RESET_B(net1670),
    .D(net1063),
    .Q(\tt6581_inst.ad_pack[19] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _9497_ (.RESET_B(net1662),
    .D(net291),
    .Q(\tt6581_inst.ad_pack[20] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _9498_ (.RESET_B(net1672),
    .D(net661),
    .Q(\tt6581_inst.ad_pack[21] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _9499_ (.RESET_B(net1666),
    .D(_0742_),
    .Q(\tt6581_inst.ad_pack[22] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _9500_ (.RESET_B(net1662),
    .D(net899),
    .Q(\tt6581_inst.ad_pack[23] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _9501_ (.RESET_B(net1659),
    .D(net916),
    .Q(\tt6581_inst.filt_f_hi[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9502_ (.RESET_B(net1661),
    .D(_0745_),
    .Q(\tt6581_inst.filt_f_hi[1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9503_ (.RESET_B(net1631),
    .D(_0746_),
    .Q(\tt6581_inst.filt_f_hi[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9504_ (.RESET_B(net1659),
    .D(net919),
    .Q(\tt6581_inst.filt_f_hi[3] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _9505_ (.RESET_B(net1661),
    .D(_0748_),
    .Q(\tt6581_inst.filt_f_hi[4] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9506_ (.RESET_B(net1631),
    .D(_0749_),
    .Q(\tt6581_inst.filt_f_hi[5] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _9507_ (.RESET_B(net1659),
    .D(_0750_),
    .Q(\tt6581_inst.filt_f_hi[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _9508_ (.RESET_B(net1660),
    .D(net794),
    .Q(\tt6581_inst.filt_f_hi[7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _9509_ (.RESET_B(net1669),
    .D(_0752_),
    .Q(\tt6581_inst.controller_inst.sr_i[16] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _9510_ (.RESET_B(net1670),
    .D(net659),
    .Q(\tt6581_inst.controller_inst.sr_i[17] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _9511_ (.RESET_B(net1669),
    .D(net884),
    .Q(\tt6581_inst.controller_inst.sr_i[18] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _9512_ (.RESET_B(net1669),
    .D(net703),
    .Q(\tt6581_inst.controller_inst.sr_i[19] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _9513_ (.RESET_B(net1663),
    .D(net778),
    .Q(\tt6581_inst.controller_inst.sr_i[20] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _9514_ (.RESET_B(net1665),
    .D(net1112),
    .Q(\tt6581_inst.controller_inst.sr_i[21] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _9515_ (.RESET_B(net1673),
    .D(_0758_),
    .Q(\tt6581_inst.controller_inst.sr_i[22] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _9516_ (.RESET_B(net1665),
    .D(net944),
    .Q(\tt6581_inst.controller_inst.sr_i[23] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _9517_ (.RESET_B(net1614),
    .D(net2),
    .Q(\tt6581_inst.spi_inst.mosi_sync[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _9518_ (.RESET_B(net1614),
    .D(net28),
    .Q(\tt6581_inst.spi_inst.mosi_sync[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _9519_ (.RESET_B(net1667),
    .D(net652),
    .Q(\tt6581_inst.filt_volume[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _9520_ (.RESET_B(net1667),
    .D(_0761_),
    .Q(\tt6581_inst.filt_volume[1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9521_ (.RESET_B(net1667),
    .D(net840),
    .Q(\tt6581_inst.filt_volume[2] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9522_ (.RESET_B(net1664),
    .D(net714),
    .Q(\tt6581_inst.filt_volume[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9523_ (.RESET_B(net1667),
    .D(_0764_),
    .Q(\tt6581_inst.filt_volume[4] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _9524_ (.RESET_B(net1667),
    .D(net780),
    .Q(\tt6581_inst.filt_volume[5] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _9525_ (.RESET_B(net1667),
    .D(net733),
    .Q(\tt6581_inst.filt_volume[6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _9526_ (.RESET_B(net1664),
    .D(net909),
    .Q(\tt6581_inst.filt_volume[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _9527_ (.RESET_B(net1618),
    .D(net807),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _9528_ (.RESET_B(net1619),
    .D(_0769_),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _9529_ (.RESET_B(net1618),
    .D(net725),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _9530_ (.RESET_B(net1614),
    .D(_0771_),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _9531_ (.RESET_B(net1613),
    .D(_0772_),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[4] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _9532_ (.RESET_B(net1613),
    .D(net975),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _9533_ (.RESET_B(net1613),
    .D(_0774_),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _9534_ (.RESET_B(net1614),
    .D(_0775_),
    .Q(\tt6581_inst.reg_file_inst.wdata_i[7] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _9535_ (.RESET_B(net1614),
    .D(net1),
    .Q(\tt6581_inst.spi_inst.cs_sync[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _9536_ (.RESET_B(net1618),
    .D(net26),
    .Q(\tt6581_inst.spi_inst.cs_sync[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _9537_ (.RESET_B(net1619),
    .D(net822),
    .Q(\tt6581_inst.reg_addr[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _9538_ (.RESET_B(net1619),
    .D(_0777_),
    .Q(\tt6581_inst.reg_addr[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _9539_ (.RESET_B(net1618),
    .D(net766),
    .Q(\tt6581_inst.reg_addr[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _9540_ (.RESET_B(net1618),
    .D(net813),
    .Q(\tt6581_inst.reg_addr[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _9541_ (.RESET_B(net1619),
    .D(net279),
    .Q(\tt6581_inst.reg_addr[4] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _9542_ (.RESET_B(net1613),
    .D(net532),
    .Q(\tt6581_inst.reg_addr[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _9543_ (.RESET_B(net1615),
    .D(net510),
    .Q(\tt6581_inst.reg_addr[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _9544_ (.RESET_B(net1674),
    .D(net179),
    .Q(\tt6581_inst.spi_inst.data_out_reg[0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _9545_ (.RESET_B(net1671),
    .D(net119),
    .Q(\tt6581_inst.spi_inst.data_out_reg[1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _9546_ (.RESET_B(net1619),
    .D(net109),
    .Q(\tt6581_inst.spi_inst.data_out_reg[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _9547_ (.RESET_B(net1671),
    .D(net95),
    .Q(\tt6581_inst.spi_inst.data_out_reg[3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _9548_ (.RESET_B(net1619),
    .D(net99),
    .Q(\tt6581_inst.spi_inst.data_out_reg[4] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _9549_ (.RESET_B(net1671),
    .D(net90),
    .Q(\tt6581_inst.spi_inst.data_out_reg[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _9550_ (.RESET_B(net1671),
    .D(net106),
    .Q(\tt6581_inst.spi_inst.data_out_reg[6] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _9551_ (.RESET_B(net1620),
    .D(net71),
    .Q(\tt6581_inst.spi_inst.data_out_reg[7] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _9552_ (.RESET_B(net1614),
    .D(_0791_),
    .Q(\tt6581_inst.reg_file_inst.we_i ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _9553_ (.RESET_B(net1619),
    .D(net139),
    .Q(\tt6581_inst.spi_inst.bit_cnt[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _9554_ (.RESET_B(net1619),
    .D(net463),
    .Q(\tt6581_inst.spi_inst.bit_cnt[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _9555_ (.RESET_B(net1620),
    .D(net578),
    .Q(\tt6581_inst.spi_inst.bit_cnt[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _9556_ (.RESET_B(net1620),
    .D(net824),
    .Q(\tt6581_inst.spi_inst.bit_cnt[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _9557_ (.RESET_B(net1614),
    .D(net3),
    .Q(\tt6581_inst.spi_inst.sclk_sync[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _9558_ (.RESET_B(net1614),
    .D(net27),
    .Q(\tt6581_inst.spi_inst.sclk_sync[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _9559_ (.RESET_B(net1618),
    .D(net35),
    .Q(\tt6581_inst.spi_inst.sclk_sync[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _9560_ (.RESET_B(net1620),
    .D(_0796_),
    .Q(\tt6581_inst.spi_inst.shift_reg[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _9561_ (.RESET_B(net1618),
    .D(_0797_),
    .Q(\tt6581_inst.spi_inst.shift_reg[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _9562_ (.RESET_B(net1618),
    .D(_0798_),
    .Q(\tt6581_inst.spi_inst.shift_reg[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _9563_ (.RESET_B(net1615),
    .D(_0799_),
    .Q(\tt6581_inst.spi_inst.shift_reg[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _9564_ (.RESET_B(net1613),
    .D(_0800_),
    .Q(\tt6581_inst.spi_inst.shift_reg[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _9565_ (.RESET_B(net1613),
    .D(net649),
    .Q(\tt6581_inst.spi_inst.shift_reg[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _9566_ (.RESET_B(net1615),
    .D(_0802_),
    .Q(\tt6581_inst.spi_inst.shift_reg[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _9567_ (.RESET_B(net1555),
    .D(_0025_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _9568_ (.RESET_B(net1560),
    .D(_0026_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _9569_ (.RESET_B(net1560),
    .D(_0027_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _9570_ (.RESET_B(net1560),
    .D(_0028_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9571_ (.RESET_B(net1560),
    .D(net68),
    .Q(\tt6581_inst.tick_gen_inst.cnt[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _9572_ (.RESET_B(net1560),
    .D(_0030_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9573_ (.RESET_B(net1560),
    .D(_0031_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9574_ (.RESET_B(net1561),
    .D(_0032_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9575_ (.RESET_B(net1562),
    .D(_0033_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _9576_ (.RESET_B(net1561),
    .D(_0034_),
    .Q(\tt6581_inst.tick_gen_inst.cnt[9] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _9577_ (.RESET_B(net1567),
    .D(net267),
    .Q(\tt6581_inst.controller_inst.sample_tick_i ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _9578_ (.RESET_B(net1644),
    .D(_0803_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _9579_ (.RESET_B(net1644),
    .D(_0804_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[5] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9580_ (.RESET_B(net1644),
    .D(_0805_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[6] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9581_ (.RESET_B(net1644),
    .D(_0806_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9582_ (.RESET_B(net1644),
    .D(_0807_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[8] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _9583_ (.RESET_B(net1653),
    .D(_0808_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[9] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _9584_ (.RESET_B(net1653),
    .D(_0809_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[10] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _9585_ (.RESET_B(net1653),
    .D(_0810_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[11] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _9586_ (.RESET_B(net1653),
    .D(_0811_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[12] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _9587_ (.RESET_B(net1653),
    .D(_0812_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[13] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9588_ (.RESET_B(net1649),
    .D(_0813_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[14] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _9589_ (.RESET_B(net1649),
    .D(_0814_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[15] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _9590_ (.RESET_B(net1651),
    .D(_0815_),
    .Q(\tt6581_inst.delta_sigma_inst.audio[16] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _9591_ (.RESET_B(net1649),
    .D(net63),
    .Q(\tt6581_inst.delta_sigma_inst.audio[17] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _9592_ (.RESET_B(net1634),
    .D(net130),
    .Q(\tt6581_inst.bypass_accum[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _9593_ (.RESET_B(net1634),
    .D(_0818_),
    .Q(\tt6581_inst.bypass_accum[1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _9594_ (.RESET_B(net1635),
    .D(net1080),
    .Q(\tt6581_inst.bypass_accum[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _9595_ (.RESET_B(net1626),
    .D(_0820_),
    .Q(\tt6581_inst.bypass_accum[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _9596_ (.RESET_B(net1627),
    .D(_0821_),
    .Q(\tt6581_inst.bypass_accum[4] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _9597_ (.RESET_B(net1627),
    .D(net1027),
    .Q(\tt6581_inst.bypass_accum[5] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _9598_ (.RESET_B(net1627),
    .D(net360),
    .Q(\tt6581_inst.bypass_accum[6] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _9599_ (.RESET_B(net1625),
    .D(_0824_),
    .Q(\tt6581_inst.bypass_accum[7] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _9600_ (.RESET_B(net1625),
    .D(net481),
    .Q(\tt6581_inst.bypass_accum[8] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _9601_ (.RESET_B(net1625),
    .D(_0826_),
    .Q(\tt6581_inst.bypass_accum[9] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _9602_ (.RESET_B(net1625),
    .D(net518),
    .Q(\tt6581_inst.bypass_accum[10] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _9603_ (.RESET_B(net1575),
    .D(net1073),
    .Q(\tt6581_inst.bypass_accum[11] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _9604_ (.RESET_B(net1625),
    .D(net487),
    .Q(\tt6581_inst.bypass_accum[12] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _9605_ (.RESET_B(net1575),
    .D(net572),
    .Q(\tt6581_inst.bypass_accum[13] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_andreasp00_5 (.L_LO(net5));
 sg13g2_tielo tt_um_andreasp00_6 (.L_LO(net6));
 sg13g2_tielo tt_um_andreasp00_7 (.L_LO(net7));
 sg13g2_tielo tt_um_andreasp00_8 (.L_LO(net8));
 sg13g2_tielo tt_um_andreasp00_9 (.L_LO(net9));
 sg13g2_tielo tt_um_andreasp00_10 (.L_LO(net10));
 sg13g2_tielo tt_um_andreasp00_11 (.L_LO(net11));
 sg13g2_tielo tt_um_andreasp00_12 (.L_LO(net12));
 sg13g2_tielo tt_um_andreasp00_13 (.L_LO(net13));
 sg13g2_tielo tt_um_andreasp00_14 (.L_LO(net14));
 sg13g2_tielo tt_um_andreasp00_15 (.L_LO(net15));
 sg13g2_tielo tt_um_andreasp00_16 (.L_LO(net16));
 sg13g2_tielo tt_um_andreasp00_17 (.L_LO(net17));
 sg13g2_tielo tt_um_andreasp00_18 (.L_LO(net18));
 sg13g2_tielo tt_um_andreasp00_19 (.L_LO(net19));
 sg13g2_tielo tt_um_andreasp00_20 (.L_LO(net20));
 sg13g2_tielo tt_um_andreasp00_21 (.L_LO(net21));
 sg13g2_tielo tt_um_andreasp00_22 (.L_LO(net22));
 sg13g2_tielo tt_um_andreasp00_23 (.L_LO(net23));
 sg13g2_tielo tt_um_andreasp00_24 (.L_LO(net24));
 sg13g2_tiehi tt_um_andreasp00_25 (.L_HI(net25));
 sg13g2_buf_1 _9628_ (.A(miso),
    .X(uio_out[2]));
 sg13g2_buf_8 _9629_ (.A(pdm),
    .X(uo_out[0]));
 sg13g2_buf_8 fanout1135 (.A(_3788_),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_8 fanout1137 (.A(_3733_),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(_3699_),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(_3699_),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(_2230_),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_8 fanout1142 (.A(_2229_),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(_2226_),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(_1882_),
    .X(net1144));
 sg13g2_buf_8 fanout1145 (.A(_1889_),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(net1147),
    .X(net1146));
 sg13g2_buf_8 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_8 fanout1148 (.A(_3965_),
    .X(net1148));
 sg13g2_buf_8 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_8 fanout1150 (.A(_3965_),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_8 fanout1152 (.A(_2065_),
    .X(net1152));
 sg13g2_buf_8 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_8 fanout1154 (.A(_2060_),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(net1157),
    .X(net1155));
 sg13g2_buf_8 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_8 fanout1157 (.A(_3335_),
    .X(net1157));
 sg13g2_buf_8 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_1 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(_3336_),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(net1163),
    .X(net1161));
 sg13g2_buf_1 fanout1162 (.A(net1163),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(_3336_),
    .X(net1163));
 sg13g2_buf_8 fanout1164 (.A(_1176_),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(_1176_),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(_1162_),
    .X(net1166));
 sg13g2_buf_8 fanout1167 (.A(_1162_),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(net1170),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(net1172),
    .X(net1170));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(_2798_),
    .X(net1172));
 sg13g2_buf_8 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_8 fanout1174 (.A(_1149_),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(net1177),
    .X(net1175));
 sg13g2_buf_1 fanout1176 (.A(net1177),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(_2796_),
    .X(net1177));
 sg13g2_buf_8 fanout1178 (.A(net1181),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_8 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_8 fanout1181 (.A(_2796_),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_8 fanout1183 (.A(_1136_),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(_1124_),
    .X(net1184));
 sg13g2_buf_8 fanout1185 (.A(_1110_),
    .X(net1185));
 sg13g2_buf_8 fanout1186 (.A(_3384_),
    .X(net1186));
 sg13g2_buf_8 fanout1187 (.A(_3364_),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(_1782_),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(_1615_),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(_1090_),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_8 fanout1194 (.A(net1198),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(net1197),
    .X(net1195));
 sg13g2_buf_1 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_2 fanout1197 (.A(net1198),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(\tt6581_inst.mult_inst.nxt_state ),
    .X(net1198));
 sg13g2_buf_8 fanout1199 (.A(_4193_),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(_4189_),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(_4184_),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(_4173_),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(_4165_),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(_4165_),
    .X(net1204));
 sg13g2_buf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(_4156_),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(_4149_),
    .X(net1207));
 sg13g2_buf_8 fanout1208 (.A(net1209),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(_3404_),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(_3404_),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(_3403_),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(_3402_),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(_3066_),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(_1617_),
    .X(net1215));
 sg13g2_buf_8 fanout1216 (.A(_1394_),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(_1387_),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(_1069_),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(_1061_),
    .X(net1219));
 sg13g2_buf_8 fanout1220 (.A(_1053_),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(net1225),
    .X(net1222));
 sg13g2_buf_8 fanout1223 (.A(net1224),
    .X(net1223));
 sg13g2_buf_8 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(_1021_),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1228),
    .X(net1226));
 sg13g2_buf_1 fanout1227 (.A(net1228),
    .X(net1227));
 sg13g2_buf_1 fanout1228 (.A(_1021_),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(net1230),
    .X(net1229));
 sg13g2_buf_2 fanout1230 (.A(net1231),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(_1021_),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(_4219_),
    .X(net1232));
 sg13g2_buf_8 fanout1233 (.A(_4219_),
    .X(net1233));
 sg13g2_buf_8 fanout1234 (.A(_4191_),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(_4188_),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(_4186_),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(_4183_),
    .X(net1237));
 sg13g2_buf_8 fanout1238 (.A(_4181_),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(_4179_),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(_4177_),
    .X(net1240));
 sg13g2_buf_8 fanout1241 (.A(_4172_),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(_4170_),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(_4164_),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(_4155_),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(_4153_),
    .X(net1245));
 sg13g2_buf_8 fanout1246 (.A(_4148_),
    .X(net1246));
 sg13g2_buf_8 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_1 fanout1248 (.A(net1249),
    .X(net1248));
 sg13g2_buf_1 fanout1249 (.A(_3355_),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(_3355_),
    .X(net1250));
 sg13g2_buf_8 fanout1251 (.A(_3349_),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(_3342_),
    .X(net1252));
 sg13g2_buf_8 fanout1253 (.A(_3340_),
    .X(net1253));
 sg13g2_buf_8 fanout1254 (.A(_2799_),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(_2799_),
    .X(net1255));
 sg13g2_buf_8 fanout1256 (.A(_2673_),
    .X(net1256));
 sg13g2_buf_8 fanout1257 (.A(_2574_),
    .X(net1257));
 sg13g2_buf_8 fanout1258 (.A(_2571_),
    .X(net1258));
 sg13g2_buf_8 fanout1259 (.A(net1260),
    .X(net1259));
 sg13g2_buf_8 fanout1260 (.A(_2562_),
    .X(net1260));
 sg13g2_buf_8 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_8 fanout1262 (.A(_2559_),
    .X(net1262));
 sg13g2_buf_8 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(_2539_),
    .X(net1264));
 sg13g2_buf_8 fanout1265 (.A(_2522_),
    .X(net1265));
 sg13g2_buf_8 fanout1266 (.A(net1267),
    .X(net1266));
 sg13g2_buf_1 fanout1267 (.A(net1268),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_1 fanout1269 (.A(_1897_),
    .X(net1269));
 sg13g2_buf_8 fanout1270 (.A(net1272),
    .X(net1270));
 sg13g2_buf_1 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(_1897_),
    .X(net1272));
 sg13g2_buf_8 fanout1273 (.A(_1397_),
    .X(net1273));
 sg13g2_buf_8 fanout1274 (.A(_1393_),
    .X(net1274));
 sg13g2_buf_8 fanout1275 (.A(_1391_),
    .X(net1275));
 sg13g2_buf_8 fanout1276 (.A(_1386_),
    .X(net1276));
 sg13g2_buf_8 fanout1277 (.A(_1384_),
    .X(net1277));
 sg13g2_buf_8 fanout1278 (.A(_1382_),
    .X(net1278));
 sg13g2_buf_8 fanout1279 (.A(_1380_),
    .X(net1279));
 sg13g2_buf_8 fanout1280 (.A(_1377_),
    .X(net1280));
 sg13g2_buf_8 fanout1281 (.A(_1071_),
    .X(net1281));
 sg13g2_buf_8 fanout1282 (.A(_1068_),
    .X(net1282));
 sg13g2_buf_8 fanout1283 (.A(_1064_),
    .X(net1283));
 sg13g2_buf_8 fanout1284 (.A(_1060_),
    .X(net1284));
 sg13g2_buf_8 fanout1285 (.A(_1058_),
    .X(net1285));
 sg13g2_buf_8 fanout1286 (.A(_1052_),
    .X(net1286));
 sg13g2_buf_8 fanout1287 (.A(net1288),
    .X(net1287));
 sg13g2_buf_1 fanout1288 (.A(net1289),
    .X(net1288));
 sg13g2_buf_1 fanout1289 (.A(net1290),
    .X(net1289));
 sg13g2_buf_1 fanout1290 (.A(_1020_),
    .X(net1290));
 sg13g2_buf_8 fanout1291 (.A(_4386_),
    .X(net1291));
 sg13g2_buf_1 fanout1292 (.A(_4386_),
    .X(net1292));
 sg13g2_buf_8 fanout1293 (.A(_4381_),
    .X(net1293));
 sg13g2_buf_8 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_8 fanout1295 (.A(_4078_),
    .X(net1295));
 sg13g2_buf_8 fanout1296 (.A(net1299),
    .X(net1296));
 sg13g2_buf_8 fanout1297 (.A(net1299),
    .X(net1297));
 sg13g2_buf_1 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_8 fanout1299 (.A(net1307),
    .X(net1299));
 sg13g2_buf_8 fanout1300 (.A(net1302),
    .X(net1300));
 sg13g2_buf_1 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_1 fanout1302 (.A(net1307),
    .X(net1302));
 sg13g2_buf_8 fanout1303 (.A(net1306),
    .X(net1303));
 sg13g2_buf_8 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_8 fanout1305 (.A(net1306),
    .X(net1305));
 sg13g2_buf_2 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_buf_8 fanout1307 (.A(_3948_),
    .X(net1307));
 sg13g2_buf_8 fanout1308 (.A(net1312),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(net1312),
    .X(net1309));
 sg13g2_buf_8 fanout1310 (.A(net1312),
    .X(net1310));
 sg13g2_buf_1 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_2 fanout1312 (.A(_3931_),
    .X(net1312));
 sg13g2_buf_8 fanout1313 (.A(net1314),
    .X(net1313));
 sg13g2_buf_2 fanout1314 (.A(_3931_),
    .X(net1314));
 sg13g2_buf_8 fanout1315 (.A(net1318),
    .X(net1315));
 sg13g2_buf_8 fanout1316 (.A(net1318),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_8 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_buf_8 fanout1319 (.A(_3931_),
    .X(net1319));
 sg13g2_buf_8 fanout1320 (.A(net1323),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(net1323),
    .X(net1321));
 sg13g2_buf_8 fanout1322 (.A(net1323),
    .X(net1322));
 sg13g2_buf_8 fanout1323 (.A(net1330),
    .X(net1323));
 sg13g2_buf_8 fanout1324 (.A(net1325),
    .X(net1324));
 sg13g2_buf_1 fanout1325 (.A(net1330),
    .X(net1325));
 sg13g2_buf_8 fanout1326 (.A(net1329),
    .X(net1326));
 sg13g2_buf_8 fanout1327 (.A(net1329),
    .X(net1327));
 sg13g2_buf_1 fanout1328 (.A(net1329),
    .X(net1328));
 sg13g2_buf_8 fanout1329 (.A(net1330),
    .X(net1329));
 sg13g2_buf_8 fanout1330 (.A(_3902_),
    .X(net1330));
 sg13g2_buf_8 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_2 fanout1332 (.A(_3333_),
    .X(net1332));
 sg13g2_buf_8 fanout1333 (.A(_3333_),
    .X(net1333));
 sg13g2_buf_8 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_8 fanout1335 (.A(net1336),
    .X(net1335));
 sg13g2_buf_8 fanout1336 (.A(_3333_),
    .X(net1336));
 sg13g2_buf_8 fanout1337 (.A(net1338),
    .X(net1337));
 sg13g2_buf_2 fanout1338 (.A(_3330_),
    .X(net1338));
 sg13g2_buf_8 fanout1339 (.A(_3330_),
    .X(net1339));
 sg13g2_buf_8 fanout1340 (.A(net1342),
    .X(net1340));
 sg13g2_buf_1 fanout1341 (.A(net1342),
    .X(net1341));
 sg13g2_buf_8 fanout1342 (.A(_3330_),
    .X(net1342));
 sg13g2_buf_8 fanout1343 (.A(_3064_),
    .X(net1343));
 sg13g2_buf_8 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_2 fanout1345 (.A(net1349),
    .X(net1345));
 sg13g2_buf_8 fanout1346 (.A(net1349),
    .X(net1346));
 sg13g2_buf_8 fanout1347 (.A(net1348),
    .X(net1347));
 sg13g2_buf_8 fanout1348 (.A(net1349),
    .X(net1348));
 sg13g2_buf_8 fanout1349 (.A(_2512_),
    .X(net1349));
 sg13g2_buf_8 fanout1350 (.A(net1351),
    .X(net1350));
 sg13g2_buf_8 fanout1351 (.A(net1353),
    .X(net1351));
 sg13g2_buf_8 fanout1352 (.A(net1353),
    .X(net1352));
 sg13g2_buf_8 fanout1353 (.A(_2000_),
    .X(net1353));
 sg13g2_buf_8 fanout1354 (.A(net1355),
    .X(net1354));
 sg13g2_buf_8 fanout1355 (.A(net1357),
    .X(net1355));
 sg13g2_buf_8 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_8 fanout1357 (.A(_1998_),
    .X(net1357));
 sg13g2_buf_8 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_8 fanout1359 (.A(net1361),
    .X(net1359));
 sg13g2_buf_8 fanout1360 (.A(net1361),
    .X(net1360));
 sg13g2_buf_8 fanout1361 (.A(_1895_),
    .X(net1361));
 sg13g2_buf_8 fanout1362 (.A(_2661_),
    .X(net1362));
 sg13g2_buf_8 fanout1363 (.A(_2661_),
    .X(net1363));
 sg13g2_buf_8 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_8 fanout1365 (.A(net1366),
    .X(net1365));
 sg13g2_buf_8 fanout1366 (.A(net1369),
    .X(net1366));
 sg13g2_buf_8 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_8 fanout1368 (.A(net1369),
    .X(net1368));
 sg13g2_buf_8 fanout1369 (.A(_1533_),
    .X(net1369));
 sg13g2_buf_8 fanout1370 (.A(net1372),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(net1372),
    .X(net1371));
 sg13g2_buf_8 fanout1372 (.A(_1533_),
    .X(net1372));
 sg13g2_buf_8 fanout1373 (.A(_1532_),
    .X(net1373));
 sg13g2_buf_8 fanout1374 (.A(_1532_),
    .X(net1374));
 sg13g2_buf_8 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_8 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_8 fanout1377 (.A(net1384),
    .X(net1377));
 sg13g2_buf_8 fanout1378 (.A(net1384),
    .X(net1378));
 sg13g2_buf_8 fanout1379 (.A(net1384),
    .X(net1379));
 sg13g2_buf_8 fanout1380 (.A(net1382),
    .X(net1380));
 sg13g2_buf_1 fanout1381 (.A(net1382),
    .X(net1381));
 sg13g2_buf_8 fanout1382 (.A(net1383),
    .X(net1382));
 sg13g2_buf_8 fanout1383 (.A(net1384),
    .X(net1383));
 sg13g2_buf_8 fanout1384 (.A(_1044_),
    .X(net1384));
 sg13g2_buf_8 fanout1385 (.A(net1387),
    .X(net1385));
 sg13g2_buf_1 fanout1386 (.A(net1387),
    .X(net1386));
 sg13g2_buf_8 fanout1387 (.A(net1389),
    .X(net1387));
 sg13g2_buf_8 fanout1388 (.A(net1389),
    .X(net1388));
 sg13g2_buf_8 fanout1389 (.A(net1392),
    .X(net1389));
 sg13g2_buf_8 fanout1390 (.A(net1391),
    .X(net1390));
 sg13g2_buf_8 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_8 fanout1392 (.A(_1043_),
    .X(net1392));
 sg13g2_buf_8 fanout1393 (.A(net1396),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(net1396),
    .X(net1394));
 sg13g2_buf_8 fanout1395 (.A(net1396),
    .X(net1395));
 sg13g2_buf_8 fanout1396 (.A(_1042_),
    .X(net1396));
 sg13g2_buf_8 fanout1397 (.A(net1398),
    .X(net1397));
 sg13g2_buf_8 fanout1398 (.A(net1399),
    .X(net1398));
 sg13g2_buf_8 fanout1399 (.A(_1042_),
    .X(net1399));
 sg13g2_buf_8 fanout1400 (.A(net1401),
    .X(net1400));
 sg13g2_buf_8 fanout1401 (.A(net1405),
    .X(net1401));
 sg13g2_buf_8 fanout1402 (.A(net1403),
    .X(net1402));
 sg13g2_buf_8 fanout1403 (.A(net1405),
    .X(net1403));
 sg13g2_buf_8 fanout1404 (.A(net1405),
    .X(net1404));
 sg13g2_buf_8 fanout1405 (.A(_1042_),
    .X(net1405));
 sg13g2_buf_8 fanout1406 (.A(net1409),
    .X(net1406));
 sg13g2_buf_8 fanout1407 (.A(net1409),
    .X(net1407));
 sg13g2_buf_8 fanout1408 (.A(net1409),
    .X(net1408));
 sg13g2_buf_8 fanout1409 (.A(net1412),
    .X(net1409));
 sg13g2_buf_8 fanout1410 (.A(net1411),
    .X(net1410));
 sg13g2_buf_8 fanout1411 (.A(net1412),
    .X(net1411));
 sg13g2_buf_8 fanout1412 (.A(net1414),
    .X(net1412));
 sg13g2_buf_8 fanout1413 (.A(net1414),
    .X(net1413));
 sg13g2_buf_8 fanout1414 (.A(_1016_),
    .X(net1414));
 sg13g2_buf_8 fanout1415 (.A(net1416),
    .X(net1415));
 sg13g2_buf_8 fanout1416 (.A(_1016_),
    .X(net1416));
 sg13g2_buf_8 fanout1417 (.A(net1426),
    .X(net1417));
 sg13g2_buf_8 fanout1418 (.A(net1426),
    .X(net1418));
 sg13g2_buf_8 fanout1419 (.A(net1420),
    .X(net1419));
 sg13g2_buf_8 fanout1420 (.A(net1426),
    .X(net1420));
 sg13g2_buf_8 fanout1421 (.A(net1425),
    .X(net1421));
 sg13g2_buf_2 fanout1422 (.A(net1425),
    .X(net1422));
 sg13g2_buf_8 fanout1423 (.A(net1424),
    .X(net1423));
 sg13g2_buf_8 fanout1424 (.A(net1425),
    .X(net1424));
 sg13g2_buf_8 fanout1425 (.A(net1426),
    .X(net1425));
 sg13g2_buf_8 fanout1426 (.A(_1015_),
    .X(net1426));
 sg13g2_buf_8 fanout1427 (.A(net1428),
    .X(net1427));
 sg13g2_buf_8 fanout1428 (.A(_1004_),
    .X(net1428));
 sg13g2_buf_8 fanout1429 (.A(net1430),
    .X(net1429));
 sg13g2_buf_8 fanout1430 (.A(_1004_),
    .X(net1430));
 sg13g2_buf_8 fanout1431 (.A(_1001_),
    .X(net1431));
 sg13g2_buf_8 fanout1432 (.A(net1433),
    .X(net1432));
 sg13g2_buf_8 fanout1433 (.A(_0998_),
    .X(net1433));
 sg13g2_buf_8 fanout1434 (.A(net1437),
    .X(net1434));
 sg13g2_buf_8 fanout1435 (.A(net1437),
    .X(net1435));
 sg13g2_buf_2 fanout1436 (.A(net1437),
    .X(net1436));
 sg13g2_buf_8 fanout1437 (.A(_0917_),
    .X(net1437));
 sg13g2_buf_8 fanout1438 (.A(net1439),
    .X(net1438));
 sg13g2_buf_8 fanout1439 (.A(net1440),
    .X(net1439));
 sg13g2_buf_8 fanout1440 (.A(net1441),
    .X(net1440));
 sg13g2_buf_8 fanout1441 (.A(_0888_),
    .X(net1441));
 sg13g2_buf_8 fanout1442 (.A(net1443),
    .X(net1442));
 sg13g2_buf_8 fanout1443 (.A(_0888_),
    .X(net1443));
 sg13g2_buf_8 fanout1444 (.A(_0888_),
    .X(net1444));
 sg13g2_buf_8 fanout1445 (.A(net1704),
    .X(net1445));
 sg13g2_buf_8 fanout1446 (.A(net1700),
    .X(net1446));
 sg13g2_buf_8 fanout1447 (.A(net1448),
    .X(net1447));
 sg13g2_buf_8 fanout1448 (.A(\tt6581_inst.reg_file_inst.we_i ),
    .X(net1448));
 sg13g2_buf_8 fanout1449 (.A(net1450),
    .X(net1449));
 sg13g2_buf_8 fanout1450 (.A(net900),
    .X(net1450));
 sg13g2_buf_8 fanout1451 (.A(net1452),
    .X(net1451));
 sg13g2_buf_8 fanout1452 (.A(net821),
    .X(net1452));
 sg13g2_buf_8 fanout1453 (.A(net1454),
    .X(net1453));
 sg13g2_buf_8 fanout1454 (.A(net961),
    .X(net1454));
 sg13g2_buf_8 fanout1455 (.A(net961),
    .X(net1455));
 sg13g2_buf_1 fanout1456 (.A(net961),
    .X(net1456));
 sg13g2_buf_8 fanout1457 (.A(net1458),
    .X(net1457));
 sg13g2_buf_8 fanout1458 (.A(net1461),
    .X(net1458));
 sg13g2_buf_8 fanout1459 (.A(net1460),
    .X(net1459));
 sg13g2_buf_8 fanout1460 (.A(net1461),
    .X(net1460));
 sg13g2_buf_8 fanout1461 (.A(net939),
    .X(net1461));
 sg13g2_buf_8 fanout1462 (.A(net1463),
    .X(net1462));
 sg13g2_buf_8 fanout1463 (.A(\tt6581_inst.reg_file_inst.wdata_i[5] ),
    .X(net1463));
 sg13g2_buf_8 fanout1464 (.A(net1465),
    .X(net1464));
 sg13g2_buf_8 fanout1465 (.A(\tt6581_inst.reg_file_inst.wdata_i[5] ),
    .X(net1465));
 sg13g2_buf_8 fanout1466 (.A(net1467),
    .X(net1466));
 sg13g2_buf_8 fanout1467 (.A(net1036),
    .X(net1467));
 sg13g2_buf_8 fanout1468 (.A(net1470),
    .X(net1468));
 sg13g2_buf_1 fanout1469 (.A(net1470),
    .X(net1469));
 sg13g2_buf_8 fanout1470 (.A(net1036),
    .X(net1470));
 sg13g2_buf_8 fanout1471 (.A(net1475),
    .X(net1471));
 sg13g2_buf_1 fanout1472 (.A(net1475),
    .X(net1472));
 sg13g2_buf_8 fanout1473 (.A(net1474),
    .X(net1473));
 sg13g2_buf_8 fanout1474 (.A(net1475),
    .X(net1474));
 sg13g2_buf_8 fanout1475 (.A(\tt6581_inst.reg_file_inst.wdata_i[3] ),
    .X(net1475));
 sg13g2_buf_8 fanout1476 (.A(net1477),
    .X(net1476));
 sg13g2_buf_8 fanout1477 (.A(net1480),
    .X(net1477));
 sg13g2_buf_8 fanout1478 (.A(net1479),
    .X(net1478));
 sg13g2_buf_8 fanout1479 (.A(net1480),
    .X(net1479));
 sg13g2_buf_8 fanout1480 (.A(\tt6581_inst.reg_file_inst.wdata_i[2] ),
    .X(net1480));
 sg13g2_buf_8 fanout1481 (.A(net1482),
    .X(net1481));
 sg13g2_buf_8 fanout1482 (.A(net792),
    .X(net1482));
 sg13g2_buf_8 fanout1483 (.A(net792),
    .X(net1483));
 sg13g2_buf_8 fanout1484 (.A(net792),
    .X(net1484));
 sg13g2_buf_8 fanout1485 (.A(\tt6581_inst.reg_file_inst.wdata_i[0] ),
    .X(net1485));
 sg13g2_buf_8 fanout1486 (.A(\tt6581_inst.reg_file_inst.wdata_i[0] ),
    .X(net1486));
 sg13g2_buf_8 fanout1487 (.A(net1488),
    .X(net1487));
 sg13g2_buf_8 fanout1488 (.A(\tt6581_inst.reg_file_inst.wdata_i[0] ),
    .X(net1488));
 sg13g2_buf_8 fanout1489 (.A(net1490),
    .X(net1489));
 sg13g2_buf_8 fanout1490 (.A(net1491),
    .X(net1490));
 sg13g2_buf_8 fanout1491 (.A(\tt6581_inst.controller_inst.mult_in_mux_o[2] ),
    .X(net1491));
 sg13g2_buf_8 fanout1492 (.A(net1493),
    .X(net1492));
 sg13g2_buf_8 fanout1493 (.A(\tt6581_inst.controller_inst.mult_in_mux_o[1] ),
    .X(net1493));
 sg13g2_buf_8 fanout1494 (.A(_0113_),
    .X(net1494));
 sg13g2_buf_8 fanout1495 (.A(net1497),
    .X(net1495));
 sg13g2_buf_8 fanout1496 (.A(net1497),
    .X(net1496));
 sg13g2_buf_8 fanout1497 (.A(\tt6581_inst.filter_accum[13] ),
    .X(net1497));
 sg13g2_buf_8 fanout1498 (.A(net1499),
    .X(net1498));
 sg13g2_buf_8 fanout1499 (.A(net62),
    .X(net1499));
 sg13g2_buf_8 fanout1500 (.A(net1504),
    .X(net1500));
 sg13g2_buf_8 fanout1501 (.A(net1502),
    .X(net1501));
 sg13g2_buf_8 fanout1502 (.A(net1503),
    .X(net1502));
 sg13g2_buf_8 fanout1503 (.A(net1504),
    .X(net1503));
 sg13g2_buf_8 fanout1504 (.A(\tt6581_inst.mult_inst.neg_result ),
    .X(net1504));
 sg13g2_buf_8 fanout1505 (.A(net1692),
    .X(net1505));
 sg13g2_buf_8 fanout1506 (.A(net1691),
    .X(net1506));
 sg13g2_buf_8 fanout1507 (.A(net1134),
    .X(net1507));
 sg13g2_buf_8 fanout1508 (.A(net1696),
    .X(net1508));
 sg13g2_buf_8 fanout1509 (.A(net1511),
    .X(net1509));
 sg13g2_buf_2 fanout1510 (.A(net1511),
    .X(net1510));
 sg13g2_buf_8 fanout1511 (.A(net1512),
    .X(net1511));
 sg13g2_buf_8 fanout1512 (.A(net1702),
    .X(net1512));
 sg13g2_buf_8 fanout1513 (.A(net1515),
    .X(net1513));
 sg13g2_buf_1 fanout1514 (.A(net1515),
    .X(net1514));
 sg13g2_buf_8 fanout1515 (.A(net1703),
    .X(net1515));
 sg13g2_buf_8 fanout1516 (.A(net1517),
    .X(net1516));
 sg13g2_buf_8 fanout1517 (.A(net1518),
    .X(net1517));
 sg13g2_buf_8 fanout1518 (.A(net1523),
    .X(net1518));
 sg13g2_buf_8 fanout1519 (.A(net1520),
    .X(net1519));
 sg13g2_buf_2 fanout1520 (.A(net1521),
    .X(net1520));
 sg13g2_buf_8 fanout1521 (.A(net1522),
    .X(net1521));
 sg13g2_buf_8 fanout1522 (.A(net1523),
    .X(net1522));
 sg13g2_buf_8 fanout1523 (.A(net1701),
    .X(net1523));
 sg13g2_buf_8 fanout1524 (.A(net1525),
    .X(net1524));
 sg13g2_buf_8 fanout1525 (.A(net1526),
    .X(net1525));
 sg13g2_buf_8 fanout1526 (.A(net220),
    .X(net1526));
 sg13g2_buf_8 fanout1527 (.A(net1528),
    .X(net1527));
 sg13g2_buf_8 fanout1528 (.A(net1529),
    .X(net1528));
 sg13g2_buf_8 fanout1529 (.A(\tt6581_inst.svf_inst.cur_state[5] ),
    .X(net1529));
 sg13g2_buf_8 fanout1530 (.A(net1531),
    .X(net1530));
 sg13g2_buf_8 fanout1531 (.A(net1699),
    .X(net1531));
 sg13g2_buf_8 fanout1532 (.A(net1533),
    .X(net1532));
 sg13g2_buf_8 fanout1533 (.A(\tt6581_inst.svf_inst.cur_state[2] ),
    .X(net1533));
 sg13g2_buf_8 fanout1534 (.A(net1535),
    .X(net1534));
 sg13g2_buf_8 fanout1535 (.A(net205),
    .X(net1535));
 sg13g2_buf_8 fanout1536 (.A(net1695),
    .X(net1536));
 sg13g2_buf_8 fanout1537 (.A(net1538),
    .X(net1537));
 sg13g2_buf_8 fanout1538 (.A(net1543),
    .X(net1538));
 sg13g2_buf_8 fanout1539 (.A(net1543),
    .X(net1539));
 sg13g2_buf_1 fanout1540 (.A(net1543),
    .X(net1540));
 sg13g2_buf_8 fanout1541 (.A(net1543),
    .X(net1541));
 sg13g2_buf_8 fanout1542 (.A(net1543),
    .X(net1542));
 sg13g2_buf_8 fanout1543 (.A(\tt6581_inst.mult_inst.cur_state ),
    .X(net1543));
 sg13g2_buf_8 fanout1544 (.A(net453),
    .X(net1544));
 sg13g2_buf_8 fanout1545 (.A(net569),
    .X(net1545));
 sg13g2_buf_8 fanout1546 (.A(net1547),
    .X(net1546));
 sg13g2_buf_8 fanout1547 (.A(net1548),
    .X(net1547));
 sg13g2_buf_8 fanout1548 (.A(net1552),
    .X(net1548));
 sg13g2_buf_8 fanout1549 (.A(net1552),
    .X(net1549));
 sg13g2_buf_8 fanout1550 (.A(net1552),
    .X(net1550));
 sg13g2_buf_8 fanout1551 (.A(net1552),
    .X(net1551));
 sg13g2_buf_8 fanout1552 (.A(net195),
    .X(net1552));
 sg13g2_buf_8 fanout1553 (.A(net1557),
    .X(net1553));
 sg13g2_buf_8 fanout1554 (.A(net1557),
    .X(net1554));
 sg13g2_buf_8 fanout1555 (.A(net1557),
    .X(net1555));
 sg13g2_buf_1 fanout1556 (.A(net1557),
    .X(net1556));
 sg13g2_buf_8 fanout1557 (.A(net1571),
    .X(net1557));
 sg13g2_buf_8 fanout1558 (.A(net1571),
    .X(net1558));
 sg13g2_buf_8 fanout1559 (.A(net1571),
    .X(net1559));
 sg13g2_buf_8 fanout1560 (.A(net1561),
    .X(net1560));
 sg13g2_buf_8 fanout1561 (.A(net1570),
    .X(net1561));
 sg13g2_buf_2 fanout1562 (.A(net1570),
    .X(net1562));
 sg13g2_buf_8 fanout1563 (.A(net1565),
    .X(net1563));
 sg13g2_buf_8 fanout1564 (.A(net1565),
    .X(net1564));
 sg13g2_buf_8 fanout1565 (.A(net1570),
    .X(net1565));
 sg13g2_buf_8 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_8 fanout1567 (.A(net1570),
    .X(net1567));
 sg13g2_buf_8 fanout1568 (.A(net1570),
    .X(net1568));
 sg13g2_buf_2 fanout1569 (.A(net1570),
    .X(net1569));
 sg13g2_buf_8 fanout1570 (.A(net1571),
    .X(net1570));
 sg13g2_buf_8 fanout1571 (.A(net1690),
    .X(net1571));
 sg13g2_buf_8 fanout1572 (.A(net1573),
    .X(net1572));
 sg13g2_buf_8 fanout1573 (.A(net1584),
    .X(net1573));
 sg13g2_buf_8 fanout1574 (.A(net1576),
    .X(net1574));
 sg13g2_buf_8 fanout1575 (.A(net1576),
    .X(net1575));
 sg13g2_buf_8 fanout1576 (.A(net1584),
    .X(net1576));
 sg13g2_buf_8 fanout1577 (.A(net1580),
    .X(net1577));
 sg13g2_buf_2 fanout1578 (.A(net1580),
    .X(net1578));
 sg13g2_buf_8 fanout1579 (.A(net1580),
    .X(net1579));
 sg13g2_buf_8 fanout1580 (.A(net1584),
    .X(net1580));
 sg13g2_buf_8 fanout1581 (.A(net1583),
    .X(net1581));
 sg13g2_buf_1 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_8 fanout1583 (.A(net1584),
    .X(net1583));
 sg13g2_buf_8 fanout1584 (.A(net1690),
    .X(net1584));
 sg13g2_buf_8 fanout1585 (.A(net1587),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(net1587),
    .X(net1586));
 sg13g2_buf_8 fanout1587 (.A(net1590),
    .X(net1587));
 sg13g2_buf_8 fanout1588 (.A(net1589),
    .X(net1588));
 sg13g2_buf_8 fanout1589 (.A(net1590),
    .X(net1589));
 sg13g2_buf_8 fanout1590 (.A(net1623),
    .X(net1590));
 sg13g2_buf_8 fanout1591 (.A(net1592),
    .X(net1591));
 sg13g2_buf_8 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_8 fanout1593 (.A(net1623),
    .X(net1593));
 sg13g2_buf_8 fanout1594 (.A(net1596),
    .X(net1594));
 sg13g2_buf_8 fanout1595 (.A(net1596),
    .X(net1595));
 sg13g2_buf_8 fanout1596 (.A(net1597),
    .X(net1596));
 sg13g2_buf_8 fanout1597 (.A(net1601),
    .X(net1597));
 sg13g2_buf_8 fanout1598 (.A(net1599),
    .X(net1598));
 sg13g2_buf_8 fanout1599 (.A(net1601),
    .X(net1599));
 sg13g2_buf_8 fanout1600 (.A(net1601),
    .X(net1600));
 sg13g2_buf_8 fanout1601 (.A(net1623),
    .X(net1601));
 sg13g2_buf_8 fanout1602 (.A(net1605),
    .X(net1602));
 sg13g2_buf_8 fanout1603 (.A(net1604),
    .X(net1603));
 sg13g2_buf_8 fanout1604 (.A(net1605),
    .X(net1604));
 sg13g2_buf_8 fanout1605 (.A(net1622),
    .X(net1605));
 sg13g2_buf_8 fanout1606 (.A(net1608),
    .X(net1606));
 sg13g2_buf_1 fanout1607 (.A(net1608),
    .X(net1607));
 sg13g2_buf_8 fanout1608 (.A(net1622),
    .X(net1608));
 sg13g2_buf_8 fanout1609 (.A(net1610),
    .X(net1609));
 sg13g2_buf_8 fanout1610 (.A(net1622),
    .X(net1610));
 sg13g2_buf_8 fanout1611 (.A(net1621),
    .X(net1611));
 sg13g2_buf_8 fanout1612 (.A(net1621),
    .X(net1612));
 sg13g2_buf_8 fanout1613 (.A(net1615),
    .X(net1613));
 sg13g2_buf_8 fanout1614 (.A(net1615),
    .X(net1614));
 sg13g2_buf_8 fanout1615 (.A(net1621),
    .X(net1615));
 sg13g2_buf_8 fanout1616 (.A(net1617),
    .X(net1616));
 sg13g2_buf_8 fanout1617 (.A(net1621),
    .X(net1617));
 sg13g2_buf_8 fanout1618 (.A(net1620),
    .X(net1618));
 sg13g2_buf_8 fanout1619 (.A(net1620),
    .X(net1619));
 sg13g2_buf_8 fanout1620 (.A(net1621),
    .X(net1620));
 sg13g2_buf_8 fanout1621 (.A(net1622),
    .X(net1621));
 sg13g2_buf_8 fanout1622 (.A(net1623),
    .X(net1622));
 sg13g2_buf_8 fanout1623 (.A(net1690),
    .X(net1623));
 sg13g2_buf_8 fanout1624 (.A(net1625),
    .X(net1624));
 sg13g2_buf_8 fanout1625 (.A(net1628),
    .X(net1625));
 sg13g2_buf_8 fanout1626 (.A(net1628),
    .X(net1626));
 sg13g2_buf_8 fanout1627 (.A(net1628),
    .X(net1627));
 sg13g2_buf_8 fanout1628 (.A(net1639),
    .X(net1628));
 sg13g2_buf_8 fanout1629 (.A(net1633),
    .X(net1629));
 sg13g2_buf_8 fanout1630 (.A(net1633),
    .X(net1630));
 sg13g2_buf_8 fanout1631 (.A(net1633),
    .X(net1631));
 sg13g2_buf_2 fanout1632 (.A(net1633),
    .X(net1632));
 sg13g2_buf_8 fanout1633 (.A(net1639),
    .X(net1633));
 sg13g2_buf_8 fanout1634 (.A(net1635),
    .X(net1634));
 sg13g2_buf_8 fanout1635 (.A(net1639),
    .X(net1635));
 sg13g2_buf_8 fanout1636 (.A(net1638),
    .X(net1636));
 sg13g2_buf_8 fanout1637 (.A(net1638),
    .X(net1637));
 sg13g2_buf_8 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_8 fanout1639 (.A(net1658),
    .X(net1639));
 sg13g2_buf_8 fanout1640 (.A(net1642),
    .X(net1640));
 sg13g2_buf_8 fanout1641 (.A(net1642),
    .X(net1641));
 sg13g2_buf_8 fanout1642 (.A(net1647),
    .X(net1642));
 sg13g2_buf_8 fanout1643 (.A(net1646),
    .X(net1643));
 sg13g2_buf_8 fanout1644 (.A(net1646),
    .X(net1644));
 sg13g2_buf_8 fanout1645 (.A(net1646),
    .X(net1645));
 sg13g2_buf_8 fanout1646 (.A(net1647),
    .X(net1646));
 sg13g2_buf_8 fanout1647 (.A(net1658),
    .X(net1647));
 sg13g2_buf_8 fanout1648 (.A(net1652),
    .X(net1648));
 sg13g2_buf_8 fanout1649 (.A(net1652),
    .X(net1649));
 sg13g2_buf_8 fanout1650 (.A(net1651),
    .X(net1650));
 sg13g2_buf_8 fanout1651 (.A(net1652),
    .X(net1651));
 sg13g2_buf_8 fanout1652 (.A(net1658),
    .X(net1652));
 sg13g2_buf_8 fanout1653 (.A(net1657),
    .X(net1653));
 sg13g2_buf_8 fanout1654 (.A(net1657),
    .X(net1654));
 sg13g2_buf_8 fanout1655 (.A(net1657),
    .X(net1655));
 sg13g2_buf_1 fanout1656 (.A(net1657),
    .X(net1656));
 sg13g2_buf_8 fanout1657 (.A(net1658),
    .X(net1657));
 sg13g2_buf_8 fanout1658 (.A(net1689),
    .X(net1658));
 sg13g2_buf_8 fanout1659 (.A(net1661),
    .X(net1659));
 sg13g2_buf_2 fanout1660 (.A(net1661),
    .X(net1660));
 sg13g2_buf_8 fanout1661 (.A(net1664),
    .X(net1661));
 sg13g2_buf_8 fanout1662 (.A(net1663),
    .X(net1662));
 sg13g2_buf_8 fanout1663 (.A(net1664),
    .X(net1663));
 sg13g2_buf_8 fanout1664 (.A(net1674),
    .X(net1664));
 sg13g2_buf_8 fanout1665 (.A(net1668),
    .X(net1665));
 sg13g2_buf_8 fanout1666 (.A(net1668),
    .X(net1666));
 sg13g2_buf_8 fanout1667 (.A(net1674),
    .X(net1667));
 sg13g2_buf_8 fanout1668 (.A(net1674),
    .X(net1668));
 sg13g2_buf_8 fanout1669 (.A(net1671),
    .X(net1669));
 sg13g2_buf_8 fanout1670 (.A(net1671),
    .X(net1670));
 sg13g2_buf_8 fanout1671 (.A(net1674),
    .X(net1671));
 sg13g2_buf_8 fanout1672 (.A(net1673),
    .X(net1672));
 sg13g2_buf_8 fanout1673 (.A(net1674),
    .X(net1673));
 sg13g2_buf_8 fanout1674 (.A(net1689),
    .X(net1674));
 sg13g2_buf_8 fanout1675 (.A(net1681),
    .X(net1675));
 sg13g2_buf_2 fanout1676 (.A(net1681),
    .X(net1676));
 sg13g2_buf_8 fanout1677 (.A(net1679),
    .X(net1677));
 sg13g2_buf_8 fanout1678 (.A(net1679),
    .X(net1678));
 sg13g2_buf_8 fanout1679 (.A(net1680),
    .X(net1679));
 sg13g2_buf_8 fanout1680 (.A(net1681),
    .X(net1680));
 sg13g2_buf_8 fanout1681 (.A(net1689),
    .X(net1681));
 sg13g2_buf_8 fanout1682 (.A(net1684),
    .X(net1682));
 sg13g2_buf_2 fanout1683 (.A(net1684),
    .X(net1683));
 sg13g2_buf_8 fanout1684 (.A(net1688),
    .X(net1684));
 sg13g2_buf_8 fanout1685 (.A(net1688),
    .X(net1685));
 sg13g2_buf_8 fanout1686 (.A(net1688),
    .X(net1686));
 sg13g2_buf_8 fanout1687 (.A(net1688),
    .X(net1687));
 sg13g2_buf_8 fanout1688 (.A(net1689),
    .X(net1688));
 sg13g2_buf_8 fanout1689 (.A(net1690),
    .X(net1689));
 sg13g2_buf_8 fanout1690 (.A(rst_n),
    .X(net1690));
 sg13g2_buf_1 input1 (.A(uio_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[3]),
    .X(net3));
 sg13g2_tielo tt_um_andreasp00_4 (.L_LO(net4));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_leaf_107_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_109_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_101_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_103_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_104_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_105_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_106_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_100_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_43_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_90_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_91_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_92_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_93_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_leaf_94_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_leaf_95_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_97_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_leaf_99_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_83_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_84_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_88_clk));
 sg13g2_inv_8 clkload31 (.A(clknet_leaf_89_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_78_clk));
 sg13g2_buf_8 clkload33 (.A(clknet_leaf_79_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_80_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_81_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_82_clk));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_70_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_54_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_56_clk));
 sg13g2_inv_4 clkload41 (.A(clknet_leaf_62_clk));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_66_clk));
 sg13g2_inv_1 clkload43 (.A(clknet_leaf_57_clk));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_60_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\tt6581_inst.spi_inst.cs_sync[0] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold2 (.A(\tt6581_inst.spi_inst.sclk_sync[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold3 (.A(\tt6581_inst.spi_inst.mosi_sync[0] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold4 (.A(\tt6581_inst.controller_inst.cur_state[6] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold5 (.A(\tt6581_inst.controller_inst.cur_state[9] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold6 (.A(\tt6581_inst.controller_inst.cur_state[4] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold7 (.A(\tt6581_inst.controller_inst.cur_state[5] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold8 (.A(\tt6581_inst.controller_inst.cur_state[1] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold9 (.A(\tt6581_inst.controller_inst.cur_state[8] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold10 (.A(\tt6581_inst.spi_inst.sclk_sync[1] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0036_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0114_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0039_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0006_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold15 (.A(\tt6581_inst.controller_inst.voice_start_o ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold16 (.A(\tt6581_inst.multi_voice_inst.nxt_state[0] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold17 (.A(\tt6581_inst.controller_inst.filt_ready_i ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0115_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold19 (.A(\tt6581_inst.delta_sigma_inst.cnt[0] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0020_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold21 (.A(\tt6581_inst.tick_gen_inst.cnt[0] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold22 (.A(\tt6581_inst.multi_voice_inst.cur_state[1] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold23 (.A(\tt6581_inst.multi_voice_inst.nxt_state[1] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold24 (.A(\tt6581_inst.svf_inst.cur_state[3] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0008_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold26 (.A(\tt6581_inst.svf_inst.cur_state[8] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0005_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold28 (.A(\tt6581_inst.svf_inst.cur_state[1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0007_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold30 (.A(\tt6581_inst.controller_inst.cur_state[2] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0010_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold32 (.A(\tt6581_inst.controller_inst.cur_state[3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0011_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold34 (.A(\tt6581_inst.controller_inst.voice_ready_i ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold35 (.A(\tt6581_inst.controller_inst.cur_state[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0001_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold37 (.A(\tt6581_inst.audio_valid ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0816_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold39 (.A(\tt6581_inst.controller_inst.cur_state[10] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold40 (.A(\tt6581_inst.mult_inst.iter[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0298_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold42 (.A(\tt6581_inst.tick_gen_inst.cnt[4] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0029_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold44 (.A(\tt6581_inst.spi_inst.data_out_reg[7] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold45 (.A(_4348_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0790_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold47 (.A(\tt6581_inst.controller_inst.mult_start_o ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold48 (.A(\tt6581_inst.mult_inst.b_reg[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0348_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold50 (.A(\tt6581_inst.mult_inst.b_reg[6] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0346_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold52 (.A(\tt6581_inst.envelope_inst.cur_state[0] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0003_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold54 (.A(\tt6581_inst.mult_inst.b_reg[13] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0353_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold56 (.A(\tt6581_inst.tick_gen_inst.cnt[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold57 (.A(\tt6581_inst.mult_inst.b_reg[11] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0351_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold59 (.A(\tt6581_inst.mult_inst.b_reg[5] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0345_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold61 (.A(\tt6581_inst.mult_inst.b_reg[2] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0342_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold63 (.A(\tt6581_inst.spi_inst.data_out_reg[5] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold64 (.A(_4306_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0788_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold66 (.A(\tt6581_inst.svf_inst.reg_band[23] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0443_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold68 (.A(\tt6581_inst.spi_inst.data_out_reg[3] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold69 (.A(_4263_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0786_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold71 (.A(\tt6581_inst.mult_inst.b_reg[7] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold72 (.A(\tt6581_inst.spi_inst.data_out_reg[4] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold73 (.A(_4284_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0787_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold75 (.A(\tt6581_inst.mult_inst.b_reg[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0344_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold77 (.A(\tt6581_inst.mult_inst.b_reg[1] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0341_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold79 (.A(\tt6581_inst.spi_inst.data_out_reg[6] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold80 (.A(_4327_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0789_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold82 (.A(\tt6581_inst.spi_inst.data_out_reg[2] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold83 (.A(_4242_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0785_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold85 (.A(\tt6581_inst.mult_inst.b_reg[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0349_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold87 (.A(\tt6581_inst.delta_sigma_inst.cnt[2] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0023_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold89 (.A(\tt6581_inst.envelope_inst.cur_state[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold90 (.A(\tt6581_inst.mult_inst.b_reg[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0343_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold92 (.A(\tt6581_inst.spi_inst.data_out_reg[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold93 (.A(_4221_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0784_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold95 (.A(\tt6581_inst.controller_inst.env_start_o ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold96 (.A(\tt6581_inst.envelope_inst.vol_regs[1][14] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold97 (.A(\tt6581_inst.envelope_inst.vol_regs[2][10] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold98 (.A(\tt6581_inst.svf_inst.reg_band[0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold99 (.A(\tt6581_inst.accum_rst ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0648_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold101 (.A(\tt6581_inst.envelope_inst.vol_regs[2][23] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold102 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][12] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold103 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][15] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold104 (.A(\tt6581_inst.bypass_accum[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0817_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold106 (.A(\tt6581_inst.envelope_inst.vol_regs[1][10] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0037_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0338_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold109 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][5] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold110 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][13] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold111 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[1][1] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0647_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold113 (.A(\tt6581_inst.spi_inst.bit_cnt[0] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0792_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold115 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][14] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold116 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[2][1] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0671_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0042_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0470_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold120 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][11] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold121 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][11] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold122 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[0][1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0645_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold124 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold125 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][17] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold126 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][6] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold127 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold128 (.A(\tt6581_inst.envelope_inst.vol_regs[1][0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold129 (.A(\tt6581_inst.envelope_inst.vol_regs[0][9] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold130 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][8] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold131 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][8] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold132 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][4] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold133 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][12] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold134 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][3] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold135 (.A(\tt6581_inst.envelope_inst.vol_regs[2][14] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold136 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][10] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold137 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][14] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold138 (.A(\tt6581_inst.envelope_inst.vol_regs[0][0] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold139 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][17] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold140 (.A(\tt6581_inst.envelope_inst.vol_regs[1][22] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][10] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold142 (.A(\tt6581_inst.control_pack[14] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold143 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][8] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold144 (.A(\tt6581_inst.mult_inst.iter[0] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold145 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][4] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold146 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][11] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0090_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold148 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][15] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold149 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][15] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold150 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0043_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold152 (.A(\tt6581_inst.spi_inst.data_out_reg[0] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold153 (.A(_4198_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0783_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold155 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][17] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0092_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0623_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold158 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][6] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold159 (.A(\tt6581_inst.envelope_inst.vol_regs[1][9] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold160 (.A(\tt6581_inst.envelope_inst.vol_regs[0][23] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold161 (.A(\tt6581_inst.envelope_inst.vol_regs[2][0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold162 (.A(\tt6581_inst.delta_sigma_inst.e1[18] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0293_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold164 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold165 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][7] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold166 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][7] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold167 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold168 (.A(\tt6581_inst.envelope_inst.vol_regs[1][12] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold169 (.A(\tt6581_inst.envelope_inst.vol_regs[0][22] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold170 (.A(\tt6581_inst.delta_sigma_inst.en ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold171 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][9] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold172 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][7] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0108_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold174 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][2] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0069_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0600_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold177 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][5] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0061_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold179 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][5] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold180 (.A(\tt6581_inst.svf_inst.cur_state[2] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold181 (.A(\tt6581_inst.mult_inst.a_reg[5] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0304_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0041_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold184 (.A(\tt6581_inst.mult_inst.a_reg[18] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0317_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold186 (.A(\tt6581_inst.mult_inst.accum[38] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0394_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold188 (.A(\tt6581_inst.svf_inst.cur_state[10] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold189 (.A(\tt6581_inst.envelope_inst.vol_regs[0][10] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold190 (.A(\tt6581_inst.envelope_inst.vol_regs[1][23] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold191 (.A(\tt6581_inst.delta_sigma_inst.e2[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0256_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0038_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold194 (.A(\tt6581_inst.envelope_inst.vol_regs[2][22] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold195 (.A(\tt6581_inst.svf_inst.cur_state[6] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold196 (.A(\tt6581_inst.envelope_inst.vol_regs[0][14] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold197 (.A(\tt6581_inst.envelope_inst.vol_regs[1][16] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold198 (.A(\tt6581_inst.envelope_inst.vol_regs[2][4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold199 (.A(\tt6581_inst.mult_inst.a_reg[4] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0303_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold201 (.A(\tt6581_inst.mult_inst.b_reg[10] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold202 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][12] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold203 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][9] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold204 (.A(\tt6581_inst.mult_inst.b_reg[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold205 (.A(\tt6581_inst.control_pack[15] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0228_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold207 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][13] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold208 (.A(\tt6581_inst.envelope_inst.vol_regs[0][6] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold209 (.A(\tt6581_inst.controller_inst.pw_hi_i[10] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0239_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold211 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold212 (.A(\tt6581_inst.mult_inst.b_reg[14] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0354_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold214 (.A(\tt6581_inst.mult_inst.b_reg[15] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0355_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0067_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold217 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][1] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold218 (.A(\tt6581_inst.mult_inst.a_reg[20] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0319_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold220 (.A(\tt6581_inst.spi_inst.shift_reg[6] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold221 (.A(_3067_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0395_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold223 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][4] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold224 (.A(\tt6581_inst.envelope_inst.vol_regs[1][4] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold225 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][9] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold226 (.A(\tt6581_inst.mult_inst.b_reg[12] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold227 (.A(\tt6581_inst.mult_inst.a_reg[22] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0321_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0085_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold230 (.A(\tt6581_inst.mult_inst.accum[6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0362_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold232 (.A(\tt6581_inst.envelope_inst.vol_regs[0][16] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold233 (.A(\tt6581_inst.envelope_inst.vol_regs[1][6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold234 (.A(\tt6581_inst.mult_inst.a_reg[38] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold235 (.A(_2511_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold236 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][14] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold237 (.A(\tt6581_inst.controller_inst.freq_lo_i[8] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0149_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold239 (.A(\tt6581_inst.envelope_inst.vol_regs[0][12] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold240 (.A(\tt6581_inst.envelope_inst.vol_regs[1][17] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold241 (.A(\tt6581_inst.tick_gen_inst.cnt[3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0035_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold243 (.A(\tt6581_inst.envelope_inst.vol_regs[1][8] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold244 (.A(\tt6581_inst.controller_inst.pw_hi_i[8] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0237_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold246 (.A(\tt6581_inst.mult_inst.a_reg[7] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0306_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold248 (.A(\tt6581_inst.mult_inst.a_reg[3] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0302_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold250 (.A(\tt6581_inst.mult_inst.accum[4] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0360_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold252 (.A(\tt6581_inst.spi_inst.shift_reg[3] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold253 (.A(_4194_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0780_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold255 (.A(\tt6581_inst.delta_sigma_inst.e1[9] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0089_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold257 (.A(\tt6581_inst.envelope_inst.vol_regs[2][20] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0040_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0444_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold260 (.A(\tt6581_inst.delta_sigma_inst.e1[11] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold261 (.A(\tt6581_inst.envelope_inst.vol_regs[1][20] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold262 (.A(\tt6581_inst.envelope_inst.vol_regs[2][1] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold263 (.A(\tt6581_inst.controller_inst.pw_hi_i[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0251_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold265 (.A(\tt6581_inst.ad_pack[20] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0740_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0068_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0079_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0048_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0098_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0101_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold272 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][16] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold273 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][0] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold274 (.A(\tt6581_inst.envelope_inst.vol_regs[0][8] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0109_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold276 (.A(\tt6581_inst.envelope_inst.vol_regs[1][18] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0082_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold278 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][16] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold279 (.A(\tt6581_inst.envelope_inst.vol_regs[2][13] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0087_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0066_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold282 (.A(\tt6581_inst.mult_inst.accum[2] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0358_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold284 (.A(\tt6581_inst.envelope_inst.vol_regs[1][19] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold285 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[1][0] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0095_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0073_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold288 (.A(\tt6581_inst.controller_inst.pw_hi_i[15] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0244_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0100_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold291 (.A(\tt6581_inst.envelope_inst.vol_regs[2][21] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0058_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold293 (.A(\tt6581_inst.controller_inst.pw_hi_i[22] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold294 (.A(\tt6581_inst.controller_inst.pw_hi_i[23] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0719_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0091_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold297 (.A(\tt6581_inst.filt_en_mode[6] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0104_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold299 (.A(\tt6581_inst.envelope_inst.vol_regs[2][7] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold300 (.A(\tt6581_inst.envelope_inst.vol_regs[0][11] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0055_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold302 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][13] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold303 (.A(\tt6581_inst.envelope_inst.vol_regs[0][20] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0065_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold305 (.A(\tt6581_inst.envelope_inst.vol_regs[0][2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold306 (.A(\tt6581_inst.envelope_inst.vol_regs[2][8] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold307 (.A(\tt6581_inst.envelope_inst.vol_regs[0][15] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold308 (.A(\tt6581_inst.envelope_inst.vol_regs[2][16] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0070_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold310 (.A(\tt6581_inst.controller_inst.pw_hi_i[13] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0054_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold312 (.A(\tt6581_inst.svf_inst.reg_band[2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0105_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold314 (.A(\tt6581_inst.envelope_inst.vol_regs[2][5] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold315 (.A(\tt6581_inst.multi_voice_inst.phase_regs[2][0] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0053_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0062_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold318 (.A(\tt6581_inst.envelope_inst.vol_regs[1][1] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0060_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0051_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold321 (.A(\tt6581_inst.envelope_inst.vol_regs[2][15] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0112_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0071_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0052_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0078_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold326 (.A(\tt6581_inst.envelope_inst.vol_regs[2][3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0097_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold328 (.A(\tt6581_inst.envelope_inst.vol_regs[0][3] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0111_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0083_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold331 (.A(\tt6581_inst.envelope_inst.vol_regs[1][5] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold332 (.A(\tt6581_inst.filt_en_mode[7] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0669_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold334 (.A(\tt6581_inst.bypass_accum[6] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0823_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold336 (.A(\tt6581_inst.controller_inst.pw_hi_i[21] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0107_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0103_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0081_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold340 (.A(\tt6581_inst.envelope_inst.vol_regs[0][18] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold341 (.A(\tt6581_inst.controller_inst.pw_lo_i[22] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0710_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold343 (.A(\tt6581_inst.mult_inst.a_reg[17] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0316_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold345 (.A(\tt6581_inst.envelope_inst.vol_regs[1][15] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold346 (.A(\tt6581_inst.svf_inst.reg_band[4] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0424_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0047_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold349 (.A(\tt6581_inst.controller_inst.pw_hi_i[12] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0241_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0093_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold352 (.A(\tt6581_inst.envelope_inst.vol_regs[2][17] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold353 (.A(\tt6581_inst.envelope_inst.vol_regs[2][9] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold354 (.A(\tt6581_inst.envelope_inst.vol_regs[2][12] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold355 (.A(\tt6581_inst.mult_inst.accum[36] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0392_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0046_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold358 (.A(\tt6581_inst.svf_inst.reg_low[0] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0106_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0074_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold361 (.A(\tt6581_inst.control_pack[3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0064_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold363 (.A(\tt6581_inst.envelope_inst.vol_regs[1][13] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold364 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[2][0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold365 (.A(\tt6581_inst.envelope_inst.vol_regs[1][7] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold366 (.A(\tt6581_inst.controller_inst.pw_hi_i[7] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0252_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold368 (.A(\tt6581_inst.envelope_inst.vol_regs[2][18] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold369 (.A(\tt6581_inst.controller_inst.freq_hi_i[18] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold370 (.A(\tt6581_inst.envelope_inst.vol_regs[2][6] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0072_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold372 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0088_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold374 (.A(\tt6581_inst.bypass_accum[7] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold375 (.A(_4416_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0057_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold377 (.A(\tt6581_inst.envelope_inst.vol_regs[0][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold378 (.A(\tt6581_inst.envelope_inst.vol_regs[2][11] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0056_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0102_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold381 (.A(\tt6581_inst.control_pack[11] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0224_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0077_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold384 (.A(\tt6581_inst.envelope_inst.vol_regs[0][5] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold385 (.A(\tt6581_inst.envelope_inst.vol_regs[1][21] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold386 (.A(\tt6581_inst.envelope_inst.vol_regs[1][11] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0076_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0080_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0063_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0045_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0086_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold392 (.A(\tt6581_inst.envelope_inst.vol_regs[1][2] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0099_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold394 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][16] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0044_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0096_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold397 (.A(\tt6581_inst.envelope_inst.vol_regs[0][7] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold398 (.A(\tt6581_inst.envelope_inst.vol_regs[0][21] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold399 (.A(\tt6581_inst.delta_sigma_inst.e2[17] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0292_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0094_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold402 (.A(\tt6581_inst.envelope_inst.vol_regs[0][13] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold403 (.A(\tt6581_inst.envelope_inst.vol_regs[0][17] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold404 (.A(\tt6581_inst.envelope_inst.vol_regs[2][2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold405 (.A(\tt6581_inst.svf_inst.reg_band[7] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0427_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold407 (.A(\tt6581_inst.mult_inst.accum[1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0357_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0050_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold410 (.A(\tt6581_inst.mult_inst.accum[0] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold411 (.A(_2797_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0356_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold413 (.A(\tt6581_inst.envelope_inst.vol_regs[1][3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold414 (.A(\tt6581_inst.controller_inst.freq_hi_i[14] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold415 (.A(\tt6581_inst.envelope_inst.vol_regs[2][19] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0110_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold417 (.A(\tt6581_inst.mult_inst.accum[3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0359_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0084_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold420 (.A(\tt6581_inst.multi_voice_inst.phase_regs[0][10] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold421 (.A(\tt6581_inst.delta_sigma_inst.audio[6] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold422 (.A(\tt6581_inst.controller_inst.freq_hi_i[19] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0691_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold424 (.A(\tt6581_inst.envelope_inst.vol_regs[0][1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0049_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold426 (.A(\tt6581_inst.controller_inst.pw_hi_i[5] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0250_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold428 (.A(\tt6581_inst.controller_inst.cur_voice[1] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold429 (.A(\tt6581_inst.controller_inst.freq_hi_i[17] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0689_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0075_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold432 (.A(\tt6581_inst.multi_voice_inst.phase_regs[1][0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold433 (.A(\tt6581_inst.delta_sigma_inst.audio[5] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold434 (.A(\tt6581_inst.envelope_inst.vol_regs[0][19] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold435 (.A(\tt6581_inst.control_pack[10] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0223_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold437 (.A(\tt6581_inst.spi_inst.bit_cnt[1] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0793_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold439 (.A(\tt6581_inst.delta_sigma_inst.e1[7] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold440 (.A(\tt6581_inst.mult_inst.accum[15] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0371_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold442 (.A(\tt6581_inst.control_pack[19] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold443 (.A(\tt6581_inst.tick_gen_inst.cnt[5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold444 (.A(_1031_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold445 (.A(\tt6581_inst.delta_sigma_inst.e1[15] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold446 (.A(\tt6581_inst.delta_sigma_inst.e1[1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0257_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0059_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold449 (.A(\tt6581_inst.filter_accum[6] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold450 (.A(_4106_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0654_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold452 (.A(\tt6581_inst.mult_inst.a_reg[24] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold453 (.A(_2497_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold454 (.A(\tt6581_inst.delta_sigma_inst.e1[5] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold455 (.A(\tt6581_inst.bypass_accum[8] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0825_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold457 (.A(\tt6581_inst.mult_inst.a_reg[32] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold458 (.A(_2505_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold459 (.A(\tt6581_inst.mult_inst.a_reg[35] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold460 (.A(_2508_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold461 (.A(\tt6581_inst.bypass_accum[12] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0829_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold463 (.A(\tt6581_inst.delta_sigma_inst.e1[0] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold464 (.A(\tt6581_inst.controller_inst.pw_hi_i[4] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0249_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold466 (.A(\tt6581_inst.mult_inst.accum[12] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0368_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold468 (.A(\tt6581_inst.controller_inst.freq_hi_i[16] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0688_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold470 (.A(\tt6581_inst.mult_inst.accum[22] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0378_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold472 (.A(\tt6581_inst.controller_inst.pw_hi_i[20] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0716_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold474 (.A(\tt6581_inst.svf_inst.hp_node[16] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold475 (.A(\tt6581_inst.svf_inst.hp_node[22] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0187_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold477 (.A(\tt6581_inst.tick_gen_inst.cnt[6] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold478 (.A(_1033_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold479 (.A(\tt6581_inst.controller_inst.pw_hi_i[1] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0246_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold481 (.A(\tt6581_inst.controller_inst.pw_hi_i[14] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold482 (.A(\tt6581_inst.multi_voice_inst.phase_last_msb[0][0] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold483 (.A(\tt6581_inst.mult_inst.a_reg[36] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold484 (.A(\tt6581_inst.reg_addr[6] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0782_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold486 (.A(\tt6581_inst.mult_inst.a_reg[33] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold487 (.A(\tt6581_inst.controller_inst.pw_lo_i[13] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0122_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold489 (.A(\tt6581_inst.delta_sigma_inst.e1[17] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold490 (.A(\tt6581_inst.delta_sigma_inst.e1[13] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold491 (.A(\tt6581_inst.svf_inst.hp_node[14] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold492 (.A(\tt6581_inst.bypass_accum[10] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0827_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold494 (.A(\tt6581_inst.mult_inst.a_reg[29] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold495 (.A(_2502_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold496 (.A(\tt6581_inst.controller_inst.freq_lo_i[22] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0686_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold498 (.A(\tt6581_inst.controller_inst.pw_lo_i[7] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0132_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold500 (.A(\tt6581_inst.mult_inst.a_reg[25] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold501 (.A(\tt6581_inst.tick_gen_inst.cnt[7] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold502 (.A(\tt6581_inst.controller_inst.freq_lo_i[20] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0684_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold504 (.A(\tt6581_inst.mult_inst.a_reg[11] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0310_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold506 (.A(\tt6581_inst.reg_addr[5] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0781_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold508 (.A(\tt6581_inst.mult_inst.a_reg[37] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold509 (.A(\tt6581_inst.ad_pack[6] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold510 (.A(\tt6581_inst.svf_inst.hp_node[23] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold511 (.A(\tt6581_inst.svf_inst.reg_band[17] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0437_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold513 (.A(\tt6581_inst.mult_inst.a_reg[30] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold514 (.A(\tt6581_inst.controller_inst.freq_hi_i[15] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0140_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold516 (.A(\tt6581_inst.mult_inst.a_reg[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0301_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold518 (.A(\tt6581_inst.filter_accum[7] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold519 (.A(_4112_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold520 (.A(\tt6581_inst.tick_gen_inst.cnt[8] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold521 (.A(\tt6581_inst.controller_inst.freq_lo_i[18] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0682_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold523 (.A(\tt6581_inst.controller_inst.pw_lo_i[20] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0708_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold525 (.A(\tt6581_inst.mult_inst.a_reg[21] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold526 (.A(\tt6581_inst.controller_inst.freq_hi_i[6] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0147_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold528 (.A(\tt6581_inst.mult_inst.a_reg[10] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0309_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold530 (.A(\tt6581_inst.mult_inst.a_reg[34] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold531 (.A(\tt6581_inst.mult_inst.accum[9] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0365_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold533 (.A(\tt6581_inst.controller_inst.pw_lo_i[3] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold534 (.A(\tt6581_inst.svf_inst.hp_node[20] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold535 (.A(\tt6581_inst.svf_inst.reg_band[3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold536 (.A(_3224_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0423_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold538 (.A(\tt6581_inst.controller_inst.freq_lo_i[17] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold539 (.A(_0681_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold540 (.A(\tt6581_inst.control_pack[16] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold541 (.A(\tt6581_inst.delta_sigma_inst.e1[2] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold542 (.A(\tt6581_inst.controller_inst.pw_hi_i[9] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0238_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold544 (.A(\tt6581_inst.controller_inst.cur_voice[0] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0254_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold546 (.A(\tt6581_inst.bypass_accum[13] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0830_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold548 (.A(\tt6581_inst.mult_inst.accum[29] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0385_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold550 (.A(\tt6581_inst.controller_inst.freq_hi_i[7] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0148_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold552 (.A(\tt6581_inst.spi_inst.bit_cnt[2] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0794_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold554 (.A(\tt6581_inst.mult_inst.a_reg[13] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0312_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold556 (.A(\tt6581_inst.controller_inst.freq_hi_i[11] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0136_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold558 (.A(\tt6581_inst.mult_inst.a_reg[27] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold559 (.A(_2500_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold560 (.A(\tt6581_inst.control_pack[6] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0235_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold562 (.A(\tt6581_inst.controller_inst.pw_hi_i[19] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold563 (.A(_0715_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold564 (.A(\tt6581_inst.mult_inst.accum[20] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold565 (.A(\tt6581_inst.control_pack[18] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold566 (.A(\tt6581_inst.control_pack[5] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0234_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold568 (.A(\tt6581_inst.controller_inst.filt_en_i[0] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0665_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold570 (.A(\tt6581_inst.controller_inst.pw_lo_i[11] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0120_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold572 (.A(\tt6581_inst.svf_inst.hp_node[2] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0167_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold574 (.A(\tt6581_inst.controller_inst.sr_i[16] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold575 (.A(\tt6581_inst.controller_inst.pw_lo_i[15] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0124_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold577 (.A(\tt6581_inst.control_pack[2] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold578 (.A(\tt6581_inst.delta_sigma_inst.e2[7] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold579 (.A(\tt6581_inst.filt_q_hi[0] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0696_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold581 (.A(\tt6581_inst.mult_inst.accum[28] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0384_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold583 (.A(\tt6581_inst.filter_accum[8] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold584 (.A(_4117_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold585 (.A(\tt6581_inst.mult_inst.accum[30] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0386_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold587 (.A(\tt6581_inst.control_pack[22] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0726_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold589 (.A(\tt6581_inst.controller_inst.pw_lo_i[16] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0704_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold591 (.A(\tt6581_inst.control_pack[20] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0724_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold593 (.A(\tt6581_inst.controller_inst.freq_hi_i[2] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold594 (.A(\tt6581_inst.controller_inst.freq_hi_i[13] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0138_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold596 (.A(\tt6581_inst.controller_inst.freq_hi_i[1] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0142_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold598 (.A(\tt6581_inst.filt_q_hi[3] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0699_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold600 (.A(\tt6581_inst.control_pack[7] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold601 (.A(_0236_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold602 (.A(\tt6581_inst.mult_inst.a_reg[26] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold603 (.A(\tt6581_inst.controller_inst.freq_hi_i[3] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0144_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold605 (.A(\tt6581_inst.mult_inst.a_reg[19] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold606 (.A(\tt6581_inst.bypass_accum[1] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold607 (.A(\tt6581_inst.filt_q_hi[6] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold608 (.A(\tt6581_inst.controller_inst.freq_lo_i[4] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0161_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold610 (.A(\tt6581_inst.filt_f_lo[6] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold611 (.A(\tt6581_inst.delta_sigma_inst.cnt[1] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold612 (.A(\tt6581_inst.ad_pack[7] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold613 (.A(_0220_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold614 (.A(\tt6581_inst.controller_inst.pw_lo_i[14] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold615 (.A(\tt6581_inst.svf_inst.hp_node[0] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0165_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold617 (.A(\tt6581_inst.svf_inst.reg_band[12] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold618 (.A(_3273_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0432_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold620 (.A(\tt6581_inst.filter_accum[10] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold621 (.A(_4126_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0658_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold623 (.A(\tt6581_inst.spi_inst.shift_reg[5] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0801_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold625 (.A(\tt6581_inst.controller_inst.pw_lo_i[18] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold626 (.A(\tt6581_inst.filt_volume[0] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold627 (.A(_0760_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold628 (.A(\tt6581_inst.controller_inst.pw_lo_i[21] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0709_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold630 (.A(\tt6581_inst.controller_inst.pw_lo_i[19] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold631 (.A(\tt6581_inst.delta_sigma_inst.e1[14] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold632 (.A(\tt6581_inst.delta_sigma_inst.e2[2] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold633 (.A(\tt6581_inst.controller_inst.sr_i[17] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0753_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold635 (.A(\tt6581_inst.ad_pack[21] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold636 (.A(_0741_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold637 (.A(\tt6581_inst.mult_inst.accum[21] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold638 (.A(\tt6581_inst.filt_q_lo[0] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold639 (.A(\tt6581_inst.ad_pack[4] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold640 (.A(_0217_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold641 (.A(\tt6581_inst.delta_sigma_inst.audio[7] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold642 (.A(\tt6581_inst.delta_sigma_inst.e2[6] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0281_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold644 (.A(\tt6581_inst.controller_inst.freq_lo_i[21] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0685_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold646 (.A(\tt6581_inst.controller_inst.freq_hi_i[10] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold647 (.A(\tt6581_inst.delta_sigma_inst.e2[12] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0287_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold649 (.A(\tt6581_inst.mult_inst.a_reg[12] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold650 (.A(\tt6581_inst.delta_sigma_inst.e2[11] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold651 (.A(\tt6581_inst.controller_inst.freq_lo_i[6] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold652 (.A(_0163_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold653 (.A(\tt6581_inst.controller_inst.sr_i[12] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold654 (.A(_0201_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold655 (.A(\tt6581_inst.ad_pack[8] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold656 (.A(\tt6581_inst.controller_inst.pw_lo_i[23] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold657 (.A(_0711_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold658 (.A(\tt6581_inst.filt_q_hi[7] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold659 (.A(_0703_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold660 (.A(\tt6581_inst.delta_sigma_inst.audio[8] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold661 (.A(\tt6581_inst.delta_sigma_inst.e2[8] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0283_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold663 (.A(\tt6581_inst.control_pack[4] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0233_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold665 (.A(\tt6581_inst.mult_inst.accum[14] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0370_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold667 (.A(\tt6581_inst.ad_pack[5] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold668 (.A(_0218_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold669 (.A(\tt6581_inst.svf_inst.hp_node[18] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold670 (.A(\tt6581_inst.mult_inst.a_reg[28] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold671 (.A(\tt6581_inst.controller_inst.freq_lo_i[2] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold672 (.A(\tt6581_inst.controller_inst.freq_lo_i[14] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold673 (.A(_0155_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold674 (.A(\tt6581_inst.filt_f_hi[4] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold675 (.A(\tt6581_inst.controller_inst.pw_lo_i[12] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold676 (.A(_0121_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold677 (.A(\tt6581_inst.controller_inst.sr_i[19] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold678 (.A(_0755_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold679 (.A(\tt6581_inst.filt_f_lo[4] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0676_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold681 (.A(\tt6581_inst.mult_inst.accum[35] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0391_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold683 (.A(\tt6581_inst.controller_inst.freq_hi_i[0] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0141_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold685 (.A(\tt6581_inst.svf_inst.hp_node[5] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold686 (.A(\tt6581_inst.delta_sigma_inst.e2[3] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold687 (.A(_0278_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold688 (.A(\tt6581_inst.filt_volume[3] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0763_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold690 (.A(\tt6581_inst.svf_inst.hp_node[6] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold691 (.A(_1146_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold692 (.A(_0171_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold693 (.A(\tt6581_inst.controller_inst.freq_lo_i[23] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0687_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold695 (.A(\tt6581_inst.svf_inst.hp_node[12] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold696 (.A(_1236_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold697 (.A(_0177_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold698 (.A(\tt6581_inst.mult_inst.accum[34] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold699 (.A(\tt6581_inst.spi_inst.shift_reg[1] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold700 (.A(_0770_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold701 (.A(\tt6581_inst.filt_q_hi[5] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold702 (.A(\tt6581_inst.svf_inst.reg_band[11] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold703 (.A(_3262_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold704 (.A(_0431_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold705 (.A(\tt6581_inst.filt_q_lo[7] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0735_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold707 (.A(\tt6581_inst.filt_volume[6] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold708 (.A(_0766_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold709 (.A(\tt6581_inst.controller_inst.freq_lo_i[13] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0154_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold711 (.A(\tt6581_inst.filt_f_hi[6] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold712 (.A(\tt6581_inst.control_pack[1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0230_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold714 (.A(\tt6581_inst.controller_inst.freq_hi_i[9] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold715 (.A(_0134_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold716 (.A(\tt6581_inst.controller_inst.sr_i[8] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold717 (.A(\tt6581_inst.filt_q_hi[1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold718 (.A(_0697_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold719 (.A(\tt6581_inst.controller_inst.pw_lo_i[9] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0118_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold721 (.A(\tt6581_inst.controller_inst.freq_lo_i[11] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold722 (.A(\tt6581_inst.svf_inst.hp_node[4] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold723 (.A(_1118_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold724 (.A(_0169_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold725 (.A(\tt6581_inst.control_pack[23] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold726 (.A(\tt6581_inst.ad_pack[12] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold727 (.A(_0209_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold728 (.A(\tt6581_inst.controller_inst.freq_lo_i[15] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold729 (.A(_0156_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold730 (.A(\tt6581_inst.mult_inst.a_reg[6] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold731 (.A(\tt6581_inst.controller_inst.freq_lo_i[1] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold732 (.A(_0158_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold733 (.A(pdm),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold734 (.A(\tt6581_inst.controller_inst.sample_tick_i ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold735 (.A(\tt6581_inst.ad_pack[11] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold736 (.A(_0208_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold737 (.A(\tt6581_inst.delta_sigma_inst.e1[3] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold738 (.A(_0259_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold739 (.A(\tt6581_inst.controller_inst.filt_en_i[2] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold740 (.A(\tt6581_inst.reg_addr[2] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold741 (.A(_0778_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold742 (.A(\tt6581_inst.delta_sigma_inst.audio[14] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold743 (.A(\tt6581_inst.controller_inst.pw_lo_i[6] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold744 (.A(\tt6581_inst.filt_q_lo[1] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold745 (.A(_0729_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold746 (.A(\tt6581_inst.spi_inst.shift_reg[2] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold747 (.A(\tt6581_inst.filt_f_lo[1] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold748 (.A(_0673_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold749 (.A(\tt6581_inst.control_pack[8] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold750 (.A(_0221_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold751 (.A(\tt6581_inst.mult_inst.a_reg[23] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold752 (.A(\tt6581_inst.controller_inst.sr_i[20] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold753 (.A(_0756_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold754 (.A(\tt6581_inst.filt_volume[5] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold755 (.A(_0765_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold756 (.A(\tt6581_inst.delta_sigma_inst.e2[1] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold757 (.A(\tt6581_inst.filt_q_hi[4] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold758 (.A(\tt6581_inst.spi_inst.shift_reg[0] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold759 (.A(\tt6581_inst.ad_pack[22] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold760 (.A(\tt6581_inst.controller_inst.freq_hi_i[8] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold761 (.A(_0133_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold762 (.A(\tt6581_inst.control_pack[9] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold763 (.A(_0222_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold764 (.A(\tt6581_inst.svf_inst.reg_band[16] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold765 (.A(_0436_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold766 (.A(\tt6581_inst.delta_sigma_inst.e1[16] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold767 (.A(\tt6581_inst.reg_file_inst.wdata_i[1] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold768 (.A(\tt6581_inst.filt_f_hi[7] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold769 (.A(_0751_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold770 (.A(\tt6581_inst.filt_f_lo[3] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold771 (.A(_0675_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold772 (.A(\tt6581_inst.controller_inst.freq_lo_i[5] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0162_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold774 (.A(\tt6581_inst.controller_inst.freq_lo_i[0] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold775 (.A(_0157_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold776 (.A(\tt6581_inst.delta_sigma_inst.e2[9] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold777 (.A(\tt6581_inst.svf_inst.hp_node[21] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold778 (.A(\tt6581_inst.mult_inst.a_reg[8] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold779 (.A(\tt6581_inst.filt_q_lo[6] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold780 (.A(\tt6581_inst.controller_inst.sr_i[9] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold781 (.A(\tt6581_inst.spi_inst.mosi_sync[1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold782 (.A(_0768_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold783 (.A(\tt6581_inst.controller_inst.freq_lo_i[10] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold784 (.A(_0151_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold785 (.A(\tt6581_inst.filt_f_lo[5] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold786 (.A(_0677_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold787 (.A(\tt6581_inst.reg_addr[3] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold788 (.A(_0779_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold789 (.A(\tt6581_inst.controller_inst.freq_lo_i[3] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold790 (.A(\tt6581_inst.delta_sigma_inst.audio[9] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold791 (.A(\tt6581_inst.mult_inst.a_reg[31] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold792 (.A(\tt6581_inst.mult_inst.a_reg[0] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold793 (.A(\tt6581_inst.svf_inst.reg_band[9] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold794 (.A(_3255_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold795 (.A(_0429_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold796 (.A(\tt6581_inst.reg_addr[0] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold797 (.A(_0776_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold798 (.A(\tt6581_inst.spi_inst.bit_cnt[3] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold799 (.A(_0795_),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold800 (.A(\tt6581_inst.tick_gen_inst.cnt[9] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold801 (.A(\tt6581_inst.spi_inst.cs_sync[1] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold802 (.A(\tt6581_inst.svf_inst.reg_band[1] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold803 (.A(_3207_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold804 (.A(_0421_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold805 (.A(\tt6581_inst.controller_inst.pw_lo_i[10] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold806 (.A(\tt6581_inst.controller_inst.pw_hi_i[3] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold807 (.A(\tt6581_inst.delta_sigma_inst.audio[11] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold808 (.A(\tt6581_inst.filt_q_lo[3] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold809 (.A(_0731_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold810 (.A(\tt6581_inst.controller_inst.freq_hi_i[4] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold811 (.A(_0145_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold812 (.A(\tt6581_inst.controller_inst.freq_hi_i[23] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold813 (.A(\tt6581_inst.delta_sigma_inst.e1[10] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold814 (.A(\tt6581_inst.filt_volume[2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold815 (.A(_0762_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold816 (.A(\tt6581_inst.mult_inst.accum[19] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold817 (.A(_0375_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold818 (.A(\tt6581_inst.filt_q_hi[2] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold819 (.A(\tt6581_inst.ad_pack[9] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold820 (.A(\tt6581_inst.spi_inst.sclk_sync[2] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold821 (.A(\tt6581_inst.filt_volume[1] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold822 (.A(\tt6581_inst.svf_inst.hp_node[7] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold823 (.A(_1158_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold824 (.A(_0172_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold825 (.A(\tt6581_inst.delta_sigma_inst.audio[16] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold826 (.A(\tt6581_inst.svf_inst.hp_node[17] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold827 (.A(\tt6581_inst.control_pack[0] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold828 (.A(_0229_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold829 (.A(\tt6581_inst.svf_inst.reg_band[5] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold830 (.A(_3231_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold831 (.A(_0425_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold832 (.A(\tt6581_inst.ad_pack[16] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold833 (.A(_0736_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold834 (.A(\tt6581_inst.filt_q_lo[4] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold835 (.A(\tt6581_inst.controller_inst.sr_i[5] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold836 (.A(_0194_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold837 (.A(\tt6581_inst.svf_inst.reg_band[14] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold838 (.A(_0434_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold839 (.A(\tt6581_inst.svf_inst.hp_node[8] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold840 (.A(_1172_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold841 (.A(_0173_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold842 (.A(\tt6581_inst.control_pack[12] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold843 (.A(_0225_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold844 (.A(\tt6581_inst.delta_sigma_inst.e1[6] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold845 (.A(\tt6581_inst.delta_sigma_inst.e2[14] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold846 (.A(\tt6581_inst.mult_inst.a_reg[9] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold847 (.A(_0308_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold848 (.A(\tt6581_inst.controller_inst.filt_en_i[1] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold849 (.A(_0666_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold850 (.A(\tt6581_inst.delta_sigma_inst.e2[15] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold851 (.A(\tt6581_inst.svf_inst.reg_band[15] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold852 (.A(_0435_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold853 (.A(\tt6581_inst.controller_inst.pw_hi_i[0] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold854 (.A(_0245_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold855 (.A(\tt6581_inst.svf_inst.reg_band[8] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold856 (.A(\tt6581_inst.mult_inst.iter[2] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold857 (.A(_1594_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold858 (.A(\tt6581_inst.controller_inst.sr_i[18] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold859 (.A(_0754_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold860 (.A(\tt6581_inst.controller_inst.pw_hi_i[17] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold861 (.A(\tt6581_inst.controller_inst.freq_lo_i[16] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold862 (.A(_0680_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold863 (.A(\tt6581_inst.controller_inst.pw_hi_i[18] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold864 (.A(\tt6581_inst.delta_sigma_inst.e2[16] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold865 (.A(\tt6581_inst.filt_f_lo[0] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold866 (.A(_0672_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold867 (.A(\tt6581_inst.svf_inst.hp_node[13] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold868 (.A(_0178_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold869 (.A(\tt6581_inst.controller_inst.freq_hi_i[22] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold870 (.A(_0694_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold871 (.A(\tt6581_inst.controller_inst.pw_hi_i[16] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold872 (.A(_0712_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold873 (.A(\tt6581_inst.ad_pack[23] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold874 (.A(_0743_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold875 (.A(\tt6581_inst.reg_addr[1] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold876 (.A(\tt6581_inst.delta_sigma_inst.e1[8] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold877 (.A(\tt6581_inst.filt_f_hi[1] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold878 (.A(\tt6581_inst.controller_inst.pw_hi_i[11] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold879 (.A(_0240_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold880 (.A(\tt6581_inst.control_pack[17] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold881 (.A(\tt6581_inst.controller_inst.sr_i[11] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold882 (.A(_0200_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold883 (.A(\tt6581_inst.filt_volume[7] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold884 (.A(_0767_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold885 (.A(\tt6581_inst.delta_sigma_inst.e2[10] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold886 (.A(\tt6581_inst.ad_pack[0] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold887 (.A(\tt6581_inst.svf_inst.reg_band[10] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold888 (.A(_3261_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold889 (.A(_0430_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold890 (.A(\tt6581_inst.filt_f_hi[0] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold891 (.A(_0744_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold892 (.A(\tt6581_inst.delta_sigma_inst.audio[15] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold893 (.A(\tt6581_inst.filt_f_hi[3] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold894 (.A(_0747_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold895 (.A(\tt6581_inst.svf_inst.reg_band[21] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold896 (.A(_3321_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold897 (.A(_0441_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold898 (.A(\tt6581_inst.filt_f_hi[5] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold899 (.A(\tt6581_inst.filt_f_lo[2] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold900 (.A(_0674_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold901 (.A(\tt6581_inst.controller_inst.freq_hi_i[5] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold902 (.A(_0146_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold903 (.A(\tt6581_inst.delta_sigma_inst.audio[10] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold904 (.A(\tt6581_inst.controller_inst.freq_lo_i[12] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold905 (.A(_0153_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold906 (.A(\tt6581_inst.ad_pack[10] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold907 (.A(_0207_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold908 (.A(\tt6581_inst.controller_inst.sr_i[0] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold909 (.A(\tt6581_inst.control_pack[13] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold910 (.A(_0226_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold911 (.A(\tt6581_inst.controller_inst.pw_lo_i[2] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold912 (.A(\tt6581_inst.svf_inst.reg_band[13] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold913 (.A(_0433_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold914 (.A(\tt6581_inst.reg_file_inst.wdata_i[6] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold915 (.A(\tt6581_inst.controller_inst.sr_i[15] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold916 (.A(_0204_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold917 (.A(\tt6581_inst.delta_sigma_inst.audio[12] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold918 (.A(\tt6581_inst.controller_inst.sr_i[23] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold919 (.A(_0759_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold920 (.A(\tt6581_inst.delta_sigma_inst.e2[5] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold921 (.A(\tt6581_inst.controller_inst.pw_hi_i[2] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold922 (.A(\tt6581_inst.delta_sigma_inst.e2[13] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold923 (.A(\tt6581_inst.controller_inst.sr_i[7] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold924 (.A(_0196_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold925 (.A(\tt6581_inst.ad_pack[13] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold926 (.A(_0210_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold927 (.A(\tt6581_inst.controller_inst.pw_lo_i[5] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold928 (.A(_0130_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold929 (.A(\tt6581_inst.controller_inst.sr_i[6] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold930 (.A(\tt6581_inst.filter_accum[1] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold931 (.A(_0649_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold932 (.A(\tt6581_inst.svf_inst.hp_node[10] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold933 (.A(_1196_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold934 (.A(_0175_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold935 (.A(\tt6581_inst.delta_sigma_inst.e1[4] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold936 (.A(\tt6581_inst.reg_file_inst.wdata_i[7] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold937 (.A(\tt6581_inst.controller_inst.sr_i[14] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold938 (.A(\tt6581_inst.mult_inst.a_reg[14] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold939 (.A(\tt6581_inst.delta_sigma_inst.audio[4] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold940 (.A(\tt6581_inst.filt_en_mode[2] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold941 (.A(\tt6581_inst.ad_pack[1] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold942 (.A(\tt6581_inst.mult_inst.iter[3] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold943 (.A(_1596_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold944 (.A(\tt6581_inst.filt_f_lo[7] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold945 (.A(\tt6581_inst.delta_sigma_inst.e2[4] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold946 (.A(\tt6581_inst.svf_inst.reg_low[4] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold947 (.A(\tt6581_inst.mult_inst.a_reg[1] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold948 (.A(_0300_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold949 (.A(\tt6581_inst.spi_inst.shift_reg[4] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold950 (.A(_0773_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold951 (.A(\tt6581_inst.mult_inst.accum[5] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold952 (.A(\tt6581_inst.mult_inst.accum[7] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold953 (.A(\tt6581_inst.filt_f_hi[2] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold954 (.A(\tt6581_inst.delta_sigma_inst.e1[12] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold955 (.A(\tt6581_inst.ad_pack[17] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold956 (.A(\tt6581_inst.control_pack[21] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold957 (.A(_0725_),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold958 (.A(\tt6581_inst.controller_inst.sr_i[22] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold959 (.A(\tt6581_inst.filt_volume[4] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold960 (.A(\tt6581_inst.ad_pack[18] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold961 (.A(_0738_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold962 (.A(\tt6581_inst.controller_inst.freq_hi_i[12] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold963 (.A(_0137_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold964 (.A(\tt6581_inst.spi_inst.is_write_cmd ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold965 (.A(\tt6581_inst.controller_inst.pw_lo_i[1] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold966 (.A(\tt6581_inst.svf_inst.reg_low[2] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold967 (.A(\tt6581_inst.controller_inst.freq_hi_i[21] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold968 (.A(_0693_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold969 (.A(\tt6581_inst.controller_inst.pw_lo_i[4] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold970 (.A(_0129_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold971 (.A(\tt6581_inst.svf_inst.hp_node[1] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold972 (.A(\tt6581_inst.mult_inst.accum[33] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold973 (.A(_0389_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold974 (.A(\tt6581_inst.controller_inst.freq_lo_i[9] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold975 (.A(\tt6581_inst.filt_q_lo[5] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold976 (.A(\tt6581_inst.svf_inst.reg_band[6] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold977 (.A(\tt6581_inst.svf_inst.hp_node[11] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold978 (.A(\tt6581_inst.filt_q_lo[2] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold979 (.A(_0730_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold980 (.A(\tt6581_inst.bypass_accum[3] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold981 (.A(_4399_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold982 (.A(\tt6581_inst.controller_inst.sr_i[13] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold983 (.A(\tt6581_inst.svf_inst.hp_node[9] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold984 (.A(_1184_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold985 (.A(_0174_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold986 (.A(\tt6581_inst.filter_accum[2] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold987 (.A(_0650_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold988 (.A(\tt6581_inst.controller_inst.sr_i[10] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold989 (.A(_0199_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold990 (.A(\tt6581_inst.mult_inst.a_reg[15] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold991 (.A(_0314_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold992 (.A(\tt6581_inst.controller_inst.freq_lo_i[19] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold993 (.A(_0683_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold994 (.A(\tt6581_inst.filter_accum[12] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold995 (.A(_0660_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold996 (.A(\tt6581_inst.svf_inst.reg_band[18] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold997 (.A(\tt6581_inst.controller_inst.freq_hi_i[20] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold998 (.A(_0692_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold999 (.A(\tt6581_inst.svf_inst.reg_low[23] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold1000 (.A(_0419_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\tt6581_inst.bypass_accum[5] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold1002 (.A(_0822_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\tt6581_inst.controller_inst.pw_lo_i[0] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold1004 (.A(_0125_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\tt6581_inst.delta_sigma_inst.audio[13] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\tt6581_inst.controller_inst.pw_lo_i[17] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\tt6581_inst.mult_inst.accum[37] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\tt6581_inst.ad_pack[15] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\tt6581_inst.svf_inst.reg_low[17] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold1010 (.A(_0413_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\tt6581_inst.reg_file_inst.wdata_i[4] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\tt6581_inst.controller_inst.sr_i[1] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\tt6581_inst.filter_accum[3] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_4095_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\tt6581_inst.tick_gen_inst.cnt[2] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\tt6581_inst.svf_inst.reg_low[13] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_3142_),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_0409_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\tt6581_inst.svf_inst.reg_low[21] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_0417_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\tt6581_inst.controller_inst.pw_lo_i[8] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_0117_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\tt6581_inst.bypass_accum[4] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\tt6581_inst.svf_inst.reg_band[20] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_0440_),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\tt6581_inst.ad_pack[3] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_0216_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\tt6581_inst.filt_en_mode[1] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\tt6581_inst.filter_accum[5] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_0653_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\tt6581_inst.ad_pack[2] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_0215_),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\tt6581_inst.ad_pack[14] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\tt6581_inst.svf_inst.reg_band[19] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\tt6581_inst.mult_inst.a_reg[16] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\tt6581_inst.svf_inst.reg_low[18] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\tt6581_inst.ad_pack[19] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_0739_),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\tt6581_inst.mult_inst.accum[18] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\tt6581_inst.svf_inst.reg_low[16] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\tt6581_inst.controller_inst.sr_i[2] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_0191_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\tt6581_inst.bypass_accum[9] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\tt6581_inst.mult_inst.iter[1] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\tt6581_inst.controller_inst.freq_lo_i[7] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\tt6581_inst.mult_inst.accum[25] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\tt6581_inst.bypass_accum[11] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_0828_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\tt6581_inst.mult_inst.accum[11] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_0367_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\tt6581_inst.svf_inst.reg_low[11] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_3130_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_0407_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\tt6581_inst.bypass_accum[2] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_0819_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\tt6581_inst.svf_inst.reg_low[22] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_0418_),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\tt6581_inst.mult_inst.accum[31] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_0387_),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\tt6581_inst.controller_inst.sr_i[4] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\tt6581_inst.multi_voice_inst.cur_state[0] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\tt6581_inst.filter_accum[4] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_4100_),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\tt6581_inst.svf_inst.reg_band[22] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\tt6581_inst.mult_inst.accum[27] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_0383_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\tt6581_inst.controller_inst.sr_i[3] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_0192_),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\tt6581_inst.svf_inst.hp_node[15] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_0180_),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\tt6581_inst.mult_inst.accum[32] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold1072 (.A(_3022_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\tt6581_inst.mult_inst.accum[26] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\tt6581_inst.mult_inst.accum[17] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_0373_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\tt6581_inst.svf_inst.reg_low[19] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold1077 (.A(_0415_),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\tt6581_inst.svf_inst.reg_low[15] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold1079 (.A(_0411_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\tt6581_inst.svf_inst.hp_node[3] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\tt6581_inst.svf_inst.hp_node[19] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\tt6581_inst.tick_gen_inst.cnt[2] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\tt6581_inst.filter_accum[11] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_0659_),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\tt6581_inst.mult_inst.accum[13] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\tt6581_inst.controller_inst.sr_i[21] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_0757_),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\tt6581_inst.svf_inst.reg_low[20] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold1089 (.A(_0416_),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\tt6581_inst.svf_inst.reg_low[7] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\tt6581_inst.svf_inst.reg_low[12] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_0408_),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\tt6581_inst.svf_inst.reg_low[10] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold1094 (.A(_0406_),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\tt6581_inst.filter_accum[9] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_0657_),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\tt6581_inst.mult_inst.accum[24] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\tt6581_inst.filt_en_mode[0] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_0662_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\tt6581_inst.mult_inst.accum[23] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_2953_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\tt6581_inst.mult_inst.accum[8] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\tt6581_inst.svf_inst.reg_low[8] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_0404_),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\tt6581_inst.filter_accum[13] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_0661_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\tt6581_inst.svf_inst.reg_low[14] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\tt6581_inst.mult_inst.accum[16] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\tt6581_inst.svf_inst.reg_low[3] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\tt6581_inst.svf_inst.reg_low[5] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\tt6581_inst.svf_inst.reg_low[9] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_3118_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold1113 (.A(_0405_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\tt6581_inst.mult_inst.accum[10] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\tt6581_inst.svf_inst.reg_low[1] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_0397_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\tt6581_inst.svf_inst.reg_low[6] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\tt6581_inst.svf_inst.cur_state[5] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\tt6581_inst.reg_file_inst.we_i ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\tt6581_inst.svf_inst.cur_state[7] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\tt6581_inst.svf_inst.cur_state[9] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\tt6581_inst.svf_inst.cur_state[9] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\tt6581_inst.reg_file_inst.we_i ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\tt6581_inst.mult_inst.accum[9] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\tt6581_inst.svf_inst.reg_band[1] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_0111_),
    .X(net1707));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_36 ();
 sg13g2_fill_1 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_54 ();
 sg13g2_fill_2 FILLER_0_59 ();
 sg13g2_fill_1 FILLER_0_76 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_4 FILLER_0_171 ();
 sg13g2_decap_4 FILLER_0_179 ();
 sg13g2_fill_2 FILLER_0_183 ();
 sg13g2_decap_4 FILLER_0_197 ();
 sg13g2_fill_1 FILLER_0_237 ();
 sg13g2_fill_1 FILLER_0_394 ();
 sg13g2_fill_2 FILLER_0_431 ();
 sg13g2_fill_1 FILLER_0_433 ();
 sg13g2_fill_1 FILLER_0_466 ();
 sg13g2_fill_2 FILLER_0_517 ();
 sg13g2_fill_2 FILLER_0_528 ();
 sg13g2_fill_1 FILLER_0_530 ();
 sg13g2_fill_2 FILLER_0_549 ();
 sg13g2_decap_4 FILLER_0_590 ();
 sg13g2_fill_1 FILLER_0_594 ();
 sg13g2_fill_1 FILLER_0_683 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_fill_2 FILLER_0_859 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_22 ();
 sg13g2_fill_2 FILLER_1_52 ();
 sg13g2_fill_2 FILLER_1_73 ();
 sg13g2_fill_2 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_152 ();
 sg13g2_fill_2 FILLER_1_161 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_fill_1 FILLER_1_177 ();
 sg13g2_fill_2 FILLER_1_192 ();
 sg13g2_fill_2 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_209 ();
 sg13g2_fill_1 FILLER_1_246 ();
 sg13g2_fill_2 FILLER_1_252 ();
 sg13g2_fill_1 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_269 ();
 sg13g2_fill_1 FILLER_1_271 ();
 sg13g2_fill_1 FILLER_1_440 ();
 sg13g2_fill_2 FILLER_1_455 ();
 sg13g2_fill_1 FILLER_1_484 ();
 sg13g2_fill_1 FILLER_1_595 ();
 sg13g2_fill_2 FILLER_1_619 ();
 sg13g2_fill_1 FILLER_1_635 ();
 sg13g2_fill_1 FILLER_1_655 ();
 sg13g2_fill_2 FILLER_1_665 ();
 sg13g2_decap_4 FILLER_1_731 ();
 sg13g2_fill_2 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_755 ();
 sg13g2_decap_8 FILLER_1_762 ();
 sg13g2_decap_8 FILLER_1_769 ();
 sg13g2_decap_8 FILLER_1_776 ();
 sg13g2_decap_8 FILLER_1_783 ();
 sg13g2_fill_1 FILLER_1_790 ();
 sg13g2_decap_8 FILLER_1_799 ();
 sg13g2_decap_8 FILLER_1_806 ();
 sg13g2_decap_8 FILLER_1_813 ();
 sg13g2_decap_8 FILLER_1_820 ();
 sg13g2_decap_8 FILLER_1_827 ();
 sg13g2_decap_8 FILLER_1_834 ();
 sg13g2_decap_8 FILLER_1_841 ();
 sg13g2_decap_8 FILLER_1_848 ();
 sg13g2_decap_8 FILLER_1_855 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_85 ();
 sg13g2_fill_2 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_246 ();
 sg13g2_fill_2 FILLER_2_293 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_fill_1 FILLER_2_313 ();
 sg13g2_fill_1 FILLER_2_412 ();
 sg13g2_fill_1 FILLER_2_423 ();
 sg13g2_fill_1 FILLER_2_492 ();
 sg13g2_fill_1 FILLER_2_498 ();
 sg13g2_fill_2 FILLER_2_525 ();
 sg13g2_fill_1 FILLER_2_527 ();
 sg13g2_fill_1 FILLER_2_581 ();
 sg13g2_fill_1 FILLER_2_636 ();
 sg13g2_fill_2 FILLER_2_660 ();
 sg13g2_fill_1 FILLER_2_662 ();
 sg13g2_fill_2 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_fill_2 FILLER_2_777 ();
 sg13g2_fill_1 FILLER_2_779 ();
 sg13g2_fill_2 FILLER_2_788 ();
 sg13g2_fill_2 FILLER_2_798 ();
 sg13g2_fill_1 FILLER_2_800 ();
 sg13g2_fill_2 FILLER_2_809 ();
 sg13g2_fill_1 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_fill_2 FILLER_2_859 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_98 ();
 sg13g2_fill_1 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_157 ();
 sg13g2_fill_1 FILLER_3_237 ();
 sg13g2_fill_2 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_283 ();
 sg13g2_fill_2 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_318 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_fill_2 FILLER_3_382 ();
 sg13g2_fill_2 FILLER_3_392 ();
 sg13g2_fill_1 FILLER_3_437 ();
 sg13g2_fill_1 FILLER_3_464 ();
 sg13g2_fill_2 FILLER_3_491 ();
 sg13g2_fill_1 FILLER_3_537 ();
 sg13g2_fill_1 FILLER_3_574 ();
 sg13g2_fill_1 FILLER_3_589 ();
 sg13g2_fill_1 FILLER_3_630 ();
 sg13g2_fill_2 FILLER_3_636 ();
 sg13g2_fill_1 FILLER_3_648 ();
 sg13g2_fill_1 FILLER_3_671 ();
 sg13g2_fill_1 FILLER_3_681 ();
 sg13g2_fill_1 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_4 FILLER_3_767 ();
 sg13g2_fill_2 FILLER_3_779 ();
 sg13g2_fill_1 FILLER_3_781 ();
 sg13g2_fill_2 FILLER_3_800 ();
 sg13g2_fill_1 FILLER_3_802 ();
 sg13g2_fill_2 FILLER_3_819 ();
 sg13g2_fill_1 FILLER_3_825 ();
 sg13g2_decap_8 FILLER_3_839 ();
 sg13g2_decap_8 FILLER_3_846 ();
 sg13g2_decap_8 FILLER_3_853 ();
 sg13g2_fill_2 FILLER_3_860 ();
 sg13g2_fill_1 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_76 ();
 sg13g2_fill_2 FILLER_4_161 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_183 ();
 sg13g2_fill_1 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_211 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_fill_2 FILLER_4_284 ();
 sg13g2_fill_1 FILLER_4_286 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_fill_2 FILLER_4_370 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_fill_1 FILLER_4_487 ();
 sg13g2_fill_2 FILLER_4_509 ();
 sg13g2_fill_2 FILLER_4_541 ();
 sg13g2_fill_1 FILLER_4_543 ();
 sg13g2_fill_1 FILLER_4_577 ();
 sg13g2_fill_1 FILLER_4_706 ();
 sg13g2_fill_1 FILLER_4_728 ();
 sg13g2_fill_1 FILLER_4_750 ();
 sg13g2_fill_2 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_211 ();
 sg13g2_fill_2 FILLER_5_238 ();
 sg13g2_decap_4 FILLER_5_265 ();
 sg13g2_decap_4 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_277 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_363 ();
 sg13g2_fill_2 FILLER_5_405 ();
 sg13g2_fill_1 FILLER_5_407 ();
 sg13g2_fill_1 FILLER_5_417 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_fill_2 FILLER_5_434 ();
 sg13g2_fill_1 FILLER_5_579 ();
 sg13g2_fill_1 FILLER_5_602 ();
 sg13g2_fill_2 FILLER_5_664 ();
 sg13g2_fill_1 FILLER_5_666 ();
 sg13g2_fill_1 FILLER_5_695 ();
 sg13g2_fill_1 FILLER_5_724 ();
 sg13g2_fill_2 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_790 ();
 sg13g2_fill_1 FILLER_5_827 ();
 sg13g2_fill_1 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_855 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_1 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_297 ();
 sg13g2_fill_1 FILLER_6_299 ();
 sg13g2_fill_1 FILLER_6_348 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_387 ();
 sg13g2_fill_2 FILLER_6_419 ();
 sg13g2_fill_1 FILLER_6_421 ();
 sg13g2_fill_1 FILLER_6_436 ();
 sg13g2_fill_2 FILLER_6_495 ();
 sg13g2_fill_1 FILLER_6_530 ();
 sg13g2_fill_1 FILLER_6_556 ();
 sg13g2_fill_2 FILLER_6_659 ();
 sg13g2_fill_1 FILLER_6_661 ();
 sg13g2_fill_1 FILLER_6_708 ();
 sg13g2_fill_2 FILLER_6_798 ();
 sg13g2_fill_1 FILLER_6_800 ();
 sg13g2_fill_2 FILLER_6_859 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_fill_1 FILLER_7_75 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_446 ();
 sg13g2_fill_2 FILLER_7_491 ();
 sg13g2_fill_2 FILLER_7_511 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_fill_2 FILLER_7_604 ();
 sg13g2_fill_1 FILLER_7_606 ();
 sg13g2_fill_2 FILLER_7_691 ();
 sg13g2_fill_2 FILLER_7_734 ();
 sg13g2_fill_2 FILLER_7_773 ();
 sg13g2_fill_1 FILLER_7_775 ();
 sg13g2_fill_2 FILLER_7_859 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_fill_1 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_76 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_fill_2 FILLER_8_125 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_fill_2 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_fill_2 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_266 ();
 sg13g2_decap_4 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_2 FILLER_8_411 ();
 sg13g2_fill_1 FILLER_8_413 ();
 sg13g2_fill_2 FILLER_8_423 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_fill_1 FILLER_8_505 ();
 sg13g2_fill_1 FILLER_8_547 ();
 sg13g2_fill_2 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_fill_2 FILLER_8_589 ();
 sg13g2_fill_1 FILLER_8_591 ();
 sg13g2_fill_2 FILLER_8_631 ();
 sg13g2_fill_1 FILLER_8_662 ();
 sg13g2_fill_1 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_2 FILLER_9_181 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_376 ();
 sg13g2_fill_2 FILLER_9_410 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_fill_1 FILLER_9_432 ();
 sg13g2_fill_2 FILLER_9_461 ();
 sg13g2_fill_1 FILLER_9_482 ();
 sg13g2_fill_1 FILLER_9_498 ();
 sg13g2_fill_2 FILLER_9_601 ();
 sg13g2_fill_1 FILLER_9_603 ();
 sg13g2_fill_2 FILLER_9_616 ();
 sg13g2_fill_2 FILLER_9_635 ();
 sg13g2_fill_2 FILLER_9_665 ();
 sg13g2_fill_2 FILLER_9_722 ();
 sg13g2_fill_2 FILLER_9_797 ();
 sg13g2_fill_2 FILLER_9_812 ();
 sg13g2_fill_2 FILLER_9_822 ();
 sg13g2_fill_1 FILLER_9_824 ();
 sg13g2_fill_1 FILLER_9_848 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_81 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_167 ();
 sg13g2_fill_1 FILLER_10_197 ();
 sg13g2_fill_2 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_4 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_325 ();
 sg13g2_fill_1 FILLER_10_345 ();
 sg13g2_fill_2 FILLER_10_387 ();
 sg13g2_fill_1 FILLER_10_447 ();
 sg13g2_fill_1 FILLER_10_466 ();
 sg13g2_fill_1 FILLER_10_480 ();
 sg13g2_fill_1 FILLER_10_489 ();
 sg13g2_fill_2 FILLER_10_587 ();
 sg13g2_fill_1 FILLER_10_614 ();
 sg13g2_fill_2 FILLER_10_631 ();
 sg13g2_fill_2 FILLER_10_646 ();
 sg13g2_fill_1 FILLER_10_684 ();
 sg13g2_fill_1 FILLER_10_727 ();
 sg13g2_fill_2 FILLER_10_734 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_2 FILLER_11_256 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_391 ();
 sg13g2_fill_2 FILLER_11_409 ();
 sg13g2_fill_1 FILLER_11_411 ();
 sg13g2_fill_1 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_502 ();
 sg13g2_fill_2 FILLER_11_548 ();
 sg13g2_fill_2 FILLER_11_567 ();
 sg13g2_fill_2 FILLER_11_631 ();
 sg13g2_fill_2 FILLER_11_645 ();
 sg13g2_fill_2 FILLER_11_661 ();
 sg13g2_fill_2 FILLER_11_710 ();
 sg13g2_fill_1 FILLER_11_767 ();
 sg13g2_fill_2 FILLER_11_777 ();
 sg13g2_fill_2 FILLER_11_859 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_30 ();
 sg13g2_fill_2 FILLER_12_74 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_393 ();
 sg13g2_fill_2 FILLER_12_419 ();
 sg13g2_fill_1 FILLER_12_546 ();
 sg13g2_fill_2 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_628 ();
 sg13g2_fill_1 FILLER_12_779 ();
 sg13g2_fill_2 FILLER_12_831 ();
 sg13g2_fill_1 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_fill_1 FILLER_13_286 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_419 ();
 sg13g2_fill_1 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_453 ();
 sg13g2_fill_2 FILLER_13_511 ();
 sg13g2_fill_1 FILLER_13_532 ();
 sg13g2_fill_1 FILLER_13_550 ();
 sg13g2_fill_2 FILLER_13_577 ();
 sg13g2_fill_1 FILLER_13_658 ();
 sg13g2_fill_1 FILLER_13_786 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_decap_4 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_472 ();
 sg13g2_fill_1 FILLER_14_494 ();
 sg13g2_fill_1 FILLER_14_535 ();
 sg13g2_fill_2 FILLER_14_609 ();
 sg13g2_fill_1 FILLER_14_611 ();
 sg13g2_fill_1 FILLER_14_659 ();
 sg13g2_fill_1 FILLER_14_673 ();
 sg13g2_fill_1 FILLER_14_792 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_374 ();
 sg13g2_fill_1 FILLER_15_412 ();
 sg13g2_fill_1 FILLER_15_445 ();
 sg13g2_fill_2 FILLER_15_454 ();
 sg13g2_fill_2 FILLER_15_479 ();
 sg13g2_fill_1 FILLER_15_549 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_fill_2 FILLER_15_601 ();
 sg13g2_fill_1 FILLER_15_603 ();
 sg13g2_fill_2 FILLER_15_652 ();
 sg13g2_fill_1 FILLER_15_654 ();
 sg13g2_fill_1 FILLER_15_740 ();
 sg13g2_fill_1 FILLER_15_759 ();
 sg13g2_fill_1 FILLER_15_801 ();
 sg13g2_fill_2 FILLER_15_823 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_29 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_16_410 ();
 sg13g2_fill_2 FILLER_16_439 ();
 sg13g2_fill_1 FILLER_16_497 ();
 sg13g2_fill_2 FILLER_16_533 ();
 sg13g2_fill_2 FILLER_16_616 ();
 sg13g2_fill_1 FILLER_16_683 ();
 sg13g2_fill_2 FILLER_16_699 ();
 sg13g2_fill_1 FILLER_16_790 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_421 ();
 sg13g2_fill_1 FILLER_17_449 ();
 sg13g2_fill_2 FILLER_17_459 ();
 sg13g2_fill_2 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_561 ();
 sg13g2_fill_2 FILLER_17_644 ();
 sg13g2_fill_2 FILLER_17_660 ();
 sg13g2_fill_1 FILLER_17_662 ();
 sg13g2_fill_2 FILLER_17_681 ();
 sg13g2_fill_2 FILLER_17_691 ();
 sg13g2_fill_1 FILLER_17_701 ();
 sg13g2_fill_1 FILLER_17_754 ();
 sg13g2_fill_2 FILLER_17_860 ();
 sg13g2_fill_2 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_343 ();
 sg13g2_decap_4 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_431 ();
 sg13g2_fill_1 FILLER_18_503 ();
 sg13g2_fill_2 FILLER_18_541 ();
 sg13g2_fill_1 FILLER_18_543 ();
 sg13g2_fill_2 FILLER_18_570 ();
 sg13g2_fill_1 FILLER_18_572 ();
 sg13g2_fill_2 FILLER_18_626 ();
 sg13g2_fill_1 FILLER_18_639 ();
 sg13g2_fill_1 FILLER_18_672 ();
 sg13g2_fill_2 FILLER_18_817 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_1 FILLER_19_445 ();
 sg13g2_fill_2 FILLER_19_457 ();
 sg13g2_fill_2 FILLER_19_485 ();
 sg13g2_fill_1 FILLER_19_487 ();
 sg13g2_fill_1 FILLER_19_534 ();
 sg13g2_fill_2 FILLER_19_589 ();
 sg13g2_fill_1 FILLER_19_591 ();
 sg13g2_fill_2 FILLER_19_630 ();
 sg13g2_fill_2 FILLER_19_658 ();
 sg13g2_fill_2 FILLER_19_733 ();
 sg13g2_fill_1 FILLER_19_788 ();
 sg13g2_fill_2 FILLER_19_807 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_410 ();
 sg13g2_fill_1 FILLER_20_412 ();
 sg13g2_decap_4 FILLER_20_426 ();
 sg13g2_fill_2 FILLER_20_444 ();
 sg13g2_fill_1 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_452 ();
 sg13g2_fill_2 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_508 ();
 sg13g2_fill_1 FILLER_20_510 ();
 sg13g2_fill_1 FILLER_20_533 ();
 sg13g2_fill_2 FILLER_20_553 ();
 sg13g2_fill_2 FILLER_20_632 ();
 sg13g2_fill_1 FILLER_20_634 ();
 sg13g2_fill_2 FILLER_20_661 ();
 sg13g2_fill_2 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_756 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_384 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_fill_1 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_440 ();
 sg13g2_fill_1 FILLER_21_463 ();
 sg13g2_fill_2 FILLER_21_512 ();
 sg13g2_fill_1 FILLER_21_543 ();
 sg13g2_fill_1 FILLER_21_558 ();
 sg13g2_fill_2 FILLER_21_611 ();
 sg13g2_fill_2 FILLER_21_647 ();
 sg13g2_fill_1 FILLER_21_649 ();
 sg13g2_fill_2 FILLER_21_726 ();
 sg13g2_fill_1 FILLER_21_808 ();
 sg13g2_fill_1 FILLER_21_833 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_fill_2 FILLER_22_452 ();
 sg13g2_fill_1 FILLER_22_454 ();
 sg13g2_fill_1 FILLER_22_500 ();
 sg13g2_fill_1 FILLER_22_526 ();
 sg13g2_fill_1 FILLER_22_563 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_fill_1 FILLER_22_642 ();
 sg13g2_fill_2 FILLER_22_661 ();
 sg13g2_fill_2 FILLER_22_677 ();
 sg13g2_fill_2 FILLER_22_715 ();
 sg13g2_fill_1 FILLER_22_717 ();
 sg13g2_fill_2 FILLER_22_734 ();
 sg13g2_fill_2 FILLER_22_769 ();
 sg13g2_fill_1 FILLER_22_771 ();
 sg13g2_fill_2 FILLER_22_822 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_fill_1 FILLER_23_27 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_449 ();
 sg13g2_fill_2 FILLER_23_522 ();
 sg13g2_fill_2 FILLER_23_536 ();
 sg13g2_fill_2 FILLER_23_543 ();
 sg13g2_fill_1 FILLER_23_545 ();
 sg13g2_fill_2 FILLER_23_556 ();
 sg13g2_fill_2 FILLER_23_566 ();
 sg13g2_fill_1 FILLER_23_617 ();
 sg13g2_fill_2 FILLER_23_646 ();
 sg13g2_fill_1 FILLER_23_667 ();
 sg13g2_fill_1 FILLER_23_789 ();
 sg13g2_fill_2 FILLER_23_825 ();
 sg13g2_fill_1 FILLER_23_846 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_414 ();
 sg13g2_fill_1 FILLER_24_416 ();
 sg13g2_fill_2 FILLER_24_438 ();
 sg13g2_fill_2 FILLER_24_452 ();
 sg13g2_fill_2 FILLER_24_467 ();
 sg13g2_fill_1 FILLER_24_469 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_decap_4 FILLER_24_523 ();
 sg13g2_fill_2 FILLER_24_527 ();
 sg13g2_fill_2 FILLER_24_591 ();
 sg13g2_fill_1 FILLER_24_620 ();
 sg13g2_fill_2 FILLER_24_634 ();
 sg13g2_fill_2 FILLER_24_683 ();
 sg13g2_fill_1 FILLER_24_685 ();
 sg13g2_fill_2 FILLER_24_696 ();
 sg13g2_fill_2 FILLER_24_703 ();
 sg13g2_fill_1 FILLER_24_719 ();
 sg13g2_fill_2 FILLER_24_764 ();
 sg13g2_fill_1 FILLER_24_766 ();
 sg13g2_fill_2 FILLER_24_784 ();
 sg13g2_fill_1 FILLER_24_799 ();
 sg13g2_fill_1 FILLER_24_818 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_465 ();
 sg13g2_fill_2 FILLER_25_626 ();
 sg13g2_fill_1 FILLER_25_628 ();
 sg13g2_fill_2 FILLER_25_668 ();
 sg13g2_fill_1 FILLER_25_670 ();
 sg13g2_fill_2 FILLER_25_692 ();
 sg13g2_fill_2 FILLER_25_823 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_391 ();
 sg13g2_fill_2 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_26_448 ();
 sg13g2_fill_1 FILLER_26_450 ();
 sg13g2_decap_4 FILLER_26_512 ();
 sg13g2_fill_2 FILLER_26_555 ();
 sg13g2_fill_1 FILLER_26_601 ();
 sg13g2_fill_1 FILLER_26_640 ();
 sg13g2_fill_2 FILLER_26_649 ();
 sg13g2_fill_1 FILLER_26_651 ();
 sg13g2_fill_2 FILLER_26_683 ();
 sg13g2_fill_1 FILLER_26_717 ();
 sg13g2_fill_2 FILLER_26_787 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_406 ();
 sg13g2_fill_2 FILLER_27_471 ();
 sg13g2_fill_1 FILLER_27_543 ();
 sg13g2_fill_2 FILLER_27_573 ();
 sg13g2_fill_1 FILLER_27_602 ();
 sg13g2_fill_1 FILLER_27_645 ();
 sg13g2_fill_2 FILLER_27_679 ();
 sg13g2_fill_2 FILLER_27_709 ();
 sg13g2_fill_2 FILLER_27_721 ();
 sg13g2_fill_1 FILLER_27_783 ();
 sg13g2_fill_2 FILLER_27_859 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_259 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_1 FILLER_28_452 ();
 sg13g2_fill_1 FILLER_28_486 ();
 sg13g2_fill_2 FILLER_28_515 ();
 sg13g2_fill_2 FILLER_28_591 ();
 sg13g2_fill_1 FILLER_28_593 ();
 sg13g2_fill_2 FILLER_28_667 ();
 sg13g2_fill_1 FILLER_28_706 ();
 sg13g2_fill_1 FILLER_28_735 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_fill_2 FILLER_28_781 ();
 sg13g2_fill_2 FILLER_28_791 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_434 ();
 sg13g2_fill_2 FILLER_29_571 ();
 sg13g2_fill_2 FILLER_29_601 ();
 sg13g2_fill_1 FILLER_29_603 ();
 sg13g2_fill_1 FILLER_29_647 ();
 sg13g2_fill_2 FILLER_29_735 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_2 FILLER_30_437 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_fill_2 FILLER_30_471 ();
 sg13g2_fill_2 FILLER_30_489 ();
 sg13g2_fill_2 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_573 ();
 sg13g2_fill_2 FILLER_30_644 ();
 sg13g2_fill_1 FILLER_30_719 ();
 sg13g2_fill_2 FILLER_30_800 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_414 ();
 sg13g2_fill_1 FILLER_31_433 ();
 sg13g2_fill_1 FILLER_31_475 ();
 sg13g2_fill_2 FILLER_31_555 ();
 sg13g2_fill_1 FILLER_31_684 ();
 sg13g2_fill_2 FILLER_31_806 ();
 sg13g2_fill_1 FILLER_31_813 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_fill_1 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_450 ();
 sg13g2_fill_1 FILLER_32_471 ();
 sg13g2_fill_2 FILLER_32_627 ();
 sg13g2_fill_1 FILLER_32_645 ();
 sg13g2_fill_2 FILLER_32_779 ();
 sg13g2_fill_1 FILLER_32_798 ();
 sg13g2_fill_1 FILLER_32_812 ();
 sg13g2_fill_2 FILLER_32_826 ();
 sg13g2_fill_1 FILLER_32_842 ();
 sg13g2_fill_1 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_491 ();
 sg13g2_fill_2 FILLER_33_512 ();
 sg13g2_fill_2 FILLER_33_597 ();
 sg13g2_fill_2 FILLER_33_681 ();
 sg13g2_fill_1 FILLER_33_737 ();
 sg13g2_fill_2 FILLER_33_775 ();
 sg13g2_fill_1 FILLER_33_777 ();
 sg13g2_fill_2 FILLER_33_800 ();
 sg13g2_fill_1 FILLER_33_833 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_546 ();
 sg13g2_fill_1 FILLER_34_574 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_fill_1 FILLER_34_617 ();
 sg13g2_fill_1 FILLER_34_659 ();
 sg13g2_fill_2 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_787 ();
 sg13g2_fill_1 FILLER_34_818 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_491 ();
 sg13g2_fill_1 FILLER_35_493 ();
 sg13g2_fill_2 FILLER_35_602 ();
 sg13g2_fill_2 FILLER_35_693 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_432 ();
 sg13g2_fill_2 FILLER_36_470 ();
 sg13g2_fill_1 FILLER_36_490 ();
 sg13g2_fill_1 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_635 ();
 sg13g2_fill_2 FILLER_36_664 ();
 sg13g2_fill_1 FILLER_36_713 ();
 sg13g2_fill_1 FILLER_36_723 ();
 sg13g2_fill_2 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_767 ();
 sg13g2_fill_1 FILLER_36_808 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_fill_2 FILLER_37_440 ();
 sg13g2_fill_1 FILLER_37_442 ();
 sg13g2_fill_2 FILLER_37_519 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_1 FILLER_37_608 ();
 sg13g2_fill_1 FILLER_37_768 ();
 sg13g2_fill_1 FILLER_37_823 ();
 sg13g2_fill_2 FILLER_37_838 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_61 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_417 ();
 sg13g2_fill_2 FILLER_38_432 ();
 sg13g2_fill_1 FILLER_38_434 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_fill_2 FILLER_38_467 ();
 sg13g2_fill_1 FILLER_38_469 ();
 sg13g2_fill_2 FILLER_38_568 ();
 sg13g2_fill_1 FILLER_38_583 ();
 sg13g2_fill_2 FILLER_38_633 ();
 sg13g2_fill_1 FILLER_38_716 ();
 sg13g2_fill_2 FILLER_38_762 ();
 sg13g2_fill_1 FILLER_38_801 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_79 ();
 sg13g2_fill_2 FILLER_39_96 ();
 sg13g2_fill_1 FILLER_39_229 ();
 sg13g2_fill_2 FILLER_39_251 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_1 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_378 ();
 sg13g2_fill_2 FILLER_39_443 ();
 sg13g2_fill_1 FILLER_39_445 ();
 sg13g2_fill_1 FILLER_39_472 ();
 sg13g2_fill_2 FILLER_39_487 ();
 sg13g2_fill_2 FILLER_39_498 ();
 sg13g2_fill_1 FILLER_39_518 ();
 sg13g2_fill_2 FILLER_39_542 ();
 sg13g2_fill_1 FILLER_39_544 ();
 sg13g2_fill_1 FILLER_39_568 ();
 sg13g2_fill_1 FILLER_39_579 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_fill_2 FILLER_39_808 ();
 sg13g2_decap_4 FILLER_39_814 ();
 sg13g2_fill_2 FILLER_39_818 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_fill_2 FILLER_39_830 ();
 sg13g2_fill_2 FILLER_39_850 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_113 ();
 sg13g2_fill_1 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_221 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_429 ();
 sg13g2_fill_1 FILLER_40_431 ();
 sg13g2_fill_1 FILLER_40_464 ();
 sg13g2_fill_2 FILLER_40_475 ();
 sg13g2_fill_1 FILLER_40_477 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_489 ();
 sg13g2_fill_2 FILLER_40_516 ();
 sg13g2_fill_2 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_591 ();
 sg13g2_fill_2 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_696 ();
 sg13g2_decap_4 FILLER_40_795 ();
 sg13g2_fill_1 FILLER_40_799 ();
 sg13g2_decap_4 FILLER_40_806 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_fill_1 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_fill_2 FILLER_40_859 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_fill_2 FILLER_41_29 ();
 sg13g2_fill_2 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_107 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_187 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_fill_2 FILLER_41_229 ();
 sg13g2_fill_1 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_243 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_fill_2 FILLER_41_411 ();
 sg13g2_fill_1 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_494 ();
 sg13g2_fill_1 FILLER_41_547 ();
 sg13g2_fill_2 FILLER_41_655 ();
 sg13g2_fill_1 FILLER_41_700 ();
 sg13g2_fill_2 FILLER_41_735 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_2 FILLER_42_74 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_fill_1 FILLER_42_176 ();
 sg13g2_fill_2 FILLER_42_200 ();
 sg13g2_fill_2 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_249 ();
 sg13g2_fill_1 FILLER_42_269 ();
 sg13g2_fill_2 FILLER_42_346 ();
 sg13g2_fill_2 FILLER_42_380 ();
 sg13g2_decap_4 FILLER_42_419 ();
 sg13g2_fill_1 FILLER_42_442 ();
 sg13g2_fill_2 FILLER_42_487 ();
 sg13g2_fill_2 FILLER_42_526 ();
 sg13g2_fill_1 FILLER_42_528 ();
 sg13g2_fill_1 FILLER_42_573 ();
 sg13g2_fill_2 FILLER_42_594 ();
 sg13g2_fill_1 FILLER_42_613 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_fill_1 FILLER_42_777 ();
 sg13g2_fill_2 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_849 ();
 sg13g2_decap_4 FILLER_42_856 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_1 FILLER_43_62 ();
 sg13g2_fill_2 FILLER_43_113 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_236 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_fill_1 FILLER_43_482 ();
 sg13g2_fill_2 FILLER_43_534 ();
 sg13g2_fill_1 FILLER_43_555 ();
 sg13g2_fill_2 FILLER_43_667 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_744 ();
 sg13g2_fill_1 FILLER_43_773 ();
 sg13g2_fill_2 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_fill_2 FILLER_44_55 ();
 sg13g2_fill_1 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_215 ();
 sg13g2_fill_1 FILLER_44_275 ();
 sg13g2_fill_2 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_384 ();
 sg13g2_fill_1 FILLER_44_419 ();
 sg13g2_fill_1 FILLER_44_476 ();
 sg13g2_fill_1 FILLER_44_487 ();
 sg13g2_fill_1 FILLER_44_498 ();
 sg13g2_fill_1 FILLER_44_527 ();
 sg13g2_fill_1 FILLER_44_573 ();
 sg13g2_fill_2 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_857 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_1 FILLER_45_135 ();
 sg13g2_fill_2 FILLER_45_171 ();
 sg13g2_fill_2 FILLER_45_191 ();
 sg13g2_fill_2 FILLER_45_241 ();
 sg13g2_fill_2 FILLER_45_284 ();
 sg13g2_fill_2 FILLER_45_412 ();
 sg13g2_fill_1 FILLER_45_414 ();
 sg13g2_fill_1 FILLER_45_425 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_fill_1 FILLER_45_545 ();
 sg13g2_fill_1 FILLER_45_733 ();
 sg13g2_fill_2 FILLER_45_761 ();
 sg13g2_fill_1 FILLER_45_763 ();
 sg13g2_fill_2 FILLER_45_804 ();
 sg13g2_fill_1 FILLER_45_820 ();
 sg13g2_decap_4 FILLER_45_848 ();
 sg13g2_fill_1 FILLER_45_852 ();
 sg13g2_fill_1 FILLER_46_41 ();
 sg13g2_fill_1 FILLER_46_106 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_2 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_fill_2 FILLER_46_299 ();
 sg13g2_fill_2 FILLER_46_331 ();
 sg13g2_fill_1 FILLER_46_421 ();
 sg13g2_fill_2 FILLER_46_431 ();
 sg13g2_fill_1 FILLER_46_433 ();
 sg13g2_fill_2 FILLER_46_505 ();
 sg13g2_fill_1 FILLER_46_507 ();
 sg13g2_fill_1 FILLER_46_527 ();
 sg13g2_fill_2 FILLER_46_644 ();
 sg13g2_fill_1 FILLER_46_674 ();
 sg13g2_fill_2 FILLER_46_693 ();
 sg13g2_fill_2 FILLER_46_775 ();
 sg13g2_fill_1 FILLER_46_777 ();
 sg13g2_fill_2 FILLER_46_791 ();
 sg13g2_fill_2 FILLER_46_806 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_47 ();
 sg13g2_fill_1 FILLER_47_53 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_fill_1 FILLER_47_187 ();
 sg13g2_fill_1 FILLER_47_303 ();
 sg13g2_fill_2 FILLER_47_392 ();
 sg13g2_fill_2 FILLER_47_446 ();
 sg13g2_fill_1 FILLER_47_448 ();
 sg13g2_fill_2 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_628 ();
 sg13g2_fill_1 FILLER_47_719 ();
 sg13g2_fill_1 FILLER_47_734 ();
 sg13g2_decap_4 FILLER_47_761 ();
 sg13g2_fill_1 FILLER_47_765 ();
 sg13g2_fill_1 FILLER_47_802 ();
 sg13g2_fill_2 FILLER_47_830 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_fill_2 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_336 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_415 ();
 sg13g2_fill_2 FILLER_48_432 ();
 sg13g2_fill_1 FILLER_48_434 ();
 sg13g2_fill_1 FILLER_48_463 ();
 sg13g2_fill_1 FILLER_48_508 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_fill_1 FILLER_48_662 ();
 sg13g2_fill_1 FILLER_48_711 ();
 sg13g2_fill_2 FILLER_48_737 ();
 sg13g2_fill_1 FILLER_48_739 ();
 sg13g2_fill_2 FILLER_48_777 ();
 sg13g2_fill_1 FILLER_48_796 ();
 sg13g2_fill_1 FILLER_49_27 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_fill_1 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_346 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_376 ();
 sg13g2_fill_1 FILLER_49_405 ();
 sg13g2_fill_1 FILLER_49_561 ();
 sg13g2_fill_1 FILLER_49_630 ();
 sg13g2_fill_2 FILLER_49_657 ();
 sg13g2_decap_4 FILLER_49_744 ();
 sg13g2_fill_1 FILLER_49_762 ();
 sg13g2_fill_2 FILLER_49_781 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_1 FILLER_50_27 ();
 sg13g2_fill_2 FILLER_50_64 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_fill_2 FILLER_50_350 ();
 sg13g2_fill_1 FILLER_50_352 ();
 sg13g2_fill_2 FILLER_50_362 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_fill_2 FILLER_50_400 ();
 sg13g2_fill_1 FILLER_50_402 ();
 sg13g2_decap_4 FILLER_50_435 ();
 sg13g2_fill_2 FILLER_50_603 ();
 sg13g2_fill_2 FILLER_50_635 ();
 sg13g2_fill_2 FILLER_50_684 ();
 sg13g2_fill_1 FILLER_50_729 ();
 sg13g2_decap_4 FILLER_50_754 ();
 sg13g2_fill_1 FILLER_50_758 ();
 sg13g2_fill_1 FILLER_50_775 ();
 sg13g2_fill_2 FILLER_50_781 ();
 sg13g2_fill_2 FILLER_50_805 ();
 sg13g2_fill_1 FILLER_50_807 ();
 sg13g2_fill_1 FILLER_50_831 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_29 ();
 sg13g2_fill_2 FILLER_51_59 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_222 ();
 sg13g2_fill_2 FILLER_51_327 ();
 sg13g2_fill_1 FILLER_51_329 ();
 sg13g2_fill_1 FILLER_51_339 ();
 sg13g2_fill_2 FILLER_51_376 ();
 sg13g2_fill_2 FILLER_51_400 ();
 sg13g2_fill_1 FILLER_51_507 ();
 sg13g2_fill_2 FILLER_51_540 ();
 sg13g2_fill_1 FILLER_51_632 ();
 sg13g2_fill_2 FILLER_51_679 ();
 sg13g2_fill_2 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_759 ();
 sg13g2_fill_2 FILLER_51_783 ();
 sg13g2_fill_1 FILLER_51_785 ();
 sg13g2_fill_2 FILLER_51_796 ();
 sg13g2_fill_1 FILLER_51_807 ();
 sg13g2_fill_2 FILLER_51_851 ();
 sg13g2_fill_2 FILLER_52_27 ();
 sg13g2_fill_1 FILLER_52_71 ();
 sg13g2_fill_2 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_318 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_fill_2 FILLER_52_376 ();
 sg13g2_fill_1 FILLER_52_378 ();
 sg13g2_fill_2 FILLER_52_388 ();
 sg13g2_fill_2 FILLER_52_404 ();
 sg13g2_fill_2 FILLER_52_412 ();
 sg13g2_fill_1 FILLER_52_445 ();
 sg13g2_fill_2 FILLER_52_456 ();
 sg13g2_fill_1 FILLER_52_458 ();
 sg13g2_fill_1 FILLER_52_486 ();
 sg13g2_fill_2 FILLER_52_521 ();
 sg13g2_fill_2 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_677 ();
 sg13g2_fill_2 FILLER_52_683 ();
 sg13g2_fill_1 FILLER_52_685 ();
 sg13g2_fill_1 FILLER_52_701 ();
 sg13g2_fill_2 FILLER_52_735 ();
 sg13g2_fill_2 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_decap_4 FILLER_52_783 ();
 sg13g2_fill_1 FILLER_52_787 ();
 sg13g2_fill_1 FILLER_52_811 ();
 sg13g2_fill_2 FILLER_52_831 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_fill_2 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_139 ();
 sg13g2_decap_4 FILLER_53_423 ();
 sg13g2_fill_2 FILLER_53_546 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_fill_2 FILLER_53_581 ();
 sg13g2_fill_2 FILLER_53_627 ();
 sg13g2_fill_2 FILLER_53_680 ();
 sg13g2_fill_2 FILLER_53_696 ();
 sg13g2_fill_1 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_742 ();
 sg13g2_fill_2 FILLER_53_759 ();
 sg13g2_fill_1 FILLER_53_761 ();
 sg13g2_fill_1 FILLER_53_791 ();
 sg13g2_fill_2 FILLER_53_808 ();
 sg13g2_fill_1 FILLER_53_842 ();
 sg13g2_fill_1 FILLER_54_146 ();
 sg13g2_fill_1 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_fill_2 FILLER_54_388 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_fill_1 FILLER_54_397 ();
 sg13g2_fill_2 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_452 ();
 sg13g2_fill_1 FILLER_54_476 ();
 sg13g2_fill_1 FILLER_54_506 ();
 sg13g2_fill_1 FILLER_54_513 ();
 sg13g2_decap_4 FILLER_54_533 ();
 sg13g2_fill_1 FILLER_54_550 ();
 sg13g2_fill_2 FILLER_54_653 ();
 sg13g2_fill_1 FILLER_54_655 ();
 sg13g2_fill_2 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_714 ();
 sg13g2_fill_2 FILLER_54_721 ();
 sg13g2_fill_1 FILLER_54_723 ();
 sg13g2_fill_2 FILLER_54_732 ();
 sg13g2_fill_1 FILLER_54_734 ();
 sg13g2_decap_4 FILLER_54_760 ();
 sg13g2_fill_2 FILLER_54_784 ();
 sg13g2_fill_1 FILLER_54_786 ();
 sg13g2_fill_2 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_303 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_fill_2 FILLER_55_384 ();
 sg13g2_fill_2 FILLER_55_405 ();
 sg13g2_fill_2 FILLER_55_444 ();
 sg13g2_fill_2 FILLER_55_484 ();
 sg13g2_fill_2 FILLER_55_514 ();
 sg13g2_fill_2 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_714 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_decap_8 FILLER_55_752 ();
 sg13g2_decap_8 FILLER_55_759 ();
 sg13g2_decap_4 FILLER_55_766 ();
 sg13g2_fill_2 FILLER_55_774 ();
 sg13g2_fill_1 FILLER_55_785 ();
 sg13g2_fill_1 FILLER_55_791 ();
 sg13g2_fill_1 FILLER_55_800 ();
 sg13g2_fill_1 FILLER_55_806 ();
 sg13g2_fill_2 FILLER_56_87 ();
 sg13g2_fill_2 FILLER_56_116 ();
 sg13g2_fill_1 FILLER_56_131 ();
 sg13g2_fill_1 FILLER_56_332 ();
 sg13g2_fill_1 FILLER_56_383 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_1 FILLER_56_431 ();
 sg13g2_fill_2 FILLER_56_445 ();
 sg13g2_fill_1 FILLER_56_476 ();
 sg13g2_fill_1 FILLER_56_518 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_fill_2 FILLER_56_618 ();
 sg13g2_fill_1 FILLER_56_620 ();
 sg13g2_fill_1 FILLER_56_640 ();
 sg13g2_fill_1 FILLER_56_659 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_fill_2 FILLER_56_685 ();
 sg13g2_fill_1 FILLER_56_687 ();
 sg13g2_fill_2 FILLER_56_711 ();
 sg13g2_fill_1 FILLER_56_713 ();
 sg13g2_fill_1 FILLER_56_720 ();
 sg13g2_fill_2 FILLER_56_733 ();
 sg13g2_fill_2 FILLER_56_759 ();
 sg13g2_fill_2 FILLER_56_800 ();
 sg13g2_fill_1 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_808 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_373 ();
 sg13g2_fill_2 FILLER_57_411 ();
 sg13g2_fill_1 FILLER_57_413 ();
 sg13g2_fill_1 FILLER_57_527 ();
 sg13g2_fill_1 FILLER_57_575 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_fill_1 FILLER_57_624 ();
 sg13g2_fill_2 FILLER_57_664 ();
 sg13g2_fill_2 FILLER_57_696 ();
 sg13g2_decap_4 FILLER_57_706 ();
 sg13g2_fill_2 FILLER_57_788 ();
 sg13g2_fill_2 FILLER_57_803 ();
 sg13g2_decap_4 FILLER_57_858 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_fill_2 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_155 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_2 FILLER_58_303 ();
 sg13g2_fill_1 FILLER_58_350 ();
 sg13g2_fill_2 FILLER_58_374 ();
 sg13g2_fill_1 FILLER_58_376 ();
 sg13g2_fill_1 FILLER_58_398 ();
 sg13g2_fill_1 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_500 ();
 sg13g2_fill_1 FILLER_58_535 ();
 sg13g2_fill_2 FILLER_58_545 ();
 sg13g2_fill_2 FILLER_58_607 ();
 sg13g2_fill_1 FILLER_58_609 ();
 sg13g2_fill_2 FILLER_58_632 ();
 sg13g2_fill_1 FILLER_58_634 ();
 sg13g2_fill_1 FILLER_58_676 ();
 sg13g2_fill_1 FILLER_58_710 ();
 sg13g2_decap_4 FILLER_58_760 ();
 sg13g2_fill_1 FILLER_58_764 ();
 sg13g2_fill_2 FILLER_58_769 ();
 sg13g2_decap_4 FILLER_58_775 ();
 sg13g2_fill_2 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_804 ();
 sg13g2_fill_2 FILLER_58_812 ();
 sg13g2_fill_2 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_fill_1 FILLER_59_27 ();
 sg13g2_fill_2 FILLER_59_43 ();
 sg13g2_fill_1 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_fill_2 FILLER_59_189 ();
 sg13g2_fill_2 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_fill_1 FILLER_59_434 ();
 sg13g2_fill_1 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_648 ();
 sg13g2_fill_1 FILLER_59_662 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_fill_1 FILLER_59_702 ();
 sg13g2_decap_4 FILLER_59_725 ();
 sg13g2_fill_2 FILLER_59_729 ();
 sg13g2_decap_4 FILLER_59_735 ();
 sg13g2_fill_1 FILLER_59_745 ();
 sg13g2_decap_4 FILLER_59_758 ();
 sg13g2_fill_2 FILLER_59_797 ();
 sg13g2_fill_2 FILLER_59_815 ();
 sg13g2_fill_1 FILLER_59_833 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_1 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_124 ();
 sg13g2_fill_2 FILLER_60_205 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_248 ();
 sg13g2_fill_2 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_2 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_662 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_fill_2 FILLER_60_682 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_fill_1 FILLER_60_690 ();
 sg13g2_fill_1 FILLER_60_712 ();
 sg13g2_decap_4 FILLER_60_731 ();
 sg13g2_fill_2 FILLER_60_735 ();
 sg13g2_fill_2 FILLER_60_750 ();
 sg13g2_fill_2 FILLER_60_760 ();
 sg13g2_fill_1 FILLER_60_762 ();
 sg13g2_fill_1 FILLER_60_782 ();
 sg13g2_fill_2 FILLER_60_807 ();
 sg13g2_fill_1 FILLER_60_823 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_46 ();
 sg13g2_fill_1 FILLER_61_48 ();
 sg13g2_fill_2 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_251 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_331 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_381 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_61_431 ();
 sg13g2_fill_2 FILLER_61_472 ();
 sg13g2_fill_1 FILLER_61_545 ();
 sg13g2_fill_2 FILLER_61_646 ();
 sg13g2_fill_1 FILLER_61_648 ();
 sg13g2_fill_2 FILLER_61_663 ();
 sg13g2_fill_1 FILLER_61_683 ();
 sg13g2_fill_1 FILLER_61_705 ();
 sg13g2_fill_1 FILLER_61_734 ();
 sg13g2_fill_2 FILLER_61_741 ();
 sg13g2_fill_1 FILLER_61_743 ();
 sg13g2_decap_8 FILLER_61_756 ();
 sg13g2_fill_2 FILLER_61_772 ();
 sg13g2_fill_1 FILLER_61_774 ();
 sg13g2_fill_2 FILLER_61_829 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_fill_1 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_293 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_398 ();
 sg13g2_fill_2 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_413 ();
 sg13g2_fill_2 FILLER_62_448 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_fill_1 FILLER_62_543 ();
 sg13g2_fill_1 FILLER_62_576 ();
 sg13g2_fill_2 FILLER_62_645 ();
 sg13g2_fill_2 FILLER_62_670 ();
 sg13g2_fill_2 FILLER_62_680 ();
 sg13g2_fill_2 FILLER_62_703 ();
 sg13g2_fill_1 FILLER_62_705 ();
 sg13g2_fill_2 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_756 ();
 sg13g2_fill_1 FILLER_62_758 ();
 sg13g2_fill_1 FILLER_62_767 ();
 sg13g2_fill_1 FILLER_62_784 ();
 sg13g2_fill_1 FILLER_62_790 ();
 sg13g2_fill_1 FILLER_62_804 ();
 sg13g2_fill_1 FILLER_62_814 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_52 ();
 sg13g2_fill_2 FILLER_63_130 ();
 sg13g2_fill_2 FILLER_63_246 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_361 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_fill_1 FILLER_63_428 ();
 sg13g2_fill_2 FILLER_63_597 ();
 sg13g2_fill_2 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_fill_2 FILLER_63_669 ();
 sg13g2_fill_1 FILLER_63_671 ();
 sg13g2_fill_2 FILLER_63_685 ();
 sg13g2_fill_2 FILLER_63_715 ();
 sg13g2_fill_2 FILLER_63_739 ();
 sg13g2_fill_1 FILLER_63_762 ();
 sg13g2_decap_4 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_775 ();
 sg13g2_fill_1 FILLER_63_781 ();
 sg13g2_fill_2 FILLER_63_786 ();
 sg13g2_fill_2 FILLER_63_813 ();
 sg13g2_fill_1 FILLER_63_815 ();
 sg13g2_fill_1 FILLER_63_820 ();
 sg13g2_fill_1 FILLER_63_843 ();
 sg13g2_fill_2 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_143 ();
 sg13g2_fill_2 FILLER_64_169 ();
 sg13g2_fill_1 FILLER_64_207 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_fill_1 FILLER_64_330 ();
 sg13g2_fill_2 FILLER_64_440 ();
 sg13g2_fill_1 FILLER_64_481 ();
 sg13g2_fill_1 FILLER_64_640 ();
 sg13g2_fill_2 FILLER_64_646 ();
 sg13g2_fill_2 FILLER_64_680 ();
 sg13g2_fill_1 FILLER_64_709 ();
 sg13g2_fill_2 FILLER_64_725 ();
 sg13g2_fill_2 FILLER_64_757 ();
 sg13g2_fill_1 FILLER_64_759 ();
 sg13g2_fill_2 FILLER_64_785 ();
 sg13g2_fill_1 FILLER_64_787 ();
 sg13g2_fill_2 FILLER_64_830 ();
 sg13g2_fill_1 FILLER_64_832 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_245 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_fill_2 FILLER_65_421 ();
 sg13g2_fill_2 FILLER_65_452 ();
 sg13g2_fill_1 FILLER_65_562 ();
 sg13g2_fill_1 FILLER_65_579 ();
 sg13g2_fill_1 FILLER_65_670 ();
 sg13g2_fill_1 FILLER_65_710 ();
 sg13g2_fill_1 FILLER_65_720 ();
 sg13g2_fill_2 FILLER_65_730 ();
 sg13g2_fill_1 FILLER_65_732 ();
 sg13g2_decap_8 FILLER_65_750 ();
 sg13g2_decap_4 FILLER_65_757 ();
 sg13g2_fill_2 FILLER_65_786 ();
 sg13g2_fill_1 FILLER_65_788 ();
 sg13g2_fill_1 FILLER_65_806 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_71 ();
 sg13g2_fill_2 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_121 ();
 sg13g2_fill_2 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_443 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_480 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_630 ();
 sg13g2_fill_2 FILLER_66_725 ();
 sg13g2_fill_1 FILLER_66_735 ();
 sg13g2_decap_4 FILLER_66_749 ();
 sg13g2_fill_1 FILLER_66_753 ();
 sg13g2_fill_1 FILLER_66_762 ();
 sg13g2_decap_4 FILLER_66_783 ();
 sg13g2_fill_1 FILLER_66_787 ();
 sg13g2_fill_2 FILLER_66_802 ();
 sg13g2_fill_1 FILLER_66_804 ();
 sg13g2_fill_1 FILLER_66_829 ();
 sg13g2_decap_4 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_2 FILLER_67_45 ();
 sg13g2_fill_2 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_241 ();
 sg13g2_fill_2 FILLER_67_261 ();
 sg13g2_fill_1 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_359 ();
 sg13g2_fill_2 FILLER_67_485 ();
 sg13g2_fill_1 FILLER_67_546 ();
 sg13g2_fill_2 FILLER_67_691 ();
 sg13g2_fill_1 FILLER_67_693 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_fill_2 FILLER_67_763 ();
 sg13g2_fill_2 FILLER_67_772 ();
 sg13g2_fill_2 FILLER_67_794 ();
 sg13g2_decap_4 FILLER_67_858 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_78 ();
 sg13g2_fill_1 FILLER_68_236 ();
 sg13g2_fill_2 FILLER_68_308 ();
 sg13g2_fill_2 FILLER_68_389 ();
 sg13g2_fill_1 FILLER_68_465 ();
 sg13g2_fill_1 FILLER_68_524 ();
 sg13g2_fill_1 FILLER_68_626 ();
 sg13g2_fill_1 FILLER_68_651 ();
 sg13g2_fill_1 FILLER_68_682 ();
 sg13g2_decap_8 FILLER_68_693 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_fill_1 FILLER_68_771 ();
 sg13g2_fill_2 FILLER_68_802 ();
 sg13g2_fill_1 FILLER_68_804 ();
 sg13g2_fill_1 FILLER_68_826 ();
 sg13g2_fill_1 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_2 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_167 ();
 sg13g2_fill_1 FILLER_69_228 ();
 sg13g2_fill_2 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_fill_1 FILLER_69_345 ();
 sg13g2_fill_1 FILLER_69_428 ();
 sg13g2_fill_1 FILLER_69_453 ();
 sg13g2_fill_2 FILLER_69_607 ();
 sg13g2_fill_2 FILLER_69_671 ();
 sg13g2_fill_1 FILLER_69_673 ();
 sg13g2_fill_1 FILLER_69_682 ();
 sg13g2_fill_2 FILLER_69_693 ();
 sg13g2_fill_1 FILLER_69_752 ();
 sg13g2_decap_8 FILLER_69_757 ();
 sg13g2_fill_2 FILLER_69_764 ();
 sg13g2_fill_1 FILLER_69_766 ();
 sg13g2_fill_2 FILLER_69_776 ();
 sg13g2_fill_1 FILLER_70_36 ();
 sg13g2_fill_2 FILLER_70_64 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_239 ();
 sg13g2_fill_2 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_374 ();
 sg13g2_fill_1 FILLER_70_432 ();
 sg13g2_fill_1 FILLER_70_480 ();
 sg13g2_fill_1 FILLER_70_556 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_2 FILLER_70_672 ();
 sg13g2_decap_8 FILLER_70_679 ();
 sg13g2_decap_8 FILLER_70_686 ();
 sg13g2_fill_2 FILLER_70_693 ();
 sg13g2_fill_2 FILLER_70_711 ();
 sg13g2_fill_1 FILLER_70_713 ();
 sg13g2_fill_1 FILLER_70_749 ();
 sg13g2_decap_4 FILLER_70_849 ();
 sg13g2_fill_1 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_166 ();
 sg13g2_fill_2 FILLER_71_285 ();
 sg13g2_fill_2 FILLER_71_413 ();
 sg13g2_fill_2 FILLER_71_503 ();
 sg13g2_fill_2 FILLER_71_524 ();
 sg13g2_fill_2 FILLER_71_607 ();
 sg13g2_fill_2 FILLER_71_678 ();
 sg13g2_fill_1 FILLER_71_680 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_816 ();
 sg13g2_fill_2 FILLER_71_833 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_37 ();
 sg13g2_fill_1 FILLER_72_105 ();
 sg13g2_fill_1 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_286 ();
 sg13g2_fill_2 FILLER_72_344 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_fill_2 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_469 ();
 sg13g2_fill_1 FILLER_72_471 ();
 sg13g2_fill_2 FILLER_72_485 ();
 sg13g2_fill_1 FILLER_72_487 ();
 sg13g2_decap_4 FILLER_72_667 ();
 sg13g2_fill_1 FILLER_72_674 ();
 sg13g2_decap_8 FILLER_72_688 ();
 sg13g2_fill_2 FILLER_72_695 ();
 sg13g2_fill_2 FILLER_72_718 ();
 sg13g2_fill_1 FILLER_72_720 ();
 sg13g2_fill_2 FILLER_72_741 ();
 sg13g2_fill_1 FILLER_72_743 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_fill_2 FILLER_72_756 ();
 sg13g2_fill_1 FILLER_72_758 ();
 sg13g2_fill_1 FILLER_72_764 ();
 sg13g2_fill_2 FILLER_72_792 ();
 sg13g2_fill_1 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_833 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_76 ();
 sg13g2_fill_2 FILLER_73_225 ();
 sg13g2_fill_1 FILLER_73_255 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_fill_2 FILLER_73_515 ();
 sg13g2_fill_1 FILLER_73_517 ();
 sg13g2_fill_2 FILLER_73_570 ();
 sg13g2_fill_2 FILLER_73_589 ();
 sg13g2_fill_1 FILLER_73_722 ();
 sg13g2_fill_2 FILLER_73_744 ();
 sg13g2_fill_1 FILLER_73_746 ();
 sg13g2_fill_1 FILLER_73_779 ();
 sg13g2_fill_1 FILLER_73_829 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_26 ();
 sg13g2_fill_1 FILLER_74_46 ();
 sg13g2_fill_2 FILLER_74_225 ();
 sg13g2_fill_1 FILLER_74_339 ();
 sg13g2_fill_2 FILLER_74_363 ();
 sg13g2_fill_2 FILLER_74_392 ();
 sg13g2_fill_1 FILLER_74_434 ();
 sg13g2_fill_1 FILLER_74_518 ();
 sg13g2_fill_2 FILLER_74_570 ();
 sg13g2_decap_8 FILLER_74_585 ();
 sg13g2_decap_8 FILLER_74_592 ();
 sg13g2_decap_8 FILLER_74_599 ();
 sg13g2_decap_4 FILLER_74_606 ();
 sg13g2_fill_2 FILLER_74_610 ();
 sg13g2_fill_2 FILLER_74_615 ();
 sg13g2_fill_1 FILLER_74_709 ();
 sg13g2_decap_4 FILLER_74_756 ();
 sg13g2_fill_1 FILLER_74_760 ();
 sg13g2_fill_1 FILLER_74_806 ();
 sg13g2_fill_1 FILLER_74_829 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_4 ();
 sg13g2_fill_2 FILLER_75_43 ();
 sg13g2_fill_1 FILLER_75_45 ();
 sg13g2_fill_2 FILLER_75_50 ();
 sg13g2_fill_2 FILLER_75_80 ();
 sg13g2_fill_2 FILLER_75_109 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_313 ();
 sg13g2_fill_1 FILLER_75_362 ();
 sg13g2_fill_2 FILLER_75_450 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_fill_2 FILLER_75_536 ();
 sg13g2_decap_8 FILLER_75_574 ();
 sg13g2_decap_8 FILLER_75_581 ();
 sg13g2_decap_8 FILLER_75_588 ();
 sg13g2_decap_8 FILLER_75_595 ();
 sg13g2_decap_8 FILLER_75_602 ();
 sg13g2_decap_8 FILLER_75_609 ();
 sg13g2_decap_4 FILLER_75_616 ();
 sg13g2_fill_1 FILLER_75_620 ();
 sg13g2_decap_4 FILLER_75_725 ();
 sg13g2_fill_1 FILLER_75_729 ();
 sg13g2_fill_2 FILLER_75_792 ();
 sg13g2_fill_1 FILLER_75_794 ();
 sg13g2_fill_1 FILLER_75_808 ();
 sg13g2_fill_1 FILLER_75_831 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_7 ();
 sg13g2_fill_2 FILLER_76_11 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_fill_2 FILLER_76_47 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_2 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_438 ();
 sg13g2_fill_1 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_572 ();
 sg13g2_decap_8 FILLER_76_579 ();
 sg13g2_decap_8 FILLER_76_586 ();
 sg13g2_decap_8 FILLER_76_593 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_8 FILLER_76_607 ();
 sg13g2_decap_8 FILLER_76_614 ();
 sg13g2_decap_8 FILLER_76_621 ();
 sg13g2_decap_8 FILLER_76_628 ();
 sg13g2_fill_2 FILLER_76_635 ();
 sg13g2_decap_4 FILLER_76_646 ();
 sg13g2_fill_1 FILLER_76_650 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_fill_1 FILLER_76_666 ();
 sg13g2_fill_2 FILLER_76_679 ();
 sg13g2_fill_1 FILLER_76_681 ();
 sg13g2_fill_2 FILLER_76_692 ();
 sg13g2_decap_4 FILLER_76_721 ();
 sg13g2_fill_1 FILLER_76_725 ();
 sg13g2_fill_2 FILLER_76_792 ();
 sg13g2_decap_4 FILLER_76_821 ();
 sg13g2_fill_1 FILLER_76_825 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_18 ();
 sg13g2_fill_2 FILLER_77_40 ();
 sg13g2_fill_2 FILLER_77_217 ();
 sg13g2_fill_2 FILLER_77_317 ();
 sg13g2_fill_2 FILLER_77_390 ();
 sg13g2_fill_2 FILLER_77_478 ();
 sg13g2_fill_1 FILLER_77_480 ();
 sg13g2_decap_8 FILLER_77_569 ();
 sg13g2_decap_8 FILLER_77_576 ();
 sg13g2_decap_8 FILLER_77_583 ();
 sg13g2_decap_8 FILLER_77_590 ();
 sg13g2_decap_8 FILLER_77_597 ();
 sg13g2_decap_8 FILLER_77_604 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_fill_2 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_650 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_fill_2 FILLER_77_708 ();
 sg13g2_fill_1 FILLER_77_710 ();
 sg13g2_decap_8 FILLER_77_747 ();
 sg13g2_fill_1 FILLER_77_754 ();
 sg13g2_fill_2 FILLER_77_758 ();
 sg13g2_fill_1 FILLER_77_760 ();
 sg13g2_decap_4 FILLER_77_770 ();
 sg13g2_fill_1 FILLER_77_774 ();
 sg13g2_decap_4 FILLER_77_788 ();
 sg13g2_decap_8 FILLER_77_796 ();
 sg13g2_decap_4 FILLER_77_803 ();
 sg13g2_fill_2 FILLER_77_807 ();
 sg13g2_decap_8 FILLER_77_817 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_4 FILLER_77_831 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_58 ();
 sg13g2_fill_2 FILLER_78_110 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_559 ();
 sg13g2_decap_8 FILLER_78_566 ();
 sg13g2_decap_8 FILLER_78_573 ();
 sg13g2_decap_8 FILLER_78_580 ();
 sg13g2_decap_8 FILLER_78_587 ();
 sg13g2_decap_8 FILLER_78_594 ();
 sg13g2_decap_8 FILLER_78_601 ();
 sg13g2_decap_8 FILLER_78_608 ();
 sg13g2_decap_8 FILLER_78_615 ();
 sg13g2_decap_8 FILLER_78_622 ();
 sg13g2_decap_8 FILLER_78_629 ();
 sg13g2_decap_8 FILLER_78_636 ();
 sg13g2_decap_8 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_650 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_8 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_decap_8 FILLER_78_678 ();
 sg13g2_decap_8 FILLER_78_685 ();
 sg13g2_decap_8 FILLER_78_692 ();
 sg13g2_decap_8 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_decap_8 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_720 ();
 sg13g2_decap_8 FILLER_78_727 ();
 sg13g2_decap_8 FILLER_78_734 ();
 sg13g2_decap_8 FILLER_78_741 ();
 sg13g2_decap_8 FILLER_78_748 ();
 sg13g2_decap_8 FILLER_78_755 ();
 sg13g2_decap_8 FILLER_78_762 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_decap_8 FILLER_78_776 ();
 sg13g2_decap_8 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_790 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_decap_8 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_4 FILLER_78_832 ();
 sg13g2_fill_1 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_41 ();
 sg13g2_fill_1 FILLER_79_117 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_284 ();
 sg13g2_fill_1 FILLER_79_340 ();
 sg13g2_decap_8 FILLER_79_559 ();
 sg13g2_decap_8 FILLER_79_566 ();
 sg13g2_decap_8 FILLER_79_573 ();
 sg13g2_decap_8 FILLER_79_580 ();
 sg13g2_decap_8 FILLER_79_587 ();
 sg13g2_decap_8 FILLER_79_594 ();
 sg13g2_decap_8 FILLER_79_601 ();
 sg13g2_decap_8 FILLER_79_608 ();
 sg13g2_decap_8 FILLER_79_615 ();
 sg13g2_decap_8 FILLER_79_622 ();
 sg13g2_decap_8 FILLER_79_629 ();
 sg13g2_decap_8 FILLER_79_636 ();
 sg13g2_decap_8 FILLER_79_643 ();
 sg13g2_decap_8 FILLER_79_650 ();
 sg13g2_decap_8 FILLER_79_657 ();
 sg13g2_decap_8 FILLER_79_664 ();
 sg13g2_decap_8 FILLER_79_671 ();
 sg13g2_decap_8 FILLER_79_678 ();
 sg13g2_decap_8 FILLER_79_685 ();
 sg13g2_decap_8 FILLER_79_692 ();
 sg13g2_decap_8 FILLER_79_699 ();
 sg13g2_decap_8 FILLER_79_706 ();
 sg13g2_decap_8 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_720 ();
 sg13g2_decap_8 FILLER_79_727 ();
 sg13g2_decap_8 FILLER_79_734 ();
 sg13g2_decap_8 FILLER_79_741 ();
 sg13g2_decap_8 FILLER_79_748 ();
 sg13g2_decap_8 FILLER_79_755 ();
 sg13g2_decap_8 FILLER_79_762 ();
 sg13g2_decap_8 FILLER_79_769 ();
 sg13g2_decap_8 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_783 ();
 sg13g2_decap_8 FILLER_79_790 ();
 sg13g2_decap_8 FILLER_79_797 ();
 sg13g2_decap_8 FILLER_79_804 ();
 sg13g2_decap_8 FILLER_79_811 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_846 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_18 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_565 ();
 sg13g2_decap_8 FILLER_80_572 ();
 sg13g2_decap_8 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_586 ();
 sg13g2_decap_8 FILLER_80_593 ();
 sg13g2_decap_8 FILLER_80_600 ();
 sg13g2_decap_8 FILLER_80_607 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_628 ();
 sg13g2_decap_8 FILLER_80_635 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_decap_8 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_fill_2 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net25;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule
