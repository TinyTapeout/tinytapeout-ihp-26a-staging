module tt_um_wedgetail_tester (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire \mod_ro_128.fabric[0] ;
 wire \mod_ro_128.fabric[100] ;
 wire \mod_ro_128.fabric[101] ;
 wire \mod_ro_128.fabric[102] ;
 wire \mod_ro_128.fabric[103] ;
 wire \mod_ro_128.fabric[104] ;
 wire \mod_ro_128.fabric[105] ;
 wire \mod_ro_128.fabric[106] ;
 wire \mod_ro_128.fabric[107] ;
 wire \mod_ro_128.fabric[108] ;
 wire \mod_ro_128.fabric[109] ;
 wire \mod_ro_128.fabric[10] ;
 wire \mod_ro_128.fabric[110] ;
 wire \mod_ro_128.fabric[111] ;
 wire \mod_ro_128.fabric[112] ;
 wire \mod_ro_128.fabric[113] ;
 wire \mod_ro_128.fabric[114] ;
 wire \mod_ro_128.fabric[115] ;
 wire \mod_ro_128.fabric[116] ;
 wire \mod_ro_128.fabric[117] ;
 wire \mod_ro_128.fabric[118] ;
 wire \mod_ro_128.fabric[119] ;
 wire \mod_ro_128.fabric[11] ;
 wire \mod_ro_128.fabric[120] ;
 wire \mod_ro_128.fabric[121] ;
 wire \mod_ro_128.fabric[122] ;
 wire \mod_ro_128.fabric[123] ;
 wire \mod_ro_128.fabric[124] ;
 wire \mod_ro_128.fabric[125] ;
 wire \mod_ro_128.fabric[126] ;
 wire \mod_ro_128.fabric[127] ;
 wire \mod_ro_128.fabric[128] ;
 wire \mod_ro_128.fabric[12] ;
 wire \mod_ro_128.fabric[13] ;
 wire \mod_ro_128.fabric[14] ;
 wire \mod_ro_128.fabric[15] ;
 wire \mod_ro_128.fabric[16] ;
 wire \mod_ro_128.fabric[17] ;
 wire \mod_ro_128.fabric[18] ;
 wire \mod_ro_128.fabric[19] ;
 wire \mod_ro_128.fabric[1] ;
 wire \mod_ro_128.fabric[20] ;
 wire \mod_ro_128.fabric[21] ;
 wire \mod_ro_128.fabric[22] ;
 wire \mod_ro_128.fabric[23] ;
 wire \mod_ro_128.fabric[24] ;
 wire \mod_ro_128.fabric[25] ;
 wire \mod_ro_128.fabric[26] ;
 wire \mod_ro_128.fabric[27] ;
 wire \mod_ro_128.fabric[28] ;
 wire \mod_ro_128.fabric[29] ;
 wire \mod_ro_128.fabric[2] ;
 wire \mod_ro_128.fabric[30] ;
 wire \mod_ro_128.fabric[31] ;
 wire \mod_ro_128.fabric[32] ;
 wire \mod_ro_128.fabric[33] ;
 wire \mod_ro_128.fabric[34] ;
 wire \mod_ro_128.fabric[35] ;
 wire \mod_ro_128.fabric[36] ;
 wire \mod_ro_128.fabric[37] ;
 wire \mod_ro_128.fabric[38] ;
 wire \mod_ro_128.fabric[39] ;
 wire \mod_ro_128.fabric[3] ;
 wire \mod_ro_128.fabric[40] ;
 wire \mod_ro_128.fabric[41] ;
 wire \mod_ro_128.fabric[42] ;
 wire \mod_ro_128.fabric[43] ;
 wire \mod_ro_128.fabric[44] ;
 wire \mod_ro_128.fabric[45] ;
 wire \mod_ro_128.fabric[46] ;
 wire \mod_ro_128.fabric[47] ;
 wire \mod_ro_128.fabric[48] ;
 wire \mod_ro_128.fabric[49] ;
 wire \mod_ro_128.fabric[4] ;
 wire \mod_ro_128.fabric[50] ;
 wire \mod_ro_128.fabric[51] ;
 wire \mod_ro_128.fabric[52] ;
 wire \mod_ro_128.fabric[53] ;
 wire \mod_ro_128.fabric[54] ;
 wire \mod_ro_128.fabric[55] ;
 wire \mod_ro_128.fabric[56] ;
 wire \mod_ro_128.fabric[57] ;
 wire \mod_ro_128.fabric[58] ;
 wire \mod_ro_128.fabric[59] ;
 wire \mod_ro_128.fabric[5] ;
 wire \mod_ro_128.fabric[60] ;
 wire \mod_ro_128.fabric[61] ;
 wire \mod_ro_128.fabric[62] ;
 wire \mod_ro_128.fabric[63] ;
 wire \mod_ro_128.fabric[64] ;
 wire \mod_ro_128.fabric[65] ;
 wire \mod_ro_128.fabric[66] ;
 wire \mod_ro_128.fabric[67] ;
 wire \mod_ro_128.fabric[68] ;
 wire \mod_ro_128.fabric[69] ;
 wire \mod_ro_128.fabric[6] ;
 wire \mod_ro_128.fabric[70] ;
 wire \mod_ro_128.fabric[71] ;
 wire \mod_ro_128.fabric[72] ;
 wire \mod_ro_128.fabric[73] ;
 wire \mod_ro_128.fabric[74] ;
 wire \mod_ro_128.fabric[75] ;
 wire \mod_ro_128.fabric[76] ;
 wire \mod_ro_128.fabric[77] ;
 wire \mod_ro_128.fabric[78] ;
 wire \mod_ro_128.fabric[79] ;
 wire \mod_ro_128.fabric[7] ;
 wire \mod_ro_128.fabric[80] ;
 wire \mod_ro_128.fabric[81] ;
 wire \mod_ro_128.fabric[82] ;
 wire \mod_ro_128.fabric[83] ;
 wire \mod_ro_128.fabric[84] ;
 wire \mod_ro_128.fabric[85] ;
 wire \mod_ro_128.fabric[86] ;
 wire \mod_ro_128.fabric[87] ;
 wire \mod_ro_128.fabric[88] ;
 wire \mod_ro_128.fabric[89] ;
 wire \mod_ro_128.fabric[8] ;
 wire \mod_ro_128.fabric[90] ;
 wire \mod_ro_128.fabric[91] ;
 wire \mod_ro_128.fabric[92] ;
 wire \mod_ro_128.fabric[93] ;
 wire \mod_ro_128.fabric[94] ;
 wire \mod_ro_128.fabric[95] ;
 wire \mod_ro_128.fabric[96] ;
 wire \mod_ro_128.fabric[97] ;
 wire \mod_ro_128.fabric[98] ;
 wire \mod_ro_128.fabric[99] ;
 wire \mod_ro_128.fabric[9] ;
 wire \mod_ro_16.fabric[0] ;
 wire \mod_ro_16.fabric[10] ;
 wire \mod_ro_16.fabric[11] ;
 wire \mod_ro_16.fabric[12] ;
 wire \mod_ro_16.fabric[13] ;
 wire \mod_ro_16.fabric[14] ;
 wire \mod_ro_16.fabric[15] ;
 wire \mod_ro_16.fabric[16] ;
 wire \mod_ro_16.fabric[1] ;
 wire \mod_ro_16.fabric[2] ;
 wire \mod_ro_16.fabric[3] ;
 wire \mod_ro_16.fabric[4] ;
 wire \mod_ro_16.fabric[5] ;
 wire \mod_ro_16.fabric[6] ;
 wire \mod_ro_16.fabric[7] ;
 wire \mod_ro_16.fabric[8] ;
 wire \mod_ro_16.fabric[9] ;
 wire \mod_ro_31.fabric[0] ;
 wire \mod_ro_31.fabric[10] ;
 wire \mod_ro_31.fabric[11] ;
 wire \mod_ro_31.fabric[12] ;
 wire \mod_ro_31.fabric[13] ;
 wire \mod_ro_31.fabric[14] ;
 wire \mod_ro_31.fabric[15] ;
 wire \mod_ro_31.fabric[16] ;
 wire \mod_ro_31.fabric[17] ;
 wire \mod_ro_31.fabric[18] ;
 wire \mod_ro_31.fabric[19] ;
 wire \mod_ro_31.fabric[1] ;
 wire \mod_ro_31.fabric[20] ;
 wire \mod_ro_31.fabric[21] ;
 wire \mod_ro_31.fabric[22] ;
 wire \mod_ro_31.fabric[23] ;
 wire \mod_ro_31.fabric[24] ;
 wire \mod_ro_31.fabric[25] ;
 wire \mod_ro_31.fabric[26] ;
 wire \mod_ro_31.fabric[27] ;
 wire \mod_ro_31.fabric[28] ;
 wire \mod_ro_31.fabric[29] ;
 wire \mod_ro_31.fabric[2] ;
 wire \mod_ro_31.fabric[30] ;
 wire \mod_ro_31.fabric[31] ;
 wire \mod_ro_31.fabric[3] ;
 wire \mod_ro_31.fabric[4] ;
 wire \mod_ro_31.fabric[5] ;
 wire \mod_ro_31.fabric[6] ;
 wire \mod_ro_31.fabric[7] ;
 wire \mod_ro_31.fabric[8] ;
 wire \mod_ro_31.fabric[9] ;
 wire \mod_ro_32_1.fabric[0] ;
 wire \mod_ro_32_1.fabric[10] ;
 wire \mod_ro_32_1.fabric[11] ;
 wire \mod_ro_32_1.fabric[12] ;
 wire \mod_ro_32_1.fabric[13] ;
 wire \mod_ro_32_1.fabric[14] ;
 wire \mod_ro_32_1.fabric[15] ;
 wire \mod_ro_32_1.fabric[16] ;
 wire \mod_ro_32_1.fabric[17] ;
 wire \mod_ro_32_1.fabric[18] ;
 wire \mod_ro_32_1.fabric[19] ;
 wire \mod_ro_32_1.fabric[1] ;
 wire \mod_ro_32_1.fabric[20] ;
 wire \mod_ro_32_1.fabric[21] ;
 wire \mod_ro_32_1.fabric[22] ;
 wire \mod_ro_32_1.fabric[23] ;
 wire \mod_ro_32_1.fabric[24] ;
 wire \mod_ro_32_1.fabric[25] ;
 wire \mod_ro_32_1.fabric[26] ;
 wire \mod_ro_32_1.fabric[27] ;
 wire \mod_ro_32_1.fabric[28] ;
 wire \mod_ro_32_1.fabric[29] ;
 wire \mod_ro_32_1.fabric[2] ;
 wire \mod_ro_32_1.fabric[30] ;
 wire \mod_ro_32_1.fabric[31] ;
 wire \mod_ro_32_1.fabric[32] ;
 wire \mod_ro_32_1.fabric[3] ;
 wire \mod_ro_32_1.fabric[4] ;
 wire \mod_ro_32_1.fabric[5] ;
 wire \mod_ro_32_1.fabric[6] ;
 wire \mod_ro_32_1.fabric[7] ;
 wire \mod_ro_32_1.fabric[8] ;
 wire \mod_ro_32_1.fabric[9] ;
 wire \mod_ro_32_2.fabric[0] ;
 wire \mod_ro_32_2.fabric[10] ;
 wire \mod_ro_32_2.fabric[11] ;
 wire \mod_ro_32_2.fabric[12] ;
 wire \mod_ro_32_2.fabric[13] ;
 wire \mod_ro_32_2.fabric[14] ;
 wire \mod_ro_32_2.fabric[15] ;
 wire \mod_ro_32_2.fabric[16] ;
 wire \mod_ro_32_2.fabric[17] ;
 wire \mod_ro_32_2.fabric[18] ;
 wire \mod_ro_32_2.fabric[19] ;
 wire \mod_ro_32_2.fabric[1] ;
 wire \mod_ro_32_2.fabric[20] ;
 wire \mod_ro_32_2.fabric[21] ;
 wire \mod_ro_32_2.fabric[22] ;
 wire \mod_ro_32_2.fabric[23] ;
 wire \mod_ro_32_2.fabric[24] ;
 wire \mod_ro_32_2.fabric[25] ;
 wire \mod_ro_32_2.fabric[26] ;
 wire \mod_ro_32_2.fabric[27] ;
 wire \mod_ro_32_2.fabric[28] ;
 wire \mod_ro_32_2.fabric[29] ;
 wire \mod_ro_32_2.fabric[2] ;
 wire \mod_ro_32_2.fabric[30] ;
 wire \mod_ro_32_2.fabric[31] ;
 wire \mod_ro_32_2.fabric[32] ;
 wire \mod_ro_32_2.fabric[3] ;
 wire \mod_ro_32_2.fabric[4] ;
 wire \mod_ro_32_2.fabric[5] ;
 wire \mod_ro_32_2.fabric[6] ;
 wire \mod_ro_32_2.fabric[7] ;
 wire \mod_ro_32_2.fabric[8] ;
 wire \mod_ro_32_2.fabric[9] ;
 wire \mod_ro_32_raw.fabric[0] ;
 wire \mod_ro_32_raw.fabric[10] ;
 wire \mod_ro_32_raw.fabric[11] ;
 wire \mod_ro_32_raw.fabric[12] ;
 wire \mod_ro_32_raw.fabric[13] ;
 wire \mod_ro_32_raw.fabric[14] ;
 wire \mod_ro_32_raw.fabric[15] ;
 wire \mod_ro_32_raw.fabric[16] ;
 wire \mod_ro_32_raw.fabric[17] ;
 wire \mod_ro_32_raw.fabric[18] ;
 wire \mod_ro_32_raw.fabric[19] ;
 wire \mod_ro_32_raw.fabric[1] ;
 wire \mod_ro_32_raw.fabric[20] ;
 wire \mod_ro_32_raw.fabric[21] ;
 wire \mod_ro_32_raw.fabric[22] ;
 wire \mod_ro_32_raw.fabric[23] ;
 wire \mod_ro_32_raw.fabric[24] ;
 wire \mod_ro_32_raw.fabric[25] ;
 wire \mod_ro_32_raw.fabric[26] ;
 wire \mod_ro_32_raw.fabric[27] ;
 wire \mod_ro_32_raw.fabric[28] ;
 wire \mod_ro_32_raw.fabric[29] ;
 wire \mod_ro_32_raw.fabric[2] ;
 wire \mod_ro_32_raw.fabric[30] ;
 wire \mod_ro_32_raw.fabric[31] ;
 wire \mod_ro_32_raw.fabric[32] ;
 wire \mod_ro_32_raw.fabric[3] ;
 wire \mod_ro_32_raw.fabric[4] ;
 wire \mod_ro_32_raw.fabric[5] ;
 wire \mod_ro_32_raw.fabric[6] ;
 wire \mod_ro_32_raw.fabric[7] ;
 wire \mod_ro_32_raw.fabric[8] ;
 wire \mod_ro_32_raw.fabric[9] ;
 wire \mod_ro_64.fabric[0] ;
 wire \mod_ro_64.fabric[10] ;
 wire \mod_ro_64.fabric[11] ;
 wire \mod_ro_64.fabric[12] ;
 wire \mod_ro_64.fabric[13] ;
 wire \mod_ro_64.fabric[14] ;
 wire \mod_ro_64.fabric[15] ;
 wire \mod_ro_64.fabric[16] ;
 wire \mod_ro_64.fabric[17] ;
 wire \mod_ro_64.fabric[18] ;
 wire \mod_ro_64.fabric[19] ;
 wire \mod_ro_64.fabric[1] ;
 wire \mod_ro_64.fabric[20] ;
 wire \mod_ro_64.fabric[21] ;
 wire \mod_ro_64.fabric[22] ;
 wire \mod_ro_64.fabric[23] ;
 wire \mod_ro_64.fabric[24] ;
 wire \mod_ro_64.fabric[25] ;
 wire \mod_ro_64.fabric[26] ;
 wire \mod_ro_64.fabric[27] ;
 wire \mod_ro_64.fabric[28] ;
 wire \mod_ro_64.fabric[29] ;
 wire \mod_ro_64.fabric[2] ;
 wire \mod_ro_64.fabric[30] ;
 wire \mod_ro_64.fabric[31] ;
 wire \mod_ro_64.fabric[32] ;
 wire \mod_ro_64.fabric[33] ;
 wire \mod_ro_64.fabric[34] ;
 wire \mod_ro_64.fabric[35] ;
 wire \mod_ro_64.fabric[36] ;
 wire \mod_ro_64.fabric[37] ;
 wire \mod_ro_64.fabric[38] ;
 wire \mod_ro_64.fabric[39] ;
 wire \mod_ro_64.fabric[3] ;
 wire \mod_ro_64.fabric[40] ;
 wire \mod_ro_64.fabric[41] ;
 wire \mod_ro_64.fabric[42] ;
 wire \mod_ro_64.fabric[43] ;
 wire \mod_ro_64.fabric[44] ;
 wire \mod_ro_64.fabric[45] ;
 wire \mod_ro_64.fabric[46] ;
 wire \mod_ro_64.fabric[47] ;
 wire \mod_ro_64.fabric[48] ;
 wire \mod_ro_64.fabric[49] ;
 wire \mod_ro_64.fabric[4] ;
 wire \mod_ro_64.fabric[50] ;
 wire \mod_ro_64.fabric[51] ;
 wire \mod_ro_64.fabric[52] ;
 wire \mod_ro_64.fabric[53] ;
 wire \mod_ro_64.fabric[54] ;
 wire \mod_ro_64.fabric[55] ;
 wire \mod_ro_64.fabric[56] ;
 wire \mod_ro_64.fabric[57] ;
 wire \mod_ro_64.fabric[58] ;
 wire \mod_ro_64.fabric[59] ;
 wire \mod_ro_64.fabric[5] ;
 wire \mod_ro_64.fabric[60] ;
 wire \mod_ro_64.fabric[61] ;
 wire \mod_ro_64.fabric[62] ;
 wire \mod_ro_64.fabric[63] ;
 wire \mod_ro_64.fabric[64] ;
 wire \mod_ro_64.fabric[6] ;
 wire \mod_ro_64.fabric[7] ;
 wire \mod_ro_64.fabric[8] ;
 wire \mod_ro_64.fabric[9] ;
 wire mux_out;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;

 sg13g2_inv_1 _09_ (.Y(_00_),
    .A(net1));
 sg13g2_inv_1 _10_ (.Y(_01_),
    .A(net2));
 sg13g2_mux2_1 _11_ (.A0(\mod_ro_32_2.fabric[0] ),
    .A1(\mod_ro_31.fabric[0] ),
    .S(net3),
    .X(_02_));
 sg13g2_nand2_1 _12_ (.Y(_03_),
    .A(net1),
    .B(_02_));
 sg13g2_a21o_1 _13_ (.A2(\mod_ro_32_2.fabric[0] ),
    .A1(net3),
    .B1(\mod_ro_32_1.fabric[0] ),
    .X(_04_));
 sg13g2_a21oi_1 _14_ (.A1(_00_),
    .A2(_04_),
    .Y(_05_),
    .B1(net2));
 sg13g2_mux2_1 _15_ (.A0(\mod_ro_64.fabric[0] ),
    .A1(\mod_ro_128.fabric[0] ),
    .S(net3),
    .X(_06_));
 sg13g2_nand3b_1 _16_ (.B(net1),
    .C(\mod_ro_16.fabric[0] ),
    .Y(_07_),
    .A_N(net3));
 sg13g2_a21oi_1 _17_ (.A1(_00_),
    .A2(_06_),
    .Y(_08_),
    .B1(_01_));
 sg13g2_a22oi_1 _18_ (.Y(mux_out),
    .B1(_07_),
    .B2(_08_),
    .A2(_05_),
    .A1(_03_));
 sg13g2_tielo tt_um_wedgetail_tester_5 (.L_LO(net5));
 sg13g2_tielo tt_um_wedgetail_tester_6 (.L_LO(net6));
 sg13g2_tielo tt_um_wedgetail_tester_7 (.L_LO(net7));
 sg13g2_tielo tt_um_wedgetail_tester_8 (.L_LO(net8));
 sg13g2_tielo tt_um_wedgetail_tester_9 (.L_LO(net9));
 sg13g2_tielo tt_um_wedgetail_tester_10 (.L_LO(net10));
 sg13g2_tielo tt_um_wedgetail_tester_11 (.L_LO(net11));
 sg13g2_tielo tt_um_wedgetail_tester_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wedgetail_tester_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wedgetail_tester_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wedgetail_tester_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wedgetail_tester_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wedgetail_tester_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wedgetail_tester_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wedgetail_tester_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wedgetail_tester_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wedgetail_tester_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wedgetail_tester_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wedgetail_tester_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wedgetail_tester_24 (.L_LO(net24));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _40_ (.A(mux_out),
    .X(uo_out[0]));
 sg13g2_buf_1 _41_ (.A(clk),
    .X(uo_out[1]));
 sg13g2_buf_1 _42_ (.A(\mod_ro_32_raw.fabric[0] ),
    .X(uo_out[2]));
 sg13g2_inv_1 \mod_ro_128.feedback  (.Y(\mod_ro_128.fabric[0] ),
    .A(\mod_ro_128.fabric[128] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[0].inv  (.Y(\mod_ro_128.fabric[1] ),
    .A(\mod_ro_128.fabric[0] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[100].inv  (.Y(\mod_ro_128.fabric[101] ),
    .A(\mod_ro_128.fabric[100] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[101].inv  (.Y(\mod_ro_128.fabric[102] ),
    .A(\mod_ro_128.fabric[101] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[102].inv  (.Y(\mod_ro_128.fabric[103] ),
    .A(\mod_ro_128.fabric[102] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[103].inv  (.Y(\mod_ro_128.fabric[104] ),
    .A(\mod_ro_128.fabric[103] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[104].inv  (.Y(\mod_ro_128.fabric[105] ),
    .A(\mod_ro_128.fabric[104] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[105].inv  (.Y(\mod_ro_128.fabric[106] ),
    .A(\mod_ro_128.fabric[105] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[106].inv  (.Y(\mod_ro_128.fabric[107] ),
    .A(\mod_ro_128.fabric[106] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[107].inv  (.Y(\mod_ro_128.fabric[108] ),
    .A(\mod_ro_128.fabric[107] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[108].inv  (.Y(\mod_ro_128.fabric[109] ),
    .A(\mod_ro_128.fabric[108] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[109].inv  (.Y(\mod_ro_128.fabric[110] ),
    .A(\mod_ro_128.fabric[109] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[10].inv  (.Y(\mod_ro_128.fabric[11] ),
    .A(\mod_ro_128.fabric[10] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[110].inv  (.Y(\mod_ro_128.fabric[111] ),
    .A(\mod_ro_128.fabric[110] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[111].inv  (.Y(\mod_ro_128.fabric[112] ),
    .A(\mod_ro_128.fabric[111] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[112].inv  (.Y(\mod_ro_128.fabric[113] ),
    .A(\mod_ro_128.fabric[112] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[113].inv  (.Y(\mod_ro_128.fabric[114] ),
    .A(\mod_ro_128.fabric[113] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[114].inv  (.Y(\mod_ro_128.fabric[115] ),
    .A(\mod_ro_128.fabric[114] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[115].inv  (.Y(\mod_ro_128.fabric[116] ),
    .A(\mod_ro_128.fabric[115] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[116].inv  (.Y(\mod_ro_128.fabric[117] ),
    .A(\mod_ro_128.fabric[116] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[117].inv  (.Y(\mod_ro_128.fabric[118] ),
    .A(\mod_ro_128.fabric[117] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[118].inv  (.Y(\mod_ro_128.fabric[119] ),
    .A(\mod_ro_128.fabric[118] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[119].inv  (.Y(\mod_ro_128.fabric[120] ),
    .A(\mod_ro_128.fabric[119] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[11].inv  (.Y(\mod_ro_128.fabric[12] ),
    .A(\mod_ro_128.fabric[11] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[120].inv  (.Y(\mod_ro_128.fabric[121] ),
    .A(\mod_ro_128.fabric[120] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[121].inv  (.Y(\mod_ro_128.fabric[122] ),
    .A(\mod_ro_128.fabric[121] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[122].inv  (.Y(\mod_ro_128.fabric[123] ),
    .A(\mod_ro_128.fabric[122] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[123].inv  (.Y(\mod_ro_128.fabric[124] ),
    .A(\mod_ro_128.fabric[123] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[124].inv  (.Y(\mod_ro_128.fabric[125] ),
    .A(\mod_ro_128.fabric[124] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[125].inv  (.Y(\mod_ro_128.fabric[126] ),
    .A(\mod_ro_128.fabric[125] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[126].inv  (.Y(\mod_ro_128.fabric[127] ),
    .A(\mod_ro_128.fabric[126] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[127].inv  (.Y(\mod_ro_128.fabric[128] ),
    .A(\mod_ro_128.fabric[127] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[12].inv  (.Y(\mod_ro_128.fabric[13] ),
    .A(\mod_ro_128.fabric[12] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[13].inv  (.Y(\mod_ro_128.fabric[14] ),
    .A(\mod_ro_128.fabric[13] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[14].inv  (.Y(\mod_ro_128.fabric[15] ),
    .A(\mod_ro_128.fabric[14] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[15].inv  (.Y(\mod_ro_128.fabric[16] ),
    .A(\mod_ro_128.fabric[15] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[16].inv  (.Y(\mod_ro_128.fabric[17] ),
    .A(\mod_ro_128.fabric[16] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[17].inv  (.Y(\mod_ro_128.fabric[18] ),
    .A(\mod_ro_128.fabric[17] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[18].inv  (.Y(\mod_ro_128.fabric[19] ),
    .A(\mod_ro_128.fabric[18] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[19].inv  (.Y(\mod_ro_128.fabric[20] ),
    .A(\mod_ro_128.fabric[19] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[1].inv  (.Y(\mod_ro_128.fabric[2] ),
    .A(\mod_ro_128.fabric[1] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[20].inv  (.Y(\mod_ro_128.fabric[21] ),
    .A(\mod_ro_128.fabric[20] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[21].inv  (.Y(\mod_ro_128.fabric[22] ),
    .A(\mod_ro_128.fabric[21] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[22].inv  (.Y(\mod_ro_128.fabric[23] ),
    .A(\mod_ro_128.fabric[22] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[23].inv  (.Y(\mod_ro_128.fabric[24] ),
    .A(\mod_ro_128.fabric[23] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[24].inv  (.Y(\mod_ro_128.fabric[25] ),
    .A(\mod_ro_128.fabric[24] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[25].inv  (.Y(\mod_ro_128.fabric[26] ),
    .A(\mod_ro_128.fabric[25] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[26].inv  (.Y(\mod_ro_128.fabric[27] ),
    .A(\mod_ro_128.fabric[26] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[27].inv  (.Y(\mod_ro_128.fabric[28] ),
    .A(\mod_ro_128.fabric[27] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[28].inv  (.Y(\mod_ro_128.fabric[29] ),
    .A(\mod_ro_128.fabric[28] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[29].inv  (.Y(\mod_ro_128.fabric[30] ),
    .A(\mod_ro_128.fabric[29] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[2].inv  (.Y(\mod_ro_128.fabric[3] ),
    .A(\mod_ro_128.fabric[2] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[30].inv  (.Y(\mod_ro_128.fabric[31] ),
    .A(\mod_ro_128.fabric[30] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[31].inv  (.Y(\mod_ro_128.fabric[32] ),
    .A(\mod_ro_128.fabric[31] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[32].inv  (.Y(\mod_ro_128.fabric[33] ),
    .A(\mod_ro_128.fabric[32] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[33].inv  (.Y(\mod_ro_128.fabric[34] ),
    .A(\mod_ro_128.fabric[33] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[34].inv  (.Y(\mod_ro_128.fabric[35] ),
    .A(\mod_ro_128.fabric[34] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[35].inv  (.Y(\mod_ro_128.fabric[36] ),
    .A(\mod_ro_128.fabric[35] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[36].inv  (.Y(\mod_ro_128.fabric[37] ),
    .A(\mod_ro_128.fabric[36] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[37].inv  (.Y(\mod_ro_128.fabric[38] ),
    .A(\mod_ro_128.fabric[37] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[38].inv  (.Y(\mod_ro_128.fabric[39] ),
    .A(\mod_ro_128.fabric[38] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[39].inv  (.Y(\mod_ro_128.fabric[40] ),
    .A(\mod_ro_128.fabric[39] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[3].inv  (.Y(\mod_ro_128.fabric[4] ),
    .A(\mod_ro_128.fabric[3] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[40].inv  (.Y(\mod_ro_128.fabric[41] ),
    .A(\mod_ro_128.fabric[40] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[41].inv  (.Y(\mod_ro_128.fabric[42] ),
    .A(\mod_ro_128.fabric[41] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[42].inv  (.Y(\mod_ro_128.fabric[43] ),
    .A(\mod_ro_128.fabric[42] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[43].inv  (.Y(\mod_ro_128.fabric[44] ),
    .A(\mod_ro_128.fabric[43] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[44].inv  (.Y(\mod_ro_128.fabric[45] ),
    .A(\mod_ro_128.fabric[44] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[45].inv  (.Y(\mod_ro_128.fabric[46] ),
    .A(\mod_ro_128.fabric[45] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[46].inv  (.Y(\mod_ro_128.fabric[47] ),
    .A(\mod_ro_128.fabric[46] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[47].inv  (.Y(\mod_ro_128.fabric[48] ),
    .A(\mod_ro_128.fabric[47] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[48].inv  (.Y(\mod_ro_128.fabric[49] ),
    .A(\mod_ro_128.fabric[48] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[49].inv  (.Y(\mod_ro_128.fabric[50] ),
    .A(\mod_ro_128.fabric[49] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[4].inv  (.Y(\mod_ro_128.fabric[5] ),
    .A(\mod_ro_128.fabric[4] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[50].inv  (.Y(\mod_ro_128.fabric[51] ),
    .A(\mod_ro_128.fabric[50] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[51].inv  (.Y(\mod_ro_128.fabric[52] ),
    .A(\mod_ro_128.fabric[51] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[52].inv  (.Y(\mod_ro_128.fabric[53] ),
    .A(\mod_ro_128.fabric[52] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[53].inv  (.Y(\mod_ro_128.fabric[54] ),
    .A(\mod_ro_128.fabric[53] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[54].inv  (.Y(\mod_ro_128.fabric[55] ),
    .A(\mod_ro_128.fabric[54] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[55].inv  (.Y(\mod_ro_128.fabric[56] ),
    .A(\mod_ro_128.fabric[55] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[56].inv  (.Y(\mod_ro_128.fabric[57] ),
    .A(\mod_ro_128.fabric[56] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[57].inv  (.Y(\mod_ro_128.fabric[58] ),
    .A(\mod_ro_128.fabric[57] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[58].inv  (.Y(\mod_ro_128.fabric[59] ),
    .A(\mod_ro_128.fabric[58] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[59].inv  (.Y(\mod_ro_128.fabric[60] ),
    .A(\mod_ro_128.fabric[59] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[5].inv  (.Y(\mod_ro_128.fabric[6] ),
    .A(\mod_ro_128.fabric[5] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[60].inv  (.Y(\mod_ro_128.fabric[61] ),
    .A(\mod_ro_128.fabric[60] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[61].inv  (.Y(\mod_ro_128.fabric[62] ),
    .A(\mod_ro_128.fabric[61] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[62].inv  (.Y(\mod_ro_128.fabric[63] ),
    .A(\mod_ro_128.fabric[62] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[63].inv  (.Y(\mod_ro_128.fabric[64] ),
    .A(\mod_ro_128.fabric[63] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[64].inv  (.Y(\mod_ro_128.fabric[65] ),
    .A(\mod_ro_128.fabric[64] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[65].inv  (.Y(\mod_ro_128.fabric[66] ),
    .A(\mod_ro_128.fabric[65] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[66].inv  (.Y(\mod_ro_128.fabric[67] ),
    .A(\mod_ro_128.fabric[66] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[67].inv  (.Y(\mod_ro_128.fabric[68] ),
    .A(\mod_ro_128.fabric[67] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[68].inv  (.Y(\mod_ro_128.fabric[69] ),
    .A(\mod_ro_128.fabric[68] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[69].inv  (.Y(\mod_ro_128.fabric[70] ),
    .A(\mod_ro_128.fabric[69] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[6].inv  (.Y(\mod_ro_128.fabric[7] ),
    .A(\mod_ro_128.fabric[6] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[70].inv  (.Y(\mod_ro_128.fabric[71] ),
    .A(\mod_ro_128.fabric[70] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[71].inv  (.Y(\mod_ro_128.fabric[72] ),
    .A(\mod_ro_128.fabric[71] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[72].inv  (.Y(\mod_ro_128.fabric[73] ),
    .A(\mod_ro_128.fabric[72] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[73].inv  (.Y(\mod_ro_128.fabric[74] ),
    .A(\mod_ro_128.fabric[73] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[74].inv  (.Y(\mod_ro_128.fabric[75] ),
    .A(\mod_ro_128.fabric[74] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[75].inv  (.Y(\mod_ro_128.fabric[76] ),
    .A(\mod_ro_128.fabric[75] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[76].inv  (.Y(\mod_ro_128.fabric[77] ),
    .A(\mod_ro_128.fabric[76] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[77].inv  (.Y(\mod_ro_128.fabric[78] ),
    .A(\mod_ro_128.fabric[77] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[78].inv  (.Y(\mod_ro_128.fabric[79] ),
    .A(\mod_ro_128.fabric[78] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[79].inv  (.Y(\mod_ro_128.fabric[80] ),
    .A(\mod_ro_128.fabric[79] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[7].inv  (.Y(\mod_ro_128.fabric[8] ),
    .A(\mod_ro_128.fabric[7] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[80].inv  (.Y(\mod_ro_128.fabric[81] ),
    .A(\mod_ro_128.fabric[80] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[81].inv  (.Y(\mod_ro_128.fabric[82] ),
    .A(\mod_ro_128.fabric[81] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[82].inv  (.Y(\mod_ro_128.fabric[83] ),
    .A(\mod_ro_128.fabric[82] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[83].inv  (.Y(\mod_ro_128.fabric[84] ),
    .A(\mod_ro_128.fabric[83] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[84].inv  (.Y(\mod_ro_128.fabric[85] ),
    .A(\mod_ro_128.fabric[84] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[85].inv  (.Y(\mod_ro_128.fabric[86] ),
    .A(\mod_ro_128.fabric[85] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[86].inv  (.Y(\mod_ro_128.fabric[87] ),
    .A(\mod_ro_128.fabric[86] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[87].inv  (.Y(\mod_ro_128.fabric[88] ),
    .A(\mod_ro_128.fabric[87] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[88].inv  (.Y(\mod_ro_128.fabric[89] ),
    .A(\mod_ro_128.fabric[88] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[89].inv  (.Y(\mod_ro_128.fabric[90] ),
    .A(\mod_ro_128.fabric[89] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[8].inv  (.Y(\mod_ro_128.fabric[9] ),
    .A(\mod_ro_128.fabric[8] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[90].inv  (.Y(\mod_ro_128.fabric[91] ),
    .A(\mod_ro_128.fabric[90] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[91].inv  (.Y(\mod_ro_128.fabric[92] ),
    .A(\mod_ro_128.fabric[91] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[92].inv  (.Y(\mod_ro_128.fabric[93] ),
    .A(\mod_ro_128.fabric[92] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[93].inv  (.Y(\mod_ro_128.fabric[94] ),
    .A(\mod_ro_128.fabric[93] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[94].inv  (.Y(\mod_ro_128.fabric[95] ),
    .A(\mod_ro_128.fabric[94] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[95].inv  (.Y(\mod_ro_128.fabric[96] ),
    .A(\mod_ro_128.fabric[95] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[96].inv  (.Y(\mod_ro_128.fabric[97] ),
    .A(\mod_ro_128.fabric[96] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[97].inv  (.Y(\mod_ro_128.fabric[98] ),
    .A(\mod_ro_128.fabric[97] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[98].inv  (.Y(\mod_ro_128.fabric[99] ),
    .A(\mod_ro_128.fabric[98] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[99].inv  (.Y(\mod_ro_128.fabric[100] ),
    .A(\mod_ro_128.fabric[99] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[9].inv  (.Y(\mod_ro_128.fabric[10] ),
    .A(\mod_ro_128.fabric[9] ));
 sg13g2_inv_1 \mod_ro_16.feedback  (.Y(\mod_ro_16.fabric[0] ),
    .A(\mod_ro_16.fabric[16] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[0].inv  (.Y(\mod_ro_16.fabric[1] ),
    .A(\mod_ro_16.fabric[0] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[10].inv  (.Y(\mod_ro_16.fabric[11] ),
    .A(\mod_ro_16.fabric[10] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[11].inv  (.Y(\mod_ro_16.fabric[12] ),
    .A(\mod_ro_16.fabric[11] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[12].inv  (.Y(\mod_ro_16.fabric[13] ),
    .A(\mod_ro_16.fabric[12] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[13].inv  (.Y(\mod_ro_16.fabric[14] ),
    .A(\mod_ro_16.fabric[13] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[14].inv  (.Y(\mod_ro_16.fabric[15] ),
    .A(\mod_ro_16.fabric[14] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[15].inv  (.Y(\mod_ro_16.fabric[16] ),
    .A(\mod_ro_16.fabric[15] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[1].inv  (.Y(\mod_ro_16.fabric[2] ),
    .A(\mod_ro_16.fabric[1] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[2].inv  (.Y(\mod_ro_16.fabric[3] ),
    .A(\mod_ro_16.fabric[2] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[3].inv  (.Y(\mod_ro_16.fabric[4] ),
    .A(\mod_ro_16.fabric[3] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[4].inv  (.Y(\mod_ro_16.fabric[5] ),
    .A(\mod_ro_16.fabric[4] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[5].inv  (.Y(\mod_ro_16.fabric[6] ),
    .A(\mod_ro_16.fabric[5] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[6].inv  (.Y(\mod_ro_16.fabric[7] ),
    .A(\mod_ro_16.fabric[6] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[7].inv  (.Y(\mod_ro_16.fabric[8] ),
    .A(\mod_ro_16.fabric[7] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[8].inv  (.Y(\mod_ro_16.fabric[9] ),
    .A(\mod_ro_16.fabric[8] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[9].inv  (.Y(\mod_ro_16.fabric[10] ),
    .A(\mod_ro_16.fabric[9] ));
 sg13g2_inv_1 \mod_ro_31.feedback  (.Y(\mod_ro_31.fabric[0] ),
    .A(\mod_ro_31.fabric[31] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[0].inv  (.Y(\mod_ro_31.fabric[1] ),
    .A(\mod_ro_31.fabric[0] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[10].inv  (.Y(\mod_ro_31.fabric[11] ),
    .A(\mod_ro_31.fabric[10] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[11].inv  (.Y(\mod_ro_31.fabric[12] ),
    .A(\mod_ro_31.fabric[11] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[12].inv  (.Y(\mod_ro_31.fabric[13] ),
    .A(\mod_ro_31.fabric[12] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[13].inv  (.Y(\mod_ro_31.fabric[14] ),
    .A(\mod_ro_31.fabric[13] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[14].inv  (.Y(\mod_ro_31.fabric[15] ),
    .A(\mod_ro_31.fabric[14] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[15].inv  (.Y(\mod_ro_31.fabric[16] ),
    .A(\mod_ro_31.fabric[15] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[16].inv  (.Y(\mod_ro_31.fabric[17] ),
    .A(\mod_ro_31.fabric[16] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[17].inv  (.Y(\mod_ro_31.fabric[18] ),
    .A(\mod_ro_31.fabric[17] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[18].inv  (.Y(\mod_ro_31.fabric[19] ),
    .A(\mod_ro_31.fabric[18] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[19].inv  (.Y(\mod_ro_31.fabric[20] ),
    .A(\mod_ro_31.fabric[19] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[1].inv  (.Y(\mod_ro_31.fabric[2] ),
    .A(\mod_ro_31.fabric[1] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[20].inv  (.Y(\mod_ro_31.fabric[21] ),
    .A(\mod_ro_31.fabric[20] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[21].inv  (.Y(\mod_ro_31.fabric[22] ),
    .A(\mod_ro_31.fabric[21] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[22].inv  (.Y(\mod_ro_31.fabric[23] ),
    .A(\mod_ro_31.fabric[22] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[23].inv  (.Y(\mod_ro_31.fabric[24] ),
    .A(\mod_ro_31.fabric[23] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[24].inv  (.Y(\mod_ro_31.fabric[25] ),
    .A(\mod_ro_31.fabric[24] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[25].inv  (.Y(\mod_ro_31.fabric[26] ),
    .A(\mod_ro_31.fabric[25] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[26].inv  (.Y(\mod_ro_31.fabric[27] ),
    .A(\mod_ro_31.fabric[26] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[27].inv  (.Y(\mod_ro_31.fabric[28] ),
    .A(\mod_ro_31.fabric[27] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[28].inv  (.Y(\mod_ro_31.fabric[29] ),
    .A(\mod_ro_31.fabric[28] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[29].inv  (.Y(\mod_ro_31.fabric[30] ),
    .A(\mod_ro_31.fabric[29] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[2].inv  (.Y(\mod_ro_31.fabric[3] ),
    .A(\mod_ro_31.fabric[2] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[30].inv  (.Y(\mod_ro_31.fabric[31] ),
    .A(\mod_ro_31.fabric[30] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[3].inv  (.Y(\mod_ro_31.fabric[4] ),
    .A(\mod_ro_31.fabric[3] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[4].inv  (.Y(\mod_ro_31.fabric[5] ),
    .A(\mod_ro_31.fabric[4] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[5].inv  (.Y(\mod_ro_31.fabric[6] ),
    .A(\mod_ro_31.fabric[5] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[6].inv  (.Y(\mod_ro_31.fabric[7] ),
    .A(\mod_ro_31.fabric[6] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[7].inv  (.Y(\mod_ro_31.fabric[8] ),
    .A(\mod_ro_31.fabric[7] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[8].inv  (.Y(\mod_ro_31.fabric[9] ),
    .A(\mod_ro_31.fabric[8] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[9].inv  (.Y(\mod_ro_31.fabric[10] ),
    .A(\mod_ro_31.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_1.feedback  (.Y(\mod_ro_32_1.fabric[0] ),
    .A(\mod_ro_32_1.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[0].inv  (.Y(\mod_ro_32_1.fabric[1] ),
    .A(\mod_ro_32_1.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[10].inv  (.Y(\mod_ro_32_1.fabric[11] ),
    .A(\mod_ro_32_1.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[11].inv  (.Y(\mod_ro_32_1.fabric[12] ),
    .A(\mod_ro_32_1.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[12].inv  (.Y(\mod_ro_32_1.fabric[13] ),
    .A(\mod_ro_32_1.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[13].inv  (.Y(\mod_ro_32_1.fabric[14] ),
    .A(\mod_ro_32_1.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[14].inv  (.Y(\mod_ro_32_1.fabric[15] ),
    .A(\mod_ro_32_1.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[15].inv  (.Y(\mod_ro_32_1.fabric[16] ),
    .A(\mod_ro_32_1.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[16].inv  (.Y(\mod_ro_32_1.fabric[17] ),
    .A(\mod_ro_32_1.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[17].inv  (.Y(\mod_ro_32_1.fabric[18] ),
    .A(\mod_ro_32_1.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[18].inv  (.Y(\mod_ro_32_1.fabric[19] ),
    .A(\mod_ro_32_1.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[19].inv  (.Y(\mod_ro_32_1.fabric[20] ),
    .A(\mod_ro_32_1.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[1].inv  (.Y(\mod_ro_32_1.fabric[2] ),
    .A(\mod_ro_32_1.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[20].inv  (.Y(\mod_ro_32_1.fabric[21] ),
    .A(\mod_ro_32_1.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[21].inv  (.Y(\mod_ro_32_1.fabric[22] ),
    .A(\mod_ro_32_1.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[22].inv  (.Y(\mod_ro_32_1.fabric[23] ),
    .A(\mod_ro_32_1.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[23].inv  (.Y(\mod_ro_32_1.fabric[24] ),
    .A(\mod_ro_32_1.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[24].inv  (.Y(\mod_ro_32_1.fabric[25] ),
    .A(\mod_ro_32_1.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[25].inv  (.Y(\mod_ro_32_1.fabric[26] ),
    .A(\mod_ro_32_1.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[26].inv  (.Y(\mod_ro_32_1.fabric[27] ),
    .A(\mod_ro_32_1.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[27].inv  (.Y(\mod_ro_32_1.fabric[28] ),
    .A(\mod_ro_32_1.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[28].inv  (.Y(\mod_ro_32_1.fabric[29] ),
    .A(\mod_ro_32_1.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[29].inv  (.Y(\mod_ro_32_1.fabric[30] ),
    .A(\mod_ro_32_1.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[2].inv  (.Y(\mod_ro_32_1.fabric[3] ),
    .A(\mod_ro_32_1.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[30].inv  (.Y(\mod_ro_32_1.fabric[31] ),
    .A(\mod_ro_32_1.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[31].inv  (.Y(\mod_ro_32_1.fabric[32] ),
    .A(\mod_ro_32_1.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[3].inv  (.Y(\mod_ro_32_1.fabric[4] ),
    .A(\mod_ro_32_1.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[4].inv  (.Y(\mod_ro_32_1.fabric[5] ),
    .A(\mod_ro_32_1.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[5].inv  (.Y(\mod_ro_32_1.fabric[6] ),
    .A(\mod_ro_32_1.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[6].inv  (.Y(\mod_ro_32_1.fabric[7] ),
    .A(\mod_ro_32_1.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[7].inv  (.Y(\mod_ro_32_1.fabric[8] ),
    .A(\mod_ro_32_1.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[8].inv  (.Y(\mod_ro_32_1.fabric[9] ),
    .A(\mod_ro_32_1.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[9].inv  (.Y(\mod_ro_32_1.fabric[10] ),
    .A(\mod_ro_32_1.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_2.feedback  (.Y(\mod_ro_32_2.fabric[0] ),
    .A(\mod_ro_32_2.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[0].inv  (.Y(\mod_ro_32_2.fabric[1] ),
    .A(\mod_ro_32_2.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[10].inv  (.Y(\mod_ro_32_2.fabric[11] ),
    .A(\mod_ro_32_2.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[11].inv  (.Y(\mod_ro_32_2.fabric[12] ),
    .A(\mod_ro_32_2.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[12].inv  (.Y(\mod_ro_32_2.fabric[13] ),
    .A(\mod_ro_32_2.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[13].inv  (.Y(\mod_ro_32_2.fabric[14] ),
    .A(\mod_ro_32_2.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[14].inv  (.Y(\mod_ro_32_2.fabric[15] ),
    .A(\mod_ro_32_2.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[15].inv  (.Y(\mod_ro_32_2.fabric[16] ),
    .A(\mod_ro_32_2.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[16].inv  (.Y(\mod_ro_32_2.fabric[17] ),
    .A(\mod_ro_32_2.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[17].inv  (.Y(\mod_ro_32_2.fabric[18] ),
    .A(\mod_ro_32_2.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[18].inv  (.Y(\mod_ro_32_2.fabric[19] ),
    .A(\mod_ro_32_2.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[19].inv  (.Y(\mod_ro_32_2.fabric[20] ),
    .A(\mod_ro_32_2.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[1].inv  (.Y(\mod_ro_32_2.fabric[2] ),
    .A(\mod_ro_32_2.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[20].inv  (.Y(\mod_ro_32_2.fabric[21] ),
    .A(\mod_ro_32_2.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[21].inv  (.Y(\mod_ro_32_2.fabric[22] ),
    .A(\mod_ro_32_2.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[22].inv  (.Y(\mod_ro_32_2.fabric[23] ),
    .A(\mod_ro_32_2.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[23].inv  (.Y(\mod_ro_32_2.fabric[24] ),
    .A(\mod_ro_32_2.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[24].inv  (.Y(\mod_ro_32_2.fabric[25] ),
    .A(\mod_ro_32_2.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[25].inv  (.Y(\mod_ro_32_2.fabric[26] ),
    .A(\mod_ro_32_2.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[26].inv  (.Y(\mod_ro_32_2.fabric[27] ),
    .A(\mod_ro_32_2.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[27].inv  (.Y(\mod_ro_32_2.fabric[28] ),
    .A(\mod_ro_32_2.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[28].inv  (.Y(\mod_ro_32_2.fabric[29] ),
    .A(\mod_ro_32_2.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[29].inv  (.Y(\mod_ro_32_2.fabric[30] ),
    .A(\mod_ro_32_2.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[2].inv  (.Y(\mod_ro_32_2.fabric[3] ),
    .A(\mod_ro_32_2.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[30].inv  (.Y(\mod_ro_32_2.fabric[31] ),
    .A(\mod_ro_32_2.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[31].inv  (.Y(\mod_ro_32_2.fabric[32] ),
    .A(\mod_ro_32_2.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[3].inv  (.Y(\mod_ro_32_2.fabric[4] ),
    .A(\mod_ro_32_2.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[4].inv  (.Y(\mod_ro_32_2.fabric[5] ),
    .A(\mod_ro_32_2.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[5].inv  (.Y(\mod_ro_32_2.fabric[6] ),
    .A(\mod_ro_32_2.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[6].inv  (.Y(\mod_ro_32_2.fabric[7] ),
    .A(\mod_ro_32_2.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[7].inv  (.Y(\mod_ro_32_2.fabric[8] ),
    .A(\mod_ro_32_2.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[8].inv  (.Y(\mod_ro_32_2.fabric[9] ),
    .A(\mod_ro_32_2.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[9].inv  (.Y(\mod_ro_32_2.fabric[10] ),
    .A(\mod_ro_32_2.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_raw.feedback  (.Y(\mod_ro_32_raw.fabric[0] ),
    .A(\mod_ro_32_raw.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[0].inv  (.Y(\mod_ro_32_raw.fabric[1] ),
    .A(\mod_ro_32_raw.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[10].inv  (.Y(\mod_ro_32_raw.fabric[11] ),
    .A(\mod_ro_32_raw.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[11].inv  (.Y(\mod_ro_32_raw.fabric[12] ),
    .A(\mod_ro_32_raw.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[12].inv  (.Y(\mod_ro_32_raw.fabric[13] ),
    .A(\mod_ro_32_raw.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[13].inv  (.Y(\mod_ro_32_raw.fabric[14] ),
    .A(\mod_ro_32_raw.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[14].inv  (.Y(\mod_ro_32_raw.fabric[15] ),
    .A(\mod_ro_32_raw.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[15].inv  (.Y(\mod_ro_32_raw.fabric[16] ),
    .A(\mod_ro_32_raw.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[16].inv  (.Y(\mod_ro_32_raw.fabric[17] ),
    .A(\mod_ro_32_raw.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[17].inv  (.Y(\mod_ro_32_raw.fabric[18] ),
    .A(\mod_ro_32_raw.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[18].inv  (.Y(\mod_ro_32_raw.fabric[19] ),
    .A(\mod_ro_32_raw.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[19].inv  (.Y(\mod_ro_32_raw.fabric[20] ),
    .A(\mod_ro_32_raw.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[1].inv  (.Y(\mod_ro_32_raw.fabric[2] ),
    .A(\mod_ro_32_raw.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[20].inv  (.Y(\mod_ro_32_raw.fabric[21] ),
    .A(\mod_ro_32_raw.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[21].inv  (.Y(\mod_ro_32_raw.fabric[22] ),
    .A(\mod_ro_32_raw.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[22].inv  (.Y(\mod_ro_32_raw.fabric[23] ),
    .A(\mod_ro_32_raw.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[23].inv  (.Y(\mod_ro_32_raw.fabric[24] ),
    .A(\mod_ro_32_raw.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[24].inv  (.Y(\mod_ro_32_raw.fabric[25] ),
    .A(\mod_ro_32_raw.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[25].inv  (.Y(\mod_ro_32_raw.fabric[26] ),
    .A(\mod_ro_32_raw.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[26].inv  (.Y(\mod_ro_32_raw.fabric[27] ),
    .A(\mod_ro_32_raw.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[27].inv  (.Y(\mod_ro_32_raw.fabric[28] ),
    .A(\mod_ro_32_raw.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[28].inv  (.Y(\mod_ro_32_raw.fabric[29] ),
    .A(\mod_ro_32_raw.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[29].inv  (.Y(\mod_ro_32_raw.fabric[30] ),
    .A(\mod_ro_32_raw.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[2].inv  (.Y(\mod_ro_32_raw.fabric[3] ),
    .A(\mod_ro_32_raw.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[30].inv  (.Y(\mod_ro_32_raw.fabric[31] ),
    .A(\mod_ro_32_raw.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[31].inv  (.Y(\mod_ro_32_raw.fabric[32] ),
    .A(\mod_ro_32_raw.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[3].inv  (.Y(\mod_ro_32_raw.fabric[4] ),
    .A(\mod_ro_32_raw.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[4].inv  (.Y(\mod_ro_32_raw.fabric[5] ),
    .A(\mod_ro_32_raw.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[5].inv  (.Y(\mod_ro_32_raw.fabric[6] ),
    .A(\mod_ro_32_raw.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[6].inv  (.Y(\mod_ro_32_raw.fabric[7] ),
    .A(\mod_ro_32_raw.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[7].inv  (.Y(\mod_ro_32_raw.fabric[8] ),
    .A(\mod_ro_32_raw.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[8].inv  (.Y(\mod_ro_32_raw.fabric[9] ),
    .A(\mod_ro_32_raw.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[9].inv  (.Y(\mod_ro_32_raw.fabric[10] ),
    .A(\mod_ro_32_raw.fabric[9] ));
 sg13g2_inv_1 \mod_ro_64.feedback  (.Y(\mod_ro_64.fabric[0] ),
    .A(\mod_ro_64.fabric[64] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[0].inv  (.Y(\mod_ro_64.fabric[1] ),
    .A(\mod_ro_64.fabric[0] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[10].inv  (.Y(\mod_ro_64.fabric[11] ),
    .A(\mod_ro_64.fabric[10] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[11].inv  (.Y(\mod_ro_64.fabric[12] ),
    .A(\mod_ro_64.fabric[11] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[12].inv  (.Y(\mod_ro_64.fabric[13] ),
    .A(\mod_ro_64.fabric[12] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[13].inv  (.Y(\mod_ro_64.fabric[14] ),
    .A(\mod_ro_64.fabric[13] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[14].inv  (.Y(\mod_ro_64.fabric[15] ),
    .A(\mod_ro_64.fabric[14] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[15].inv  (.Y(\mod_ro_64.fabric[16] ),
    .A(\mod_ro_64.fabric[15] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[16].inv  (.Y(\mod_ro_64.fabric[17] ),
    .A(\mod_ro_64.fabric[16] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[17].inv  (.Y(\mod_ro_64.fabric[18] ),
    .A(\mod_ro_64.fabric[17] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[18].inv  (.Y(\mod_ro_64.fabric[19] ),
    .A(\mod_ro_64.fabric[18] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[19].inv  (.Y(\mod_ro_64.fabric[20] ),
    .A(\mod_ro_64.fabric[19] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[1].inv  (.Y(\mod_ro_64.fabric[2] ),
    .A(\mod_ro_64.fabric[1] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[20].inv  (.Y(\mod_ro_64.fabric[21] ),
    .A(\mod_ro_64.fabric[20] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[21].inv  (.Y(\mod_ro_64.fabric[22] ),
    .A(\mod_ro_64.fabric[21] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[22].inv  (.Y(\mod_ro_64.fabric[23] ),
    .A(\mod_ro_64.fabric[22] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[23].inv  (.Y(\mod_ro_64.fabric[24] ),
    .A(\mod_ro_64.fabric[23] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[24].inv  (.Y(\mod_ro_64.fabric[25] ),
    .A(\mod_ro_64.fabric[24] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[25].inv  (.Y(\mod_ro_64.fabric[26] ),
    .A(\mod_ro_64.fabric[25] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[26].inv  (.Y(\mod_ro_64.fabric[27] ),
    .A(\mod_ro_64.fabric[26] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[27].inv  (.Y(\mod_ro_64.fabric[28] ),
    .A(\mod_ro_64.fabric[27] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[28].inv  (.Y(\mod_ro_64.fabric[29] ),
    .A(\mod_ro_64.fabric[28] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[29].inv  (.Y(\mod_ro_64.fabric[30] ),
    .A(\mod_ro_64.fabric[29] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[2].inv  (.Y(\mod_ro_64.fabric[3] ),
    .A(\mod_ro_64.fabric[2] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[30].inv  (.Y(\mod_ro_64.fabric[31] ),
    .A(\mod_ro_64.fabric[30] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[31].inv  (.Y(\mod_ro_64.fabric[32] ),
    .A(\mod_ro_64.fabric[31] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[32].inv  (.Y(\mod_ro_64.fabric[33] ),
    .A(\mod_ro_64.fabric[32] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[33].inv  (.Y(\mod_ro_64.fabric[34] ),
    .A(\mod_ro_64.fabric[33] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[34].inv  (.Y(\mod_ro_64.fabric[35] ),
    .A(\mod_ro_64.fabric[34] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[35].inv  (.Y(\mod_ro_64.fabric[36] ),
    .A(\mod_ro_64.fabric[35] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[36].inv  (.Y(\mod_ro_64.fabric[37] ),
    .A(\mod_ro_64.fabric[36] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[37].inv  (.Y(\mod_ro_64.fabric[38] ),
    .A(\mod_ro_64.fabric[37] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[38].inv  (.Y(\mod_ro_64.fabric[39] ),
    .A(\mod_ro_64.fabric[38] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[39].inv  (.Y(\mod_ro_64.fabric[40] ),
    .A(\mod_ro_64.fabric[39] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[3].inv  (.Y(\mod_ro_64.fabric[4] ),
    .A(\mod_ro_64.fabric[3] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[40].inv  (.Y(\mod_ro_64.fabric[41] ),
    .A(\mod_ro_64.fabric[40] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[41].inv  (.Y(\mod_ro_64.fabric[42] ),
    .A(\mod_ro_64.fabric[41] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[42].inv  (.Y(\mod_ro_64.fabric[43] ),
    .A(\mod_ro_64.fabric[42] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[43].inv  (.Y(\mod_ro_64.fabric[44] ),
    .A(\mod_ro_64.fabric[43] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[44].inv  (.Y(\mod_ro_64.fabric[45] ),
    .A(\mod_ro_64.fabric[44] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[45].inv  (.Y(\mod_ro_64.fabric[46] ),
    .A(\mod_ro_64.fabric[45] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[46].inv  (.Y(\mod_ro_64.fabric[47] ),
    .A(\mod_ro_64.fabric[46] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[47].inv  (.Y(\mod_ro_64.fabric[48] ),
    .A(\mod_ro_64.fabric[47] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[48].inv  (.Y(\mod_ro_64.fabric[49] ),
    .A(\mod_ro_64.fabric[48] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[49].inv  (.Y(\mod_ro_64.fabric[50] ),
    .A(\mod_ro_64.fabric[49] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[4].inv  (.Y(\mod_ro_64.fabric[5] ),
    .A(\mod_ro_64.fabric[4] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[50].inv  (.Y(\mod_ro_64.fabric[51] ),
    .A(\mod_ro_64.fabric[50] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[51].inv  (.Y(\mod_ro_64.fabric[52] ),
    .A(\mod_ro_64.fabric[51] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[52].inv  (.Y(\mod_ro_64.fabric[53] ),
    .A(\mod_ro_64.fabric[52] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[53].inv  (.Y(\mod_ro_64.fabric[54] ),
    .A(\mod_ro_64.fabric[53] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[54].inv  (.Y(\mod_ro_64.fabric[55] ),
    .A(\mod_ro_64.fabric[54] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[55].inv  (.Y(\mod_ro_64.fabric[56] ),
    .A(\mod_ro_64.fabric[55] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[56].inv  (.Y(\mod_ro_64.fabric[57] ),
    .A(\mod_ro_64.fabric[56] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[57].inv  (.Y(\mod_ro_64.fabric[58] ),
    .A(\mod_ro_64.fabric[57] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[58].inv  (.Y(\mod_ro_64.fabric[59] ),
    .A(\mod_ro_64.fabric[58] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[59].inv  (.Y(\mod_ro_64.fabric[60] ),
    .A(\mod_ro_64.fabric[59] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[5].inv  (.Y(\mod_ro_64.fabric[6] ),
    .A(\mod_ro_64.fabric[5] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[60].inv  (.Y(\mod_ro_64.fabric[61] ),
    .A(\mod_ro_64.fabric[60] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[61].inv  (.Y(\mod_ro_64.fabric[62] ),
    .A(\mod_ro_64.fabric[61] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[62].inv  (.Y(\mod_ro_64.fabric[63] ),
    .A(\mod_ro_64.fabric[62] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[63].inv  (.Y(\mod_ro_64.fabric[64] ),
    .A(\mod_ro_64.fabric[63] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[6].inv  (.Y(\mod_ro_64.fabric[7] ),
    .A(\mod_ro_64.fabric[6] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[7].inv  (.Y(\mod_ro_64.fabric[8] ),
    .A(\mod_ro_64.fabric[7] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[8].inv  (.Y(\mod_ro_64.fabric[9] ),
    .A(\mod_ro_64.fabric[8] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[9].inv  (.Y(\mod_ro_64.fabric[10] ),
    .A(\mod_ro_64.fabric[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_tielo tt_um_wedgetail_tester_4 (.L_LO(net4));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_4 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_4 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_4 FILLER_28_385 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_4 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_29_379 ();
 sg13g2_decap_4 FILLER_29_393 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_decap_4 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_4 FILLER_31_273 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_decap_4 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_390 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_4 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_4 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_368 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_decap_4 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_4 FILLER_34_385 ();
 sg13g2_fill_1 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_decap_8 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_decap_4 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_decap_8 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_321 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_373 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_4 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_fill_1 FILLER_36_367 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_decap_4 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_4 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_decap_4 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_2 FILLER_38_320 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_fill_2 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule
