module tt_um_corey (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire \byte_cnt[0] ;
 wire \byte_cnt[1] ;
 wire \byte_cnt[2] ;
 wire \byte_cnt[3] ;
 wire \byte_cnt[4] ;
 wire inv_done;
 wire inv_go;
 wire \inv_result[0] ;
 wire \inv_result[100] ;
 wire \inv_result[101] ;
 wire \inv_result[102] ;
 wire \inv_result[103] ;
 wire \inv_result[104] ;
 wire \inv_result[105] ;
 wire \inv_result[106] ;
 wire \inv_result[107] ;
 wire \inv_result[108] ;
 wire \inv_result[109] ;
 wire \inv_result[10] ;
 wire \inv_result[110] ;
 wire \inv_result[111] ;
 wire \inv_result[112] ;
 wire \inv_result[113] ;
 wire \inv_result[114] ;
 wire \inv_result[115] ;
 wire \inv_result[116] ;
 wire \inv_result[117] ;
 wire \inv_result[118] ;
 wire \inv_result[119] ;
 wire \inv_result[11] ;
 wire \inv_result[120] ;
 wire \inv_result[121] ;
 wire \inv_result[122] ;
 wire \inv_result[123] ;
 wire \inv_result[124] ;
 wire \inv_result[125] ;
 wire \inv_result[126] ;
 wire \inv_result[127] ;
 wire \inv_result[128] ;
 wire \inv_result[129] ;
 wire \inv_result[12] ;
 wire \inv_result[130] ;
 wire \inv_result[131] ;
 wire \inv_result[132] ;
 wire \inv_result[133] ;
 wire \inv_result[134] ;
 wire \inv_result[135] ;
 wire \inv_result[136] ;
 wire \inv_result[137] ;
 wire \inv_result[138] ;
 wire \inv_result[139] ;
 wire \inv_result[13] ;
 wire \inv_result[140] ;
 wire \inv_result[141] ;
 wire \inv_result[142] ;
 wire \inv_result[143] ;
 wire \inv_result[144] ;
 wire \inv_result[145] ;
 wire \inv_result[146] ;
 wire \inv_result[147] ;
 wire \inv_result[148] ;
 wire \inv_result[149] ;
 wire \inv_result[14] ;
 wire \inv_result[150] ;
 wire \inv_result[151] ;
 wire \inv_result[152] ;
 wire \inv_result[153] ;
 wire \inv_result[154] ;
 wire \inv_result[155] ;
 wire \inv_result[156] ;
 wire \inv_result[157] ;
 wire \inv_result[158] ;
 wire \inv_result[159] ;
 wire \inv_result[15] ;
 wire \inv_result[160] ;
 wire \inv_result[161] ;
 wire \inv_result[162] ;
 wire \inv_result[163] ;
 wire \inv_result[164] ;
 wire \inv_result[165] ;
 wire \inv_result[166] ;
 wire \inv_result[167] ;
 wire \inv_result[168] ;
 wire \inv_result[169] ;
 wire \inv_result[16] ;
 wire \inv_result[170] ;
 wire \inv_result[171] ;
 wire \inv_result[172] ;
 wire \inv_result[173] ;
 wire \inv_result[174] ;
 wire \inv_result[175] ;
 wire \inv_result[176] ;
 wire \inv_result[177] ;
 wire \inv_result[178] ;
 wire \inv_result[179] ;
 wire \inv_result[17] ;
 wire \inv_result[180] ;
 wire \inv_result[181] ;
 wire \inv_result[182] ;
 wire \inv_result[183] ;
 wire \inv_result[184] ;
 wire \inv_result[185] ;
 wire \inv_result[186] ;
 wire \inv_result[187] ;
 wire \inv_result[188] ;
 wire \inv_result[189] ;
 wire \inv_result[18] ;
 wire \inv_result[190] ;
 wire \inv_result[191] ;
 wire \inv_result[192] ;
 wire \inv_result[193] ;
 wire \inv_result[194] ;
 wire \inv_result[195] ;
 wire \inv_result[196] ;
 wire \inv_result[197] ;
 wire \inv_result[198] ;
 wire \inv_result[199] ;
 wire \inv_result[19] ;
 wire \inv_result[1] ;
 wire \inv_result[200] ;
 wire \inv_result[201] ;
 wire \inv_result[202] ;
 wire \inv_result[203] ;
 wire \inv_result[204] ;
 wire \inv_result[205] ;
 wire \inv_result[206] ;
 wire \inv_result[207] ;
 wire \inv_result[208] ;
 wire \inv_result[209] ;
 wire \inv_result[20] ;
 wire \inv_result[210] ;
 wire \inv_result[211] ;
 wire \inv_result[212] ;
 wire \inv_result[213] ;
 wire \inv_result[214] ;
 wire \inv_result[215] ;
 wire \inv_result[216] ;
 wire \inv_result[217] ;
 wire \inv_result[218] ;
 wire \inv_result[219] ;
 wire \inv_result[21] ;
 wire \inv_result[220] ;
 wire \inv_result[221] ;
 wire \inv_result[222] ;
 wire \inv_result[223] ;
 wire \inv_result[224] ;
 wire \inv_result[225] ;
 wire \inv_result[226] ;
 wire \inv_result[227] ;
 wire \inv_result[228] ;
 wire \inv_result[229] ;
 wire \inv_result[22] ;
 wire \inv_result[230] ;
 wire \inv_result[231] ;
 wire \inv_result[232] ;
 wire \inv_result[233] ;
 wire \inv_result[234] ;
 wire \inv_result[235] ;
 wire \inv_result[236] ;
 wire \inv_result[237] ;
 wire \inv_result[238] ;
 wire \inv_result[239] ;
 wire \inv_result[23] ;
 wire \inv_result[240] ;
 wire \inv_result[241] ;
 wire \inv_result[242] ;
 wire \inv_result[243] ;
 wire \inv_result[244] ;
 wire \inv_result[245] ;
 wire \inv_result[246] ;
 wire \inv_result[247] ;
 wire \inv_result[248] ;
 wire \inv_result[249] ;
 wire \inv_result[24] ;
 wire \inv_result[250] ;
 wire \inv_result[251] ;
 wire \inv_result[252] ;
 wire \inv_result[253] ;
 wire \inv_result[254] ;
 wire \inv_result[255] ;
 wire \inv_result[25] ;
 wire \inv_result[26] ;
 wire \inv_result[27] ;
 wire \inv_result[28] ;
 wire \inv_result[29] ;
 wire \inv_result[2] ;
 wire \inv_result[30] ;
 wire \inv_result[31] ;
 wire \inv_result[32] ;
 wire \inv_result[33] ;
 wire \inv_result[34] ;
 wire \inv_result[35] ;
 wire \inv_result[36] ;
 wire \inv_result[37] ;
 wire \inv_result[38] ;
 wire \inv_result[39] ;
 wire \inv_result[3] ;
 wire \inv_result[40] ;
 wire \inv_result[41] ;
 wire \inv_result[42] ;
 wire \inv_result[43] ;
 wire \inv_result[44] ;
 wire \inv_result[45] ;
 wire \inv_result[46] ;
 wire \inv_result[47] ;
 wire \inv_result[48] ;
 wire \inv_result[49] ;
 wire \inv_result[4] ;
 wire \inv_result[50] ;
 wire \inv_result[51] ;
 wire \inv_result[52] ;
 wire \inv_result[53] ;
 wire \inv_result[54] ;
 wire \inv_result[55] ;
 wire \inv_result[56] ;
 wire \inv_result[57] ;
 wire \inv_result[58] ;
 wire \inv_result[59] ;
 wire \inv_result[5] ;
 wire \inv_result[60] ;
 wire \inv_result[61] ;
 wire \inv_result[62] ;
 wire \inv_result[63] ;
 wire \inv_result[64] ;
 wire \inv_result[65] ;
 wire \inv_result[66] ;
 wire \inv_result[67] ;
 wire \inv_result[68] ;
 wire \inv_result[69] ;
 wire \inv_result[6] ;
 wire \inv_result[70] ;
 wire \inv_result[71] ;
 wire \inv_result[72] ;
 wire \inv_result[73] ;
 wire \inv_result[74] ;
 wire \inv_result[75] ;
 wire \inv_result[76] ;
 wire \inv_result[77] ;
 wire \inv_result[78] ;
 wire \inv_result[79] ;
 wire \inv_result[7] ;
 wire \inv_result[80] ;
 wire \inv_result[81] ;
 wire \inv_result[82] ;
 wire \inv_result[83] ;
 wire \inv_result[84] ;
 wire \inv_result[85] ;
 wire \inv_result[86] ;
 wire \inv_result[87] ;
 wire \inv_result[88] ;
 wire \inv_result[89] ;
 wire \inv_result[8] ;
 wire \inv_result[90] ;
 wire \inv_result[91] ;
 wire \inv_result[92] ;
 wire \inv_result[93] ;
 wire \inv_result[94] ;
 wire \inv_result[95] ;
 wire \inv_result[96] ;
 wire \inv_result[97] ;
 wire \inv_result[98] ;
 wire \inv_result[99] ;
 wire \inv_result[9] ;
 wire rd_prev;
 wire \shift_reg[0] ;
 wire \shift_reg[100] ;
 wire \shift_reg[101] ;
 wire \shift_reg[102] ;
 wire \shift_reg[103] ;
 wire \shift_reg[104] ;
 wire \shift_reg[105] ;
 wire \shift_reg[106] ;
 wire \shift_reg[107] ;
 wire \shift_reg[108] ;
 wire \shift_reg[109] ;
 wire \shift_reg[10] ;
 wire \shift_reg[110] ;
 wire \shift_reg[111] ;
 wire \shift_reg[112] ;
 wire \shift_reg[113] ;
 wire \shift_reg[114] ;
 wire \shift_reg[115] ;
 wire \shift_reg[116] ;
 wire \shift_reg[117] ;
 wire \shift_reg[118] ;
 wire \shift_reg[119] ;
 wire \shift_reg[11] ;
 wire \shift_reg[120] ;
 wire \shift_reg[121] ;
 wire \shift_reg[122] ;
 wire \shift_reg[123] ;
 wire \shift_reg[124] ;
 wire \shift_reg[125] ;
 wire \shift_reg[126] ;
 wire \shift_reg[127] ;
 wire \shift_reg[128] ;
 wire \shift_reg[129] ;
 wire \shift_reg[12] ;
 wire \shift_reg[130] ;
 wire \shift_reg[131] ;
 wire \shift_reg[132] ;
 wire \shift_reg[133] ;
 wire \shift_reg[134] ;
 wire \shift_reg[135] ;
 wire \shift_reg[136] ;
 wire \shift_reg[137] ;
 wire \shift_reg[138] ;
 wire \shift_reg[139] ;
 wire \shift_reg[13] ;
 wire \shift_reg[140] ;
 wire \shift_reg[141] ;
 wire \shift_reg[142] ;
 wire \shift_reg[143] ;
 wire \shift_reg[144] ;
 wire \shift_reg[145] ;
 wire \shift_reg[146] ;
 wire \shift_reg[147] ;
 wire \shift_reg[148] ;
 wire \shift_reg[149] ;
 wire \shift_reg[14] ;
 wire \shift_reg[150] ;
 wire \shift_reg[151] ;
 wire \shift_reg[152] ;
 wire \shift_reg[153] ;
 wire \shift_reg[154] ;
 wire \shift_reg[155] ;
 wire \shift_reg[156] ;
 wire \shift_reg[157] ;
 wire \shift_reg[158] ;
 wire \shift_reg[159] ;
 wire \shift_reg[15] ;
 wire \shift_reg[160] ;
 wire \shift_reg[161] ;
 wire \shift_reg[162] ;
 wire \shift_reg[163] ;
 wire \shift_reg[164] ;
 wire \shift_reg[165] ;
 wire \shift_reg[166] ;
 wire \shift_reg[167] ;
 wire \shift_reg[168] ;
 wire \shift_reg[169] ;
 wire \shift_reg[16] ;
 wire \shift_reg[170] ;
 wire \shift_reg[171] ;
 wire \shift_reg[172] ;
 wire \shift_reg[173] ;
 wire \shift_reg[174] ;
 wire \shift_reg[175] ;
 wire \shift_reg[176] ;
 wire \shift_reg[177] ;
 wire \shift_reg[178] ;
 wire \shift_reg[179] ;
 wire \shift_reg[17] ;
 wire \shift_reg[180] ;
 wire \shift_reg[181] ;
 wire \shift_reg[182] ;
 wire \shift_reg[183] ;
 wire \shift_reg[184] ;
 wire \shift_reg[185] ;
 wire \shift_reg[186] ;
 wire \shift_reg[187] ;
 wire \shift_reg[188] ;
 wire \shift_reg[189] ;
 wire \shift_reg[18] ;
 wire \shift_reg[190] ;
 wire \shift_reg[191] ;
 wire \shift_reg[192] ;
 wire \shift_reg[193] ;
 wire \shift_reg[194] ;
 wire \shift_reg[195] ;
 wire \shift_reg[196] ;
 wire \shift_reg[197] ;
 wire \shift_reg[198] ;
 wire \shift_reg[199] ;
 wire \shift_reg[19] ;
 wire \shift_reg[1] ;
 wire \shift_reg[200] ;
 wire \shift_reg[201] ;
 wire \shift_reg[202] ;
 wire \shift_reg[203] ;
 wire \shift_reg[204] ;
 wire \shift_reg[205] ;
 wire \shift_reg[206] ;
 wire \shift_reg[207] ;
 wire \shift_reg[208] ;
 wire \shift_reg[209] ;
 wire \shift_reg[20] ;
 wire \shift_reg[210] ;
 wire \shift_reg[211] ;
 wire \shift_reg[212] ;
 wire \shift_reg[213] ;
 wire \shift_reg[214] ;
 wire \shift_reg[215] ;
 wire \shift_reg[216] ;
 wire \shift_reg[217] ;
 wire \shift_reg[218] ;
 wire \shift_reg[219] ;
 wire \shift_reg[21] ;
 wire \shift_reg[220] ;
 wire \shift_reg[221] ;
 wire \shift_reg[222] ;
 wire \shift_reg[223] ;
 wire \shift_reg[224] ;
 wire \shift_reg[225] ;
 wire \shift_reg[226] ;
 wire \shift_reg[227] ;
 wire \shift_reg[228] ;
 wire \shift_reg[229] ;
 wire \shift_reg[22] ;
 wire \shift_reg[230] ;
 wire \shift_reg[231] ;
 wire \shift_reg[232] ;
 wire \shift_reg[233] ;
 wire \shift_reg[234] ;
 wire \shift_reg[235] ;
 wire \shift_reg[236] ;
 wire \shift_reg[237] ;
 wire \shift_reg[238] ;
 wire \shift_reg[239] ;
 wire \shift_reg[23] ;
 wire \shift_reg[240] ;
 wire \shift_reg[241] ;
 wire \shift_reg[242] ;
 wire \shift_reg[243] ;
 wire \shift_reg[244] ;
 wire \shift_reg[245] ;
 wire \shift_reg[246] ;
 wire \shift_reg[247] ;
 wire \shift_reg[248] ;
 wire \shift_reg[249] ;
 wire \shift_reg[24] ;
 wire \shift_reg[250] ;
 wire \shift_reg[251] ;
 wire \shift_reg[252] ;
 wire \shift_reg[253] ;
 wire \shift_reg[254] ;
 wire \shift_reg[255] ;
 wire \shift_reg[25] ;
 wire \shift_reg[26] ;
 wire \shift_reg[27] ;
 wire \shift_reg[28] ;
 wire \shift_reg[29] ;
 wire \shift_reg[2] ;
 wire \shift_reg[30] ;
 wire \shift_reg[31] ;
 wire \shift_reg[32] ;
 wire \shift_reg[33] ;
 wire \shift_reg[34] ;
 wire \shift_reg[35] ;
 wire \shift_reg[36] ;
 wire \shift_reg[37] ;
 wire \shift_reg[38] ;
 wire \shift_reg[39] ;
 wire \shift_reg[3] ;
 wire \shift_reg[40] ;
 wire \shift_reg[41] ;
 wire \shift_reg[42] ;
 wire \shift_reg[43] ;
 wire \shift_reg[44] ;
 wire \shift_reg[45] ;
 wire \shift_reg[46] ;
 wire \shift_reg[47] ;
 wire \shift_reg[48] ;
 wire \shift_reg[49] ;
 wire \shift_reg[4] ;
 wire \shift_reg[50] ;
 wire \shift_reg[51] ;
 wire \shift_reg[52] ;
 wire \shift_reg[53] ;
 wire \shift_reg[54] ;
 wire \shift_reg[55] ;
 wire \shift_reg[56] ;
 wire \shift_reg[57] ;
 wire \shift_reg[58] ;
 wire \shift_reg[59] ;
 wire \shift_reg[5] ;
 wire \shift_reg[60] ;
 wire \shift_reg[61] ;
 wire \shift_reg[62] ;
 wire \shift_reg[63] ;
 wire \shift_reg[64] ;
 wire \shift_reg[65] ;
 wire \shift_reg[66] ;
 wire \shift_reg[67] ;
 wire \shift_reg[68] ;
 wire \shift_reg[69] ;
 wire \shift_reg[6] ;
 wire \shift_reg[70] ;
 wire \shift_reg[71] ;
 wire \shift_reg[72] ;
 wire \shift_reg[73] ;
 wire \shift_reg[74] ;
 wire \shift_reg[75] ;
 wire \shift_reg[76] ;
 wire \shift_reg[77] ;
 wire \shift_reg[78] ;
 wire \shift_reg[79] ;
 wire \shift_reg[7] ;
 wire \shift_reg[80] ;
 wire \shift_reg[81] ;
 wire \shift_reg[82] ;
 wire \shift_reg[83] ;
 wire \shift_reg[84] ;
 wire \shift_reg[85] ;
 wire \shift_reg[86] ;
 wire \shift_reg[87] ;
 wire \shift_reg[88] ;
 wire \shift_reg[89] ;
 wire \shift_reg[8] ;
 wire \shift_reg[90] ;
 wire \shift_reg[91] ;
 wire \shift_reg[92] ;
 wire \shift_reg[93] ;
 wire \shift_reg[94] ;
 wire \shift_reg[95] ;
 wire \shift_reg[96] ;
 wire \shift_reg[97] ;
 wire \shift_reg[98] ;
 wire \shift_reg[99] ;
 wire \shift_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \u_inv.counter[0] ;
 wire \u_inv.counter[1] ;
 wire \u_inv.counter[2] ;
 wire \u_inv.counter[3] ;
 wire \u_inv.counter[4] ;
 wire \u_inv.counter[5] ;
 wire \u_inv.counter[6] ;
 wire \u_inv.counter[7] ;
 wire \u_inv.counter[8] ;
 wire \u_inv.counter[9] ;
 wire \u_inv.d_next[0] ;
 wire \u_inv.d_next[100] ;
 wire \u_inv.d_next[101] ;
 wire \u_inv.d_next[102] ;
 wire \u_inv.d_next[103] ;
 wire \u_inv.d_next[104] ;
 wire \u_inv.d_next[105] ;
 wire \u_inv.d_next[106] ;
 wire \u_inv.d_next[107] ;
 wire \u_inv.d_next[108] ;
 wire \u_inv.d_next[109] ;
 wire \u_inv.d_next[10] ;
 wire \u_inv.d_next[110] ;
 wire \u_inv.d_next[111] ;
 wire \u_inv.d_next[112] ;
 wire \u_inv.d_next[113] ;
 wire \u_inv.d_next[114] ;
 wire \u_inv.d_next[115] ;
 wire \u_inv.d_next[116] ;
 wire \u_inv.d_next[117] ;
 wire \u_inv.d_next[118] ;
 wire \u_inv.d_next[119] ;
 wire \u_inv.d_next[11] ;
 wire \u_inv.d_next[120] ;
 wire \u_inv.d_next[121] ;
 wire \u_inv.d_next[122] ;
 wire \u_inv.d_next[123] ;
 wire \u_inv.d_next[124] ;
 wire \u_inv.d_next[125] ;
 wire \u_inv.d_next[126] ;
 wire \u_inv.d_next[127] ;
 wire \u_inv.d_next[128] ;
 wire \u_inv.d_next[129] ;
 wire \u_inv.d_next[12] ;
 wire \u_inv.d_next[130] ;
 wire \u_inv.d_next[131] ;
 wire \u_inv.d_next[132] ;
 wire \u_inv.d_next[133] ;
 wire \u_inv.d_next[134] ;
 wire \u_inv.d_next[135] ;
 wire \u_inv.d_next[136] ;
 wire \u_inv.d_next[137] ;
 wire \u_inv.d_next[138] ;
 wire \u_inv.d_next[139] ;
 wire \u_inv.d_next[13] ;
 wire \u_inv.d_next[140] ;
 wire \u_inv.d_next[141] ;
 wire \u_inv.d_next[142] ;
 wire \u_inv.d_next[143] ;
 wire \u_inv.d_next[144] ;
 wire \u_inv.d_next[145] ;
 wire \u_inv.d_next[146] ;
 wire \u_inv.d_next[147] ;
 wire \u_inv.d_next[148] ;
 wire \u_inv.d_next[149] ;
 wire \u_inv.d_next[14] ;
 wire \u_inv.d_next[150] ;
 wire \u_inv.d_next[151] ;
 wire \u_inv.d_next[152] ;
 wire \u_inv.d_next[153] ;
 wire \u_inv.d_next[154] ;
 wire \u_inv.d_next[155] ;
 wire \u_inv.d_next[156] ;
 wire \u_inv.d_next[157] ;
 wire \u_inv.d_next[158] ;
 wire \u_inv.d_next[159] ;
 wire \u_inv.d_next[15] ;
 wire \u_inv.d_next[160] ;
 wire \u_inv.d_next[161] ;
 wire \u_inv.d_next[162] ;
 wire \u_inv.d_next[163] ;
 wire \u_inv.d_next[164] ;
 wire \u_inv.d_next[165] ;
 wire \u_inv.d_next[166] ;
 wire \u_inv.d_next[167] ;
 wire \u_inv.d_next[168] ;
 wire \u_inv.d_next[169] ;
 wire \u_inv.d_next[16] ;
 wire \u_inv.d_next[170] ;
 wire \u_inv.d_next[171] ;
 wire \u_inv.d_next[172] ;
 wire \u_inv.d_next[173] ;
 wire \u_inv.d_next[174] ;
 wire \u_inv.d_next[175] ;
 wire \u_inv.d_next[176] ;
 wire \u_inv.d_next[177] ;
 wire \u_inv.d_next[178] ;
 wire \u_inv.d_next[179] ;
 wire \u_inv.d_next[17] ;
 wire \u_inv.d_next[180] ;
 wire \u_inv.d_next[181] ;
 wire \u_inv.d_next[182] ;
 wire \u_inv.d_next[183] ;
 wire \u_inv.d_next[184] ;
 wire \u_inv.d_next[185] ;
 wire \u_inv.d_next[186] ;
 wire \u_inv.d_next[187] ;
 wire \u_inv.d_next[188] ;
 wire \u_inv.d_next[189] ;
 wire \u_inv.d_next[18] ;
 wire \u_inv.d_next[190] ;
 wire \u_inv.d_next[191] ;
 wire \u_inv.d_next[192] ;
 wire \u_inv.d_next[193] ;
 wire \u_inv.d_next[194] ;
 wire \u_inv.d_next[195] ;
 wire \u_inv.d_next[196] ;
 wire \u_inv.d_next[197] ;
 wire \u_inv.d_next[198] ;
 wire \u_inv.d_next[199] ;
 wire \u_inv.d_next[19] ;
 wire \u_inv.d_next[1] ;
 wire \u_inv.d_next[200] ;
 wire \u_inv.d_next[201] ;
 wire \u_inv.d_next[202] ;
 wire \u_inv.d_next[203] ;
 wire \u_inv.d_next[204] ;
 wire \u_inv.d_next[205] ;
 wire \u_inv.d_next[206] ;
 wire \u_inv.d_next[207] ;
 wire \u_inv.d_next[208] ;
 wire \u_inv.d_next[209] ;
 wire \u_inv.d_next[20] ;
 wire \u_inv.d_next[210] ;
 wire \u_inv.d_next[211] ;
 wire \u_inv.d_next[212] ;
 wire \u_inv.d_next[213] ;
 wire \u_inv.d_next[214] ;
 wire \u_inv.d_next[215] ;
 wire \u_inv.d_next[216] ;
 wire \u_inv.d_next[217] ;
 wire \u_inv.d_next[218] ;
 wire \u_inv.d_next[219] ;
 wire \u_inv.d_next[21] ;
 wire \u_inv.d_next[220] ;
 wire \u_inv.d_next[221] ;
 wire \u_inv.d_next[222] ;
 wire \u_inv.d_next[223] ;
 wire \u_inv.d_next[224] ;
 wire \u_inv.d_next[225] ;
 wire \u_inv.d_next[226] ;
 wire \u_inv.d_next[227] ;
 wire \u_inv.d_next[228] ;
 wire \u_inv.d_next[229] ;
 wire \u_inv.d_next[22] ;
 wire \u_inv.d_next[230] ;
 wire \u_inv.d_next[231] ;
 wire \u_inv.d_next[232] ;
 wire \u_inv.d_next[233] ;
 wire \u_inv.d_next[234] ;
 wire \u_inv.d_next[235] ;
 wire \u_inv.d_next[236] ;
 wire \u_inv.d_next[237] ;
 wire \u_inv.d_next[238] ;
 wire \u_inv.d_next[239] ;
 wire \u_inv.d_next[23] ;
 wire \u_inv.d_next[240] ;
 wire \u_inv.d_next[241] ;
 wire \u_inv.d_next[242] ;
 wire \u_inv.d_next[243] ;
 wire \u_inv.d_next[244] ;
 wire \u_inv.d_next[245] ;
 wire \u_inv.d_next[246] ;
 wire \u_inv.d_next[247] ;
 wire \u_inv.d_next[248] ;
 wire \u_inv.d_next[249] ;
 wire \u_inv.d_next[24] ;
 wire \u_inv.d_next[250] ;
 wire \u_inv.d_next[251] ;
 wire \u_inv.d_next[252] ;
 wire \u_inv.d_next[253] ;
 wire \u_inv.d_next[254] ;
 wire \u_inv.d_next[255] ;
 wire \u_inv.d_next[256] ;
 wire \u_inv.d_next[25] ;
 wire \u_inv.d_next[26] ;
 wire \u_inv.d_next[27] ;
 wire \u_inv.d_next[28] ;
 wire \u_inv.d_next[29] ;
 wire \u_inv.d_next[2] ;
 wire \u_inv.d_next[30] ;
 wire \u_inv.d_next[31] ;
 wire \u_inv.d_next[32] ;
 wire \u_inv.d_next[33] ;
 wire \u_inv.d_next[34] ;
 wire \u_inv.d_next[35] ;
 wire \u_inv.d_next[36] ;
 wire \u_inv.d_next[37] ;
 wire \u_inv.d_next[38] ;
 wire \u_inv.d_next[39] ;
 wire \u_inv.d_next[3] ;
 wire \u_inv.d_next[40] ;
 wire \u_inv.d_next[41] ;
 wire \u_inv.d_next[42] ;
 wire \u_inv.d_next[43] ;
 wire \u_inv.d_next[44] ;
 wire \u_inv.d_next[45] ;
 wire \u_inv.d_next[46] ;
 wire \u_inv.d_next[47] ;
 wire \u_inv.d_next[48] ;
 wire \u_inv.d_next[49] ;
 wire \u_inv.d_next[4] ;
 wire \u_inv.d_next[50] ;
 wire \u_inv.d_next[51] ;
 wire \u_inv.d_next[52] ;
 wire \u_inv.d_next[53] ;
 wire \u_inv.d_next[54] ;
 wire \u_inv.d_next[55] ;
 wire \u_inv.d_next[56] ;
 wire \u_inv.d_next[57] ;
 wire \u_inv.d_next[58] ;
 wire \u_inv.d_next[59] ;
 wire \u_inv.d_next[5] ;
 wire \u_inv.d_next[60] ;
 wire \u_inv.d_next[61] ;
 wire \u_inv.d_next[62] ;
 wire \u_inv.d_next[63] ;
 wire \u_inv.d_next[64] ;
 wire \u_inv.d_next[65] ;
 wire \u_inv.d_next[66] ;
 wire \u_inv.d_next[67] ;
 wire \u_inv.d_next[68] ;
 wire \u_inv.d_next[69] ;
 wire \u_inv.d_next[6] ;
 wire \u_inv.d_next[70] ;
 wire \u_inv.d_next[71] ;
 wire \u_inv.d_next[72] ;
 wire \u_inv.d_next[73] ;
 wire \u_inv.d_next[74] ;
 wire \u_inv.d_next[75] ;
 wire \u_inv.d_next[76] ;
 wire \u_inv.d_next[77] ;
 wire \u_inv.d_next[78] ;
 wire \u_inv.d_next[79] ;
 wire \u_inv.d_next[7] ;
 wire \u_inv.d_next[80] ;
 wire \u_inv.d_next[81] ;
 wire \u_inv.d_next[82] ;
 wire \u_inv.d_next[83] ;
 wire \u_inv.d_next[84] ;
 wire \u_inv.d_next[85] ;
 wire \u_inv.d_next[86] ;
 wire \u_inv.d_next[87] ;
 wire \u_inv.d_next[88] ;
 wire \u_inv.d_next[89] ;
 wire \u_inv.d_next[8] ;
 wire \u_inv.d_next[90] ;
 wire \u_inv.d_next[91] ;
 wire \u_inv.d_next[92] ;
 wire \u_inv.d_next[93] ;
 wire \u_inv.d_next[94] ;
 wire \u_inv.d_next[95] ;
 wire \u_inv.d_next[96] ;
 wire \u_inv.d_next[97] ;
 wire \u_inv.d_next[98] ;
 wire \u_inv.d_next[99] ;
 wire \u_inv.d_next[9] ;
 wire \u_inv.d_reg[0] ;
 wire \u_inv.d_reg[100] ;
 wire \u_inv.d_reg[101] ;
 wire \u_inv.d_reg[102] ;
 wire \u_inv.d_reg[103] ;
 wire \u_inv.d_reg[104] ;
 wire \u_inv.d_reg[105] ;
 wire \u_inv.d_reg[106] ;
 wire \u_inv.d_reg[107] ;
 wire \u_inv.d_reg[108] ;
 wire \u_inv.d_reg[109] ;
 wire \u_inv.d_reg[10] ;
 wire \u_inv.d_reg[110] ;
 wire \u_inv.d_reg[111] ;
 wire \u_inv.d_reg[112] ;
 wire \u_inv.d_reg[113] ;
 wire \u_inv.d_reg[114] ;
 wire \u_inv.d_reg[115] ;
 wire \u_inv.d_reg[116] ;
 wire \u_inv.d_reg[117] ;
 wire \u_inv.d_reg[118] ;
 wire \u_inv.d_reg[119] ;
 wire \u_inv.d_reg[11] ;
 wire \u_inv.d_reg[120] ;
 wire \u_inv.d_reg[121] ;
 wire \u_inv.d_reg[122] ;
 wire \u_inv.d_reg[123] ;
 wire \u_inv.d_reg[124] ;
 wire \u_inv.d_reg[125] ;
 wire \u_inv.d_reg[126] ;
 wire \u_inv.d_reg[127] ;
 wire \u_inv.d_reg[128] ;
 wire \u_inv.d_reg[129] ;
 wire \u_inv.d_reg[12] ;
 wire \u_inv.d_reg[130] ;
 wire \u_inv.d_reg[131] ;
 wire \u_inv.d_reg[132] ;
 wire \u_inv.d_reg[133] ;
 wire \u_inv.d_reg[134] ;
 wire \u_inv.d_reg[135] ;
 wire \u_inv.d_reg[136] ;
 wire \u_inv.d_reg[137] ;
 wire \u_inv.d_reg[138] ;
 wire \u_inv.d_reg[139] ;
 wire \u_inv.d_reg[13] ;
 wire \u_inv.d_reg[140] ;
 wire \u_inv.d_reg[141] ;
 wire \u_inv.d_reg[142] ;
 wire \u_inv.d_reg[143] ;
 wire \u_inv.d_reg[144] ;
 wire \u_inv.d_reg[145] ;
 wire \u_inv.d_reg[146] ;
 wire \u_inv.d_reg[147] ;
 wire \u_inv.d_reg[148] ;
 wire \u_inv.d_reg[149] ;
 wire \u_inv.d_reg[14] ;
 wire \u_inv.d_reg[150] ;
 wire \u_inv.d_reg[151] ;
 wire \u_inv.d_reg[152] ;
 wire \u_inv.d_reg[153] ;
 wire \u_inv.d_reg[154] ;
 wire \u_inv.d_reg[155] ;
 wire \u_inv.d_reg[156] ;
 wire \u_inv.d_reg[157] ;
 wire \u_inv.d_reg[158] ;
 wire \u_inv.d_reg[159] ;
 wire \u_inv.d_reg[15] ;
 wire \u_inv.d_reg[160] ;
 wire \u_inv.d_reg[161] ;
 wire \u_inv.d_reg[162] ;
 wire \u_inv.d_reg[163] ;
 wire \u_inv.d_reg[164] ;
 wire \u_inv.d_reg[165] ;
 wire \u_inv.d_reg[166] ;
 wire \u_inv.d_reg[167] ;
 wire \u_inv.d_reg[168] ;
 wire \u_inv.d_reg[169] ;
 wire \u_inv.d_reg[16] ;
 wire \u_inv.d_reg[170] ;
 wire \u_inv.d_reg[171] ;
 wire \u_inv.d_reg[172] ;
 wire \u_inv.d_reg[173] ;
 wire \u_inv.d_reg[174] ;
 wire \u_inv.d_reg[175] ;
 wire \u_inv.d_reg[176] ;
 wire \u_inv.d_reg[177] ;
 wire \u_inv.d_reg[178] ;
 wire \u_inv.d_reg[179] ;
 wire \u_inv.d_reg[17] ;
 wire \u_inv.d_reg[180] ;
 wire \u_inv.d_reg[181] ;
 wire \u_inv.d_reg[182] ;
 wire \u_inv.d_reg[183] ;
 wire \u_inv.d_reg[184] ;
 wire \u_inv.d_reg[185] ;
 wire \u_inv.d_reg[186] ;
 wire \u_inv.d_reg[187] ;
 wire \u_inv.d_reg[188] ;
 wire \u_inv.d_reg[189] ;
 wire \u_inv.d_reg[18] ;
 wire \u_inv.d_reg[190] ;
 wire \u_inv.d_reg[191] ;
 wire \u_inv.d_reg[192] ;
 wire \u_inv.d_reg[193] ;
 wire \u_inv.d_reg[194] ;
 wire \u_inv.d_reg[195] ;
 wire \u_inv.d_reg[196] ;
 wire \u_inv.d_reg[197] ;
 wire \u_inv.d_reg[198] ;
 wire \u_inv.d_reg[199] ;
 wire \u_inv.d_reg[19] ;
 wire \u_inv.d_reg[1] ;
 wire \u_inv.d_reg[200] ;
 wire \u_inv.d_reg[201] ;
 wire \u_inv.d_reg[202] ;
 wire \u_inv.d_reg[203] ;
 wire \u_inv.d_reg[204] ;
 wire \u_inv.d_reg[205] ;
 wire \u_inv.d_reg[206] ;
 wire \u_inv.d_reg[207] ;
 wire \u_inv.d_reg[208] ;
 wire \u_inv.d_reg[209] ;
 wire \u_inv.d_reg[20] ;
 wire \u_inv.d_reg[210] ;
 wire \u_inv.d_reg[211] ;
 wire \u_inv.d_reg[212] ;
 wire \u_inv.d_reg[213] ;
 wire \u_inv.d_reg[214] ;
 wire \u_inv.d_reg[215] ;
 wire \u_inv.d_reg[216] ;
 wire \u_inv.d_reg[217] ;
 wire \u_inv.d_reg[218] ;
 wire \u_inv.d_reg[219] ;
 wire \u_inv.d_reg[21] ;
 wire \u_inv.d_reg[220] ;
 wire \u_inv.d_reg[221] ;
 wire \u_inv.d_reg[222] ;
 wire \u_inv.d_reg[223] ;
 wire \u_inv.d_reg[224] ;
 wire \u_inv.d_reg[225] ;
 wire \u_inv.d_reg[226] ;
 wire \u_inv.d_reg[227] ;
 wire \u_inv.d_reg[228] ;
 wire \u_inv.d_reg[229] ;
 wire \u_inv.d_reg[22] ;
 wire \u_inv.d_reg[230] ;
 wire \u_inv.d_reg[231] ;
 wire \u_inv.d_reg[232] ;
 wire \u_inv.d_reg[233] ;
 wire \u_inv.d_reg[234] ;
 wire \u_inv.d_reg[235] ;
 wire \u_inv.d_reg[236] ;
 wire \u_inv.d_reg[237] ;
 wire \u_inv.d_reg[238] ;
 wire \u_inv.d_reg[239] ;
 wire \u_inv.d_reg[23] ;
 wire \u_inv.d_reg[240] ;
 wire \u_inv.d_reg[241] ;
 wire \u_inv.d_reg[242] ;
 wire \u_inv.d_reg[243] ;
 wire \u_inv.d_reg[244] ;
 wire \u_inv.d_reg[245] ;
 wire \u_inv.d_reg[246] ;
 wire \u_inv.d_reg[247] ;
 wire \u_inv.d_reg[248] ;
 wire \u_inv.d_reg[249] ;
 wire \u_inv.d_reg[24] ;
 wire \u_inv.d_reg[250] ;
 wire \u_inv.d_reg[251] ;
 wire \u_inv.d_reg[252] ;
 wire \u_inv.d_reg[253] ;
 wire \u_inv.d_reg[254] ;
 wire \u_inv.d_reg[255] ;
 wire \u_inv.d_reg[256] ;
 wire \u_inv.d_reg[25] ;
 wire \u_inv.d_reg[26] ;
 wire \u_inv.d_reg[27] ;
 wire \u_inv.d_reg[28] ;
 wire \u_inv.d_reg[29] ;
 wire \u_inv.d_reg[2] ;
 wire \u_inv.d_reg[30] ;
 wire \u_inv.d_reg[31] ;
 wire \u_inv.d_reg[32] ;
 wire \u_inv.d_reg[33] ;
 wire \u_inv.d_reg[34] ;
 wire \u_inv.d_reg[35] ;
 wire \u_inv.d_reg[36] ;
 wire \u_inv.d_reg[37] ;
 wire \u_inv.d_reg[38] ;
 wire \u_inv.d_reg[39] ;
 wire \u_inv.d_reg[3] ;
 wire \u_inv.d_reg[40] ;
 wire \u_inv.d_reg[41] ;
 wire \u_inv.d_reg[42] ;
 wire \u_inv.d_reg[43] ;
 wire \u_inv.d_reg[44] ;
 wire \u_inv.d_reg[45] ;
 wire \u_inv.d_reg[46] ;
 wire \u_inv.d_reg[47] ;
 wire \u_inv.d_reg[48] ;
 wire \u_inv.d_reg[49] ;
 wire \u_inv.d_reg[4] ;
 wire \u_inv.d_reg[50] ;
 wire \u_inv.d_reg[51] ;
 wire \u_inv.d_reg[52] ;
 wire \u_inv.d_reg[53] ;
 wire \u_inv.d_reg[54] ;
 wire \u_inv.d_reg[55] ;
 wire \u_inv.d_reg[56] ;
 wire \u_inv.d_reg[57] ;
 wire \u_inv.d_reg[58] ;
 wire \u_inv.d_reg[59] ;
 wire \u_inv.d_reg[5] ;
 wire \u_inv.d_reg[60] ;
 wire \u_inv.d_reg[61] ;
 wire \u_inv.d_reg[62] ;
 wire \u_inv.d_reg[63] ;
 wire \u_inv.d_reg[64] ;
 wire \u_inv.d_reg[65] ;
 wire \u_inv.d_reg[66] ;
 wire \u_inv.d_reg[67] ;
 wire \u_inv.d_reg[68] ;
 wire \u_inv.d_reg[69] ;
 wire \u_inv.d_reg[6] ;
 wire \u_inv.d_reg[70] ;
 wire \u_inv.d_reg[71] ;
 wire \u_inv.d_reg[72] ;
 wire \u_inv.d_reg[73] ;
 wire \u_inv.d_reg[74] ;
 wire \u_inv.d_reg[75] ;
 wire \u_inv.d_reg[76] ;
 wire \u_inv.d_reg[77] ;
 wire \u_inv.d_reg[78] ;
 wire \u_inv.d_reg[79] ;
 wire \u_inv.d_reg[7] ;
 wire \u_inv.d_reg[80] ;
 wire \u_inv.d_reg[81] ;
 wire \u_inv.d_reg[82] ;
 wire \u_inv.d_reg[83] ;
 wire \u_inv.d_reg[84] ;
 wire \u_inv.d_reg[85] ;
 wire \u_inv.d_reg[86] ;
 wire \u_inv.d_reg[87] ;
 wire \u_inv.d_reg[88] ;
 wire \u_inv.d_reg[89] ;
 wire \u_inv.d_reg[8] ;
 wire \u_inv.d_reg[90] ;
 wire \u_inv.d_reg[91] ;
 wire \u_inv.d_reg[92] ;
 wire \u_inv.d_reg[93] ;
 wire \u_inv.d_reg[94] ;
 wire \u_inv.d_reg[95] ;
 wire \u_inv.d_reg[96] ;
 wire \u_inv.d_reg[97] ;
 wire \u_inv.d_reg[98] ;
 wire \u_inv.d_reg[99] ;
 wire \u_inv.d_reg[9] ;
 wire \u_inv.delta_reg[0] ;
 wire \u_inv.delta_reg[1] ;
 wire \u_inv.delta_reg[2] ;
 wire \u_inv.delta_reg[3] ;
 wire \u_inv.delta_reg[4] ;
 wire \u_inv.delta_reg[5] ;
 wire \u_inv.delta_reg[6] ;
 wire \u_inv.delta_reg[7] ;
 wire \u_inv.delta_reg[8] ;
 wire \u_inv.delta_reg[9] ;
 wire \u_inv.f_next[0] ;
 wire \u_inv.f_next[100] ;
 wire \u_inv.f_next[101] ;
 wire \u_inv.f_next[102] ;
 wire \u_inv.f_next[103] ;
 wire \u_inv.f_next[104] ;
 wire \u_inv.f_next[105] ;
 wire \u_inv.f_next[106] ;
 wire \u_inv.f_next[107] ;
 wire \u_inv.f_next[108] ;
 wire \u_inv.f_next[109] ;
 wire \u_inv.f_next[10] ;
 wire \u_inv.f_next[110] ;
 wire \u_inv.f_next[111] ;
 wire \u_inv.f_next[112] ;
 wire \u_inv.f_next[113] ;
 wire \u_inv.f_next[114] ;
 wire \u_inv.f_next[115] ;
 wire \u_inv.f_next[116] ;
 wire \u_inv.f_next[117] ;
 wire \u_inv.f_next[118] ;
 wire \u_inv.f_next[119] ;
 wire \u_inv.f_next[11] ;
 wire \u_inv.f_next[120] ;
 wire \u_inv.f_next[121] ;
 wire \u_inv.f_next[122] ;
 wire \u_inv.f_next[123] ;
 wire \u_inv.f_next[124] ;
 wire \u_inv.f_next[125] ;
 wire \u_inv.f_next[126] ;
 wire \u_inv.f_next[127] ;
 wire \u_inv.f_next[128] ;
 wire \u_inv.f_next[129] ;
 wire \u_inv.f_next[12] ;
 wire \u_inv.f_next[130] ;
 wire \u_inv.f_next[131] ;
 wire \u_inv.f_next[132] ;
 wire \u_inv.f_next[133] ;
 wire \u_inv.f_next[134] ;
 wire \u_inv.f_next[135] ;
 wire \u_inv.f_next[136] ;
 wire \u_inv.f_next[137] ;
 wire \u_inv.f_next[138] ;
 wire \u_inv.f_next[139] ;
 wire \u_inv.f_next[13] ;
 wire \u_inv.f_next[140] ;
 wire \u_inv.f_next[141] ;
 wire \u_inv.f_next[142] ;
 wire \u_inv.f_next[143] ;
 wire \u_inv.f_next[144] ;
 wire \u_inv.f_next[145] ;
 wire \u_inv.f_next[146] ;
 wire \u_inv.f_next[147] ;
 wire \u_inv.f_next[148] ;
 wire \u_inv.f_next[149] ;
 wire \u_inv.f_next[14] ;
 wire \u_inv.f_next[150] ;
 wire \u_inv.f_next[151] ;
 wire \u_inv.f_next[152] ;
 wire \u_inv.f_next[153] ;
 wire \u_inv.f_next[154] ;
 wire \u_inv.f_next[155] ;
 wire \u_inv.f_next[156] ;
 wire \u_inv.f_next[157] ;
 wire \u_inv.f_next[158] ;
 wire \u_inv.f_next[159] ;
 wire \u_inv.f_next[15] ;
 wire \u_inv.f_next[160] ;
 wire \u_inv.f_next[161] ;
 wire \u_inv.f_next[162] ;
 wire \u_inv.f_next[163] ;
 wire \u_inv.f_next[164] ;
 wire \u_inv.f_next[165] ;
 wire \u_inv.f_next[166] ;
 wire \u_inv.f_next[167] ;
 wire \u_inv.f_next[168] ;
 wire \u_inv.f_next[169] ;
 wire \u_inv.f_next[16] ;
 wire \u_inv.f_next[170] ;
 wire \u_inv.f_next[171] ;
 wire \u_inv.f_next[172] ;
 wire \u_inv.f_next[173] ;
 wire \u_inv.f_next[174] ;
 wire \u_inv.f_next[175] ;
 wire \u_inv.f_next[176] ;
 wire \u_inv.f_next[177] ;
 wire \u_inv.f_next[178] ;
 wire \u_inv.f_next[179] ;
 wire \u_inv.f_next[17] ;
 wire \u_inv.f_next[180] ;
 wire \u_inv.f_next[181] ;
 wire \u_inv.f_next[182] ;
 wire \u_inv.f_next[183] ;
 wire \u_inv.f_next[184] ;
 wire \u_inv.f_next[185] ;
 wire \u_inv.f_next[186] ;
 wire \u_inv.f_next[187] ;
 wire \u_inv.f_next[188] ;
 wire \u_inv.f_next[189] ;
 wire \u_inv.f_next[18] ;
 wire \u_inv.f_next[190] ;
 wire \u_inv.f_next[191] ;
 wire \u_inv.f_next[192] ;
 wire \u_inv.f_next[193] ;
 wire \u_inv.f_next[194] ;
 wire \u_inv.f_next[195] ;
 wire \u_inv.f_next[196] ;
 wire \u_inv.f_next[197] ;
 wire \u_inv.f_next[198] ;
 wire \u_inv.f_next[199] ;
 wire \u_inv.f_next[19] ;
 wire \u_inv.f_next[1] ;
 wire \u_inv.f_next[200] ;
 wire \u_inv.f_next[201] ;
 wire \u_inv.f_next[202] ;
 wire \u_inv.f_next[203] ;
 wire \u_inv.f_next[204] ;
 wire \u_inv.f_next[205] ;
 wire \u_inv.f_next[206] ;
 wire \u_inv.f_next[207] ;
 wire \u_inv.f_next[208] ;
 wire \u_inv.f_next[209] ;
 wire \u_inv.f_next[20] ;
 wire \u_inv.f_next[210] ;
 wire \u_inv.f_next[211] ;
 wire \u_inv.f_next[212] ;
 wire \u_inv.f_next[213] ;
 wire \u_inv.f_next[214] ;
 wire \u_inv.f_next[215] ;
 wire \u_inv.f_next[216] ;
 wire \u_inv.f_next[217] ;
 wire \u_inv.f_next[218] ;
 wire \u_inv.f_next[219] ;
 wire \u_inv.f_next[21] ;
 wire \u_inv.f_next[220] ;
 wire \u_inv.f_next[221] ;
 wire \u_inv.f_next[222] ;
 wire \u_inv.f_next[223] ;
 wire \u_inv.f_next[224] ;
 wire \u_inv.f_next[225] ;
 wire \u_inv.f_next[226] ;
 wire \u_inv.f_next[227] ;
 wire \u_inv.f_next[228] ;
 wire \u_inv.f_next[229] ;
 wire \u_inv.f_next[22] ;
 wire \u_inv.f_next[230] ;
 wire \u_inv.f_next[231] ;
 wire \u_inv.f_next[232] ;
 wire \u_inv.f_next[233] ;
 wire \u_inv.f_next[234] ;
 wire \u_inv.f_next[235] ;
 wire \u_inv.f_next[236] ;
 wire \u_inv.f_next[237] ;
 wire \u_inv.f_next[238] ;
 wire \u_inv.f_next[239] ;
 wire \u_inv.f_next[23] ;
 wire \u_inv.f_next[240] ;
 wire \u_inv.f_next[241] ;
 wire \u_inv.f_next[242] ;
 wire \u_inv.f_next[243] ;
 wire \u_inv.f_next[244] ;
 wire \u_inv.f_next[245] ;
 wire \u_inv.f_next[246] ;
 wire \u_inv.f_next[247] ;
 wire \u_inv.f_next[248] ;
 wire \u_inv.f_next[249] ;
 wire \u_inv.f_next[24] ;
 wire \u_inv.f_next[250] ;
 wire \u_inv.f_next[251] ;
 wire \u_inv.f_next[252] ;
 wire \u_inv.f_next[253] ;
 wire \u_inv.f_next[254] ;
 wire \u_inv.f_next[255] ;
 wire \u_inv.f_next[256] ;
 wire \u_inv.f_next[25] ;
 wire \u_inv.f_next[26] ;
 wire \u_inv.f_next[27] ;
 wire \u_inv.f_next[28] ;
 wire \u_inv.f_next[29] ;
 wire \u_inv.f_next[2] ;
 wire \u_inv.f_next[30] ;
 wire \u_inv.f_next[31] ;
 wire \u_inv.f_next[32] ;
 wire \u_inv.f_next[33] ;
 wire \u_inv.f_next[34] ;
 wire \u_inv.f_next[35] ;
 wire \u_inv.f_next[36] ;
 wire \u_inv.f_next[37] ;
 wire \u_inv.f_next[38] ;
 wire \u_inv.f_next[39] ;
 wire \u_inv.f_next[3] ;
 wire \u_inv.f_next[40] ;
 wire \u_inv.f_next[41] ;
 wire \u_inv.f_next[42] ;
 wire \u_inv.f_next[43] ;
 wire \u_inv.f_next[44] ;
 wire \u_inv.f_next[45] ;
 wire \u_inv.f_next[46] ;
 wire \u_inv.f_next[47] ;
 wire \u_inv.f_next[48] ;
 wire \u_inv.f_next[49] ;
 wire \u_inv.f_next[4] ;
 wire \u_inv.f_next[50] ;
 wire \u_inv.f_next[51] ;
 wire \u_inv.f_next[52] ;
 wire \u_inv.f_next[53] ;
 wire \u_inv.f_next[54] ;
 wire \u_inv.f_next[55] ;
 wire \u_inv.f_next[56] ;
 wire \u_inv.f_next[57] ;
 wire \u_inv.f_next[58] ;
 wire \u_inv.f_next[59] ;
 wire \u_inv.f_next[5] ;
 wire \u_inv.f_next[60] ;
 wire \u_inv.f_next[61] ;
 wire \u_inv.f_next[62] ;
 wire \u_inv.f_next[63] ;
 wire \u_inv.f_next[64] ;
 wire \u_inv.f_next[65] ;
 wire \u_inv.f_next[66] ;
 wire \u_inv.f_next[67] ;
 wire \u_inv.f_next[68] ;
 wire \u_inv.f_next[69] ;
 wire \u_inv.f_next[6] ;
 wire \u_inv.f_next[70] ;
 wire \u_inv.f_next[71] ;
 wire \u_inv.f_next[72] ;
 wire \u_inv.f_next[73] ;
 wire \u_inv.f_next[74] ;
 wire \u_inv.f_next[75] ;
 wire \u_inv.f_next[76] ;
 wire \u_inv.f_next[77] ;
 wire \u_inv.f_next[78] ;
 wire \u_inv.f_next[79] ;
 wire \u_inv.f_next[7] ;
 wire \u_inv.f_next[80] ;
 wire \u_inv.f_next[81] ;
 wire \u_inv.f_next[82] ;
 wire \u_inv.f_next[83] ;
 wire \u_inv.f_next[84] ;
 wire \u_inv.f_next[85] ;
 wire \u_inv.f_next[86] ;
 wire \u_inv.f_next[87] ;
 wire \u_inv.f_next[88] ;
 wire \u_inv.f_next[89] ;
 wire \u_inv.f_next[8] ;
 wire \u_inv.f_next[90] ;
 wire \u_inv.f_next[91] ;
 wire \u_inv.f_next[92] ;
 wire \u_inv.f_next[93] ;
 wire \u_inv.f_next[94] ;
 wire \u_inv.f_next[95] ;
 wire \u_inv.f_next[96] ;
 wire \u_inv.f_next[97] ;
 wire \u_inv.f_next[98] ;
 wire \u_inv.f_next[99] ;
 wire \u_inv.f_next[9] ;
 wire \u_inv.f_reg[0] ;
 wire \u_inv.f_reg[100] ;
 wire \u_inv.f_reg[101] ;
 wire \u_inv.f_reg[102] ;
 wire \u_inv.f_reg[103] ;
 wire \u_inv.f_reg[104] ;
 wire \u_inv.f_reg[105] ;
 wire \u_inv.f_reg[106] ;
 wire \u_inv.f_reg[107] ;
 wire \u_inv.f_reg[108] ;
 wire \u_inv.f_reg[109] ;
 wire \u_inv.f_reg[10] ;
 wire \u_inv.f_reg[110] ;
 wire \u_inv.f_reg[111] ;
 wire \u_inv.f_reg[112] ;
 wire \u_inv.f_reg[113] ;
 wire \u_inv.f_reg[114] ;
 wire \u_inv.f_reg[115] ;
 wire \u_inv.f_reg[116] ;
 wire \u_inv.f_reg[117] ;
 wire \u_inv.f_reg[118] ;
 wire \u_inv.f_reg[119] ;
 wire \u_inv.f_reg[11] ;
 wire \u_inv.f_reg[120] ;
 wire \u_inv.f_reg[121] ;
 wire \u_inv.f_reg[122] ;
 wire \u_inv.f_reg[123] ;
 wire \u_inv.f_reg[124] ;
 wire \u_inv.f_reg[125] ;
 wire \u_inv.f_reg[126] ;
 wire \u_inv.f_reg[127] ;
 wire \u_inv.f_reg[128] ;
 wire \u_inv.f_reg[129] ;
 wire \u_inv.f_reg[12] ;
 wire \u_inv.f_reg[130] ;
 wire \u_inv.f_reg[131] ;
 wire \u_inv.f_reg[132] ;
 wire \u_inv.f_reg[133] ;
 wire \u_inv.f_reg[134] ;
 wire \u_inv.f_reg[135] ;
 wire \u_inv.f_reg[136] ;
 wire \u_inv.f_reg[137] ;
 wire \u_inv.f_reg[138] ;
 wire \u_inv.f_reg[139] ;
 wire \u_inv.f_reg[13] ;
 wire \u_inv.f_reg[140] ;
 wire \u_inv.f_reg[141] ;
 wire \u_inv.f_reg[142] ;
 wire \u_inv.f_reg[143] ;
 wire \u_inv.f_reg[144] ;
 wire \u_inv.f_reg[145] ;
 wire \u_inv.f_reg[146] ;
 wire \u_inv.f_reg[147] ;
 wire \u_inv.f_reg[148] ;
 wire \u_inv.f_reg[149] ;
 wire \u_inv.f_reg[14] ;
 wire \u_inv.f_reg[150] ;
 wire \u_inv.f_reg[151] ;
 wire \u_inv.f_reg[152] ;
 wire \u_inv.f_reg[153] ;
 wire \u_inv.f_reg[154] ;
 wire \u_inv.f_reg[155] ;
 wire \u_inv.f_reg[156] ;
 wire \u_inv.f_reg[157] ;
 wire \u_inv.f_reg[158] ;
 wire \u_inv.f_reg[159] ;
 wire \u_inv.f_reg[15] ;
 wire \u_inv.f_reg[160] ;
 wire \u_inv.f_reg[161] ;
 wire \u_inv.f_reg[162] ;
 wire \u_inv.f_reg[163] ;
 wire \u_inv.f_reg[164] ;
 wire \u_inv.f_reg[165] ;
 wire \u_inv.f_reg[166] ;
 wire \u_inv.f_reg[167] ;
 wire \u_inv.f_reg[168] ;
 wire \u_inv.f_reg[169] ;
 wire \u_inv.f_reg[16] ;
 wire \u_inv.f_reg[170] ;
 wire \u_inv.f_reg[171] ;
 wire \u_inv.f_reg[172] ;
 wire \u_inv.f_reg[173] ;
 wire \u_inv.f_reg[174] ;
 wire \u_inv.f_reg[175] ;
 wire \u_inv.f_reg[176] ;
 wire \u_inv.f_reg[177] ;
 wire \u_inv.f_reg[178] ;
 wire \u_inv.f_reg[179] ;
 wire \u_inv.f_reg[17] ;
 wire \u_inv.f_reg[180] ;
 wire \u_inv.f_reg[181] ;
 wire \u_inv.f_reg[182] ;
 wire \u_inv.f_reg[183] ;
 wire \u_inv.f_reg[184] ;
 wire \u_inv.f_reg[185] ;
 wire \u_inv.f_reg[186] ;
 wire \u_inv.f_reg[187] ;
 wire \u_inv.f_reg[188] ;
 wire \u_inv.f_reg[189] ;
 wire \u_inv.f_reg[18] ;
 wire \u_inv.f_reg[190] ;
 wire \u_inv.f_reg[191] ;
 wire \u_inv.f_reg[192] ;
 wire \u_inv.f_reg[193] ;
 wire \u_inv.f_reg[194] ;
 wire \u_inv.f_reg[195] ;
 wire \u_inv.f_reg[196] ;
 wire \u_inv.f_reg[197] ;
 wire \u_inv.f_reg[198] ;
 wire \u_inv.f_reg[199] ;
 wire \u_inv.f_reg[19] ;
 wire \u_inv.f_reg[1] ;
 wire \u_inv.f_reg[200] ;
 wire \u_inv.f_reg[201] ;
 wire \u_inv.f_reg[202] ;
 wire \u_inv.f_reg[203] ;
 wire \u_inv.f_reg[204] ;
 wire \u_inv.f_reg[205] ;
 wire \u_inv.f_reg[206] ;
 wire \u_inv.f_reg[207] ;
 wire \u_inv.f_reg[208] ;
 wire \u_inv.f_reg[209] ;
 wire \u_inv.f_reg[20] ;
 wire \u_inv.f_reg[210] ;
 wire \u_inv.f_reg[211] ;
 wire \u_inv.f_reg[212] ;
 wire \u_inv.f_reg[213] ;
 wire \u_inv.f_reg[214] ;
 wire \u_inv.f_reg[215] ;
 wire \u_inv.f_reg[216] ;
 wire \u_inv.f_reg[217] ;
 wire \u_inv.f_reg[218] ;
 wire \u_inv.f_reg[219] ;
 wire \u_inv.f_reg[21] ;
 wire \u_inv.f_reg[220] ;
 wire \u_inv.f_reg[221] ;
 wire \u_inv.f_reg[222] ;
 wire \u_inv.f_reg[223] ;
 wire \u_inv.f_reg[224] ;
 wire \u_inv.f_reg[225] ;
 wire \u_inv.f_reg[226] ;
 wire \u_inv.f_reg[227] ;
 wire \u_inv.f_reg[228] ;
 wire \u_inv.f_reg[229] ;
 wire \u_inv.f_reg[22] ;
 wire \u_inv.f_reg[230] ;
 wire \u_inv.f_reg[231] ;
 wire \u_inv.f_reg[232] ;
 wire \u_inv.f_reg[233] ;
 wire \u_inv.f_reg[234] ;
 wire \u_inv.f_reg[235] ;
 wire \u_inv.f_reg[236] ;
 wire \u_inv.f_reg[237] ;
 wire \u_inv.f_reg[238] ;
 wire \u_inv.f_reg[239] ;
 wire \u_inv.f_reg[23] ;
 wire \u_inv.f_reg[240] ;
 wire \u_inv.f_reg[241] ;
 wire \u_inv.f_reg[242] ;
 wire \u_inv.f_reg[243] ;
 wire \u_inv.f_reg[244] ;
 wire \u_inv.f_reg[245] ;
 wire \u_inv.f_reg[246] ;
 wire \u_inv.f_reg[247] ;
 wire \u_inv.f_reg[248] ;
 wire \u_inv.f_reg[249] ;
 wire \u_inv.f_reg[24] ;
 wire \u_inv.f_reg[250] ;
 wire \u_inv.f_reg[251] ;
 wire \u_inv.f_reg[252] ;
 wire \u_inv.f_reg[253] ;
 wire \u_inv.f_reg[254] ;
 wire \u_inv.f_reg[255] ;
 wire \u_inv.f_reg[256] ;
 wire \u_inv.f_reg[25] ;
 wire \u_inv.f_reg[26] ;
 wire \u_inv.f_reg[27] ;
 wire \u_inv.f_reg[28] ;
 wire \u_inv.f_reg[29] ;
 wire \u_inv.f_reg[2] ;
 wire \u_inv.f_reg[30] ;
 wire \u_inv.f_reg[31] ;
 wire \u_inv.f_reg[32] ;
 wire \u_inv.f_reg[33] ;
 wire \u_inv.f_reg[34] ;
 wire \u_inv.f_reg[35] ;
 wire \u_inv.f_reg[36] ;
 wire \u_inv.f_reg[37] ;
 wire \u_inv.f_reg[38] ;
 wire \u_inv.f_reg[39] ;
 wire \u_inv.f_reg[3] ;
 wire \u_inv.f_reg[40] ;
 wire \u_inv.f_reg[41] ;
 wire \u_inv.f_reg[42] ;
 wire \u_inv.f_reg[43] ;
 wire \u_inv.f_reg[44] ;
 wire \u_inv.f_reg[45] ;
 wire \u_inv.f_reg[46] ;
 wire \u_inv.f_reg[47] ;
 wire \u_inv.f_reg[48] ;
 wire \u_inv.f_reg[49] ;
 wire \u_inv.f_reg[4] ;
 wire \u_inv.f_reg[50] ;
 wire \u_inv.f_reg[51] ;
 wire \u_inv.f_reg[52] ;
 wire \u_inv.f_reg[53] ;
 wire \u_inv.f_reg[54] ;
 wire \u_inv.f_reg[55] ;
 wire \u_inv.f_reg[56] ;
 wire \u_inv.f_reg[57] ;
 wire \u_inv.f_reg[58] ;
 wire \u_inv.f_reg[59] ;
 wire \u_inv.f_reg[5] ;
 wire \u_inv.f_reg[60] ;
 wire \u_inv.f_reg[61] ;
 wire \u_inv.f_reg[62] ;
 wire \u_inv.f_reg[63] ;
 wire \u_inv.f_reg[64] ;
 wire \u_inv.f_reg[65] ;
 wire \u_inv.f_reg[66] ;
 wire \u_inv.f_reg[67] ;
 wire \u_inv.f_reg[68] ;
 wire \u_inv.f_reg[69] ;
 wire \u_inv.f_reg[6] ;
 wire \u_inv.f_reg[70] ;
 wire \u_inv.f_reg[71] ;
 wire \u_inv.f_reg[72] ;
 wire \u_inv.f_reg[73] ;
 wire \u_inv.f_reg[74] ;
 wire \u_inv.f_reg[75] ;
 wire \u_inv.f_reg[76] ;
 wire \u_inv.f_reg[77] ;
 wire \u_inv.f_reg[78] ;
 wire \u_inv.f_reg[79] ;
 wire \u_inv.f_reg[7] ;
 wire \u_inv.f_reg[80] ;
 wire \u_inv.f_reg[81] ;
 wire \u_inv.f_reg[82] ;
 wire \u_inv.f_reg[83] ;
 wire \u_inv.f_reg[84] ;
 wire \u_inv.f_reg[85] ;
 wire \u_inv.f_reg[86] ;
 wire \u_inv.f_reg[87] ;
 wire \u_inv.f_reg[88] ;
 wire \u_inv.f_reg[89] ;
 wire \u_inv.f_reg[8] ;
 wire \u_inv.f_reg[90] ;
 wire \u_inv.f_reg[91] ;
 wire \u_inv.f_reg[92] ;
 wire \u_inv.f_reg[93] ;
 wire \u_inv.f_reg[94] ;
 wire \u_inv.f_reg[95] ;
 wire \u_inv.f_reg[96] ;
 wire \u_inv.f_reg[97] ;
 wire \u_inv.f_reg[98] ;
 wire \u_inv.f_reg[99] ;
 wire \u_inv.f_reg[9] ;
 wire \u_inv.input_reg[0] ;
 wire \u_inv.input_reg[100] ;
 wire \u_inv.input_reg[101] ;
 wire \u_inv.input_reg[102] ;
 wire \u_inv.input_reg[103] ;
 wire \u_inv.input_reg[104] ;
 wire \u_inv.input_reg[105] ;
 wire \u_inv.input_reg[106] ;
 wire \u_inv.input_reg[107] ;
 wire \u_inv.input_reg[108] ;
 wire \u_inv.input_reg[109] ;
 wire \u_inv.input_reg[10] ;
 wire \u_inv.input_reg[110] ;
 wire \u_inv.input_reg[111] ;
 wire \u_inv.input_reg[112] ;
 wire \u_inv.input_reg[113] ;
 wire \u_inv.input_reg[114] ;
 wire \u_inv.input_reg[115] ;
 wire \u_inv.input_reg[116] ;
 wire \u_inv.input_reg[117] ;
 wire \u_inv.input_reg[118] ;
 wire \u_inv.input_reg[119] ;
 wire \u_inv.input_reg[11] ;
 wire \u_inv.input_reg[120] ;
 wire \u_inv.input_reg[121] ;
 wire \u_inv.input_reg[122] ;
 wire \u_inv.input_reg[123] ;
 wire \u_inv.input_reg[124] ;
 wire \u_inv.input_reg[125] ;
 wire \u_inv.input_reg[126] ;
 wire \u_inv.input_reg[127] ;
 wire \u_inv.input_reg[128] ;
 wire \u_inv.input_reg[129] ;
 wire \u_inv.input_reg[12] ;
 wire \u_inv.input_reg[130] ;
 wire \u_inv.input_reg[131] ;
 wire \u_inv.input_reg[132] ;
 wire \u_inv.input_reg[133] ;
 wire \u_inv.input_reg[134] ;
 wire \u_inv.input_reg[135] ;
 wire \u_inv.input_reg[136] ;
 wire \u_inv.input_reg[137] ;
 wire \u_inv.input_reg[138] ;
 wire \u_inv.input_reg[139] ;
 wire \u_inv.input_reg[13] ;
 wire \u_inv.input_reg[140] ;
 wire \u_inv.input_reg[141] ;
 wire \u_inv.input_reg[142] ;
 wire \u_inv.input_reg[143] ;
 wire \u_inv.input_reg[144] ;
 wire \u_inv.input_reg[145] ;
 wire \u_inv.input_reg[146] ;
 wire \u_inv.input_reg[147] ;
 wire \u_inv.input_reg[148] ;
 wire \u_inv.input_reg[149] ;
 wire \u_inv.input_reg[14] ;
 wire \u_inv.input_reg[150] ;
 wire \u_inv.input_reg[151] ;
 wire \u_inv.input_reg[152] ;
 wire \u_inv.input_reg[153] ;
 wire \u_inv.input_reg[154] ;
 wire \u_inv.input_reg[155] ;
 wire \u_inv.input_reg[156] ;
 wire \u_inv.input_reg[157] ;
 wire \u_inv.input_reg[158] ;
 wire \u_inv.input_reg[159] ;
 wire \u_inv.input_reg[15] ;
 wire \u_inv.input_reg[160] ;
 wire \u_inv.input_reg[161] ;
 wire \u_inv.input_reg[162] ;
 wire \u_inv.input_reg[163] ;
 wire \u_inv.input_reg[164] ;
 wire \u_inv.input_reg[165] ;
 wire \u_inv.input_reg[166] ;
 wire \u_inv.input_reg[167] ;
 wire \u_inv.input_reg[168] ;
 wire \u_inv.input_reg[169] ;
 wire \u_inv.input_reg[16] ;
 wire \u_inv.input_reg[170] ;
 wire \u_inv.input_reg[171] ;
 wire \u_inv.input_reg[172] ;
 wire \u_inv.input_reg[173] ;
 wire \u_inv.input_reg[174] ;
 wire \u_inv.input_reg[175] ;
 wire \u_inv.input_reg[176] ;
 wire \u_inv.input_reg[177] ;
 wire \u_inv.input_reg[178] ;
 wire \u_inv.input_reg[179] ;
 wire \u_inv.input_reg[17] ;
 wire \u_inv.input_reg[180] ;
 wire \u_inv.input_reg[181] ;
 wire \u_inv.input_reg[182] ;
 wire \u_inv.input_reg[183] ;
 wire \u_inv.input_reg[184] ;
 wire \u_inv.input_reg[185] ;
 wire \u_inv.input_reg[186] ;
 wire \u_inv.input_reg[187] ;
 wire \u_inv.input_reg[188] ;
 wire \u_inv.input_reg[189] ;
 wire \u_inv.input_reg[18] ;
 wire \u_inv.input_reg[190] ;
 wire \u_inv.input_reg[191] ;
 wire \u_inv.input_reg[192] ;
 wire \u_inv.input_reg[193] ;
 wire \u_inv.input_reg[194] ;
 wire \u_inv.input_reg[195] ;
 wire \u_inv.input_reg[196] ;
 wire \u_inv.input_reg[197] ;
 wire \u_inv.input_reg[198] ;
 wire \u_inv.input_reg[199] ;
 wire \u_inv.input_reg[19] ;
 wire \u_inv.input_reg[1] ;
 wire \u_inv.input_reg[200] ;
 wire \u_inv.input_reg[201] ;
 wire \u_inv.input_reg[202] ;
 wire \u_inv.input_reg[203] ;
 wire \u_inv.input_reg[204] ;
 wire \u_inv.input_reg[205] ;
 wire \u_inv.input_reg[206] ;
 wire \u_inv.input_reg[207] ;
 wire \u_inv.input_reg[208] ;
 wire \u_inv.input_reg[209] ;
 wire \u_inv.input_reg[20] ;
 wire \u_inv.input_reg[210] ;
 wire \u_inv.input_reg[211] ;
 wire \u_inv.input_reg[212] ;
 wire \u_inv.input_reg[213] ;
 wire \u_inv.input_reg[214] ;
 wire \u_inv.input_reg[215] ;
 wire \u_inv.input_reg[216] ;
 wire \u_inv.input_reg[217] ;
 wire \u_inv.input_reg[218] ;
 wire \u_inv.input_reg[219] ;
 wire \u_inv.input_reg[21] ;
 wire \u_inv.input_reg[220] ;
 wire \u_inv.input_reg[221] ;
 wire \u_inv.input_reg[222] ;
 wire \u_inv.input_reg[223] ;
 wire \u_inv.input_reg[224] ;
 wire \u_inv.input_reg[225] ;
 wire \u_inv.input_reg[226] ;
 wire \u_inv.input_reg[227] ;
 wire \u_inv.input_reg[228] ;
 wire \u_inv.input_reg[229] ;
 wire \u_inv.input_reg[22] ;
 wire \u_inv.input_reg[230] ;
 wire \u_inv.input_reg[231] ;
 wire \u_inv.input_reg[232] ;
 wire \u_inv.input_reg[233] ;
 wire \u_inv.input_reg[234] ;
 wire \u_inv.input_reg[235] ;
 wire \u_inv.input_reg[236] ;
 wire \u_inv.input_reg[237] ;
 wire \u_inv.input_reg[238] ;
 wire \u_inv.input_reg[239] ;
 wire \u_inv.input_reg[23] ;
 wire \u_inv.input_reg[240] ;
 wire \u_inv.input_reg[241] ;
 wire \u_inv.input_reg[242] ;
 wire \u_inv.input_reg[243] ;
 wire \u_inv.input_reg[244] ;
 wire \u_inv.input_reg[245] ;
 wire \u_inv.input_reg[246] ;
 wire \u_inv.input_reg[247] ;
 wire \u_inv.input_reg[248] ;
 wire \u_inv.input_reg[249] ;
 wire \u_inv.input_reg[24] ;
 wire \u_inv.input_reg[250] ;
 wire \u_inv.input_reg[251] ;
 wire \u_inv.input_reg[252] ;
 wire \u_inv.input_reg[253] ;
 wire \u_inv.input_reg[254] ;
 wire \u_inv.input_reg[255] ;
 wire \u_inv.input_reg[25] ;
 wire \u_inv.input_reg[26] ;
 wire \u_inv.input_reg[27] ;
 wire \u_inv.input_reg[28] ;
 wire \u_inv.input_reg[29] ;
 wire \u_inv.input_reg[2] ;
 wire \u_inv.input_reg[30] ;
 wire \u_inv.input_reg[31] ;
 wire \u_inv.input_reg[32] ;
 wire \u_inv.input_reg[33] ;
 wire \u_inv.input_reg[34] ;
 wire \u_inv.input_reg[35] ;
 wire \u_inv.input_reg[36] ;
 wire \u_inv.input_reg[37] ;
 wire \u_inv.input_reg[38] ;
 wire \u_inv.input_reg[39] ;
 wire \u_inv.input_reg[3] ;
 wire \u_inv.input_reg[40] ;
 wire \u_inv.input_reg[41] ;
 wire \u_inv.input_reg[42] ;
 wire \u_inv.input_reg[43] ;
 wire \u_inv.input_reg[44] ;
 wire \u_inv.input_reg[45] ;
 wire \u_inv.input_reg[46] ;
 wire \u_inv.input_reg[47] ;
 wire \u_inv.input_reg[48] ;
 wire \u_inv.input_reg[49] ;
 wire \u_inv.input_reg[4] ;
 wire \u_inv.input_reg[50] ;
 wire \u_inv.input_reg[51] ;
 wire \u_inv.input_reg[52] ;
 wire \u_inv.input_reg[53] ;
 wire \u_inv.input_reg[54] ;
 wire \u_inv.input_reg[55] ;
 wire \u_inv.input_reg[56] ;
 wire \u_inv.input_reg[57] ;
 wire \u_inv.input_reg[58] ;
 wire \u_inv.input_reg[59] ;
 wire \u_inv.input_reg[5] ;
 wire \u_inv.input_reg[60] ;
 wire \u_inv.input_reg[61] ;
 wire \u_inv.input_reg[62] ;
 wire \u_inv.input_reg[63] ;
 wire \u_inv.input_reg[64] ;
 wire \u_inv.input_reg[65] ;
 wire \u_inv.input_reg[66] ;
 wire \u_inv.input_reg[67] ;
 wire \u_inv.input_reg[68] ;
 wire \u_inv.input_reg[69] ;
 wire \u_inv.input_reg[6] ;
 wire \u_inv.input_reg[70] ;
 wire \u_inv.input_reg[71] ;
 wire \u_inv.input_reg[72] ;
 wire \u_inv.input_reg[73] ;
 wire \u_inv.input_reg[74] ;
 wire \u_inv.input_reg[75] ;
 wire \u_inv.input_reg[76] ;
 wire \u_inv.input_reg[77] ;
 wire \u_inv.input_reg[78] ;
 wire \u_inv.input_reg[79] ;
 wire \u_inv.input_reg[7] ;
 wire \u_inv.input_reg[80] ;
 wire \u_inv.input_reg[81] ;
 wire \u_inv.input_reg[82] ;
 wire \u_inv.input_reg[83] ;
 wire \u_inv.input_reg[84] ;
 wire \u_inv.input_reg[85] ;
 wire \u_inv.input_reg[86] ;
 wire \u_inv.input_reg[87] ;
 wire \u_inv.input_reg[88] ;
 wire \u_inv.input_reg[89] ;
 wire \u_inv.input_reg[8] ;
 wire \u_inv.input_reg[90] ;
 wire \u_inv.input_reg[91] ;
 wire \u_inv.input_reg[92] ;
 wire \u_inv.input_reg[93] ;
 wire \u_inv.input_reg[94] ;
 wire \u_inv.input_reg[95] ;
 wire \u_inv.input_reg[96] ;
 wire \u_inv.input_reg[97] ;
 wire \u_inv.input_reg[98] ;
 wire \u_inv.input_reg[99] ;
 wire \u_inv.input_reg[9] ;
 wire \u_inv.input_valid ;
 wire \u_inv.load_input ;
 wire \u_inv.state[0] ;
 wire \u_inv.state[1] ;
 wire net1062;
 wire clknet_leaf_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire wr_prev;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire [0:0] _17369_;

 sg13g2_inv_1 _17370_ (.Y(_10326_),
    .A(net2530));
 sg13g2_inv_1 _17371_ (.Y(_10327_),
    .A(net2535));
 sg13g2_inv_2 _17372_ (.Y(_10328_),
    .A(net2340));
 sg13g2_inv_1 _17373_ (.Y(_10329_),
    .A(net2244));
 sg13g2_inv_1 _17374_ (.Y(_10330_),
    .A(net3282));
 sg13g2_inv_1 _17375_ (.Y(_10331_),
    .A(net3180));
 sg13g2_inv_1 _17376_ (.Y(_10332_),
    .A(\u_inv.f_next[249] ));
 sg13g2_inv_1 _17377_ (.Y(_10333_),
    .A(net2890));
 sg13g2_inv_1 _17378_ (.Y(_10334_),
    .A(net2336));
 sg13g2_inv_1 _17379_ (.Y(_10335_),
    .A(net1661));
 sg13g2_inv_1 _17380_ (.Y(_10336_),
    .A(net2197));
 sg13g2_inv_2 _17381_ (.Y(_10337_),
    .A(net1439));
 sg13g2_inv_1 _17382_ (.Y(_10338_),
    .A(net2181));
 sg13g2_inv_1 _17383_ (.Y(_10339_),
    .A(net1826));
 sg13g2_inv_1 _17384_ (.Y(_10340_),
    .A(net3309));
 sg13g2_inv_1 _17385_ (.Y(_10341_),
    .A(net2696));
 sg13g2_inv_2 _17386_ (.Y(_10342_),
    .A(net2764));
 sg13g2_inv_1 _17387_ (.Y(_10343_),
    .A(net3232));
 sg13g2_inv_1 _17388_ (.Y(_10344_),
    .A(net1967));
 sg13g2_inv_1 _17389_ (.Y(_10345_),
    .A(net1625));
 sg13g2_inv_2 _17390_ (.Y(_10346_),
    .A(net2347));
 sg13g2_inv_1 _17391_ (.Y(_10347_),
    .A(net1412));
 sg13g2_inv_2 _17392_ (.Y(_10348_),
    .A(net2193));
 sg13g2_inv_1 _17393_ (.Y(_10349_),
    .A(net2947));
 sg13g2_inv_1 _17394_ (.Y(_10350_),
    .A(net3249));
 sg13g2_inv_1 _17395_ (.Y(_10351_),
    .A(net3263));
 sg13g2_inv_1 _17396_ (.Y(_10352_),
    .A(net2212));
 sg13g2_inv_1 _17397_ (.Y(_10353_),
    .A(net3277));
 sg13g2_inv_1 _17398_ (.Y(_10354_),
    .A(net4954));
 sg13g2_inv_1 _17399_ (.Y(_10355_),
    .A(\u_inv.f_next[226] ));
 sg13g2_inv_1 _17400_ (.Y(_10356_),
    .A(net2266));
 sg13g2_inv_1 _17401_ (.Y(_10357_),
    .A(net2049));
 sg13g2_inv_2 _17402_ (.Y(_10358_),
    .A(net2338));
 sg13g2_inv_1 _17403_ (.Y(_10359_),
    .A(net1463));
 sg13g2_inv_1 _17404_ (.Y(_10360_),
    .A(net2277));
 sg13g2_inv_1 _17405_ (.Y(_10361_),
    .A(net1709));
 sg13g2_inv_1 _17406_ (.Y(_10362_),
    .A(net2236));
 sg13g2_inv_1 _17407_ (.Y(_10363_),
    .A(net2109));
 sg13g2_inv_1 _17408_ (.Y(_10364_),
    .A(net2258));
 sg13g2_inv_1 _17409_ (.Y(_10365_),
    .A(net2195));
 sg13g2_inv_2 _17410_ (.Y(_10366_),
    .A(net2124));
 sg13g2_inv_1 _17411_ (.Y(_10367_),
    .A(net1696));
 sg13g2_inv_2 _17412_ (.Y(_10368_),
    .A(net2477));
 sg13g2_inv_1 _17413_ (.Y(_10369_),
    .A(net2983));
 sg13g2_inv_2 _17414_ (.Y(_10370_),
    .A(net2832));
 sg13g2_inv_1 _17415_ (.Y(_10371_),
    .A(net2206));
 sg13g2_inv_1 _17416_ (.Y(_10372_),
    .A(net2549));
 sg13g2_inv_1 _17417_ (.Y(_10373_),
    .A(net2482));
 sg13g2_inv_1 _17418_ (.Y(_10374_),
    .A(net2177));
 sg13g2_inv_1 _17419_ (.Y(_10375_),
    .A(net2664));
 sg13g2_inv_1 _17420_ (.Y(_10376_),
    .A(net2943));
 sg13g2_inv_2 _17421_ (.Y(_10377_),
    .A(net2809));
 sg13g2_inv_1 _17422_ (.Y(_10378_),
    .A(net4953));
 sg13g2_inv_1 _17423_ (.Y(_10379_),
    .A(net1959));
 sg13g2_inv_1 _17424_ (.Y(_10380_),
    .A(net1992));
 sg13g2_inv_1 _17425_ (.Y(_10381_),
    .A(net2509));
 sg13g2_inv_1 _17426_ (.Y(_10382_),
    .A(net3304));
 sg13g2_inv_1 _17427_ (.Y(_10383_),
    .A(net1627));
 sg13g2_inv_1 _17428_ (.Y(_10384_),
    .A(net1704));
 sg13g2_inv_1 _17429_ (.Y(_10385_),
    .A(net1770));
 sg13g2_inv_2 _17430_ (.Y(_10386_),
    .A(net2440));
 sg13g2_inv_2 _17431_ (.Y(_10387_),
    .A(net3005));
 sg13g2_inv_1 _17432_ (.Y(_10388_),
    .A(net2771));
 sg13g2_inv_1 _17433_ (.Y(_10389_),
    .A(net2242));
 sg13g2_inv_2 _17434_ (.Y(_10390_),
    .A(net3276));
 sg13g2_inv_1 _17435_ (.Y(_10391_),
    .A(net2316));
 sg13g2_inv_1 _17436_ (.Y(_10392_),
    .A(net2129));
 sg13g2_inv_1 _17437_ (.Y(_10393_),
    .A(net2188));
 sg13g2_inv_1 _17438_ (.Y(_10394_),
    .A(net2984));
 sg13g2_inv_1 _17439_ (.Y(_10395_),
    .A(net3265));
 sg13g2_inv_1 _17440_ (.Y(_10396_),
    .A(net2175));
 sg13g2_inv_1 _17441_ (.Y(_10397_),
    .A(net2151));
 sg13g2_inv_1 _17442_ (.Y(_10398_),
    .A(net2366));
 sg13g2_inv_1 _17443_ (.Y(_10399_),
    .A(net2791));
 sg13g2_inv_1 _17444_ (.Y(_10400_),
    .A(net2616));
 sg13g2_inv_2 _17445_ (.Y(_10401_),
    .A(net2497));
 sg13g2_inv_1 _17446_ (.Y(_10402_),
    .A(\u_inv.f_next[179] ));
 sg13g2_inv_1 _17447_ (.Y(_10403_),
    .A(net3295));
 sg13g2_inv_1 _17448_ (.Y(_10404_),
    .A(net2231));
 sg13g2_inv_1 _17449_ (.Y(_10405_),
    .A(net2044));
 sg13g2_inv_1 _17450_ (.Y(_10406_),
    .A(net2191));
 sg13g2_inv_1 _17451_ (.Y(_10407_),
    .A(net2630));
 sg13g2_inv_2 _17452_ (.Y(_10408_),
    .A(net2202));
 sg13g2_inv_1 _17453_ (.Y(_10409_),
    .A(\u_inv.f_next[172] ));
 sg13g2_inv_2 _17454_ (.Y(_10410_),
    .A(net2784));
 sg13g2_inv_2 _17455_ (.Y(_10411_),
    .A(net3137));
 sg13g2_inv_1 _17456_ (.Y(_10412_),
    .A(net2083));
 sg13g2_inv_1 _17457_ (.Y(_10413_),
    .A(net2818));
 sg13g2_inv_2 _17458_ (.Y(_10414_),
    .A(net2504));
 sg13g2_inv_1 _17459_ (.Y(_10415_),
    .A(\u_inv.f_next[166] ));
 sg13g2_inv_1 _17460_ (.Y(_10416_),
    .A(net2854));
 sg13g2_inv_1 _17461_ (.Y(_10417_),
    .A(net2256));
 sg13g2_inv_1 _17462_ (.Y(_10418_),
    .A(net1908));
 sg13g2_inv_1 _17463_ (.Y(_10419_),
    .A(net1772));
 sg13g2_inv_1 _17464_ (.Y(_10420_),
    .A(net2140));
 sg13g2_inv_1 _17465_ (.Y(_10421_),
    .A(net3271));
 sg13g2_inv_2 _17466_ (.Y(_10422_),
    .A(\u_inv.f_next[159] ));
 sg13g2_inv_1 _17467_ (.Y(_10423_),
    .A(net1475));
 sg13g2_inv_1 _17468_ (.Y(_10424_),
    .A(net3028));
 sg13g2_inv_1 _17469_ (.Y(_10425_),
    .A(net1748));
 sg13g2_inv_1 _17470_ (.Y(_10426_),
    .A(net3199));
 sg13g2_inv_2 _17471_ (.Y(_10427_),
    .A(net2411));
 sg13g2_inv_1 _17472_ (.Y(_10428_),
    .A(net2878));
 sg13g2_inv_2 _17473_ (.Y(_10429_),
    .A(net2334));
 sg13g2_inv_1 _17474_ (.Y(_10430_),
    .A(net3042));
 sg13g2_inv_1 _17475_ (.Y(_10431_),
    .A(net3093));
 sg13g2_inv_2 _17476_ (.Y(_10432_),
    .A(net2792));
 sg13g2_inv_1 _17477_ (.Y(_10433_),
    .A(net3242));
 sg13g2_inv_1 _17478_ (.Y(_10434_),
    .A(net3018));
 sg13g2_inv_1 _17479_ (.Y(_10435_),
    .A(net3305));
 sg13g2_inv_1 _17480_ (.Y(_10436_),
    .A(\u_inv.f_next[145] ));
 sg13g2_inv_1 _17481_ (.Y(_10437_),
    .A(net2073));
 sg13g2_inv_1 _17482_ (.Y(_10438_),
    .A(net2419));
 sg13g2_inv_1 _17483_ (.Y(_10439_),
    .A(net2799));
 sg13g2_inv_2 _17484_ (.Y(_10440_),
    .A(net2406));
 sg13g2_inv_1 _17485_ (.Y(_10441_),
    .A(net1728));
 sg13g2_inv_1 _17486_ (.Y(_10442_),
    .A(net3141));
 sg13g2_inv_1 _17487_ (.Y(_10443_),
    .A(\u_inv.f_next[138] ));
 sg13g2_inv_1 _17488_ (.Y(_10444_),
    .A(net2332));
 sg13g2_inv_1 _17489_ (.Y(_10445_),
    .A(net3283));
 sg13g2_inv_1 _17490_ (.Y(_10446_),
    .A(net2868));
 sg13g2_inv_1 _17491_ (.Y(_10447_),
    .A(net2618));
 sg13g2_inv_1 _17492_ (.Y(_10448_),
    .A(net2400));
 sg13g2_inv_1 _17493_ (.Y(_10449_),
    .A(net2097));
 sg13g2_inv_1 _17494_ (.Y(_10450_),
    .A(net2720));
 sg13g2_inv_1 _17495_ (.Y(_10451_),
    .A(net3279));
 sg13g2_inv_1 _17496_ (.Y(_10452_),
    .A(net1878));
 sg13g2_inv_1 _17497_ (.Y(_10453_),
    .A(net2561));
 sg13g2_inv_2 _17498_ (.Y(_10454_),
    .A(net2545));
 sg13g2_inv_1 _17499_ (.Y(_10455_),
    .A(net2821));
 sg13g2_inv_2 _17500_ (.Y(_10456_),
    .A(net2171));
 sg13g2_inv_1 _17501_ (.Y(_10457_),
    .A(net1558));
 sg13g2_inv_2 _17502_ (.Y(_10458_),
    .A(net2884));
 sg13g2_inv_1 _17503_ (.Y(_10459_),
    .A(net2164));
 sg13g2_inv_2 _17504_ (.Y(_10460_),
    .A(net2420));
 sg13g2_inv_1 _17505_ (.Y(_10461_),
    .A(net3299));
 sg13g2_inv_1 _17506_ (.Y(_10462_),
    .A(\u_inv.f_next[119] ));
 sg13g2_inv_1 _17507_ (.Y(_10463_),
    .A(net3140));
 sg13g2_inv_1 _17508_ (.Y(_10464_),
    .A(net2989));
 sg13g2_inv_2 _17509_ (.Y(_10465_),
    .A(net2223));
 sg13g2_inv_1 _17510_ (.Y(_10466_),
    .A(net2997));
 sg13g2_inv_1 _17511_ (.Y(_10467_),
    .A(net2404));
 sg13g2_inv_1 _17512_ (.Y(_10468_),
    .A(net2661));
 sg13g2_inv_1 _17513_ (.Y(_10469_),
    .A(net1527));
 sg13g2_inv_1 _17514_ (.Y(_10470_),
    .A(net2148));
 sg13g2_inv_1 _17515_ (.Y(_10471_),
    .A(net2100));
 sg13g2_inv_1 _17516_ (.Y(_10472_),
    .A(net2526));
 sg13g2_inv_2 _17517_ (.Y(_10473_),
    .A(net2778));
 sg13g2_inv_2 _17518_ (.Y(_10474_),
    .A(net2585));
 sg13g2_inv_1 _17519_ (.Y(_10475_),
    .A(net3284));
 sg13g2_inv_1 _17520_ (.Y(_10476_),
    .A(net4957));
 sg13g2_inv_1 _17521_ (.Y(_10477_),
    .A(net3162));
 sg13g2_inv_1 _17522_ (.Y(_10478_),
    .A(net2328));
 sg13g2_inv_1 _17523_ (.Y(_10479_),
    .A(net3221));
 sg13g2_inv_1 _17524_ (.Y(_10480_),
    .A(net2018));
 sg13g2_inv_1 _17525_ (.Y(_10481_),
    .A(net3083));
 sg13g2_inv_1 _17526_ (.Y(_10482_),
    .A(net1761));
 sg13g2_inv_1 _17527_ (.Y(_10483_),
    .A(net2086));
 sg13g2_inv_1 _17528_ (.Y(_10484_),
    .A(net3204));
 sg13g2_inv_2 _17529_ (.Y(_10485_),
    .A(net2499));
 sg13g2_inv_2 _17530_ (.Y(_10486_),
    .A(net2380));
 sg13g2_inv_1 _17531_ (.Y(_10487_),
    .A(net1799));
 sg13g2_inv_1 _17532_ (.Y(_10488_),
    .A(net2842));
 sg13g2_inv_1 _17533_ (.Y(_10489_),
    .A(net2353));
 sg13g2_inv_1 _17534_ (.Y(_10490_),
    .A(net2940));
 sg13g2_inv_1 _17535_ (.Y(_10491_),
    .A(net3111));
 sg13g2_inv_1 _17536_ (.Y(_10492_),
    .A(net2865));
 sg13g2_inv_1 _17537_ (.Y(_10493_),
    .A(net3245));
 sg13g2_inv_1 _17538_ (.Y(_10494_),
    .A(\u_inv.f_next[87] ));
 sg13g2_inv_1 _17539_ (.Y(_10495_),
    .A(net3227));
 sg13g2_inv_1 _17540_ (.Y(_10496_),
    .A(net3156));
 sg13g2_inv_1 _17541_ (.Y(_10497_),
    .A(net3153));
 sg13g2_inv_1 _17542_ (.Y(_10498_),
    .A(net3084));
 sg13g2_inv_1 _17543_ (.Y(_10499_),
    .A(net2382));
 sg13g2_inv_1 _17544_ (.Y(_10500_),
    .A(\u_inv.f_next[81] ));
 sg13g2_inv_1 _17545_ (.Y(_10501_),
    .A(net3071));
 sg13g2_inv_1 _17546_ (.Y(_10502_),
    .A(net2568));
 sg13g2_inv_2 _17547_ (.Y(_10503_),
    .A(net2271));
 sg13g2_inv_1 _17548_ (.Y(_10504_),
    .A(net2769));
 sg13g2_inv_1 _17549_ (.Y(_10505_),
    .A(net3037));
 sg13g2_inv_1 _17550_ (.Y(_10506_),
    .A(net2979));
 sg13g2_inv_2 _17551_ (.Y(_10507_),
    .A(net2571));
 sg13g2_inv_1 _17552_ (.Y(_10508_),
    .A(net2308));
 sg13g2_inv_1 _17553_ (.Y(_10509_),
    .A(net2067));
 sg13g2_inv_2 _17554_ (.Y(_10510_),
    .A(net2317));
 sg13g2_inv_1 _17555_ (.Y(_10511_),
    .A(net1539));
 sg13g2_inv_2 _17556_ (.Y(_10512_),
    .A(net2554));
 sg13g2_inv_1 _17557_ (.Y(_10513_),
    .A(net2060));
 sg13g2_inv_1 _17558_ (.Y(_10514_),
    .A(net2349));
 sg13g2_inv_2 _17559_ (.Y(_10515_),
    .A(net2217));
 sg13g2_inv_1 _17560_ (.Y(_10516_),
    .A(net2051));
 sg13g2_inv_1 _17561_ (.Y(_10517_),
    .A(net2147));
 sg13g2_inv_1 _17562_ (.Y(_10518_),
    .A(net3301));
 sg13g2_inv_1 _17563_ (.Y(_10519_),
    .A(net1969));
 sg13g2_inv_1 _17564_ (.Y(_10520_),
    .A(\u_inv.f_next[61] ));
 sg13g2_inv_1 _17565_ (.Y(_10521_),
    .A(net3124));
 sg13g2_inv_1 _17566_ (.Y(_10522_),
    .A(\u_inv.f_next[59] ));
 sg13g2_inv_1 _17567_ (.Y(_10523_),
    .A(net3248));
 sg13g2_inv_1 _17568_ (.Y(_10524_),
    .A(net3178));
 sg13g2_inv_1 _17569_ (.Y(_10525_),
    .A(net2689));
 sg13g2_inv_2 _17570_ (.Y(_10526_),
    .A(net2313));
 sg13g2_inv_2 _17571_ (.Y(_10527_),
    .A(net3169));
 sg13g2_inv_1 _17572_ (.Y(_10528_),
    .A(net2857));
 sg13g2_inv_1 _17573_ (.Y(_10529_),
    .A(net2402));
 sg13g2_inv_1 _17574_ (.Y(_10530_),
    .A(net2702));
 sg13g2_inv_1 _17575_ (.Y(_10531_),
    .A(net2234));
 sg13g2_inv_1 _17576_ (.Y(_10532_),
    .A(net3015));
 sg13g2_inv_2 _17577_ (.Y(_10533_),
    .A(net2485));
 sg13g2_inv_1 _17578_ (.Y(_10534_),
    .A(\u_inv.f_next[47] ));
 sg13g2_inv_1 _17579_ (.Y(_10535_),
    .A(net2831));
 sg13g2_inv_1 _17580_ (.Y(_10536_),
    .A(net2593));
 sg13g2_inv_2 _17581_ (.Y(_10537_),
    .A(net3013));
 sg13g2_inv_1 _17582_ (.Y(_10538_),
    .A(net3306));
 sg13g2_inv_1 _17583_ (.Y(_10539_),
    .A(net2306));
 sg13g2_inv_1 _17584_ (.Y(_10540_),
    .A(net1905));
 sg13g2_inv_1 _17585_ (.Y(_10541_),
    .A(net2156));
 sg13g2_inv_2 _17586_ (.Y(_10542_),
    .A(net2513));
 sg13g2_inv_2 _17587_ (.Y(_10543_),
    .A(net2610));
 sg13g2_inv_2 _17588_ (.Y(_10544_),
    .A(net2937));
 sg13g2_inv_1 _17589_ (.Y(_10545_),
    .A(net2077));
 sg13g2_inv_1 _17590_ (.Y(_10546_),
    .A(net2801));
 sg13g2_inv_2 _17591_ (.Y(_10547_),
    .A(net2896));
 sg13g2_inv_1 _17592_ (.Y(_10548_),
    .A(net3228));
 sg13g2_inv_1 _17593_ (.Y(_10549_),
    .A(net2280));
 sg13g2_inv_2 _17594_ (.Y(_10550_),
    .A(net2712));
 sg13g2_inv_1 _17595_ (.Y(_10551_),
    .A(net3308));
 sg13g2_inv_1 _17596_ (.Y(_10552_),
    .A(net3119));
 sg13g2_inv_2 _17597_ (.Y(_10553_),
    .A(net3209));
 sg13g2_inv_1 _17598_ (.Y(_10554_),
    .A(net3133));
 sg13g2_inv_1 _17599_ (.Y(_10555_),
    .A(net3246));
 sg13g2_inv_2 _17600_ (.Y(_10556_),
    .A(net2722));
 sg13g2_inv_1 _17601_ (.Y(_10557_),
    .A(net1754));
 sg13g2_inv_2 _17602_ (.Y(_10558_),
    .A(net2430));
 sg13g2_inv_2 _17603_ (.Y(_10559_),
    .A(net2643));
 sg13g2_inv_2 _17604_ (.Y(_10560_),
    .A(net2250));
 sg13g2_inv_1 _17605_ (.Y(_10561_),
    .A(\u_inv.f_next[20] ));
 sg13g2_inv_1 _17606_ (.Y(_10562_),
    .A(net2812));
 sg13g2_inv_1 _17607_ (.Y(_10563_),
    .A(net2290));
 sg13g2_inv_1 _17608_ (.Y(_10564_),
    .A(net1744));
 sg13g2_inv_1 _17609_ (.Y(_10565_),
    .A(net3189));
 sg13g2_inv_1 _17610_ (.Y(_10566_),
    .A(\u_inv.f_next[15] ));
 sg13g2_inv_1 _17611_ (.Y(_10567_),
    .A(net3297));
 sg13g2_inv_1 _17612_ (.Y(_10568_),
    .A(net4958));
 sg13g2_inv_1 _17613_ (.Y(_10569_),
    .A(net2528));
 sg13g2_inv_1 _17614_ (.Y(_10570_),
    .A(net3044));
 sg13g2_inv_2 _17615_ (.Y(_10571_),
    .A(net2601));
 sg13g2_inv_1 _17616_ (.Y(_10572_),
    .A(net2143));
 sg13g2_inv_1 _17617_ (.Y(_10573_),
    .A(net2122));
 sg13g2_inv_1 _17618_ (.Y(_10574_),
    .A(net2186));
 sg13g2_inv_1 _17619_ (.Y(_10575_),
    .A(\u_inv.f_next[2] ));
 sg13g2_inv_1 _17620_ (.Y(_10576_),
    .A(net3290));
 sg13g2_inv_8 _17621_ (.Y(_10577_),
    .A(net4685));
 sg13g2_inv_1 _17622_ (.Y(_10578_),
    .A(net2275));
 sg13g2_inv_1 _17623_ (.Y(_10579_),
    .A(\u_inv.d_next[231] ));
 sg13g2_inv_1 _17624_ (.Y(_10580_),
    .A(\u_inv.d_next[223] ));
 sg13g2_inv_1 _17625_ (.Y(_10581_),
    .A(net2013));
 sg13g2_inv_1 _17626_ (.Y(_10582_),
    .A(net2931));
 sg13g2_inv_1 _17627_ (.Y(_10583_),
    .A(net2967));
 sg13g2_inv_1 _17628_ (.Y(_10584_),
    .A(net2913));
 sg13g2_inv_1 _17629_ (.Y(_10585_),
    .A(net2998));
 sg13g2_inv_1 _17630_ (.Y(_10586_),
    .A(net2762));
 sg13g2_inv_1 _17631_ (.Y(_10587_),
    .A(net2454));
 sg13g2_inv_1 _17632_ (.Y(_10588_),
    .A(\u_inv.d_next[191] ));
 sg13g2_inv_1 _17633_ (.Y(_10589_),
    .A(net2297));
 sg13g2_inv_1 _17634_ (.Y(_10590_),
    .A(net2672));
 sg13g2_inv_2 _17635_ (.Y(_10591_),
    .A(net2273));
 sg13g2_inv_1 _17636_ (.Y(_10592_),
    .A(net2392));
 sg13g2_inv_1 _17637_ (.Y(_10593_),
    .A(net2342));
 sg13g2_inv_2 _17638_ (.Y(_10594_),
    .A(net3164));
 sg13g2_inv_1 _17639_ (.Y(_10595_),
    .A(net2906));
 sg13g2_inv_1 _17640_ (.Y(_10596_),
    .A(net2269));
 sg13g2_inv_1 _17641_ (.Y(_10597_),
    .A(net2311));
 sg13g2_inv_1 _17642_ (.Y(_10598_),
    .A(net3106));
 sg13g2_inv_1 _17643_ (.Y(_10599_),
    .A(net2364));
 sg13g2_inv_1 _17644_ (.Y(_10600_),
    .A(net2924));
 sg13g2_inv_1 _17645_ (.Y(_10601_),
    .A(net2489));
 sg13g2_inv_1 _17646_ (.Y(_10602_),
    .A(\u_inv.d_next[121] ));
 sg13g2_inv_1 _17647_ (.Y(_10603_),
    .A(\u_inv.d_next[114] ));
 sg13g2_inv_1 _17648_ (.Y(_10604_),
    .A(net2976));
 sg13g2_inv_1 _17649_ (.Y(_10605_),
    .A(net3293));
 sg13g2_inv_1 _17650_ (.Y(_10606_),
    .A(net2806));
 sg13g2_inv_1 _17651_ (.Y(_10607_),
    .A(\u_inv.d_next[103] ));
 sg13g2_inv_1 _17652_ (.Y(_10608_),
    .A(net2263));
 sg13g2_inv_1 _17653_ (.Y(_10609_),
    .A(net3020));
 sg13g2_inv_1 _17654_ (.Y(_10610_),
    .A(net2524));
 sg13g2_inv_1 _17655_ (.Y(_10611_),
    .A(net2647));
 sg13g2_inv_1 _17656_ (.Y(_10612_),
    .A(net2991));
 sg13g2_inv_1 _17657_ (.Y(_10613_),
    .A(net2625));
 sg13g2_inv_1 _17658_ (.Y(_10614_),
    .A(net3038));
 sg13g2_inv_1 _17659_ (.Y(_10615_),
    .A(\u_inv.d_next[47] ));
 sg13g2_inv_1 _17660_ (.Y(_10616_),
    .A(net2957));
 sg13g2_inv_1 _17661_ (.Y(_10617_),
    .A(\u_inv.d_next[31] ));
 sg13g2_inv_1 _17662_ (.Y(_10618_),
    .A(net2649));
 sg13g2_inv_1 _17663_ (.Y(_10619_),
    .A(\u_inv.d_next[19] ));
 sg13g2_inv_1 _17664_ (.Y(_10620_),
    .A(\u_inv.d_next[14] ));
 sg13g2_inv_1 _17665_ (.Y(_10621_),
    .A(\u_inv.d_next[9] ));
 sg13g2_inv_1 _17666_ (.Y(_10622_),
    .A(net2547));
 sg13g2_inv_1 _17667_ (.Y(_10623_),
    .A(net2558));
 sg13g2_inv_1 _17668_ (.Y(_10624_),
    .A(net2479));
 sg13g2_inv_8 _17669_ (.Y(_10625_),
    .A(net4612));
 sg13g2_inv_1 _17670_ (.Y(_10626_),
    .A(net2883));
 sg13g2_inv_1 _17671_ (.Y(_10627_),
    .A(\u_inv.input_valid ));
 sg13g2_inv_1 _17672_ (.Y(_10628_),
    .A(net1603));
 sg13g2_inv_1 _17673_ (.Y(_10629_),
    .A(\u_inv.delta_reg[4] ));
 sg13g2_inv_1 _17674_ (.Y(_10630_),
    .A(net1680));
 sg13g2_inv_1 _17675_ (.Y(_10631_),
    .A(net3160));
 sg13g2_inv_1 _17676_ (.Y(_10632_),
    .A(inv_go));
 sg13g2_inv_1 _17677_ (.Y(_10633_),
    .A(net1631));
 sg13g2_inv_8 _17678_ (.Y(_10634_),
    .A(net4729));
 sg13g2_inv_1 _17679_ (.Y(_10635_),
    .A(net2996));
 sg13g2_inv_1 _17680_ (.Y(_10636_),
    .A(\u_inv.f_reg[254] ));
 sg13g2_inv_1 _17681_ (.Y(_10637_),
    .A(\u_inv.f_reg[253] ));
 sg13g2_inv_1 _17682_ (.Y(_10638_),
    .A(net2322));
 sg13g2_inv_1 _17683_ (.Y(_10639_),
    .A(net3075));
 sg13g2_inv_1 _17684_ (.Y(_10640_),
    .A(net2427));
 sg13g2_inv_1 _17685_ (.Y(_10641_),
    .A(net3091));
 sg13g2_inv_1 _17686_ (.Y(_10642_),
    .A(net2903));
 sg13g2_inv_1 _17687_ (.Y(_10643_),
    .A(net2880));
 sg13g2_inv_1 _17688_ (.Y(_10644_),
    .A(net2226));
 sg13g2_inv_1 _17689_ (.Y(_10645_),
    .A(net2653));
 sg13g2_inv_1 _17690_ (.Y(_10646_),
    .A(net2024));
 sg13g2_inv_1 _17691_ (.Y(_10647_),
    .A(net2886));
 sg13g2_inv_1 _17692_ (.Y(_10648_),
    .A(net2379));
 sg13g2_inv_1 _17693_ (.Y(_10649_),
    .A(net3184));
 sg13g2_inv_1 _17694_ (.Y(_10650_),
    .A(net3177));
 sg13g2_inv_1 _17695_ (.Y(_10651_),
    .A(\u_inv.f_reg[239] ));
 sg13g2_inv_1 _17696_ (.Y(_10652_),
    .A(net2145));
 sg13g2_inv_1 _17697_ (.Y(_10653_),
    .A(net2688));
 sg13g2_inv_1 _17698_ (.Y(_10654_),
    .A(net2090));
 sg13g2_inv_1 _17699_ (.Y(_10655_),
    .A(\u_inv.f_reg[235] ));
 sg13g2_inv_1 _17700_ (.Y(_10656_),
    .A(net1971));
 sg13g2_inv_1 _17701_ (.Y(_10657_),
    .A(net2749));
 sg13g2_inv_1 _17702_ (.Y(_10658_),
    .A(net2681));
 sg13g2_inv_1 _17703_ (.Y(_10659_),
    .A(\u_inv.f_reg[231] ));
 sg13g2_inv_1 _17704_ (.Y(_10660_),
    .A(net2964));
 sg13g2_inv_1 _17705_ (.Y(_10661_),
    .A(net2861));
 sg13g2_inv_1 _17706_ (.Y(_10662_),
    .A(\u_inv.f_reg[228] ));
 sg13g2_inv_1 _17707_ (.Y(_10663_),
    .A(net3193));
 sg13g2_inv_1 _17708_ (.Y(_10664_),
    .A(net2361));
 sg13g2_inv_2 _17709_ (.Y(_10665_),
    .A(net2417));
 sg13g2_inv_1 _17710_ (.Y(_10666_),
    .A(net2523));
 sg13g2_inv_1 _17711_ (.Y(_10667_),
    .A(\u_inv.f_reg[223] ));
 sg13g2_inv_1 _17712_ (.Y(_10668_),
    .A(net1867));
 sg13g2_inv_1 _17713_ (.Y(_10669_),
    .A(net3003));
 sg13g2_inv_1 _17714_ (.Y(_10670_),
    .A(net2544));
 sg13g2_inv_1 _17715_ (.Y(_10671_),
    .A(net2444));
 sg13g2_inv_1 _17716_ (.Y(_10672_),
    .A(net2676));
 sg13g2_inv_2 _17717_ (.Y(_10673_),
    .A(net2495));
 sg13g2_inv_1 _17718_ (.Y(_10674_),
    .A(net2446));
 sg13g2_inv_1 _17719_ (.Y(_10675_),
    .A(net2484));
 sg13g2_inv_1 _17720_ (.Y(_10676_),
    .A(net2115));
 sg13g2_inv_1 _17721_ (.Y(_10677_),
    .A(\u_inv.f_reg[213] ));
 sg13g2_inv_1 _17722_ (.Y(_10678_),
    .A(net2320));
 sg13g2_inv_1 _17723_ (.Y(_10679_),
    .A(\u_inv.f_reg[211] ));
 sg13g2_inv_1 _17724_ (.Y(_10680_),
    .A(net2370));
 sg13g2_inv_1 _17725_ (.Y(_10681_),
    .A(net2839));
 sg13g2_inv_1 _17726_ (.Y(_10682_),
    .A(\u_inv.f_reg[208] ));
 sg13g2_inv_1 _17727_ (.Y(_10683_),
    .A(net3050));
 sg13g2_inv_1 _17728_ (.Y(_10684_),
    .A(net3270));
 sg13g2_inv_1 _17729_ (.Y(_10685_),
    .A(\u_inv.f_reg[205] ));
 sg13g2_inv_1 _17730_ (.Y(_10686_),
    .A(net2254));
 sg13g2_inv_1 _17731_ (.Y(_10687_),
    .A(net3259));
 sg13g2_inv_1 _17732_ (.Y(_10688_),
    .A(net2211));
 sg13g2_inv_1 _17733_ (.Y(_10689_),
    .A(net2438));
 sg13g2_inv_1 _17734_ (.Y(_10690_),
    .A(net2566));
 sg13g2_inv_1 _17735_ (.Y(_10691_),
    .A(net2677));
 sg13g2_inv_1 _17736_ (.Y(_10692_),
    .A(net2410));
 sg13g2_inv_1 _17737_ (.Y(_10693_),
    .A(net2646));
 sg13g2_inv_1 _17738_ (.Y(_10694_),
    .A(net2464));
 sg13g2_inv_1 _17739_ (.Y(_10695_),
    .A(\u_inv.f_reg[195] ));
 sg13g2_inv_1 _17740_ (.Y(_10696_),
    .A(net2358));
 sg13g2_inv_1 _17741_ (.Y(_10697_),
    .A(\u_inv.f_reg[193] ));
 sg13g2_inv_1 _17742_ (.Y(_10698_),
    .A(net3012));
 sg13g2_inv_1 _17743_ (.Y(_10699_),
    .A(net2575));
 sg13g2_inv_1 _17744_ (.Y(_10700_),
    .A(net2325));
 sg13g2_inv_1 _17745_ (.Y(_10701_),
    .A(net3006));
 sg13g2_inv_1 _17746_ (.Y(_10702_),
    .A(net2995));
 sg13g2_inv_1 _17747_ (.Y(_10703_),
    .A(net3116));
 sg13g2_inv_1 _17748_ (.Y(_10704_),
    .A(net1941));
 sg13g2_inv_1 _17749_ (.Y(_10705_),
    .A(net2475));
 sg13g2_inv_1 _17750_ (.Y(_10706_),
    .A(net2633));
 sg13g2_inv_1 _17751_ (.Y(_10707_),
    .A(net2928));
 sg13g2_inv_1 _17752_ (.Y(_10708_),
    .A(net2916));
 sg13g2_inv_1 _17753_ (.Y(_10709_),
    .A(\u_inv.f_reg[181] ));
 sg13g2_inv_1 _17754_ (.Y(_10710_),
    .A(\u_inv.f_reg[180] ));
 sg13g2_inv_1 _17755_ (.Y(_10711_),
    .A(net2471));
 sg13g2_inv_1 _17756_ (.Y(_10712_),
    .A(net2247));
 sg13g2_inv_1 _17757_ (.Y(_10713_),
    .A(net2709));
 sg13g2_inv_1 _17758_ (.Y(_10714_),
    .A(net2726));
 sg13g2_inv_1 _17759_ (.Y(_10715_),
    .A(net2591));
 sg13g2_inv_1 _17760_ (.Y(_10716_),
    .A(net2603));
 sg13g2_inv_1 _17761_ (.Y(_10717_),
    .A(\u_inv.f_reg[173] ));
 sg13g2_inv_1 _17762_ (.Y(_10718_),
    .A(net2287));
 sg13g2_inv_1 _17763_ (.Y(_10719_),
    .A(\u_inv.f_reg[171] ));
 sg13g2_inv_1 _17764_ (.Y(_10720_),
    .A(net2750));
 sg13g2_inv_1 _17765_ (.Y(_10721_),
    .A(net3128));
 sg13g2_inv_1 _17766_ (.Y(_10722_),
    .A(net2950));
 sg13g2_inv_1 _17767_ (.Y(_10723_),
    .A(\u_inv.f_reg[167] ));
 sg13g2_inv_1 _17768_ (.Y(_10724_),
    .A(net2002));
 sg13g2_inv_1 _17769_ (.Y(_10725_),
    .A(net3251));
 sg13g2_inv_1 _17770_ (.Y(_10726_),
    .A(net3280));
 sg13g2_inv_1 _17771_ (.Y(_10727_),
    .A(net2715));
 sg13g2_inv_1 _17772_ (.Y(_10728_),
    .A(net1926));
 sg13g2_inv_1 _17773_ (.Y(_10729_),
    .A(net3187));
 sg13g2_inv_1 _17774_ (.Y(_10730_),
    .A(net2434));
 sg13g2_inv_1 _17775_ (.Y(_10731_),
    .A(net1956));
 sg13g2_inv_1 _17776_ (.Y(_10732_),
    .A(net1924));
 sg13g2_inv_1 _17777_ (.Y(_10733_),
    .A(\u_inv.f_reg[157] ));
 sg13g2_inv_1 _17778_ (.Y(_10734_),
    .A(net2301));
 sg13g2_inv_1 _17779_ (.Y(_10735_),
    .A(net2827));
 sg13g2_inv_1 _17780_ (.Y(_10736_),
    .A(\u_inv.f_reg[154] ));
 sg13g2_inv_1 _17781_ (.Y(_10737_),
    .A(net3102));
 sg13g2_inv_1 _17782_ (.Y(_10738_),
    .A(\u_inv.f_reg[152] ));
 sg13g2_inv_1 _17783_ (.Y(_10739_),
    .A(\u_inv.f_reg[151] ));
 sg13g2_inv_1 _17784_ (.Y(_10740_),
    .A(net3077));
 sg13g2_inv_1 _17785_ (.Y(_10741_),
    .A(\u_inv.f_reg[149] ));
 sg13g2_inv_1 _17786_ (.Y(_10742_),
    .A(net3296));
 sg13g2_inv_1 _17787_ (.Y(_10743_),
    .A(\u_inv.f_reg[147] ));
 sg13g2_inv_1 _17788_ (.Y(_10744_),
    .A(net3100));
 sg13g2_inv_1 _17789_ (.Y(_10745_),
    .A(net2683));
 sg13g2_inv_1 _17790_ (.Y(_10746_),
    .A(net2278));
 sg13g2_inv_1 _17791_ (.Y(_10747_),
    .A(net2629));
 sg13g2_inv_1 _17792_ (.Y(_10748_),
    .A(net2860));
 sg13g2_inv_1 _17793_ (.Y(_10749_),
    .A(\u_inv.f_reg[141] ));
 sg13g2_inv_1 _17794_ (.Y(_10750_),
    .A(net3145));
 sg13g2_inv_1 _17795_ (.Y(_10751_),
    .A(\u_inv.f_reg[139] ));
 sg13g2_inv_1 _17796_ (.Y(_10752_),
    .A(net2167));
 sg13g2_inv_1 _17797_ (.Y(_10753_),
    .A(net2396));
 sg13g2_inv_1 _17798_ (.Y(_10754_),
    .A(net2158));
 sg13g2_inv_1 _17799_ (.Y(_10755_),
    .A(net3103));
 sg13g2_inv_1 _17800_ (.Y(_10756_),
    .A(net2975));
 sg13g2_inv_1 _17801_ (.Y(_10757_),
    .A(net2915));
 sg13g2_inv_1 _17802_ (.Y(_10758_),
    .A(net2282));
 sg13g2_inv_1 _17803_ (.Y(_10759_),
    .A(net3183));
 sg13g2_inv_1 _17804_ (.Y(_10760_),
    .A(net2813));
 sg13g2_inv_1 _17805_ (.Y(_10761_),
    .A(net2487));
 sg13g2_inv_1 _17806_ (.Y(_10762_),
    .A(net2590));
 sg13g2_inv_1 _17807_ (.Y(_10763_),
    .A(\u_inv.f_reg[127] ));
 sg13g2_inv_1 _17808_ (.Y(_10764_),
    .A(net2102));
 sg13g2_inv_1 _17809_ (.Y(_10765_),
    .A(\u_inv.f_reg[125] ));
 sg13g2_inv_1 _17810_ (.Y(_10766_),
    .A(net2592));
 sg13g2_inv_1 _17811_ (.Y(_10767_),
    .A(\u_inv.f_reg[123] ));
 sg13g2_inv_1 _17812_ (.Y(_10768_),
    .A(net2219));
 sg13g2_inv_1 _17813_ (.Y(_10769_),
    .A(\u_inv.f_reg[121] ));
 sg13g2_inv_1 _17814_ (.Y(_10770_),
    .A(net2386));
 sg13g2_inv_1 _17815_ (.Y(_10771_),
    .A(net2469));
 sg13g2_inv_1 _17816_ (.Y(_10772_),
    .A(net2034));
 sg13g2_inv_1 _17817_ (.Y(_10773_),
    .A(net3109));
 sg13g2_inv_1 _17818_ (.Y(_10774_),
    .A(\u_inv.f_reg[116] ));
 sg13g2_inv_1 _17819_ (.Y(_10775_),
    .A(net3063));
 sg13g2_inv_1 _17820_ (.Y(_10776_),
    .A(\u_inv.f_reg[114] ));
 sg13g2_inv_1 _17821_ (.Y(_10777_),
    .A(net2736));
 sg13g2_inv_1 _17822_ (.Y(_10778_),
    .A(net2620));
 sg13g2_inv_1 _17823_ (.Y(_10779_),
    .A(\u_inv.f_reg[111] ));
 sg13g2_inv_1 _17824_ (.Y(_10780_),
    .A(net2779));
 sg13g2_inv_1 _17825_ (.Y(_10781_),
    .A(\u_inv.f_reg[109] ));
 sg13g2_inv_1 _17826_ (.Y(_10782_),
    .A(net2414));
 sg13g2_inv_1 _17827_ (.Y(_10783_),
    .A(\u_inv.f_reg[107] ));
 sg13g2_inv_1 _17828_ (.Y(_10784_),
    .A(net2372));
 sg13g2_inv_2 _17829_ (.Y(_10785_),
    .A(net2985));
 sg13g2_inv_1 _17830_ (.Y(_10786_),
    .A(net2595));
 sg13g2_inv_1 _17831_ (.Y(_10787_),
    .A(net3110));
 sg13g2_inv_1 _17832_ (.Y(_10788_),
    .A(net1976));
 sg13g2_inv_1 _17833_ (.Y(_10789_),
    .A(net2691));
 sg13g2_inv_1 _17834_ (.Y(_10790_),
    .A(net2887));
 sg13g2_inv_1 _17835_ (.Y(_10791_),
    .A(net2589));
 sg13g2_inv_1 _17836_ (.Y(_10792_),
    .A(net2324));
 sg13g2_inv_1 _17837_ (.Y(_10793_),
    .A(net2686));
 sg13g2_inv_1 _17838_ (.Y(_10794_),
    .A(\u_inv.f_reg[96] ));
 sg13g2_inv_1 _17839_ (.Y(_10795_),
    .A(\u_inv.f_reg[95] ));
 sg13g2_inv_1 _17840_ (.Y(_10796_),
    .A(net2169));
 sg13g2_inv_1 _17841_ (.Y(_10797_),
    .A(\u_inv.f_reg[93] ));
 sg13g2_inv_1 _17842_ (.Y(_10798_),
    .A(net2409));
 sg13g2_inv_1 _17843_ (.Y(_10799_),
    .A(net2942));
 sg13g2_inv_1 _17844_ (.Y(_10800_),
    .A(net2521));
 sg13g2_inv_1 _17845_ (.Y(_10801_),
    .A(\u_inv.f_reg[89] ));
 sg13g2_inv_2 _17846_ (.Y(_10802_),
    .A(net2377));
 sg13g2_inv_1 _17847_ (.Y(_10803_),
    .A(net2741));
 sg13g2_inv_1 _17848_ (.Y(_10804_),
    .A(net1900));
 sg13g2_inv_1 _17849_ (.Y(_10805_),
    .A(\u_inv.f_reg[85] ));
 sg13g2_inv_1 _17850_ (.Y(_10806_),
    .A(net2532));
 sg13g2_inv_1 _17851_ (.Y(_10807_),
    .A(net3186));
 sg13g2_inv_1 _17852_ (.Y(_10808_),
    .A(\u_inv.f_reg[82] ));
 sg13g2_inv_1 _17853_ (.Y(_10809_),
    .A(net2141));
 sg13g2_inv_1 _17854_ (.Y(_10810_),
    .A(\u_inv.f_reg[80] ));
 sg13g2_inv_1 _17855_ (.Y(_10811_),
    .A(\u_inv.f_reg[79] ));
 sg13g2_inv_1 _17856_ (.Y(_10812_),
    .A(\u_inv.f_reg[78] ));
 sg13g2_inv_1 _17857_ (.Y(_10813_),
    .A(\u_inv.f_reg[77] ));
 sg13g2_inv_1 _17858_ (.Y(_10814_),
    .A(net2302));
 sg13g2_inv_1 _17859_ (.Y(_10815_),
    .A(\u_inv.f_reg[75] ));
 sg13g2_inv_1 _17860_ (.Y(_10816_),
    .A(\u_inv.f_reg[74] ));
 sg13g2_inv_2 _17861_ (.Y(_10817_),
    .A(net2397));
 sg13g2_inv_1 _17862_ (.Y(_10818_),
    .A(net2553));
 sg13g2_inv_1 _17863_ (.Y(_10819_),
    .A(\u_inv.f_reg[71] ));
 sg13g2_inv_1 _17864_ (.Y(_10820_),
    .A(net1903));
 sg13g2_inv_1 _17865_ (.Y(_10821_),
    .A(\u_inv.f_reg[69] ));
 sg13g2_inv_1 _17866_ (.Y(_10822_),
    .A(net2707));
 sg13g2_inv_1 _17867_ (.Y(_10823_),
    .A(\u_inv.f_reg[67] ));
 sg13g2_inv_1 _17868_ (.Y(_10824_),
    .A(\u_inv.f_reg[66] ));
 sg13g2_inv_1 _17869_ (.Y(_10825_),
    .A(net2279));
 sg13g2_inv_1 _17870_ (.Y(_10826_),
    .A(net2660));
 sg13g2_inv_1 _17871_ (.Y(_10827_),
    .A(net3129));
 sg13g2_inv_1 _17872_ (.Y(_10828_),
    .A(net2941));
 sg13g2_inv_1 _17873_ (.Y(_10829_),
    .A(net2473));
 sg13g2_inv_1 _17874_ (.Y(_10830_),
    .A(net2355));
 sg13g2_inv_1 _17875_ (.Y(_10831_),
    .A(net2639));
 sg13g2_inv_1 _17876_ (.Y(_10832_),
    .A(net2199));
 sg13g2_inv_1 _17877_ (.Y(_10833_),
    .A(\u_inv.f_reg[57] ));
 sg13g2_inv_1 _17878_ (.Y(_10834_),
    .A(net3011));
 sg13g2_inv_1 _17879_ (.Y(_10835_),
    .A(\u_inv.f_reg[55] ));
 sg13g2_inv_1 _17880_ (.Y(_10836_),
    .A(net2551));
 sg13g2_inv_1 _17881_ (.Y(_10837_),
    .A(net3054));
 sg13g2_inv_1 _17882_ (.Y(_10838_),
    .A(net2755));
 sg13g2_inv_1 _17883_ (.Y(_10839_),
    .A(net2754));
 sg13g2_inv_1 _17884_ (.Y(_10840_),
    .A(net2293));
 sg13g2_inv_1 _17885_ (.Y(_10841_),
    .A(net2261));
 sg13g2_inv_1 _17886_ (.Y(_10842_),
    .A(\u_inv.f_reg[48] ));
 sg13g2_inv_1 _17887_ (.Y(_10843_),
    .A(net2920));
 sg13g2_inv_1 _17888_ (.Y(_10844_),
    .A(net2456));
 sg13g2_inv_1 _17889_ (.Y(_10845_),
    .A(\u_inv.f_reg[45] ));
 sg13g2_inv_1 _17890_ (.Y(_10846_),
    .A(net2259));
 sg13g2_inv_1 _17891_ (.Y(_10847_),
    .A(net3253));
 sg13g2_inv_1 _17892_ (.Y(_10848_),
    .A(net2466));
 sg13g2_inv_1 _17893_ (.Y(_10849_),
    .A(net2634));
 sg13g2_inv_1 _17894_ (.Y(_10850_),
    .A(net2285));
 sg13g2_inv_1 _17895_ (.Y(_10851_),
    .A(\u_inv.f_reg[39] ));
 sg13g2_inv_2 _17896_ (.Y(_10852_),
    .A(net2153));
 sg13g2_inv_1 _17897_ (.Y(_10853_),
    .A(net2502));
 sg13g2_inv_1 _17898_ (.Y(_10854_),
    .A(net2969));
 sg13g2_inv_1 _17899_ (.Y(_10855_),
    .A(\u_inv.f_reg[35] ));
 sg13g2_inv_1 _17900_ (.Y(_10856_),
    .A(net2710));
 sg13g2_inv_1 _17901_ (.Y(_10857_),
    .A(net2091));
 sg13g2_inv_1 _17902_ (.Y(_10858_),
    .A(\u_inv.f_reg[31] ));
 sg13g2_inv_1 _17903_ (.Y(_10859_),
    .A(net2578));
 sg13g2_inv_1 _17904_ (.Y(_10860_),
    .A(net3200));
 sg13g2_inv_1 _17905_ (.Y(_10861_),
    .A(net2517));
 sg13g2_inv_1 _17906_ (.Y(_10862_),
    .A(\u_inv.f_reg[27] ));
 sg13g2_inv_1 _17907_ (.Y(_10863_),
    .A(net2679));
 sg13g2_inv_1 _17908_ (.Y(_10864_),
    .A(net2974));
 sg13g2_inv_1 _17909_ (.Y(_10865_),
    .A(net2729));
 sg13g2_inv_1 _17910_ (.Y(_10866_),
    .A(\u_inv.f_reg[23] ));
 sg13g2_inv_1 _17911_ (.Y(_10867_),
    .A(net2227));
 sg13g2_inv_1 _17912_ (.Y(_10868_),
    .A(\u_inv.f_reg[21] ));
 sg13g2_inv_1 _17913_ (.Y(_10869_),
    .A(net2587));
 sg13g2_inv_1 _17914_ (.Y(_10870_),
    .A(net2047));
 sg13g2_inv_1 _17915_ (.Y(_10871_),
    .A(\u_inv.f_reg[18] ));
 sg13g2_inv_1 _17916_ (.Y(_10872_),
    .A(net2636));
 sg13g2_inv_1 _17917_ (.Y(_10873_),
    .A(net2718));
 sg13g2_inv_1 _17918_ (.Y(_10874_),
    .A(net2295));
 sg13g2_inv_1 _17919_ (.Y(_10875_),
    .A(net3088));
 sg13g2_inv_1 _17920_ (.Y(_10876_),
    .A(net2573));
 sg13g2_inv_1 _17921_ (.Y(_10877_),
    .A(net3121));
 sg13g2_inv_1 _17922_ (.Y(_10878_),
    .A(net3261));
 sg13g2_inv_1 _17923_ (.Y(_10879_),
    .A(\u_inv.f_reg[10] ));
 sg13g2_inv_1 _17924_ (.Y(_10880_),
    .A(\u_inv.f_reg[5] ));
 sg13g2_inv_1 _17925_ (.Y(_10881_),
    .A(\u_inv.f_reg[3] ));
 sg13g2_inv_1 _17926_ (.Y(_10882_),
    .A(net1984));
 sg13g2_inv_1 _17927_ (.Y(_10883_),
    .A(net2583));
 sg13g2_inv_1 _17928_ (.Y(_10884_),
    .A(\u_inv.d_reg[252] ));
 sg13g2_inv_1 _17929_ (.Y(_10885_),
    .A(\u_inv.d_reg[245] ));
 sg13g2_inv_2 _17930_ (.Y(_10886_),
    .A(\u_inv.d_reg[238] ));
 sg13g2_inv_1 _17931_ (.Y(_10887_),
    .A(\u_inv.d_reg[232] ));
 sg13g2_inv_4 _17932_ (.A(\u_inv.d_reg[223] ),
    .Y(_10888_));
 sg13g2_inv_4 _17933_ (.A(\u_inv.d_reg[222] ),
    .Y(_10889_));
 sg13g2_inv_1 _17934_ (.Y(_10890_),
    .A(\u_inv.d_reg[220] ));
 sg13g2_inv_2 _17935_ (.Y(_10891_),
    .A(\u_inv.d_reg[217] ));
 sg13g2_inv_2 _17936_ (.Y(_10892_),
    .A(\u_inv.d_reg[216] ));
 sg13g2_inv_1 _17937_ (.Y(_10893_),
    .A(\u_inv.d_reg[213] ));
 sg13g2_inv_2 _17938_ (.Y(_10894_),
    .A(\u_inv.d_reg[211] ));
 sg13g2_inv_2 _17939_ (.Y(_10895_),
    .A(\u_inv.d_reg[210] ));
 sg13g2_inv_2 _17940_ (.Y(_10896_),
    .A(\u_inv.d_reg[201] ));
 sg13g2_inv_1 _17941_ (.Y(_10897_),
    .A(\u_inv.d_reg[195] ));
 sg13g2_inv_2 _17942_ (.Y(_10898_),
    .A(\u_inv.d_reg[194] ));
 sg13g2_inv_1 _17943_ (.Y(_10899_),
    .A(\u_inv.d_reg[189] ));
 sg13g2_inv_1 _17944_ (.Y(_10900_),
    .A(\u_inv.d_reg[188] ));
 sg13g2_inv_1 _17945_ (.Y(_10901_),
    .A(\u_inv.d_reg[185] ));
 sg13g2_inv_1 _17946_ (.Y(_10902_),
    .A(\u_inv.d_reg[183] ));
 sg13g2_inv_2 _17947_ (.Y(_10903_),
    .A(\u_inv.d_reg[182] ));
 sg13g2_inv_1 _17948_ (.Y(_10904_),
    .A(\u_inv.d_reg[181] ));
 sg13g2_inv_1 _17949_ (.Y(_10905_),
    .A(\u_inv.d_reg[179] ));
 sg13g2_inv_1 _17950_ (.Y(_10906_),
    .A(\u_inv.d_reg[173] ));
 sg13g2_inv_1 _17951_ (.Y(_10907_),
    .A(\u_inv.d_reg[172] ));
 sg13g2_inv_2 _17952_ (.Y(_10908_),
    .A(\u_inv.d_reg[171] ));
 sg13g2_inv_2 _17953_ (.Y(_10909_),
    .A(\u_inv.d_reg[169] ));
 sg13g2_inv_1 _17954_ (.Y(_10910_),
    .A(\u_inv.d_reg[168] ));
 sg13g2_inv_2 _17955_ (.Y(_10911_),
    .A(\u_inv.d_reg[166] ));
 sg13g2_inv_1 _17956_ (.Y(_10912_),
    .A(\u_inv.d_reg[163] ));
 sg13g2_inv_1 _17957_ (.Y(_10913_),
    .A(\u_inv.d_reg[159] ));
 sg13g2_inv_1 _17958_ (.Y(_10914_),
    .A(\u_inv.d_reg[157] ));
 sg13g2_inv_2 _17959_ (.Y(_10915_),
    .A(\u_inv.d_reg[155] ));
 sg13g2_inv_1 _17960_ (.Y(_10916_),
    .A(\u_inv.d_reg[151] ));
 sg13g2_inv_2 _17961_ (.Y(_10917_),
    .A(\u_inv.d_reg[142] ));
 sg13g2_inv_2 _17962_ (.Y(_10918_),
    .A(\u_inv.d_reg[135] ));
 sg13g2_inv_1 _17963_ (.Y(_10919_),
    .A(net4779));
 sg13g2_inv_1 _17964_ (.Y(_10920_),
    .A(\u_inv.d_reg[127] ));
 sg13g2_inv_1 _17965_ (.Y(_10921_),
    .A(\u_inv.d_reg[121] ));
 sg13g2_inv_2 _17966_ (.Y(_10922_),
    .A(\u_inv.d_reg[111] ));
 sg13g2_inv_1 _17967_ (.Y(_10923_),
    .A(\u_inv.d_reg[109] ));
 sg13g2_inv_1 _17968_ (.Y(_10924_),
    .A(\u_inv.d_reg[105] ));
 sg13g2_inv_2 _17969_ (.Y(_10925_),
    .A(\u_inv.d_reg[103] ));
 sg13g2_inv_1 _17970_ (.Y(_10926_),
    .A(\u_inv.d_reg[98] ));
 sg13g2_inv_2 _17971_ (.Y(_10927_),
    .A(\u_inv.d_reg[95] ));
 sg13g2_inv_1 _17972_ (.Y(_10928_),
    .A(\u_inv.d_reg[90] ));
 sg13g2_inv_1 _17973_ (.Y(_10929_),
    .A(\u_inv.d_reg[85] ));
 sg13g2_inv_1 _17974_ (.Y(_10930_),
    .A(net4782));
 sg13g2_inv_1 _17975_ (.Y(_10931_),
    .A(\u_inv.d_reg[75] ));
 sg13g2_inv_2 _17976_ (.Y(_10932_),
    .A(\u_inv.d_reg[69] ));
 sg13g2_inv_1 _17977_ (.Y(_10933_),
    .A(\u_inv.d_reg[67] ));
 sg13g2_inv_2 _17978_ (.Y(_10934_),
    .A(\u_inv.d_reg[61] ));
 sg13g2_inv_1 _17979_ (.Y(_10935_),
    .A(\u_inv.d_reg[58] ));
 sg13g2_inv_1 _17980_ (.Y(_10936_),
    .A(\u_inv.d_reg[57] ));
 sg13g2_inv_1 _17981_ (.Y(_10937_),
    .A(\u_inv.d_reg[53] ));
 sg13g2_inv_2 _17982_ (.Y(_10938_),
    .A(\u_inv.d_reg[52] ));
 sg13g2_inv_1 _17983_ (.Y(_10939_),
    .A(\u_inv.d_reg[51] ));
 sg13g2_inv_1 _17984_ (.Y(_10940_),
    .A(\u_inv.d_reg[50] ));
 sg13g2_inv_1 _17985_ (.Y(_10941_),
    .A(\u_inv.d_reg[49] ));
 sg13g2_inv_1 _17986_ (.Y(_10942_),
    .A(\u_inv.d_reg[47] ));
 sg13g2_inv_1 _17987_ (.Y(_10943_),
    .A(\u_inv.d_reg[46] ));
 sg13g2_inv_1 _17988_ (.Y(_10944_),
    .A(\u_inv.d_reg[41] ));
 sg13g2_inv_1 _17989_ (.Y(_10945_),
    .A(\u_inv.d_reg[34] ));
 sg13g2_inv_2 _17990_ (.Y(_10946_),
    .A(\u_inv.d_reg[31] ));
 sg13g2_inv_2 _17991_ (.Y(_10947_),
    .A(\u_inv.d_reg[30] ));
 sg13g2_inv_1 _17992_ (.Y(_10948_),
    .A(\u_inv.d_reg[29] ));
 sg13g2_inv_1 _17993_ (.Y(_10949_),
    .A(\u_inv.d_reg[24] ));
 sg13g2_inv_1 _17994_ (.Y(_10950_),
    .A(net4791));
 sg13g2_inv_1 _17995_ (.Y(_10951_),
    .A(\u_inv.d_reg[16] ));
 sg13g2_inv_2 _17996_ (.Y(_10952_),
    .A(\u_inv.d_reg[15] ));
 sg13g2_inv_2 _17997_ (.Y(_10953_),
    .A(\u_inv.d_reg[14] ));
 sg13g2_inv_1 _17998_ (.Y(_10954_),
    .A(\u_inv.d_reg[12] ));
 sg13g2_inv_2 _17999_ (.Y(_10955_),
    .A(\u_inv.d_reg[9] ));
 sg13g2_inv_2 _18000_ (.Y(_10956_),
    .A(\u_inv.d_reg[8] ));
 sg13g2_inv_1 _18001_ (.Y(_10957_),
    .A(net1621));
 sg13g2_inv_1 _18002_ (.Y(_10958_),
    .A(net1811));
 sg13g2_inv_1 _18003_ (.Y(_10959_),
    .A(net1683));
 sg13g2_inv_1 _18004_ (.Y(_10960_),
    .A(net1758));
 sg13g2_inv_1 _18005_ (.Y(_10961_),
    .A(net1722));
 sg13g2_inv_1 _18006_ (.Y(_10962_),
    .A(net1695));
 sg13g2_inv_1 _18007_ (.Y(_10963_),
    .A(net1814));
 sg13g2_inv_1 _18008_ (.Y(_10964_),
    .A(net1720));
 sg13g2_inv_1 _18009_ (.Y(_10965_),
    .A(net1718));
 sg13g2_inv_1 _18010_ (.Y(_10966_),
    .A(net1750));
 sg13g2_inv_1 _18011_ (.Y(_10967_),
    .A(net1725));
 sg13g2_inv_1 _18012_ (.Y(_10968_),
    .A(net1801));
 sg13g2_inv_1 _18013_ (.Y(_10969_),
    .A(net1813));
 sg13g2_inv_1 _18014_ (.Y(_10970_),
    .A(net1715));
 sg13g2_inv_1 _18015_ (.Y(_10971_),
    .A(net1708));
 sg13g2_inv_1 _18016_ (.Y(_10972_),
    .A(net1974));
 sg13g2_inv_1 _18017_ (.Y(_10973_),
    .A(net1682));
 sg13g2_inv_1 _18018_ (.Y(_10974_),
    .A(net1888));
 sg13g2_inv_1 _18019_ (.Y(_10975_),
    .A(net2031));
 sg13g2_inv_1 _18020_ (.Y(_10976_),
    .A(net1894));
 sg13g2_inv_1 _18021_ (.Y(_10977_),
    .A(net2654));
 sg13g2_inv_1 _18022_ (.Y(_10978_),
    .A(net1740));
 sg13g2_inv_1 _18023_ (.Y(_10979_),
    .A(net2463));
 sg13g2_inv_1 _18024_ (.Y(_10980_),
    .A(net2016));
 sg13g2_inv_1 _18025_ (.Y(_10981_),
    .A(net2488));
 sg13g2_inv_1 _18026_ (.Y(_10982_),
    .A(net2006));
 sg13g2_inv_1 _18027_ (.Y(_10983_),
    .A(net1742));
 sg13g2_inv_1 _18028_ (.Y(_10984_),
    .A(net1732));
 sg13g2_inv_1 _18029_ (.Y(_10985_),
    .A(net1172));
 sg13g2_inv_1 _18030_ (.Y(_10986_),
    .A(net1893));
 sg13g2_inv_1 _18031_ (.Y(_10987_),
    .A(net1690));
 sg13g2_inv_1 _18032_ (.Y(_10988_),
    .A(net1491));
 sg13g2_inv_2 _18033_ (.Y(_10989_),
    .A(net1369));
 sg13g2_inv_1 _18034_ (.Y(_10990_),
    .A(net1850));
 sg13g2_inv_1 _18035_ (.Y(_10991_),
    .A(net1829));
 sg13g2_inv_2 _18036_ (.Y(_10992_),
    .A(net1169));
 sg13g2_inv_2 _18037_ (.Y(_10993_),
    .A(net1347));
 sg13g2_inv_2 _18038_ (.Y(_10994_),
    .A(net1190));
 sg13g2_inv_1 _18039_ (.Y(_10995_),
    .A(net1582));
 sg13g2_inv_2 _18040_ (.Y(_10996_),
    .A(net1509));
 sg13g2_inv_1 _18041_ (.Y(_10997_),
    .A(net1515));
 sg13g2_inv_1 _18042_ (.Y(_10998_),
    .A(net1505));
 sg13g2_inv_1 _18043_ (.Y(_10999_),
    .A(net1624));
 sg13g2_inv_1 _18044_ (.Y(_11000_),
    .A(net1245));
 sg13g2_inv_1 _18045_ (.Y(_11001_),
    .A(net1768));
 sg13g2_inv_1 _18046_ (.Y(_11002_),
    .A(net1298));
 sg13g2_inv_1 _18047_ (.Y(_11003_),
    .A(net1954));
 sg13g2_inv_2 _18048_ (.Y(_11004_),
    .A(net1264));
 sg13g2_inv_1 _18049_ (.Y(_11005_),
    .A(net1325));
 sg13g2_inv_2 _18050_ (.Y(_11006_),
    .A(net1367));
 sg13g2_inv_1 _18051_ (.Y(_11007_),
    .A(net1671));
 sg13g2_inv_2 _18052_ (.Y(_11008_),
    .A(net2418));
 sg13g2_inv_2 _18053_ (.Y(_11009_),
    .A(net1666));
 sg13g2_inv_1 _18054_ (.Y(_11010_),
    .A(net1746));
 sg13g2_inv_1 _18055_ (.Y(_11011_),
    .A(net1314));
 sg13g2_inv_1 _18056_ (.Y(_11012_),
    .A(net1279));
 sg13g2_inv_2 _18057_ (.Y(_11013_),
    .A(net1271));
 sg13g2_inv_1 _18058_ (.Y(_11014_),
    .A(net1246));
 sg13g2_inv_1 _18059_ (.Y(_11015_),
    .A(net2017));
 sg13g2_inv_1 _18060_ (.Y(_11016_),
    .A(net1738));
 sg13g2_inv_1 _18061_ (.Y(_11017_),
    .A(net1931));
 sg13g2_inv_1 _18062_ (.Y(_11018_),
    .A(net1655));
 sg13g2_inv_1 _18063_ (.Y(_11019_),
    .A(net1140));
 sg13g2_inv_1 _18064_ (.Y(_11020_),
    .A(net1881));
 sg13g2_inv_1 _18065_ (.Y(_11021_),
    .A(net1186));
 sg13g2_inv_1 _18066_ (.Y(_11022_),
    .A(net2208));
 sg13g2_inv_1 _18067_ (.Y(_11023_),
    .A(net1391));
 sg13g2_inv_1 _18068_ (.Y(_11024_),
    .A(net1516));
 sg13g2_inv_1 _18069_ (.Y(_11025_),
    .A(net1175));
 sg13g2_inv_1 _18070_ (.Y(_11026_),
    .A(net1401));
 sg13g2_inv_1 _18071_ (.Y(_11027_),
    .A(net1131));
 sg13g2_inv_1 _18072_ (.Y(_11028_),
    .A(net1561));
 sg13g2_inv_1 _18073_ (.Y(_11029_),
    .A(net1171));
 sg13g2_inv_1 _18074_ (.Y(_11030_),
    .A(net1114));
 sg13g2_inv_1 _18075_ (.Y(_11031_),
    .A(net1382));
 sg13g2_inv_1 _18076_ (.Y(_11032_),
    .A(net1079));
 sg13g2_inv_1 _18077_ (.Y(_11033_),
    .A(net1159));
 sg13g2_inv_2 _18078_ (.Y(_11034_),
    .A(net1569));
 sg13g2_inv_2 _18079_ (.Y(_11035_),
    .A(net1608));
 sg13g2_inv_2 _18080_ (.Y(_11036_),
    .A(net1237));
 sg13g2_inv_2 _18081_ (.Y(_11037_),
    .A(net1225));
 sg13g2_inv_2 _18082_ (.Y(_11038_),
    .A(net1142));
 sg13g2_inv_2 _18083_ (.Y(_11039_),
    .A(net1452));
 sg13g2_inv_2 _18084_ (.Y(_11040_),
    .A(net1438));
 sg13g2_nor2_2 _18085_ (.A(net2883),
    .B(net2072),
    .Y(uio_out[0]));
 sg13g2_nor2b_2 _18086_ (.A(\state[0] ),
    .B_N(\state[1] ),
    .Y(uio_out[1]));
 sg13g2_nor2_2 _18087_ (.A(_10626_),
    .B(\state[1] ),
    .Y(_11041_));
 sg13g2_nand2b_2 _18088_ (.Y(_11042_),
    .B(\state[0] ),
    .A_N(\state[1] ));
 sg13g2_nand2_2 _18089_ (.Y(_11043_),
    .A(net2221),
    .B(net4453));
 sg13g2_nand3_1 _18090_ (.B(net3298),
    .C(net4453),
    .A(\u_inv.state[1] ),
    .Y(_11044_));
 sg13g2_nand3_1 _18091_ (.B(net4964),
    .C(_11044_),
    .A(net4511),
    .Y(_11045_));
 sg13g2_inv_2 _18092_ (.Y(_17369_[0]),
    .A(net4965));
 sg13g2_nand2_2 _18093_ (.Y(_11046_),
    .A(net4511),
    .B(net2836));
 sg13g2_nand2_1 _18094_ (.Y(_00001_),
    .A(_11043_),
    .B(_11046_));
 sg13g2_and3_1 _18095_ (.X(_11047_),
    .A(net1294),
    .B(net1069),
    .C(net2011));
 sg13g2_nand3_1 _18096_ (.B(net1102),
    .C(_11047_),
    .A(net1215),
    .Y(_11048_));
 sg13g2_nand2b_2 _18097_ (.Y(_11049_),
    .B(net9),
    .A_N(net1533));
 sg13g2_nor2_2 _18098_ (.A(net4966),
    .B(_11049_),
    .Y(_11050_));
 sg13g2_nor3_1 _18099_ (.A(\state[0] ),
    .B(\state[1] ),
    .C(_11049_),
    .Y(_11051_));
 sg13g2_nor2b_1 _18100_ (.A(net1216),
    .B_N(_11051_),
    .Y(_00000_));
 sg13g2_a21oi_1 _18101_ (.A1(_10627_),
    .A2(_10632_),
    .Y(_00002_),
    .B1(net1063));
 sg13g2_nor2_1 _18102_ (.A(net2072),
    .B(net2221),
    .Y(_11052_));
 sg13g2_nor2_1 _18103_ (.A(uio_out[0]),
    .B(_11052_),
    .Y(_11053_));
 sg13g2_a221oi_1 _18104_ (.B2(_10626_),
    .C1(_11053_),
    .B1(_11049_),
    .A1(uio_out[0]),
    .Y(_00003_),
    .A2(net1216));
 sg13g2_a21oi_1 _18105_ (.A1(uio_out[1]),
    .A2(_11049_),
    .Y(_11054_),
    .B1(net4391));
 sg13g2_nor3_1 _18106_ (.A(uio_out[0]),
    .B(_11052_),
    .C(net1534),
    .Y(_00004_));
 sg13g2_nor2_1 _18107_ (.A(net1069),
    .B(_11050_),
    .Y(_11055_));
 sg13g2_a21oi_1 _18108_ (.A1(net1069),
    .A2(_11051_),
    .Y(_00005_),
    .B1(_11055_));
 sg13g2_and3_1 _18109_ (.X(_11056_),
    .A(net1294),
    .B(net1069),
    .C(_11050_));
 sg13g2_a21oi_1 _18110_ (.A1(net1069),
    .A2(_11050_),
    .Y(_11057_),
    .B1(net1294));
 sg13g2_and2_1 _18111_ (.A(net2072),
    .B(_11050_),
    .X(_11058_));
 sg13g2_nor3_1 _18112_ (.A(_11056_),
    .B(net1295),
    .C(_11058_),
    .Y(_00006_));
 sg13g2_xnor2_1 _18113_ (.Y(_11059_),
    .A(net2011),
    .B(_11056_));
 sg13g2_nor2_1 _18114_ (.A(_11058_),
    .B(_11059_),
    .Y(_00007_));
 sg13g2_and3_1 _18115_ (.X(_11060_),
    .A(net1102),
    .B(_11047_),
    .C(_11050_));
 sg13g2_a21oi_1 _18116_ (.A1(_11047_),
    .A2(_11051_),
    .Y(_11061_),
    .B1(net1102));
 sg13g2_nor3_1 _18117_ (.A(_11058_),
    .B(_11060_),
    .C(net1103),
    .Y(_00008_));
 sg13g2_xnor2_1 _18118_ (.Y(_11062_),
    .A(net1215),
    .B(_11060_));
 sg13g2_nor2_1 _18119_ (.A(_11058_),
    .B(_11062_),
    .Y(_00009_));
 sg13g2_nor2_2 _18120_ (.A(net4511),
    .B(\u_inv.state[1] ),
    .Y(_11063_));
 sg13g2_nand2b_1 _18121_ (.Y(_11064_),
    .B(net4601),
    .A_N(\u_inv.state[1] ));
 sg13g2_nand2_2 _18122_ (.Y(_11065_),
    .A(_11045_),
    .B(net4435));
 sg13g2_and2_1 _18123_ (.A(net4811),
    .B(_11065_),
    .X(_11066_));
 sg13g2_nand2_1 _18124_ (.Y(_11067_),
    .A(net4812),
    .B(_11065_));
 sg13g2_o21ai_1 _18125_ (.B1(net4000),
    .Y(_11068_),
    .A1(net4636),
    .A2(net4434));
 sg13g2_and2_1 _18126_ (.A(net4959),
    .B(_11068_),
    .X(_11069_));
 sg13g2_xnor2_1 _18127_ (.Y(_11070_),
    .A(\u_inv.f_next[256] ),
    .B(net4725));
 sg13g2_nand2_1 _18128_ (.Y(_11071_),
    .A(_10326_),
    .B(_10635_));
 sg13g2_xor2_1 _18129_ (.B(\u_inv.f_reg[255] ),
    .A(\u_inv.f_next[255] ),
    .X(_11072_));
 sg13g2_nand2_1 _18130_ (.Y(_11073_),
    .A(\u_inv.f_next[254] ),
    .B(_10636_));
 sg13g2_nand2_1 _18131_ (.Y(_11074_),
    .A(\u_inv.f_next[255] ),
    .B(_10635_));
 sg13g2_o21ai_1 _18132_ (.B1(_11074_),
    .Y(_11075_),
    .A1(_11072_),
    .A2(_11073_));
 sg13g2_nand2_1 _18133_ (.Y(_11076_),
    .A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ));
 sg13g2_xnor2_1 _18134_ (.Y(_11077_),
    .A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ));
 sg13g2_nor2b_1 _18135_ (.A(_11072_),
    .B_N(_11077_),
    .Y(_11078_));
 sg13g2_xor2_1 _18136_ (.B(\u_inv.f_reg[31] ),
    .A(\u_inv.f_next[31] ),
    .X(_11079_));
 sg13g2_xnor2_1 _18137_ (.Y(_11080_),
    .A(\u_inv.f_next[31] ),
    .B(\u_inv.f_reg[31] ));
 sg13g2_nand2_1 _18138_ (.Y(_11081_),
    .A(\u_inv.f_next[30] ),
    .B(\u_inv.f_reg[30] ));
 sg13g2_xor2_1 _18139_ (.B(\u_inv.f_reg[30] ),
    .A(\u_inv.f_next[30] ),
    .X(_11082_));
 sg13g2_xnor2_1 _18140_ (.Y(_11083_),
    .A(\u_inv.f_next[30] ),
    .B(\u_inv.f_reg[30] ));
 sg13g2_nor2_1 _18141_ (.A(_11079_),
    .B(_11082_),
    .Y(_11084_));
 sg13g2_xor2_1 _18142_ (.B(\u_inv.f_reg[29] ),
    .A(\u_inv.f_next[29] ),
    .X(_11085_));
 sg13g2_xnor2_1 _18143_ (.Y(_11086_),
    .A(\u_inv.f_next[29] ),
    .B(\u_inv.f_reg[29] ));
 sg13g2_nand2_1 _18144_ (.Y(_11087_),
    .A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ));
 sg13g2_xor2_1 _18145_ (.B(\u_inv.f_reg[28] ),
    .A(\u_inv.f_next[28] ),
    .X(_11088_));
 sg13g2_xnor2_1 _18146_ (.Y(_11089_),
    .A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ));
 sg13g2_nand3_1 _18147_ (.B(_11086_),
    .C(_11089_),
    .A(_11084_),
    .Y(_11090_));
 sg13g2_nand2_1 _18148_ (.Y(_11091_),
    .A(\u_inv.f_next[18] ),
    .B(\u_inv.f_reg[18] ));
 sg13g2_xor2_1 _18149_ (.B(\u_inv.f_reg[18] ),
    .A(\u_inv.f_next[18] ),
    .X(_11092_));
 sg13g2_inv_2 _18150_ (.Y(_11093_),
    .A(_11092_));
 sg13g2_xor2_1 _18151_ (.B(\u_inv.f_reg[17] ),
    .A(\u_inv.f_next[17] ),
    .X(_11094_));
 sg13g2_nor2_1 _18152_ (.A(\u_inv.f_next[19] ),
    .B(\u_inv.f_reg[19] ),
    .Y(_11095_));
 sg13g2_nand2_1 _18153_ (.Y(_11096_),
    .A(\u_inv.f_next[19] ),
    .B(\u_inv.f_reg[19] ));
 sg13g2_nor2b_2 _18154_ (.A(_11095_),
    .B_N(_11096_),
    .Y(_11097_));
 sg13g2_nand2b_2 _18155_ (.Y(_11098_),
    .B(_11096_),
    .A_N(_11095_));
 sg13g2_nand2_1 _18156_ (.Y(_11099_),
    .A(\u_inv.f_next[15] ),
    .B(\u_inv.f_reg[15] ));
 sg13g2_xnor2_1 _18157_ (.Y(_11100_),
    .A(\u_inv.f_next[15] ),
    .B(\u_inv.f_reg[15] ));
 sg13g2_nor2_1 _18158_ (.A(_10567_),
    .B(_10875_),
    .Y(_11101_));
 sg13g2_xor2_1 _18159_ (.B(\u_inv.f_reg[14] ),
    .A(\u_inv.f_next[14] ),
    .X(_11102_));
 sg13g2_xnor2_1 _18160_ (.Y(_11103_),
    .A(\u_inv.f_next[14] ),
    .B(\u_inv.f_reg[14] ));
 sg13g2_nor2_1 _18161_ (.A(\u_inv.f_next[13] ),
    .B(\u_inv.f_reg[13] ),
    .Y(_11104_));
 sg13g2_nand2_1 _18162_ (.Y(_11105_),
    .A(\u_inv.f_next[13] ),
    .B(\u_inv.f_reg[13] ));
 sg13g2_nand2b_2 _18163_ (.Y(_11106_),
    .B(_11105_),
    .A_N(_11104_));
 sg13g2_nand2_1 _18164_ (.Y(_11107_),
    .A(\u_inv.f_next[10] ),
    .B(\u_inv.f_reg[10] ));
 sg13g2_xor2_1 _18165_ (.B(\u_inv.f_reg[10] ),
    .A(\u_inv.f_next[10] ),
    .X(_11108_));
 sg13g2_inv_2 _18166_ (.Y(_11109_),
    .A(_11108_));
 sg13g2_nor2b_1 _18167_ (.A(\u_inv.f_reg[9] ),
    .B_N(\u_inv.f_next[9] ),
    .Y(_11110_));
 sg13g2_nor2_1 _18168_ (.A(\u_inv.f_next[9] ),
    .B(\u_inv.f_reg[9] ),
    .Y(_11111_));
 sg13g2_xor2_1 _18169_ (.B(\u_inv.f_reg[9] ),
    .A(\u_inv.f_next[9] ),
    .X(_11112_));
 sg13g2_and2_1 _18170_ (.A(\u_inv.f_next[8] ),
    .B(\u_inv.f_reg[8] ),
    .X(_11113_));
 sg13g2_xor2_1 _18171_ (.B(\u_inv.f_reg[8] ),
    .A(\u_inv.f_next[8] ),
    .X(_11114_));
 sg13g2_nand2b_1 _18172_ (.Y(_11115_),
    .B(\u_inv.f_next[7] ),
    .A_N(\u_inv.f_reg[7] ));
 sg13g2_nand2_1 _18173_ (.Y(_11116_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_xnor2_1 _18174_ (.Y(_11117_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_nor2_1 _18175_ (.A(_10572_),
    .B(\u_inv.f_reg[6] ),
    .Y(_11118_));
 sg13g2_xor2_1 _18176_ (.B(\u_inv.f_reg[6] ),
    .A(\u_inv.f_next[6] ),
    .X(_11119_));
 sg13g2_nand2_1 _18177_ (.Y(_11120_),
    .A(\u_inv.f_next[5] ),
    .B(_10880_));
 sg13g2_nand2_1 _18178_ (.Y(_11121_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_xnor2_1 _18179_ (.Y(_11122_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_nor2b_1 _18180_ (.A(\u_inv.f_reg[4] ),
    .B_N(\u_inv.f_next[4] ),
    .Y(_11123_));
 sg13g2_xor2_1 _18181_ (.B(\u_inv.f_reg[4] ),
    .A(\u_inv.f_next[4] ),
    .X(_11124_));
 sg13g2_nand2_1 _18182_ (.Y(_11125_),
    .A(\u_inv.f_next[3] ),
    .B(_10881_));
 sg13g2_nand2_1 _18183_ (.Y(_11126_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_xnor2_1 _18184_ (.Y(_11127_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_nor2_1 _18185_ (.A(_10575_),
    .B(\u_inv.f_reg[2] ),
    .Y(_11128_));
 sg13g2_nand2_1 _18186_ (.Y(_11129_),
    .A(\u_inv.f_next[2] ),
    .B(\u_inv.f_reg[2] ));
 sg13g2_inv_1 _18187_ (.Y(_11130_),
    .A(_11129_));
 sg13g2_or2_1 _18188_ (.X(_11131_),
    .B(\u_inv.f_reg[2] ),
    .A(\u_inv.f_next[2] ));
 sg13g2_and2_1 _18189_ (.A(_11129_),
    .B(_11131_),
    .X(_11132_));
 sg13g2_nor2b_1 _18190_ (.A(\u_inv.f_next[1] ),
    .B_N(\u_inv.f_reg[1] ),
    .Y(_11133_));
 sg13g2_nand2b_1 _18191_ (.Y(_11134_),
    .B(\u_inv.f_next[1] ),
    .A_N(\u_inv.f_reg[1] ));
 sg13g2_nor2b_1 _18192_ (.A(net4638),
    .B_N(\u_inv.f_reg[0] ),
    .Y(_11135_));
 sg13g2_a21oi_1 _18193_ (.A1(_11134_),
    .A2(_11135_),
    .Y(_11136_),
    .B1(_11133_));
 sg13g2_a221oi_1 _18194_ (.B2(_11135_),
    .C1(_11133_),
    .B1(_11134_),
    .A1(_11129_),
    .Y(_11137_),
    .A2(_11131_));
 sg13g2_o21ai_1 _18195_ (.B1(_11127_),
    .Y(_11138_),
    .A1(_11128_),
    .A2(_11137_));
 sg13g2_a21oi_1 _18196_ (.A1(_11125_),
    .A2(_11138_),
    .Y(_11139_),
    .B1(_11124_));
 sg13g2_o21ai_1 _18197_ (.B1(_11122_),
    .Y(_11140_),
    .A1(_11123_),
    .A2(_11139_));
 sg13g2_a21oi_1 _18198_ (.A1(_11120_),
    .A2(_11140_),
    .Y(_11141_),
    .B1(_11119_));
 sg13g2_o21ai_1 _18199_ (.B1(_11117_),
    .Y(_11142_),
    .A1(_11118_),
    .A2(_11141_));
 sg13g2_a21o_1 _18200_ (.A2(_11142_),
    .A1(_11115_),
    .B1(_11114_),
    .X(_11143_));
 sg13g2_nand2b_1 _18201_ (.Y(_11144_),
    .B(\u_inv.f_next[8] ),
    .A_N(\u_inv.f_reg[8] ));
 sg13g2_a21oi_1 _18202_ (.A1(_11143_),
    .A2(_11144_),
    .Y(_11145_),
    .B1(_11112_));
 sg13g2_o21ai_1 _18203_ (.B1(_11109_),
    .Y(_11146_),
    .A1(_11110_),
    .A2(_11145_));
 sg13g2_inv_1 _18204_ (.Y(_11147_),
    .A(_11146_));
 sg13g2_o21ai_1 _18205_ (.B1(_11146_),
    .Y(_11148_),
    .A1(_10571_),
    .A2(\u_inv.f_reg[10] ));
 sg13g2_a22oi_1 _18206_ (.Y(_11149_),
    .B1(_10879_),
    .B2(\u_inv.f_next[10] ),
    .A2(_10878_),
    .A1(\u_inv.f_next[11] ));
 sg13g2_nand2_1 _18207_ (.Y(_11150_),
    .A(_11146_),
    .B(_11149_));
 sg13g2_o21ai_1 _18208_ (.B1(_11150_),
    .Y(_11151_),
    .A1(\u_inv.f_next[11] ),
    .A2(_10878_));
 sg13g2_nand2_1 _18209_ (.Y(_11152_),
    .A(\u_inv.f_next[12] ),
    .B(\u_inv.f_reg[12] ));
 sg13g2_xor2_1 _18210_ (.B(\u_inv.f_reg[12] ),
    .A(\u_inv.f_next[12] ),
    .X(_11153_));
 sg13g2_xnor2_1 _18211_ (.Y(_11154_),
    .A(\u_inv.f_next[12] ),
    .B(\u_inv.f_reg[12] ));
 sg13g2_nand2b_1 _18212_ (.Y(_11155_),
    .B(_11154_),
    .A_N(_11151_));
 sg13g2_nand2b_1 _18213_ (.Y(_11156_),
    .B(_11106_),
    .A_N(_11155_));
 sg13g2_nand4_1 _18214_ (.B(_11103_),
    .C(_11106_),
    .A(_11100_),
    .Y(_11157_),
    .D(_11154_));
 sg13g2_a221oi_1 _18215_ (.B2(_11149_),
    .C1(_11157_),
    .B1(_11146_),
    .A1(_10570_),
    .Y(_11158_),
    .A2(\u_inv.f_reg[11] ));
 sg13g2_nand2_1 _18216_ (.Y(_11159_),
    .A(\u_inv.f_next[14] ),
    .B(_10875_));
 sg13g2_nand2_1 _18217_ (.Y(_11160_),
    .A(\u_inv.f_next[13] ),
    .B(_10876_));
 sg13g2_nand3_1 _18218_ (.B(_10877_),
    .C(_11106_),
    .A(\u_inv.f_next[12] ),
    .Y(_11161_));
 sg13g2_and2_1 _18219_ (.A(_11160_),
    .B(_11161_),
    .X(_11162_));
 sg13g2_o21ai_1 _18220_ (.B1(_11159_),
    .Y(_11163_),
    .A1(_11102_),
    .A2(_11162_));
 sg13g2_nand2_1 _18221_ (.Y(_11164_),
    .A(_11100_),
    .B(_11163_));
 sg13g2_o21ai_1 _18222_ (.B1(_11164_),
    .Y(_11165_),
    .A1(_10566_),
    .A2(\u_inv.f_reg[15] ));
 sg13g2_nor2_1 _18223_ (.A(_11158_),
    .B(_11165_),
    .Y(_11166_));
 sg13g2_nor2_1 _18224_ (.A(_10565_),
    .B(_10873_),
    .Y(_11167_));
 sg13g2_xor2_1 _18225_ (.B(\u_inv.f_reg[16] ),
    .A(\u_inv.f_next[16] ),
    .X(_11168_));
 sg13g2_nor2_1 _18226_ (.A(_11166_),
    .B(_11168_),
    .Y(_11169_));
 sg13g2_inv_1 _18227_ (.Y(_11170_),
    .A(_11169_));
 sg13g2_nor4_1 _18228_ (.A(_11092_),
    .B(_11094_),
    .C(_11097_),
    .D(_11168_),
    .Y(_11171_));
 sg13g2_o21ai_1 _18229_ (.B1(_11171_),
    .Y(_11172_),
    .A1(_11158_),
    .A2(_11165_));
 sg13g2_nor2_1 _18230_ (.A(_10562_),
    .B(\u_inv.f_reg[19] ),
    .Y(_11173_));
 sg13g2_nand2_1 _18231_ (.Y(_11174_),
    .A(\u_inv.f_next[18] ),
    .B(_10871_));
 sg13g2_nor2_1 _18232_ (.A(_10564_),
    .B(\u_inv.f_reg[17] ),
    .Y(_11175_));
 sg13g2_nand2_1 _18233_ (.Y(_11176_),
    .A(\u_inv.f_next[16] ),
    .B(_10873_));
 sg13g2_nor2_1 _18234_ (.A(_11094_),
    .B(_11176_),
    .Y(_11177_));
 sg13g2_o21ai_1 _18235_ (.B1(_11093_),
    .Y(_11178_),
    .A1(_11175_),
    .A2(_11177_));
 sg13g2_nand2_1 _18236_ (.Y(_11179_),
    .A(_11174_),
    .B(_11178_));
 sg13g2_a21oi_1 _18237_ (.A1(_11098_),
    .A2(_11179_),
    .Y(_11180_),
    .B1(_11173_));
 sg13g2_nand2_1 _18238_ (.Y(_11181_),
    .A(\u_inv.f_next[20] ),
    .B(\u_inv.f_reg[20] ));
 sg13g2_xor2_1 _18239_ (.B(\u_inv.f_reg[20] ),
    .A(\u_inv.f_next[20] ),
    .X(_11182_));
 sg13g2_xnor2_1 _18240_ (.Y(_11183_),
    .A(\u_inv.f_next[20] ),
    .B(\u_inv.f_reg[20] ));
 sg13g2_a21oi_1 _18241_ (.A1(_11172_),
    .A2(_11180_),
    .Y(_11184_),
    .B1(_11182_));
 sg13g2_nand2_1 _18242_ (.Y(_11185_),
    .A(\u_inv.f_next[22] ),
    .B(\u_inv.f_reg[22] ));
 sg13g2_xor2_1 _18243_ (.B(\u_inv.f_reg[22] ),
    .A(\u_inv.f_next[22] ),
    .X(_11186_));
 sg13g2_xnor2_1 _18244_ (.Y(_11187_),
    .A(\u_inv.f_next[21] ),
    .B(\u_inv.f_reg[21] ));
 sg13g2_xor2_1 _18245_ (.B(\u_inv.f_reg[23] ),
    .A(\u_inv.f_next[23] ),
    .X(_11188_));
 sg13g2_inv_1 _18246_ (.Y(_11189_),
    .A(_11188_));
 sg13g2_nor2_1 _18247_ (.A(_11186_),
    .B(_11188_),
    .Y(_11190_));
 sg13g2_nand3_1 _18248_ (.B(_11187_),
    .C(_11190_),
    .A(_11183_),
    .Y(_11191_));
 sg13g2_a21o_1 _18249_ (.A2(_11180_),
    .A1(_11172_),
    .B1(_11191_),
    .X(_11192_));
 sg13g2_nor2_1 _18250_ (.A(_10558_),
    .B(\u_inv.f_reg[23] ),
    .Y(_11193_));
 sg13g2_nor2_1 _18251_ (.A(_10559_),
    .B(\u_inv.f_reg[22] ),
    .Y(_11194_));
 sg13g2_nand2_1 _18252_ (.Y(_11195_),
    .A(\u_inv.f_next[21] ),
    .B(_10868_));
 sg13g2_nor2_1 _18253_ (.A(_10561_),
    .B(\u_inv.f_reg[20] ),
    .Y(_11196_));
 sg13g2_nand2_1 _18254_ (.Y(_11197_),
    .A(_11187_),
    .B(_11196_));
 sg13g2_nand2_1 _18255_ (.Y(_11198_),
    .A(_11195_),
    .B(_11197_));
 sg13g2_a221oi_1 _18256_ (.B2(_11190_),
    .C1(_11193_),
    .B1(_11198_),
    .A1(_11189_),
    .Y(_11199_),
    .A2(_11194_));
 sg13g2_and2_1 _18257_ (.A(_11192_),
    .B(_11199_),
    .X(_11200_));
 sg13g2_xnor2_1 _18258_ (.Y(_11201_),
    .A(\u_inv.f_next[24] ),
    .B(\u_inv.f_reg[24] ));
 sg13g2_inv_1 _18259_ (.Y(_11202_),
    .A(_11201_));
 sg13g2_xor2_1 _18260_ (.B(\u_inv.f_reg[25] ),
    .A(\u_inv.f_next[25] ),
    .X(_11203_));
 sg13g2_xnor2_1 _18261_ (.Y(_11204_),
    .A(\u_inv.f_next[25] ),
    .B(\u_inv.f_reg[25] ));
 sg13g2_nor2_1 _18262_ (.A(_10555_),
    .B(_10863_),
    .Y(_11205_));
 sg13g2_xnor2_1 _18263_ (.Y(_11206_),
    .A(\u_inv.f_next[26] ),
    .B(\u_inv.f_reg[26] ));
 sg13g2_inv_2 _18264_ (.Y(_11207_),
    .A(_11206_));
 sg13g2_xor2_1 _18265_ (.B(\u_inv.f_reg[27] ),
    .A(\u_inv.f_next[27] ),
    .X(_11208_));
 sg13g2_nor2_1 _18266_ (.A(_11207_),
    .B(_11208_),
    .Y(_11209_));
 sg13g2_nand3_1 _18267_ (.B(_11204_),
    .C(_11209_),
    .A(_11201_),
    .Y(_11210_));
 sg13g2_nor2_1 _18268_ (.A(_11200_),
    .B(_11210_),
    .Y(_11211_));
 sg13g2_or2_1 _18269_ (.X(_11212_),
    .B(_11210_),
    .A(_11090_));
 sg13g2_a21oi_2 _18270_ (.B1(_11212_),
    .Y(_11213_),
    .A2(_11199_),
    .A1(_11192_));
 sg13g2_nand2_1 _18271_ (.Y(_11214_),
    .A(\u_inv.f_next[29] ),
    .B(_10860_));
 sg13g2_nor2_1 _18272_ (.A(_10553_),
    .B(\u_inv.f_reg[28] ),
    .Y(_11215_));
 sg13g2_nand2_1 _18273_ (.Y(_11216_),
    .A(\u_inv.f_next[24] ),
    .B(_10865_));
 sg13g2_nand2_1 _18274_ (.Y(_11217_),
    .A(\u_inv.f_next[26] ),
    .B(_10863_));
 sg13g2_nand2_1 _18275_ (.Y(_11218_),
    .A(\u_inv.f_next[27] ),
    .B(_10862_));
 sg13g2_o21ai_1 _18276_ (.B1(_11218_),
    .Y(_11219_),
    .A1(_11208_),
    .A2(_11217_));
 sg13g2_nor2_1 _18277_ (.A(_10556_),
    .B(\u_inv.f_reg[25] ),
    .Y(_11220_));
 sg13g2_nor2_1 _18278_ (.A(_11203_),
    .B(_11216_),
    .Y(_11221_));
 sg13g2_o21ai_1 _18279_ (.B1(_11209_),
    .Y(_11222_),
    .A1(_11220_),
    .A2(_11221_));
 sg13g2_nand2b_1 _18280_ (.Y(_11223_),
    .B(_11222_),
    .A_N(_11219_));
 sg13g2_a21oi_1 _18281_ (.A1(_11089_),
    .A2(_11223_),
    .Y(_11224_),
    .B1(_11215_));
 sg13g2_o21ai_1 _18282_ (.B1(_11214_),
    .Y(_11225_),
    .A1(_11085_),
    .A2(_11224_));
 sg13g2_nor2_1 _18283_ (.A(_10551_),
    .B(\u_inv.f_reg[30] ),
    .Y(_11226_));
 sg13g2_nor2_1 _18284_ (.A(_10550_),
    .B(\u_inv.f_reg[31] ),
    .Y(_11227_));
 sg13g2_a221oi_1 _18285_ (.B2(_11080_),
    .C1(_11227_),
    .B1(_11226_),
    .A1(_11084_),
    .Y(_11228_),
    .A2(_11225_));
 sg13g2_inv_1 _18286_ (.Y(_11229_),
    .A(_11228_));
 sg13g2_nand2b_2 _18287_ (.Y(_11230_),
    .B(_11228_),
    .A_N(_11213_));
 sg13g2_xor2_1 _18288_ (.B(\u_inv.f_reg[35] ),
    .A(\u_inv.f_next[35] ),
    .X(_11231_));
 sg13g2_xor2_1 _18289_ (.B(\u_inv.f_reg[34] ),
    .A(\u_inv.f_next[34] ),
    .X(_11232_));
 sg13g2_nor2_1 _18290_ (.A(_11231_),
    .B(_11232_),
    .Y(_11233_));
 sg13g2_nand2_1 _18291_ (.Y(_11234_),
    .A(\u_inv.f_next[32] ),
    .B(\u_inv.f_reg[32] ));
 sg13g2_xnor2_1 _18292_ (.Y(_11235_),
    .A(\u_inv.f_next[32] ),
    .B(\u_inv.f_reg[32] ));
 sg13g2_inv_1 _18293_ (.Y(_11236_),
    .A(_11235_));
 sg13g2_nor2_2 _18294_ (.A(\u_inv.f_next[33] ),
    .B(\u_inv.f_reg[33] ),
    .Y(_11237_));
 sg13g2_nand2_1 _18295_ (.Y(_11238_),
    .A(\u_inv.f_next[33] ),
    .B(\u_inv.f_reg[33] ));
 sg13g2_nor2b_2 _18296_ (.A(_11237_),
    .B_N(_11238_),
    .Y(_11239_));
 sg13g2_nand2b_1 _18297_ (.Y(_11240_),
    .B(_11238_),
    .A_N(_11237_));
 sg13g2_nor4_1 _18298_ (.A(_11231_),
    .B(_11232_),
    .C(_11236_),
    .D(_11239_),
    .Y(_11241_));
 sg13g2_xor2_1 _18299_ (.B(\u_inv.f_reg[37] ),
    .A(\u_inv.f_next[37] ),
    .X(_11242_));
 sg13g2_xor2_1 _18300_ (.B(\u_inv.f_reg[36] ),
    .A(\u_inv.f_next[36] ),
    .X(_11243_));
 sg13g2_nor2_1 _18301_ (.A(_11242_),
    .B(_11243_),
    .Y(_11244_));
 sg13g2_nand2_1 _18302_ (.Y(_11245_),
    .A(_10542_),
    .B(_10851_));
 sg13g2_nor2_1 _18303_ (.A(_10542_),
    .B(_10851_),
    .Y(_11246_));
 sg13g2_xnor2_1 _18304_ (.Y(_11247_),
    .A(\u_inv.f_next[39] ),
    .B(\u_inv.f_reg[39] ));
 sg13g2_nor2_1 _18305_ (.A(_10543_),
    .B(_10852_),
    .Y(_11248_));
 sg13g2_nand2_1 _18306_ (.Y(_11249_),
    .A(_10543_),
    .B(_10852_));
 sg13g2_nand2b_2 _18307_ (.Y(_11250_),
    .B(_11249_),
    .A_N(_11248_));
 sg13g2_and2_1 _18308_ (.A(_11247_),
    .B(_11250_),
    .X(_11251_));
 sg13g2_and3_1 _18309_ (.X(_11252_),
    .A(_11241_),
    .B(_11244_),
    .C(_11251_));
 sg13g2_o21ai_1 _18310_ (.B1(_11252_),
    .Y(_11253_),
    .A1(_11213_),
    .A2(_11229_));
 sg13g2_nand2_1 _18311_ (.Y(_11254_),
    .A(\u_inv.f_next[35] ),
    .B(_10855_));
 sg13g2_nor2_1 _18312_ (.A(_10547_),
    .B(\u_inv.f_reg[34] ),
    .Y(_11255_));
 sg13g2_nor2_1 _18313_ (.A(_10548_),
    .B(\u_inv.f_reg[33] ),
    .Y(_11256_));
 sg13g2_nand2b_1 _18314_ (.Y(_11257_),
    .B(\u_inv.f_next[32] ),
    .A_N(\u_inv.f_reg[32] ));
 sg13g2_nor2_1 _18315_ (.A(_11239_),
    .B(_11257_),
    .Y(_11258_));
 sg13g2_o21ai_1 _18316_ (.B1(_11233_),
    .Y(_11259_),
    .A1(_11256_),
    .A2(_11258_));
 sg13g2_nand2b_1 _18317_ (.Y(_11260_),
    .B(_11255_),
    .A_N(_11231_));
 sg13g2_nand3_1 _18318_ (.B(_11259_),
    .C(_11260_),
    .A(_11254_),
    .Y(_11261_));
 sg13g2_nand2_1 _18319_ (.Y(_11262_),
    .A(\u_inv.f_next[36] ),
    .B(_10854_));
 sg13g2_nor2_1 _18320_ (.A(_10544_),
    .B(\u_inv.f_reg[37] ),
    .Y(_11263_));
 sg13g2_a21oi_1 _18321_ (.A1(_11244_),
    .A2(_11261_),
    .Y(_11264_),
    .B1(_11263_));
 sg13g2_o21ai_1 _18322_ (.B1(_11264_),
    .Y(_11265_),
    .A1(_11242_),
    .A2(_11262_));
 sg13g2_nand3_1 _18323_ (.B(_10852_),
    .C(_11247_),
    .A(\u_inv.f_next[38] ),
    .Y(_11266_));
 sg13g2_o21ai_1 _18324_ (.B1(_11266_),
    .Y(_11267_),
    .A1(_10542_),
    .A2(\u_inv.f_reg[39] ));
 sg13g2_a21o_1 _18325_ (.A2(_11265_),
    .A1(_11251_),
    .B1(_11267_),
    .X(_11268_));
 sg13g2_inv_2 _18326_ (.Y(_11269_),
    .A(_11268_));
 sg13g2_nand2_1 _18327_ (.Y(_11270_),
    .A(_11253_),
    .B(_11269_));
 sg13g2_inv_1 _18328_ (.Y(_11271_),
    .A(_11270_));
 sg13g2_nand2_1 _18329_ (.Y(_11272_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_xnor2_1 _18330_ (.Y(_11273_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_inv_1 _18331_ (.Y(_11274_),
    .A(_11273_));
 sg13g2_xor2_1 _18332_ (.B(\u_inv.f_reg[43] ),
    .A(\u_inv.f_next[43] ),
    .X(_11275_));
 sg13g2_xnor2_1 _18333_ (.Y(_11276_),
    .A(\u_inv.f_next[43] ),
    .B(\u_inv.f_reg[43] ));
 sg13g2_xnor2_1 _18334_ (.Y(_11277_),
    .A(\u_inv.f_next[40] ),
    .B(\u_inv.f_reg[40] ));
 sg13g2_xnor2_1 _18335_ (.Y(_11278_),
    .A(\u_inv.f_next[41] ),
    .B(\u_inv.f_reg[41] ));
 sg13g2_inv_1 _18336_ (.Y(_11279_),
    .A(_11278_));
 sg13g2_nand4_1 _18337_ (.B(_11276_),
    .C(_11277_),
    .A(_11273_),
    .Y(_11280_),
    .D(_11278_));
 sg13g2_xnor2_1 _18338_ (.Y(_11281_),
    .A(\u_inv.f_next[45] ),
    .B(\u_inv.f_reg[45] ));
 sg13g2_xnor2_1 _18339_ (.Y(_11282_),
    .A(\u_inv.f_next[44] ),
    .B(\u_inv.f_reg[44] ));
 sg13g2_nand2_1 _18340_ (.Y(_11283_),
    .A(_11281_),
    .B(_11282_));
 sg13g2_xor2_1 _18341_ (.B(\u_inv.f_reg[47] ),
    .A(\u_inv.f_next[47] ),
    .X(_11284_));
 sg13g2_xnor2_1 _18342_ (.Y(_11285_),
    .A(\u_inv.f_next[47] ),
    .B(\u_inv.f_reg[47] ));
 sg13g2_nand2_1 _18343_ (.Y(_11286_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_xor2_1 _18344_ (.B(\u_inv.f_reg[46] ),
    .A(\u_inv.f_next[46] ),
    .X(_11287_));
 sg13g2_xnor2_1 _18345_ (.Y(_11288_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_nor4_1 _18346_ (.A(_11280_),
    .B(_11283_),
    .C(_11284_),
    .D(_11287_),
    .Y(_11289_));
 sg13g2_inv_1 _18347_ (.Y(_11290_),
    .A(_11289_));
 sg13g2_a21oi_2 _18348_ (.B1(_11290_),
    .Y(_11291_),
    .A2(_11269_),
    .A1(_11253_));
 sg13g2_nor2_1 _18349_ (.A(_10540_),
    .B(\u_inv.f_reg[41] ),
    .Y(_11292_));
 sg13g2_nor2_1 _18350_ (.A(_10541_),
    .B(\u_inv.f_reg[40] ),
    .Y(_11293_));
 sg13g2_a21oi_1 _18351_ (.A1(_11278_),
    .A2(_11293_),
    .Y(_11294_),
    .B1(_11292_));
 sg13g2_nor3_1 _18352_ (.A(_11274_),
    .B(_11275_),
    .C(_11294_),
    .Y(_11295_));
 sg13g2_nand2_1 _18353_ (.Y(_11296_),
    .A(\u_inv.f_next[42] ),
    .B(_10848_));
 sg13g2_nand2_1 _18354_ (.Y(_11297_),
    .A(\u_inv.f_next[43] ),
    .B(_10847_));
 sg13g2_o21ai_1 _18355_ (.B1(_11297_),
    .Y(_11298_),
    .A1(_11275_),
    .A2(_11296_));
 sg13g2_nor2_1 _18356_ (.A(_11295_),
    .B(_11298_),
    .Y(_11299_));
 sg13g2_nor2_1 _18357_ (.A(_10537_),
    .B(\u_inv.f_reg[44] ),
    .Y(_11300_));
 sg13g2_nand2_1 _18358_ (.Y(_11301_),
    .A(\u_inv.f_next[45] ),
    .B(_10845_));
 sg13g2_o21ai_1 _18359_ (.B1(_11301_),
    .Y(_11302_),
    .A1(_11283_),
    .A2(_11299_));
 sg13g2_a21oi_1 _18360_ (.A1(_11281_),
    .A2(_11300_),
    .Y(_11303_),
    .B1(_11302_));
 sg13g2_nor2_1 _18361_ (.A(_10535_),
    .B(\u_inv.f_reg[46] ),
    .Y(_11304_));
 sg13g2_nor2_1 _18362_ (.A(_11287_),
    .B(_11303_),
    .Y(_11305_));
 sg13g2_o21ai_1 _18363_ (.B1(_11285_),
    .Y(_11306_),
    .A1(_11304_),
    .A2(_11305_));
 sg13g2_o21ai_1 _18364_ (.B1(_11306_),
    .Y(_11307_),
    .A1(_10534_),
    .A2(\u_inv.f_reg[47] ));
 sg13g2_or2_1 _18365_ (.X(_11308_),
    .B(_11307_),
    .A(_11291_));
 sg13g2_xor2_1 _18366_ (.B(\u_inv.f_reg[63] ),
    .A(\u_inv.f_next[63] ),
    .X(_11309_));
 sg13g2_xor2_1 _18367_ (.B(\u_inv.f_reg[62] ),
    .A(\u_inv.f_next[62] ),
    .X(_11310_));
 sg13g2_nor2_1 _18368_ (.A(_11309_),
    .B(_11310_),
    .Y(_11311_));
 sg13g2_xnor2_1 _18369_ (.Y(_11312_),
    .A(\u_inv.f_next[61] ),
    .B(\u_inv.f_reg[61] ));
 sg13g2_xnor2_1 _18370_ (.Y(_11313_),
    .A(\u_inv.f_next[60] ),
    .B(\u_inv.f_reg[60] ));
 sg13g2_nand3_1 _18371_ (.B(_11312_),
    .C(_11313_),
    .A(_11311_),
    .Y(_11314_));
 sg13g2_nand2_1 _18372_ (.Y(_11315_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_xnor2_1 _18373_ (.Y(_11316_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_xor2_1 _18374_ (.B(\u_inv.f_reg[57] ),
    .A(\u_inv.f_next[57] ),
    .X(_11317_));
 sg13g2_xnor2_1 _18375_ (.Y(_11318_),
    .A(\u_inv.f_next[59] ),
    .B(\u_inv.f_reg[59] ));
 sg13g2_and2_1 _18376_ (.A(_11316_),
    .B(_11318_),
    .X(_11319_));
 sg13g2_nand2b_1 _18377_ (.Y(_11320_),
    .B(_11319_),
    .A_N(_11317_));
 sg13g2_xor2_1 _18378_ (.B(\u_inv.f_reg[56] ),
    .A(\u_inv.f_next[56] ),
    .X(_11321_));
 sg13g2_nor3_1 _18379_ (.A(_11314_),
    .B(_11320_),
    .C(_11321_),
    .Y(_11322_));
 sg13g2_xnor2_1 _18380_ (.Y(_11323_),
    .A(\u_inv.f_next[48] ),
    .B(\u_inv.f_reg[48] ));
 sg13g2_xnor2_1 _18381_ (.Y(_11324_),
    .A(\u_inv.f_next[55] ),
    .B(\u_inv.f_reg[55] ));
 sg13g2_xnor2_1 _18382_ (.Y(_11325_),
    .A(\u_inv.f_next[54] ),
    .B(\u_inv.f_reg[54] ));
 sg13g2_nand2_1 _18383_ (.Y(_11326_),
    .A(_11324_),
    .B(_11325_));
 sg13g2_xor2_1 _18384_ (.B(\u_inv.f_reg[52] ),
    .A(\u_inv.f_next[52] ),
    .X(_11327_));
 sg13g2_xor2_1 _18385_ (.B(\u_inv.f_reg[53] ),
    .A(\u_inv.f_next[53] ),
    .X(_11328_));
 sg13g2_nor3_1 _18386_ (.A(_11326_),
    .B(_11327_),
    .C(_11328_),
    .Y(_11329_));
 sg13g2_xnor2_1 _18387_ (.Y(_11330_),
    .A(\u_inv.f_next[51] ),
    .B(\u_inv.f_reg[51] ));
 sg13g2_xnor2_1 _18388_ (.Y(_11331_),
    .A(\u_inv.f_next[50] ),
    .B(\u_inv.f_reg[50] ));
 sg13g2_nor2_1 _18389_ (.A(\u_inv.f_next[49] ),
    .B(\u_inv.f_reg[49] ),
    .Y(_11332_));
 sg13g2_xnor2_1 _18390_ (.Y(_11333_),
    .A(\u_inv.f_next[49] ),
    .B(\u_inv.f_reg[49] ));
 sg13g2_and4_1 _18391_ (.A(_11323_),
    .B(_11330_),
    .C(_11331_),
    .D(_11333_),
    .X(_11334_));
 sg13g2_and2_1 _18392_ (.A(_11329_),
    .B(_11334_),
    .X(_11335_));
 sg13g2_and2_1 _18393_ (.A(_11322_),
    .B(_11335_),
    .X(_11336_));
 sg13g2_o21ai_1 _18394_ (.B1(_11336_),
    .Y(_11337_),
    .A1(_11291_),
    .A2(_11307_));
 sg13g2_nor2_1 _18395_ (.A(_10526_),
    .B(\u_inv.f_reg[55] ),
    .Y(_11338_));
 sg13g2_nor2_1 _18396_ (.A(_10528_),
    .B(\u_inv.f_reg[53] ),
    .Y(_11339_));
 sg13g2_nand2_1 _18397_ (.Y(_11340_),
    .A(\u_inv.f_next[52] ),
    .B(_10838_));
 sg13g2_nor2_1 _18398_ (.A(_11328_),
    .B(_11340_),
    .Y(_11341_));
 sg13g2_nor2_1 _18399_ (.A(_10533_),
    .B(\u_inv.f_reg[48] ),
    .Y(_11342_));
 sg13g2_nor2_1 _18400_ (.A(_10531_),
    .B(\u_inv.f_reg[50] ),
    .Y(_11343_));
 sg13g2_nor2_1 _18401_ (.A(_10532_),
    .B(\u_inv.f_reg[49] ),
    .Y(_11344_));
 sg13g2_a21o_1 _18402_ (.A2(_11342_),
    .A1(_11333_),
    .B1(_11344_),
    .X(_11345_));
 sg13g2_and2_1 _18403_ (.A(_11331_),
    .B(_11345_),
    .X(_11346_));
 sg13g2_o21ai_1 _18404_ (.B1(_11330_),
    .Y(_11347_),
    .A1(_11343_),
    .A2(_11346_));
 sg13g2_o21ai_1 _18405_ (.B1(_11347_),
    .Y(_11348_),
    .A1(_10530_),
    .A2(\u_inv.f_reg[51] ));
 sg13g2_o21ai_1 _18406_ (.B1(_11325_),
    .Y(_11349_),
    .A1(_11339_),
    .A2(_11341_));
 sg13g2_o21ai_1 _18407_ (.B1(_11349_),
    .Y(_11350_),
    .A1(_10527_),
    .A2(\u_inv.f_reg[54] ));
 sg13g2_a221oi_1 _18408_ (.B2(_11324_),
    .C1(_11338_),
    .B1(_11350_),
    .A1(_11329_),
    .Y(_11351_),
    .A2(_11348_));
 sg13g2_inv_2 _18409_ (.Y(_11352_),
    .A(_11351_));
 sg13g2_nor2_1 _18410_ (.A(_10520_),
    .B(\u_inv.f_reg[61] ),
    .Y(_11353_));
 sg13g2_nor2_1 _18411_ (.A(_10521_),
    .B(\u_inv.f_reg[60] ),
    .Y(_11354_));
 sg13g2_a21o_1 _18412_ (.A2(_11354_),
    .A1(_11312_),
    .B1(_11353_),
    .X(_11355_));
 sg13g2_nand2_1 _18413_ (.Y(_11356_),
    .A(\u_inv.f_next[62] ),
    .B(_10828_));
 sg13g2_nor2_1 _18414_ (.A(_11309_),
    .B(_11356_),
    .Y(_11357_));
 sg13g2_a221oi_1 _18415_ (.B2(_11355_),
    .C1(_11357_),
    .B1(_11311_),
    .A1(\u_inv.f_next[63] ),
    .Y(_11358_),
    .A2(_10827_));
 sg13g2_nor2_1 _18416_ (.A(_10522_),
    .B(\u_inv.f_reg[59] ),
    .Y(_11359_));
 sg13g2_nor2_1 _18417_ (.A(_10523_),
    .B(\u_inv.f_reg[58] ),
    .Y(_11360_));
 sg13g2_nand2_1 _18418_ (.Y(_11361_),
    .A(\u_inv.f_next[57] ),
    .B(_10833_));
 sg13g2_nand2_1 _18419_ (.Y(_11362_),
    .A(\u_inv.f_next[56] ),
    .B(_10834_));
 sg13g2_o21ai_1 _18420_ (.B1(_11361_),
    .Y(_11363_),
    .A1(_11317_),
    .A2(_11362_));
 sg13g2_a221oi_1 _18421_ (.B2(_11319_),
    .C1(_11359_),
    .B1(_11363_),
    .A1(_11318_),
    .Y(_11364_),
    .A2(_11360_));
 sg13g2_o21ai_1 _18422_ (.B1(_11358_),
    .Y(_11365_),
    .A1(_11314_),
    .A2(_11364_));
 sg13g2_a21oi_2 _18423_ (.B1(_11365_),
    .Y(_11366_),
    .A2(_11352_),
    .A1(_11322_));
 sg13g2_nand2_1 _18424_ (.Y(_11367_),
    .A(_11337_),
    .B(_11366_));
 sg13g2_xor2_1 _18425_ (.B(\u_inv.f_reg[75] ),
    .A(\u_inv.f_next[75] ),
    .X(_11368_));
 sg13g2_nor2_1 _18426_ (.A(_10507_),
    .B(_10816_),
    .Y(_11369_));
 sg13g2_xor2_1 _18427_ (.B(\u_inv.f_reg[74] ),
    .A(\u_inv.f_next[74] ),
    .X(_11370_));
 sg13g2_nor2_1 _18428_ (.A(_11368_),
    .B(_11370_),
    .Y(_11371_));
 sg13g2_xor2_1 _18429_ (.B(\u_inv.f_reg[72] ),
    .A(\u_inv.f_next[72] ),
    .X(_11372_));
 sg13g2_xor2_1 _18430_ (.B(\u_inv.f_reg[73] ),
    .A(\u_inv.f_next[73] ),
    .X(_11373_));
 sg13g2_or4_1 _18431_ (.A(_11368_),
    .B(_11370_),
    .C(_11372_),
    .D(_11373_),
    .X(_11374_));
 sg13g2_nand2_1 _18432_ (.Y(_11375_),
    .A(\u_inv.f_next[79] ),
    .B(\u_inv.f_reg[79] ));
 sg13g2_xnor2_1 _18433_ (.Y(_11376_),
    .A(\u_inv.f_next[79] ),
    .B(\u_inv.f_reg[79] ));
 sg13g2_nor2_1 _18434_ (.A(_10503_),
    .B(_10812_),
    .Y(_11377_));
 sg13g2_xnor2_1 _18435_ (.Y(_11378_),
    .A(\u_inv.f_next[78] ),
    .B(\u_inv.f_reg[78] ));
 sg13g2_nand2_1 _18436_ (.Y(_11379_),
    .A(_11376_),
    .B(_11378_));
 sg13g2_xnor2_1 _18437_ (.Y(_11380_),
    .A(\u_inv.f_next[77] ),
    .B(\u_inv.f_reg[77] ));
 sg13g2_nand2_1 _18438_ (.Y(_11381_),
    .A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ));
 sg13g2_xnor2_1 _18439_ (.Y(_11382_),
    .A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ));
 sg13g2_nand2_1 _18440_ (.Y(_11383_),
    .A(_11380_),
    .B(_11382_));
 sg13g2_nor3_1 _18441_ (.A(_11374_),
    .B(_11379_),
    .C(_11383_),
    .Y(_11384_));
 sg13g2_xor2_1 _18442_ (.B(\u_inv.f_reg[67] ),
    .A(\u_inv.f_next[67] ),
    .X(_11385_));
 sg13g2_nor2_1 _18443_ (.A(_10515_),
    .B(_10824_),
    .Y(_11386_));
 sg13g2_xor2_1 _18444_ (.B(\u_inv.f_reg[66] ),
    .A(\u_inv.f_next[66] ),
    .X(_11387_));
 sg13g2_nor2_1 _18445_ (.A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ),
    .Y(_11388_));
 sg13g2_nand2_1 _18446_ (.Y(_11389_),
    .A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ));
 sg13g2_nor2b_2 _18447_ (.A(_11388_),
    .B_N(_11389_),
    .Y(_11390_));
 sg13g2_nand2_1 _18448_ (.Y(_11391_),
    .A(\u_inv.f_next[64] ),
    .B(\u_inv.f_reg[64] ));
 sg13g2_xor2_1 _18449_ (.B(\u_inv.f_reg[64] ),
    .A(\u_inv.f_next[64] ),
    .X(_11392_));
 sg13g2_nor4_1 _18450_ (.A(_11385_),
    .B(_11387_),
    .C(_11390_),
    .D(_11392_),
    .Y(_11393_));
 sg13g2_xor2_1 _18451_ (.B(\u_inv.f_reg[71] ),
    .A(\u_inv.f_next[71] ),
    .X(_11394_));
 sg13g2_inv_2 _18452_ (.Y(_11395_),
    .A(_11394_));
 sg13g2_nand2_1 _18453_ (.Y(_11396_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_xnor2_1 _18454_ (.Y(_11397_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_xor2_1 _18455_ (.B(\u_inv.f_reg[69] ),
    .A(\u_inv.f_next[69] ),
    .X(_11398_));
 sg13g2_nor2_1 _18456_ (.A(_10513_),
    .B(_10822_),
    .Y(_11399_));
 sg13g2_xor2_1 _18457_ (.B(\u_inv.f_reg[68] ),
    .A(\u_inv.f_next[68] ),
    .X(_11400_));
 sg13g2_nor2_1 _18458_ (.A(_11398_),
    .B(_11400_),
    .Y(_11401_));
 sg13g2_and4_1 _18459_ (.A(_11393_),
    .B(_11395_),
    .C(_11397_),
    .D(_11401_),
    .X(_11402_));
 sg13g2_and2_1 _18460_ (.A(_11384_),
    .B(_11402_),
    .X(_11403_));
 sg13g2_inv_1 _18461_ (.Y(_11404_),
    .A(_11403_));
 sg13g2_a21oi_2 _18462_ (.B1(_11404_),
    .Y(_11405_),
    .A2(_11366_),
    .A1(_11337_));
 sg13g2_nand2_1 _18463_ (.Y(_11406_),
    .A(\u_inv.f_next[77] ),
    .B(_10813_));
 sg13g2_nor2_1 _18464_ (.A(_10505_),
    .B(\u_inv.f_reg[76] ),
    .Y(_11407_));
 sg13g2_nor2_1 _18465_ (.A(_10507_),
    .B(net3099),
    .Y(_11408_));
 sg13g2_nand2_1 _18466_ (.Y(_11409_),
    .A(\u_inv.f_next[73] ),
    .B(_10817_));
 sg13g2_nand2_1 _18467_ (.Y(_11410_),
    .A(\u_inv.f_next[72] ),
    .B(_10818_));
 sg13g2_o21ai_1 _18468_ (.B1(_11409_),
    .Y(_11411_),
    .A1(_11373_),
    .A2(_11410_));
 sg13g2_nor3_1 _18469_ (.A(_10507_),
    .B(\u_inv.f_reg[74] ),
    .C(_11368_),
    .Y(_11412_));
 sg13g2_a221oi_1 _18470_ (.B2(_11411_),
    .C1(_11412_),
    .B1(_11371_),
    .A1(\u_inv.f_next[75] ),
    .Y(_11413_),
    .A2(_10815_));
 sg13g2_o21ai_1 _18471_ (.B1(_11406_),
    .Y(_11414_),
    .A1(_11383_),
    .A2(_11413_));
 sg13g2_a21oi_1 _18472_ (.A1(_11380_),
    .A2(_11407_),
    .Y(_11415_),
    .B1(_11414_));
 sg13g2_nand2_1 _18473_ (.Y(_11416_),
    .A(\u_inv.f_next[67] ),
    .B(_10823_));
 sg13g2_nor2_1 _18474_ (.A(_10515_),
    .B(\u_inv.f_reg[66] ),
    .Y(_11417_));
 sg13g2_nor3_1 _18475_ (.A(_10517_),
    .B(\u_inv.f_reg[64] ),
    .C(_11390_),
    .Y(_11418_));
 sg13g2_a21o_1 _18476_ (.A2(_10825_),
    .A1(\u_inv.f_next[65] ),
    .B1(_11418_),
    .X(_11419_));
 sg13g2_nor2b_1 _18477_ (.A(_11387_),
    .B_N(_11419_),
    .Y(_11420_));
 sg13g2_nor2_1 _18478_ (.A(_11417_),
    .B(_11420_),
    .Y(_11421_));
 sg13g2_o21ai_1 _18479_ (.B1(_11416_),
    .Y(_11422_),
    .A1(_11385_),
    .A2(_11421_));
 sg13g2_nand2_1 _18480_ (.Y(_11423_),
    .A(\u_inv.f_next[68] ),
    .B(_10822_));
 sg13g2_nor2_1 _18481_ (.A(_10512_),
    .B(\u_inv.f_reg[69] ),
    .Y(_11424_));
 sg13g2_a21oi_1 _18482_ (.A1(_11401_),
    .A2(_11422_),
    .Y(_11425_),
    .B1(_11424_));
 sg13g2_o21ai_1 _18483_ (.B1(_11425_),
    .Y(_11426_),
    .A1(_11398_),
    .A2(_11423_));
 sg13g2_nand2_1 _18484_ (.Y(_11427_),
    .A(\u_inv.f_next[71] ),
    .B(_10819_));
 sg13g2_nor2_1 _18485_ (.A(_10511_),
    .B(\u_inv.f_reg[70] ),
    .Y(_11428_));
 sg13g2_a21oi_1 _18486_ (.A1(_11397_),
    .A2(_11426_),
    .Y(_11429_),
    .B1(_11428_));
 sg13g2_o21ai_1 _18487_ (.B1(_11427_),
    .Y(_11430_),
    .A1(_11394_),
    .A2(_11429_));
 sg13g2_nor2_1 _18488_ (.A(_10503_),
    .B(\u_inv.f_reg[78] ),
    .Y(_11431_));
 sg13g2_and2_1 _18489_ (.A(_11376_),
    .B(_11431_),
    .X(_11432_));
 sg13g2_a221oi_1 _18490_ (.B2(_11430_),
    .C1(_11432_),
    .B1(_11384_),
    .A1(\u_inv.f_next[79] ),
    .Y(_11433_),
    .A2(_10811_));
 sg13g2_o21ai_1 _18491_ (.B1(_11433_),
    .Y(_11434_),
    .A1(_11379_),
    .A2(_11415_));
 sg13g2_nor2_2 _18492_ (.A(_11405_),
    .B(_11434_),
    .Y(_11435_));
 sg13g2_xnor2_1 _18493_ (.Y(_11436_),
    .A(\u_inv.f_next[95] ),
    .B(\u_inv.f_reg[95] ));
 sg13g2_nand2_1 _18494_ (.Y(_11437_),
    .A(\u_inv.f_next[94] ),
    .B(\u_inv.f_reg[94] ));
 sg13g2_xnor2_1 _18495_ (.Y(_11438_),
    .A(\u_inv.f_next[94] ),
    .B(\u_inv.f_reg[94] ));
 sg13g2_and2_1 _18496_ (.A(_11436_),
    .B(_11438_),
    .X(_11439_));
 sg13g2_xor2_1 _18497_ (.B(\u_inv.f_reg[93] ),
    .A(\u_inv.f_next[93] ),
    .X(_11440_));
 sg13g2_nor2_1 _18498_ (.A(_10489_),
    .B(_10798_),
    .Y(_11441_));
 sg13g2_xor2_1 _18499_ (.B(\u_inv.f_reg[92] ),
    .A(\u_inv.f_next[92] ),
    .X(_11442_));
 sg13g2_nor2_1 _18500_ (.A(_11440_),
    .B(_11442_),
    .Y(_11443_));
 sg13g2_nand2_1 _18501_ (.Y(_11444_),
    .A(_11439_),
    .B(_11443_));
 sg13g2_nand2_1 _18502_ (.Y(_11445_),
    .A(\u_inv.f_next[90] ),
    .B(\u_inv.f_reg[90] ));
 sg13g2_xor2_1 _18503_ (.B(\u_inv.f_reg[90] ),
    .A(\u_inv.f_next[90] ),
    .X(_11446_));
 sg13g2_xnor2_1 _18504_ (.Y(_11447_),
    .A(\u_inv.f_next[90] ),
    .B(\u_inv.f_reg[90] ));
 sg13g2_xor2_1 _18505_ (.B(\u_inv.f_reg[89] ),
    .A(\u_inv.f_next[89] ),
    .X(_11448_));
 sg13g2_xor2_1 _18506_ (.B(\u_inv.f_reg[91] ),
    .A(\u_inv.f_next[91] ),
    .X(_11449_));
 sg13g2_nor3_1 _18507_ (.A(_11446_),
    .B(_11448_),
    .C(_11449_),
    .Y(_11450_));
 sg13g2_nor2_1 _18508_ (.A(_10493_),
    .B(_10802_),
    .Y(_11451_));
 sg13g2_xor2_1 _18509_ (.B(\u_inv.f_reg[88] ),
    .A(\u_inv.f_next[88] ),
    .X(_11452_));
 sg13g2_nor2_1 _18510_ (.A(_11444_),
    .B(_11452_),
    .Y(_11453_));
 sg13g2_nand2_1 _18511_ (.Y(_11454_),
    .A(_11450_),
    .B(_11453_));
 sg13g2_xnor2_1 _18512_ (.Y(_11455_),
    .A(\u_inv.f_next[87] ),
    .B(\u_inv.f_reg[87] ));
 sg13g2_nand2_1 _18513_ (.Y(_11456_),
    .A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ));
 sg13g2_xnor2_1 _18514_ (.Y(_11457_),
    .A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ));
 sg13g2_and2_1 _18515_ (.A(_11455_),
    .B(_11457_),
    .X(_11458_));
 sg13g2_xnor2_1 _18516_ (.Y(_11459_),
    .A(\u_inv.f_next[84] ),
    .B(\u_inv.f_reg[84] ));
 sg13g2_xor2_1 _18517_ (.B(\u_inv.f_reg[85] ),
    .A(\u_inv.f_next[85] ),
    .X(_11460_));
 sg13g2_xnor2_1 _18518_ (.Y(_11461_),
    .A(\u_inv.f_next[85] ),
    .B(\u_inv.f_reg[85] ));
 sg13g2_nand3_1 _18519_ (.B(_11459_),
    .C(_11461_),
    .A(_11458_),
    .Y(_11462_));
 sg13g2_xor2_1 _18520_ (.B(\u_inv.f_reg[83] ),
    .A(\u_inv.f_next[83] ),
    .X(_11463_));
 sg13g2_xnor2_1 _18521_ (.Y(_11464_),
    .A(\u_inv.f_next[83] ),
    .B(\u_inv.f_reg[83] ));
 sg13g2_nand2_1 _18522_ (.Y(_11465_),
    .A(\u_inv.f_next[82] ),
    .B(\u_inv.f_reg[82] ));
 sg13g2_xnor2_1 _18523_ (.Y(_11466_),
    .A(\u_inv.f_next[82] ),
    .B(\u_inv.f_reg[82] ));
 sg13g2_and2_1 _18524_ (.A(_11464_),
    .B(_11466_),
    .X(_11467_));
 sg13g2_xnor2_1 _18525_ (.Y(_11468_),
    .A(\u_inv.f_next[80] ),
    .B(\u_inv.f_reg[80] ));
 sg13g2_nand2_1 _18526_ (.Y(_11469_),
    .A(_10500_),
    .B(_10809_));
 sg13g2_nand2_1 _18527_ (.Y(_11470_),
    .A(\u_inv.f_next[81] ),
    .B(\u_inv.f_reg[81] ));
 sg13g2_and2_1 _18528_ (.A(_11469_),
    .B(_11470_),
    .X(_11471_));
 sg13g2_nand3b_1 _18529_ (.B(_11467_),
    .C(_11468_),
    .Y(_11472_),
    .A_N(_11471_));
 sg13g2_nor2_1 _18530_ (.A(_11462_),
    .B(_11472_),
    .Y(_11473_));
 sg13g2_inv_1 _18531_ (.Y(_11474_),
    .A(_11473_));
 sg13g2_nand2b_1 _18532_ (.Y(_11475_),
    .B(_11473_),
    .A_N(_11454_));
 sg13g2_inv_1 _18533_ (.Y(_11476_),
    .A(_11475_));
 sg13g2_o21ai_1 _18534_ (.B1(_11476_),
    .Y(_11477_),
    .A1(_11405_),
    .A2(_11434_));
 sg13g2_nand2_1 _18535_ (.Y(_11478_),
    .A(\u_inv.f_next[82] ),
    .B(_10808_));
 sg13g2_nor2_1 _18536_ (.A(_10500_),
    .B(\u_inv.f_reg[81] ),
    .Y(_11479_));
 sg13g2_nand2_1 _18537_ (.Y(_11480_),
    .A(\u_inv.f_next[80] ),
    .B(_10810_));
 sg13g2_nor2_1 _18538_ (.A(_11471_),
    .B(_11480_),
    .Y(_11481_));
 sg13g2_o21ai_1 _18539_ (.B1(_11466_),
    .Y(_11482_),
    .A1(_11479_),
    .A2(_11481_));
 sg13g2_a21oi_1 _18540_ (.A1(_11478_),
    .A2(_11482_),
    .Y(_11483_),
    .B1(_11463_));
 sg13g2_a21oi_1 _18541_ (.A1(\u_inv.f_next[83] ),
    .A2(_10807_),
    .Y(_11484_),
    .B1(_11483_));
 sg13g2_nand2_1 _18542_ (.Y(_11485_),
    .A(\u_inv.f_next[85] ),
    .B(_10805_));
 sg13g2_nand2_1 _18543_ (.Y(_11486_),
    .A(\u_inv.f_next[84] ),
    .B(_10806_));
 sg13g2_o21ai_1 _18544_ (.B1(_11485_),
    .Y(_11487_),
    .A1(_11460_),
    .A2(_11486_));
 sg13g2_nor2_1 _18545_ (.A(_10495_),
    .B(\u_inv.f_reg[86] ),
    .Y(_11488_));
 sg13g2_nor2_1 _18546_ (.A(_10494_),
    .B(\u_inv.f_reg[87] ),
    .Y(_11489_));
 sg13g2_a21oi_1 _18547_ (.A1(_11455_),
    .A2(_11488_),
    .Y(_11490_),
    .B1(_11489_));
 sg13g2_o21ai_1 _18548_ (.B1(_11490_),
    .Y(_11491_),
    .A1(_11462_),
    .A2(_11484_));
 sg13g2_a21oi_1 _18549_ (.A1(_11458_),
    .A2(_11487_),
    .Y(_11492_),
    .B1(_11491_));
 sg13g2_nand2_1 _18550_ (.Y(_11493_),
    .A(\u_inv.f_next[93] ),
    .B(_10797_));
 sg13g2_nor2_1 _18551_ (.A(_10489_),
    .B(\u_inv.f_reg[92] ),
    .Y(_11494_));
 sg13g2_nand2b_1 _18552_ (.Y(_11495_),
    .B(_11494_),
    .A_N(_11440_));
 sg13g2_nand2_1 _18553_ (.Y(_11496_),
    .A(_11493_),
    .B(_11495_));
 sg13g2_nor2_1 _18554_ (.A(_10487_),
    .B(\u_inv.f_reg[94] ),
    .Y(_11497_));
 sg13g2_nand2_1 _18555_ (.Y(_11498_),
    .A(\u_inv.f_next[91] ),
    .B(_10799_));
 sg13g2_nor2_1 _18556_ (.A(_10491_),
    .B(\u_inv.f_reg[90] ),
    .Y(_11499_));
 sg13g2_nand2_1 _18557_ (.Y(_11500_),
    .A(\u_inv.f_next[89] ),
    .B(_10801_));
 sg13g2_nand2_1 _18558_ (.Y(_11501_),
    .A(\u_inv.f_next[88] ),
    .B(_10802_));
 sg13g2_o21ai_1 _18559_ (.B1(_11500_),
    .Y(_11502_),
    .A1(_11448_),
    .A2(_11501_));
 sg13g2_a21oi_1 _18560_ (.A1(_11447_),
    .A2(_11502_),
    .Y(_11503_),
    .B1(_11499_));
 sg13g2_o21ai_1 _18561_ (.B1(_11498_),
    .Y(_11504_),
    .A1(_11449_),
    .A2(_11503_));
 sg13g2_nor2b_1 _18562_ (.A(_11444_),
    .B_N(_11504_),
    .Y(_11505_));
 sg13g2_a221oi_1 _18563_ (.B2(_11496_),
    .C1(_11505_),
    .B1(_11439_),
    .A1(\u_inv.f_next[95] ),
    .Y(_11506_),
    .A2(_10795_));
 sg13g2_o21ai_1 _18564_ (.B1(_11506_),
    .Y(_11507_),
    .A1(_11454_),
    .A2(_11492_));
 sg13g2_a21oi_2 _18565_ (.B1(_11507_),
    .Y(_11508_),
    .A2(_11497_),
    .A1(_11436_));
 sg13g2_nand2_2 _18566_ (.Y(_11509_),
    .A(_11477_),
    .B(_11508_));
 sg13g2_xor2_1 _18567_ (.B(\u_inv.f_reg[123] ),
    .A(\u_inv.f_next[123] ),
    .X(_11510_));
 sg13g2_xnor2_1 _18568_ (.Y(_11511_),
    .A(\u_inv.f_next[123] ),
    .B(\u_inv.f_reg[123] ));
 sg13g2_xnor2_1 _18569_ (.Y(_11512_),
    .A(\u_inv.f_next[122] ),
    .B(\u_inv.f_reg[122] ));
 sg13g2_nand2_1 _18570_ (.Y(_11513_),
    .A(\u_inv.f_next[120] ),
    .B(\u_inv.f_reg[120] ));
 sg13g2_xnor2_1 _18571_ (.Y(_11514_),
    .A(\u_inv.f_next[120] ),
    .B(\u_inv.f_reg[120] ));
 sg13g2_nand2_1 _18572_ (.Y(_11515_),
    .A(\u_inv.f_next[121] ),
    .B(\u_inv.f_reg[121] ));
 sg13g2_nor2_1 _18573_ (.A(\u_inv.f_next[121] ),
    .B(\u_inv.f_reg[121] ),
    .Y(_11516_));
 sg13g2_xor2_1 _18574_ (.B(\u_inv.f_reg[121] ),
    .A(\u_inv.f_next[121] ),
    .X(_11517_));
 sg13g2_nand3_1 _18575_ (.B(_11512_),
    .C(_11514_),
    .A(_11511_),
    .Y(_11518_));
 sg13g2_nor2_1 _18576_ (.A(_11517_),
    .B(_11518_),
    .Y(_11519_));
 sg13g2_xnor2_1 _18577_ (.Y(_11520_),
    .A(\u_inv.f_next[127] ),
    .B(\u_inv.f_reg[127] ));
 sg13g2_nand2_1 _18578_ (.Y(_11521_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_xnor2_1 _18579_ (.Y(_11522_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_and2_1 _18580_ (.A(_11520_),
    .B(_11522_),
    .X(_11523_));
 sg13g2_xor2_1 _18581_ (.B(\u_inv.f_reg[125] ),
    .A(\u_inv.f_next[125] ),
    .X(_11524_));
 sg13g2_nor2_1 _18582_ (.A(_10457_),
    .B(_10766_),
    .Y(_11525_));
 sg13g2_xor2_1 _18583_ (.B(\u_inv.f_reg[124] ),
    .A(\u_inv.f_next[124] ),
    .X(_11526_));
 sg13g2_nor2_1 _18584_ (.A(_11524_),
    .B(_11526_),
    .Y(_11527_));
 sg13g2_nand3_1 _18585_ (.B(_11523_),
    .C(_11527_),
    .A(_11519_),
    .Y(_11528_));
 sg13g2_xor2_1 _18586_ (.B(\u_inv.f_reg[115] ),
    .A(\u_inv.f_next[115] ),
    .X(_11529_));
 sg13g2_nand2_1 _18587_ (.Y(_11530_),
    .A(\u_inv.f_next[114] ),
    .B(\u_inv.f_reg[114] ));
 sg13g2_xnor2_1 _18588_ (.Y(_11531_),
    .A(\u_inv.f_next[114] ),
    .B(\u_inv.f_reg[114] ));
 sg13g2_inv_2 _18589_ (.Y(_11532_),
    .A(_11531_));
 sg13g2_nor2_1 _18590_ (.A(_10469_),
    .B(_10778_),
    .Y(_11533_));
 sg13g2_xor2_1 _18591_ (.B(\u_inv.f_reg[112] ),
    .A(\u_inv.f_next[112] ),
    .X(_11534_));
 sg13g2_xor2_1 _18592_ (.B(\u_inv.f_reg[113] ),
    .A(\u_inv.f_next[113] ),
    .X(_11535_));
 sg13g2_or4_1 _18593_ (.A(_11529_),
    .B(_11532_),
    .C(_11534_),
    .D(_11535_),
    .X(_11536_));
 sg13g2_xnor2_1 _18594_ (.Y(_11537_),
    .A(\u_inv.f_next[119] ),
    .B(\u_inv.f_reg[119] ));
 sg13g2_nand2_1 _18595_ (.Y(_11538_),
    .A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ));
 sg13g2_xnor2_1 _18596_ (.Y(_11539_),
    .A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ));
 sg13g2_and2_1 _18597_ (.A(_11537_),
    .B(_11539_),
    .X(_11540_));
 sg13g2_xnor2_1 _18598_ (.Y(_11541_),
    .A(\u_inv.f_next[117] ),
    .B(\u_inv.f_reg[117] ));
 sg13g2_nor2_1 _18599_ (.A(_10465_),
    .B(_10774_),
    .Y(_11542_));
 sg13g2_xor2_1 _18600_ (.B(\u_inv.f_reg[116] ),
    .A(\u_inv.f_next[116] ),
    .X(_11543_));
 sg13g2_xnor2_1 _18601_ (.Y(_11544_),
    .A(\u_inv.f_next[116] ),
    .B(\u_inv.f_reg[116] ));
 sg13g2_nand3_1 _18602_ (.B(_11541_),
    .C(_11544_),
    .A(_11540_),
    .Y(_11545_));
 sg13g2_or2_1 _18603_ (.X(_11546_),
    .B(_11545_),
    .A(_11536_));
 sg13g2_nor2_2 _18604_ (.A(_11528_),
    .B(_11546_),
    .Y(_11547_));
 sg13g2_nor2_1 _18605_ (.A(\u_inv.f_next[111] ),
    .B(\u_inv.f_reg[111] ),
    .Y(_11548_));
 sg13g2_nand2_1 _18606_ (.Y(_11549_),
    .A(\u_inv.f_next[111] ),
    .B(\u_inv.f_reg[111] ));
 sg13g2_nor2b_2 _18607_ (.A(_11548_),
    .B_N(_11549_),
    .Y(_11550_));
 sg13g2_nand2_1 _18608_ (.Y(_11551_),
    .A(\u_inv.f_next[110] ),
    .B(\u_inv.f_reg[110] ));
 sg13g2_xor2_1 _18609_ (.B(\u_inv.f_reg[110] ),
    .A(\u_inv.f_next[110] ),
    .X(_11552_));
 sg13g2_nor2_1 _18610_ (.A(_11550_),
    .B(_11552_),
    .Y(_11553_));
 sg13g2_xnor2_1 _18611_ (.Y(_11554_),
    .A(\u_inv.f_next[109] ),
    .B(\u_inv.f_reg[109] ));
 sg13g2_xnor2_1 _18612_ (.Y(_11555_),
    .A(\u_inv.f_next[108] ),
    .B(\u_inv.f_reg[108] ));
 sg13g2_nand3_1 _18613_ (.B(_11554_),
    .C(_11555_),
    .A(_11553_),
    .Y(_11556_));
 sg13g2_xor2_1 _18614_ (.B(\u_inv.f_reg[104] ),
    .A(\u_inv.f_next[104] ),
    .X(_11557_));
 sg13g2_xor2_1 _18615_ (.B(\u_inv.f_reg[105] ),
    .A(\u_inv.f_next[105] ),
    .X(_11558_));
 sg13g2_xnor2_1 _18616_ (.Y(_11559_),
    .A(\u_inv.f_next[105] ),
    .B(\u_inv.f_reg[105] ));
 sg13g2_xnor2_1 _18617_ (.Y(_11560_),
    .A(\u_inv.f_next[107] ),
    .B(\u_inv.f_reg[107] ));
 sg13g2_xnor2_1 _18618_ (.Y(_11561_),
    .A(\u_inv.f_next[106] ),
    .B(\u_inv.f_reg[106] ));
 sg13g2_and2_1 _18619_ (.A(_11560_),
    .B(_11561_),
    .X(_11562_));
 sg13g2_nand2_1 _18620_ (.Y(_11563_),
    .A(_11559_),
    .B(_11562_));
 sg13g2_nor3_1 _18621_ (.A(_11556_),
    .B(_11557_),
    .C(_11563_),
    .Y(_11564_));
 sg13g2_xnor2_1 _18622_ (.Y(_11565_),
    .A(\u_inv.f_next[98] ),
    .B(\u_inv.f_reg[98] ));
 sg13g2_xnor2_1 _18623_ (.Y(_11566_),
    .A(\u_inv.f_next[99] ),
    .B(\u_inv.f_reg[99] ));
 sg13g2_xnor2_1 _18624_ (.Y(_11567_),
    .A(\u_inv.f_next[96] ),
    .B(\u_inv.f_reg[96] ));
 sg13g2_nor2_1 _18625_ (.A(\u_inv.f_next[97] ),
    .B(\u_inv.f_reg[97] ),
    .Y(_11568_));
 sg13g2_xor2_1 _18626_ (.B(\u_inv.f_reg[97] ),
    .A(\u_inv.f_next[97] ),
    .X(_11569_));
 sg13g2_nand3_1 _18627_ (.B(_11566_),
    .C(_11567_),
    .A(_11565_),
    .Y(_11570_));
 sg13g2_nor2_1 _18628_ (.A(_11569_),
    .B(_11570_),
    .Y(_11571_));
 sg13g2_xnor2_1 _18629_ (.Y(_11572_),
    .A(\u_inv.f_next[101] ),
    .B(\u_inv.f_reg[101] ));
 sg13g2_inv_1 _18630_ (.Y(_11573_),
    .A(_11572_));
 sg13g2_nor2_1 _18631_ (.A(_10481_),
    .B(_10790_),
    .Y(_11574_));
 sg13g2_xor2_1 _18632_ (.B(\u_inv.f_reg[100] ),
    .A(\u_inv.f_next[100] ),
    .X(_11575_));
 sg13g2_nor2_1 _18633_ (.A(_11573_),
    .B(_11575_),
    .Y(_11576_));
 sg13g2_xor2_1 _18634_ (.B(\u_inv.f_reg[103] ),
    .A(\u_inv.f_next[103] ),
    .X(_11577_));
 sg13g2_xnor2_1 _18635_ (.Y(_11578_),
    .A(\u_inv.f_next[103] ),
    .B(\u_inv.f_reg[103] ));
 sg13g2_nand2_1 _18636_ (.Y(_11579_),
    .A(\u_inv.f_next[102] ),
    .B(\u_inv.f_reg[102] ));
 sg13g2_xnor2_1 _18637_ (.Y(_11580_),
    .A(\u_inv.f_next[102] ),
    .B(\u_inv.f_reg[102] ));
 sg13g2_and4_1 _18638_ (.A(_11571_),
    .B(_11576_),
    .C(_11578_),
    .D(_11580_),
    .X(_11581_));
 sg13g2_and2_1 _18639_ (.A(_11564_),
    .B(_11581_),
    .X(_11582_));
 sg13g2_and2_1 _18640_ (.A(_11547_),
    .B(_11582_),
    .X(_11583_));
 sg13g2_inv_1 _18641_ (.Y(_11584_),
    .A(_11583_));
 sg13g2_a21oi_2 _18642_ (.B1(_11584_),
    .Y(_11585_),
    .A2(_11508_),
    .A1(_11477_));
 sg13g2_nand2_1 _18643_ (.Y(_11586_),
    .A(\u_inv.f_next[117] ),
    .B(_10773_));
 sg13g2_nor2_1 _18644_ (.A(_10465_),
    .B(\u_inv.f_reg[116] ),
    .Y(_11587_));
 sg13g2_nand2_1 _18645_ (.Y(_11588_),
    .A(\u_inv.f_next[114] ),
    .B(_10776_));
 sg13g2_nor2_1 _18646_ (.A(_10468_),
    .B(\u_inv.f_reg[113] ),
    .Y(_11589_));
 sg13g2_nand2_1 _18647_ (.Y(_11590_),
    .A(\u_inv.f_next[112] ),
    .B(_10778_));
 sg13g2_nor2_1 _18648_ (.A(_11535_),
    .B(_11590_),
    .Y(_11591_));
 sg13g2_o21ai_1 _18649_ (.B1(_11531_),
    .Y(_11592_),
    .A1(_11589_),
    .A2(_11591_));
 sg13g2_a21oi_1 _18650_ (.A1(_11588_),
    .A2(_11592_),
    .Y(_11593_),
    .B1(_11529_));
 sg13g2_a21oi_1 _18651_ (.A1(\u_inv.f_next[115] ),
    .A2(_10775_),
    .Y(_11594_),
    .B1(_11593_));
 sg13g2_nor2_1 _18652_ (.A(_11543_),
    .B(_11594_),
    .Y(_11595_));
 sg13g2_o21ai_1 _18653_ (.B1(_11541_),
    .Y(_11596_),
    .A1(_11587_),
    .A2(_11595_));
 sg13g2_nand2_1 _18654_ (.Y(_11597_),
    .A(_11586_),
    .B(_11596_));
 sg13g2_nor2_1 _18655_ (.A(_10463_),
    .B(\u_inv.f_reg[118] ),
    .Y(_11598_));
 sg13g2_nor2_1 _18656_ (.A(_10462_),
    .B(\u_inv.f_reg[119] ),
    .Y(_11599_));
 sg13g2_a221oi_1 _18657_ (.B2(_11537_),
    .C1(_11599_),
    .B1(_11598_),
    .A1(_11540_),
    .Y(_11600_),
    .A2(_11597_));
 sg13g2_nand2_1 _18658_ (.Y(_11601_),
    .A(net3204),
    .B(_10793_));
 sg13g2_nor2_1 _18659_ (.A(_10485_),
    .B(\u_inv.f_reg[96] ),
    .Y(_11602_));
 sg13g2_nand2b_1 _18660_ (.Y(_11603_),
    .B(_11602_),
    .A_N(_11569_));
 sg13g2_nand2_1 _18661_ (.Y(_11604_),
    .A(_11601_),
    .B(_11603_));
 sg13g2_nand3_1 _18662_ (.B(_11566_),
    .C(_11604_),
    .A(_11565_),
    .Y(_11605_));
 sg13g2_nor2_1 _18663_ (.A(_10483_),
    .B(\u_inv.f_reg[98] ),
    .Y(_11606_));
 sg13g2_o21ai_1 _18664_ (.B1(_11605_),
    .Y(_11607_),
    .A1(_10482_),
    .A2(\u_inv.f_reg[99] ));
 sg13g2_a21o_1 _18665_ (.A2(_11606_),
    .A1(_11566_),
    .B1(_11607_),
    .X(_11608_));
 sg13g2_nand2_1 _18666_ (.Y(_11609_),
    .A(\u_inv.f_next[100] ),
    .B(_10790_));
 sg13g2_nor2_1 _18667_ (.A(_10480_),
    .B(\u_inv.f_reg[101] ),
    .Y(_11610_));
 sg13g2_a21oi_1 _18668_ (.A1(_11576_),
    .A2(_11608_),
    .Y(_11611_),
    .B1(_11610_));
 sg13g2_o21ai_1 _18669_ (.B1(_11611_),
    .Y(_11612_),
    .A1(_11573_),
    .A2(_11609_));
 sg13g2_nand2_1 _18670_ (.Y(_11613_),
    .A(\u_inv.f_next[103] ),
    .B(_10787_));
 sg13g2_nor2_1 _18671_ (.A(_10479_),
    .B(\u_inv.f_reg[102] ),
    .Y(_11614_));
 sg13g2_a21oi_1 _18672_ (.A1(_11580_),
    .A2(_11612_),
    .Y(_11615_),
    .B1(_11614_));
 sg13g2_o21ai_1 _18673_ (.B1(_11613_),
    .Y(_11616_),
    .A1(_11577_),
    .A2(_11615_));
 sg13g2_nand2_1 _18674_ (.Y(_11617_),
    .A(_11564_),
    .B(_11616_));
 sg13g2_nand2_1 _18675_ (.Y(_11618_),
    .A(\u_inv.f_next[109] ),
    .B(_10781_));
 sg13g2_nor2_1 _18676_ (.A(_10473_),
    .B(\u_inv.f_reg[108] ),
    .Y(_11619_));
 sg13g2_nand2_1 _18677_ (.Y(_11620_),
    .A(_11554_),
    .B(_11619_));
 sg13g2_nand2_1 _18678_ (.Y(_11621_),
    .A(_11618_),
    .B(_11620_));
 sg13g2_nand2_1 _18679_ (.Y(_11622_),
    .A(\u_inv.f_next[111] ),
    .B(_10779_));
 sg13g2_nor3_1 _18680_ (.A(_10471_),
    .B(\u_inv.f_reg[110] ),
    .C(_11550_),
    .Y(_11623_));
 sg13g2_nor2_1 _18681_ (.A(_10474_),
    .B(\u_inv.f_reg[107] ),
    .Y(_11624_));
 sg13g2_nor2_1 _18682_ (.A(_10475_),
    .B(\u_inv.f_reg[106] ),
    .Y(_11625_));
 sg13g2_nand2_1 _18683_ (.Y(_11626_),
    .A(\u_inv.f_next[105] ),
    .B(_10785_));
 sg13g2_nand2_1 _18684_ (.Y(_11627_),
    .A(\u_inv.f_next[104] ),
    .B(_10786_));
 sg13g2_o21ai_1 _18685_ (.B1(_11626_),
    .Y(_11628_),
    .A1(_11558_),
    .A2(_11627_));
 sg13g2_a221oi_1 _18686_ (.B2(_11562_),
    .C1(_11624_),
    .B1(_11628_),
    .A1(_11560_),
    .Y(_11629_),
    .A2(_11625_));
 sg13g2_or2_1 _18687_ (.X(_11630_),
    .B(_11629_),
    .A(_11556_));
 sg13g2_a21oi_1 _18688_ (.A1(_11553_),
    .A2(_11621_),
    .Y(_11631_),
    .B1(_11623_));
 sg13g2_nand4_1 _18689_ (.B(_11622_),
    .C(_11630_),
    .A(_11617_),
    .Y(_11632_),
    .D(_11631_));
 sg13g2_nand2_1 _18690_ (.Y(_11633_),
    .A(\u_inv.f_next[123] ),
    .B(_10767_));
 sg13g2_nor2_1 _18691_ (.A(_10459_),
    .B(\u_inv.f_reg[122] ),
    .Y(_11634_));
 sg13g2_nand2_1 _18692_ (.Y(_11635_),
    .A(\u_inv.f_next[121] ),
    .B(_10769_));
 sg13g2_nor2_1 _18693_ (.A(_10461_),
    .B(net2386),
    .Y(_11636_));
 sg13g2_nand2b_1 _18694_ (.Y(_11637_),
    .B(_11636_),
    .A_N(_11517_));
 sg13g2_nand2_1 _18695_ (.Y(_11638_),
    .A(_11635_),
    .B(_11637_));
 sg13g2_a21oi_1 _18696_ (.A1(_11512_),
    .A2(_11638_),
    .Y(_11639_),
    .B1(_11634_));
 sg13g2_o21ai_1 _18697_ (.B1(_11633_),
    .Y(_11640_),
    .A1(_11510_),
    .A2(_11639_));
 sg13g2_nand2_1 _18698_ (.Y(_11641_),
    .A(\u_inv.f_next[124] ),
    .B(_10766_));
 sg13g2_nor2_1 _18699_ (.A(_10456_),
    .B(\u_inv.f_reg[125] ),
    .Y(_11642_));
 sg13g2_a21oi_1 _18700_ (.A1(_11527_),
    .A2(_11640_),
    .Y(_11643_),
    .B1(_11642_));
 sg13g2_o21ai_1 _18701_ (.B1(_11643_),
    .Y(_11644_),
    .A1(_11524_),
    .A2(_11641_));
 sg13g2_nor2_1 _18702_ (.A(_10455_),
    .B(\u_inv.f_reg[126] ),
    .Y(_11645_));
 sg13g2_a22oi_1 _18703_ (.Y(_11646_),
    .B1(_11645_),
    .B2(_11520_),
    .A2(_11644_),
    .A1(_11523_));
 sg13g2_o21ai_1 _18704_ (.B1(_11646_),
    .Y(_11647_),
    .A1(_11528_),
    .A2(_11600_));
 sg13g2_a21oi_1 _18705_ (.A1(_11547_),
    .A2(_11632_),
    .Y(_11648_),
    .B1(_11647_));
 sg13g2_o21ai_1 _18706_ (.B1(_11648_),
    .Y(_11649_),
    .A1(_10454_),
    .A2(\u_inv.f_reg[127] ));
 sg13g2_nor2_2 _18707_ (.A(_11585_),
    .B(_11649_),
    .Y(_11650_));
 sg13g2_xor2_1 _18708_ (.B(\u_inv.f_reg[152] ),
    .A(\u_inv.f_next[152] ),
    .X(_11651_));
 sg13g2_xor2_1 _18709_ (.B(\u_inv.f_reg[153] ),
    .A(\u_inv.f_next[153] ),
    .X(_11652_));
 sg13g2_nor2_1 _18710_ (.A(_10427_),
    .B(_10736_),
    .Y(_11653_));
 sg13g2_xor2_1 _18711_ (.B(\u_inv.f_reg[154] ),
    .A(\u_inv.f_next[154] ),
    .X(_11654_));
 sg13g2_xor2_1 _18712_ (.B(\u_inv.f_reg[155] ),
    .A(\u_inv.f_next[155] ),
    .X(_11655_));
 sg13g2_xnor2_1 _18713_ (.Y(_11656_),
    .A(\u_inv.f_next[155] ),
    .B(\u_inv.f_reg[155] ));
 sg13g2_nor4_1 _18714_ (.A(_11651_),
    .B(_11652_),
    .C(_11654_),
    .D(_11655_),
    .Y(_11657_));
 sg13g2_inv_1 _18715_ (.Y(_11658_),
    .A(_11657_));
 sg13g2_xor2_1 _18716_ (.B(\u_inv.f_reg[149] ),
    .A(\u_inv.f_next[149] ),
    .X(_11659_));
 sg13g2_nand2_1 _18717_ (.Y(_11660_),
    .A(\u_inv.f_next[150] ),
    .B(\u_inv.f_reg[150] ));
 sg13g2_xor2_1 _18718_ (.B(\u_inv.f_reg[150] ),
    .A(\u_inv.f_next[150] ),
    .X(_11661_));
 sg13g2_xnor2_1 _18719_ (.Y(_11662_),
    .A(\u_inv.f_next[150] ),
    .B(\u_inv.f_reg[150] ));
 sg13g2_xor2_1 _18720_ (.B(\u_inv.f_reg[148] ),
    .A(\u_inv.f_next[148] ),
    .X(_11663_));
 sg13g2_xnor2_1 _18721_ (.Y(_11664_),
    .A(\u_inv.f_next[148] ),
    .B(\u_inv.f_reg[148] ));
 sg13g2_xor2_1 _18722_ (.B(\u_inv.f_reg[151] ),
    .A(\u_inv.f_next[151] ),
    .X(_11665_));
 sg13g2_nor4_1 _18723_ (.A(_11659_),
    .B(_11661_),
    .C(_11663_),
    .D(_11665_),
    .Y(_11666_));
 sg13g2_nand2_1 _18724_ (.Y(_11667_),
    .A(\u_inv.f_next[146] ),
    .B(\u_inv.f_reg[146] ));
 sg13g2_xor2_1 _18725_ (.B(\u_inv.f_reg[146] ),
    .A(\u_inv.f_next[146] ),
    .X(_11668_));
 sg13g2_xnor2_1 _18726_ (.Y(_11669_),
    .A(\u_inv.f_next[146] ),
    .B(\u_inv.f_reg[146] ));
 sg13g2_nand2_1 _18727_ (.Y(_11670_),
    .A(\u_inv.f_next[144] ),
    .B(\u_inv.f_reg[144] ));
 sg13g2_xnor2_1 _18728_ (.Y(_11671_),
    .A(\u_inv.f_next[144] ),
    .B(\u_inv.f_reg[144] ));
 sg13g2_xor2_1 _18729_ (.B(\u_inv.f_reg[147] ),
    .A(\u_inv.f_next[147] ),
    .X(_11672_));
 sg13g2_inv_1 _18730_ (.Y(_11673_),
    .A(_11672_));
 sg13g2_xnor2_1 _18731_ (.Y(_11674_),
    .A(\u_inv.f_next[145] ),
    .B(\u_inv.f_reg[145] ));
 sg13g2_nand4_1 _18732_ (.B(_11671_),
    .C(_11673_),
    .A(_11669_),
    .Y(_11675_),
    .D(_11674_));
 sg13g2_nor2_1 _18733_ (.A(\u_inv.f_next[159] ),
    .B(\u_inv.f_reg[159] ),
    .Y(_11676_));
 sg13g2_nand2_1 _18734_ (.Y(_11677_),
    .A(\u_inv.f_next[159] ),
    .B(\u_inv.f_reg[159] ));
 sg13g2_nand2b_2 _18735_ (.Y(_11678_),
    .B(_11677_),
    .A_N(_11676_));
 sg13g2_nand2_1 _18736_ (.Y(_11679_),
    .A(\u_inv.f_next[158] ),
    .B(\u_inv.f_reg[158] ));
 sg13g2_xor2_1 _18737_ (.B(\u_inv.f_reg[158] ),
    .A(\u_inv.f_next[158] ),
    .X(_11680_));
 sg13g2_inv_1 _18738_ (.Y(_11681_),
    .A(_11680_));
 sg13g2_nand2_1 _18739_ (.Y(_11682_),
    .A(_10424_),
    .B(_10733_));
 sg13g2_xnor2_1 _18740_ (.Y(_11683_),
    .A(\u_inv.f_next[157] ),
    .B(\u_inv.f_reg[157] ));
 sg13g2_xnor2_1 _18741_ (.Y(_11684_),
    .A(\u_inv.f_next[156] ),
    .B(\u_inv.f_reg[156] ));
 sg13g2_nand4_1 _18742_ (.B(_11681_),
    .C(_11683_),
    .A(_11678_),
    .Y(_11685_),
    .D(_11684_));
 sg13g2_nor3_1 _18743_ (.A(_11658_),
    .B(_11675_),
    .C(_11685_),
    .Y(_11686_));
 sg13g2_nand2_1 _18744_ (.Y(_11687_),
    .A(_11666_),
    .B(_11686_));
 sg13g2_nor2_1 _18745_ (.A(\u_inv.f_next[143] ),
    .B(\u_inv.f_reg[143] ),
    .Y(_11688_));
 sg13g2_nor2_1 _18746_ (.A(_10438_),
    .B(_10747_),
    .Y(_11689_));
 sg13g2_nand2_1 _18747_ (.Y(_11690_),
    .A(\u_inv.f_next[143] ),
    .B(\u_inv.f_reg[143] ));
 sg13g2_nor2_2 _18748_ (.A(_11688_),
    .B(_11689_),
    .Y(_11691_));
 sg13g2_nand2_1 _18749_ (.Y(_11692_),
    .A(\u_inv.f_next[142] ),
    .B(\u_inv.f_reg[142] ));
 sg13g2_xnor2_1 _18750_ (.Y(_11693_),
    .A(\u_inv.f_next[142] ),
    .B(\u_inv.f_reg[142] ));
 sg13g2_nor2b_2 _18751_ (.A(_11691_),
    .B_N(_11693_),
    .Y(_11694_));
 sg13g2_xor2_1 _18752_ (.B(\u_inv.f_reg[141] ),
    .A(\u_inv.f_next[141] ),
    .X(_11695_));
 sg13g2_xor2_1 _18753_ (.B(\u_inv.f_reg[140] ),
    .A(\u_inv.f_next[140] ),
    .X(_11696_));
 sg13g2_nor2_1 _18754_ (.A(_11695_),
    .B(_11696_),
    .Y(_11697_));
 sg13g2_nand2_1 _18755_ (.Y(_11698_),
    .A(_11694_),
    .B(_11697_));
 sg13g2_xnor2_1 _18756_ (.Y(_11699_),
    .A(\u_inv.f_next[139] ),
    .B(\u_inv.f_reg[139] ));
 sg13g2_inv_1 _18757_ (.Y(_11700_),
    .A(_11699_));
 sg13g2_nand2_1 _18758_ (.Y(_11701_),
    .A(\u_inv.f_next[138] ),
    .B(\u_inv.f_reg[138] ));
 sg13g2_xnor2_1 _18759_ (.Y(_11702_),
    .A(\u_inv.f_next[138] ),
    .B(\u_inv.f_reg[138] ));
 sg13g2_xnor2_1 _18760_ (.Y(_11703_),
    .A(\u_inv.f_next[136] ),
    .B(\u_inv.f_reg[136] ));
 sg13g2_nor2_1 _18761_ (.A(\u_inv.f_next[137] ),
    .B(\u_inv.f_reg[137] ),
    .Y(_11704_));
 sg13g2_xor2_1 _18762_ (.B(net2396),
    .A(\u_inv.f_next[137] ),
    .X(_11705_));
 sg13g2_inv_2 _18763_ (.Y(_11706_),
    .A(_11705_));
 sg13g2_and4_1 _18764_ (.A(_11699_),
    .B(_11702_),
    .C(_11703_),
    .D(_11706_),
    .X(_11707_));
 sg13g2_nand3_1 _18765_ (.B(_11697_),
    .C(_11707_),
    .A(_11694_),
    .Y(_11708_));
 sg13g2_nor2_1 _18766_ (.A(\u_inv.f_next[135] ),
    .B(\u_inv.f_reg[135] ),
    .Y(_11709_));
 sg13g2_xor2_1 _18767_ (.B(\u_inv.f_reg[135] ),
    .A(\u_inv.f_next[135] ),
    .X(_11710_));
 sg13g2_xnor2_1 _18768_ (.Y(_11711_),
    .A(\u_inv.f_next[135] ),
    .B(\u_inv.f_reg[135] ));
 sg13g2_nand2_1 _18769_ (.Y(_11712_),
    .A(\u_inv.f_next[134] ),
    .B(\u_inv.f_reg[134] ));
 sg13g2_xor2_1 _18770_ (.B(\u_inv.f_reg[134] ),
    .A(\u_inv.f_next[134] ),
    .X(_11713_));
 sg13g2_xnor2_1 _18771_ (.Y(_11714_),
    .A(\u_inv.f_next[134] ),
    .B(\u_inv.f_reg[134] ));
 sg13g2_xnor2_1 _18772_ (.Y(_11715_),
    .A(\u_inv.f_next[132] ),
    .B(\u_inv.f_reg[132] ));
 sg13g2_xor2_1 _18773_ (.B(\u_inv.f_reg[133] ),
    .A(\u_inv.f_next[133] ),
    .X(_11716_));
 sg13g2_xnor2_1 _18774_ (.Y(_11717_),
    .A(\u_inv.f_next[133] ),
    .B(\u_inv.f_reg[133] ));
 sg13g2_nand4_1 _18775_ (.B(_11714_),
    .C(_11715_),
    .A(_11711_),
    .Y(_11718_),
    .D(_11717_));
 sg13g2_xor2_1 _18776_ (.B(\u_inv.f_reg[131] ),
    .A(\u_inv.f_next[131] ),
    .X(_11719_));
 sg13g2_xnor2_1 _18777_ (.Y(_11720_),
    .A(\u_inv.f_next[131] ),
    .B(\u_inv.f_reg[131] ));
 sg13g2_nand2_1 _18778_ (.Y(_11721_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_xnor2_1 _18779_ (.Y(_11722_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_nand2_1 _18780_ (.Y(_11723_),
    .A(\u_inv.f_next[128] ),
    .B(\u_inv.f_reg[128] ));
 sg13g2_xnor2_1 _18781_ (.Y(_11724_),
    .A(\u_inv.f_next[128] ),
    .B(\u_inv.f_reg[128] ));
 sg13g2_xnor2_1 _18782_ (.Y(_11725_),
    .A(\u_inv.f_next[129] ),
    .B(\u_inv.f_reg[129] ));
 sg13g2_nand4_1 _18783_ (.B(_11722_),
    .C(_11724_),
    .A(_11720_),
    .Y(_11726_),
    .D(_11725_));
 sg13g2_or2_1 _18784_ (.X(_11727_),
    .B(_11726_),
    .A(_11718_));
 sg13g2_or2_1 _18785_ (.X(_11728_),
    .B(_11727_),
    .A(_11708_));
 sg13g2_nor2_2 _18786_ (.A(_11687_),
    .B(_11728_),
    .Y(_11729_));
 sg13g2_xor2_1 _18787_ (.B(\u_inv.f_reg[191] ),
    .A(\u_inv.f_next[191] ),
    .X(_11730_));
 sg13g2_nand2_1 _18788_ (.Y(_11731_),
    .A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ));
 sg13g2_xor2_1 _18789_ (.B(\u_inv.f_reg[190] ),
    .A(\u_inv.f_next[190] ),
    .X(_11732_));
 sg13g2_xnor2_1 _18790_ (.Y(_11733_),
    .A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ));
 sg13g2_xnor2_1 _18791_ (.Y(_11734_),
    .A(\u_inv.f_next[189] ),
    .B(\u_inv.f_reg[189] ));
 sg13g2_nor2_1 _18792_ (.A(_10393_),
    .B(_10702_),
    .Y(_11735_));
 sg13g2_xor2_1 _18793_ (.B(\u_inv.f_reg[188] ),
    .A(\u_inv.f_next[188] ),
    .X(_11736_));
 sg13g2_xnor2_1 _18794_ (.Y(_11737_),
    .A(\u_inv.f_next[188] ),
    .B(\u_inv.f_reg[188] ));
 sg13g2_nor3_1 _18795_ (.A(_11730_),
    .B(_11732_),
    .C(_11736_),
    .Y(_11738_));
 sg13g2_nand2_1 _18796_ (.Y(_11739_),
    .A(_11734_),
    .B(_11738_));
 sg13g2_xor2_1 _18797_ (.B(\u_inv.f_reg[187] ),
    .A(\u_inv.f_next[187] ),
    .X(_11740_));
 sg13g2_xnor2_1 _18798_ (.Y(_11741_),
    .A(\u_inv.f_next[187] ),
    .B(\u_inv.f_reg[187] ));
 sg13g2_nand2_1 _18799_ (.Y(_11742_),
    .A(\u_inv.f_next[186] ),
    .B(\u_inv.f_reg[186] ));
 sg13g2_xnor2_1 _18800_ (.Y(_11743_),
    .A(\u_inv.f_next[186] ),
    .B(\u_inv.f_reg[186] ));
 sg13g2_xnor2_1 _18801_ (.Y(_11744_),
    .A(\u_inv.f_next[184] ),
    .B(\u_inv.f_reg[184] ));
 sg13g2_xor2_1 _18802_ (.B(\u_inv.f_reg[185] ),
    .A(\u_inv.f_next[185] ),
    .X(_11745_));
 sg13g2_nand3_1 _18803_ (.B(_11743_),
    .C(_11744_),
    .A(_11741_),
    .Y(_11746_));
 sg13g2_nor2_1 _18804_ (.A(_11745_),
    .B(_11746_),
    .Y(_11747_));
 sg13g2_nand2b_2 _18805_ (.Y(_11748_),
    .B(_11747_),
    .A_N(_11739_));
 sg13g2_xor2_1 _18806_ (.B(\u_inv.f_reg[183] ),
    .A(\u_inv.f_next[183] ),
    .X(_11749_));
 sg13g2_xnor2_1 _18807_ (.Y(_11750_),
    .A(\u_inv.f_next[183] ),
    .B(\u_inv.f_reg[183] ));
 sg13g2_nand2_1 _18808_ (.Y(_11751_),
    .A(\u_inv.f_next[182] ),
    .B(\u_inv.f_reg[182] ));
 sg13g2_xor2_1 _18809_ (.B(\u_inv.f_reg[182] ),
    .A(\u_inv.f_next[182] ),
    .X(_11752_));
 sg13g2_xnor2_1 _18810_ (.Y(_11753_),
    .A(\u_inv.f_next[182] ),
    .B(\u_inv.f_reg[182] ));
 sg13g2_nor2_1 _18811_ (.A(_10401_),
    .B(_10710_),
    .Y(_11754_));
 sg13g2_xor2_1 _18812_ (.B(\u_inv.f_reg[180] ),
    .A(\u_inv.f_next[180] ),
    .X(_11755_));
 sg13g2_xnor2_1 _18813_ (.Y(_11756_),
    .A(\u_inv.f_next[180] ),
    .B(\u_inv.f_reg[180] ));
 sg13g2_xnor2_1 _18814_ (.Y(_11757_),
    .A(\u_inv.f_next[181] ),
    .B(\u_inv.f_reg[181] ));
 sg13g2_nand4_1 _18815_ (.B(_11753_),
    .C(_11756_),
    .A(_11750_),
    .Y(_11758_),
    .D(_11757_));
 sg13g2_xor2_1 _18816_ (.B(\u_inv.f_reg[176] ),
    .A(\u_inv.f_next[176] ),
    .X(_11759_));
 sg13g2_xor2_1 _18817_ (.B(\u_inv.f_reg[177] ),
    .A(\u_inv.f_next[177] ),
    .X(_11760_));
 sg13g2_nor2_1 _18818_ (.A(_11759_),
    .B(_11760_),
    .Y(_11761_));
 sg13g2_nand2_1 _18819_ (.Y(_11762_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_xnor2_1 _18820_ (.Y(_11763_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_xnor2_1 _18821_ (.Y(_11764_),
    .A(\u_inv.f_next[179] ),
    .B(\u_inv.f_reg[179] ));
 sg13g2_and3_1 _18822_ (.X(_11765_),
    .A(_11761_),
    .B(net4433),
    .C(_11764_));
 sg13g2_nand3_1 _18823_ (.B(net4433),
    .C(_11764_),
    .A(_11761_),
    .Y(_11766_));
 sg13g2_nor3_2 _18824_ (.A(_11748_),
    .B(_11758_),
    .C(_11766_),
    .Y(_11767_));
 sg13g2_xor2_1 _18825_ (.B(\u_inv.f_reg[175] ),
    .A(\u_inv.f_next[175] ),
    .X(_11768_));
 sg13g2_nor2_1 _18826_ (.A(_10407_),
    .B(_10716_),
    .Y(_11769_));
 sg13g2_xor2_1 _18827_ (.B(\u_inv.f_reg[174] ),
    .A(\u_inv.f_next[174] ),
    .X(_11770_));
 sg13g2_nor2_1 _18828_ (.A(_11768_),
    .B(_11770_),
    .Y(_11771_));
 sg13g2_xnor2_1 _18829_ (.Y(_11772_),
    .A(\u_inv.f_next[173] ),
    .B(\u_inv.f_reg[173] ));
 sg13g2_nand2_1 _18830_ (.Y(_11773_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_xnor2_1 _18831_ (.Y(_11774_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_nand3_1 _18832_ (.B(_11772_),
    .C(_11774_),
    .A(_11771_),
    .Y(_11775_));
 sg13g2_xor2_1 _18833_ (.B(\u_inv.f_reg[171] ),
    .A(\u_inv.f_next[171] ),
    .X(_11776_));
 sg13g2_xnor2_1 _18834_ (.Y(_11777_),
    .A(\u_inv.f_next[171] ),
    .B(\u_inv.f_reg[171] ));
 sg13g2_nor2_1 _18835_ (.A(_10411_),
    .B(_10720_),
    .Y(_11778_));
 sg13g2_xor2_1 _18836_ (.B(\u_inv.f_reg[170] ),
    .A(\u_inv.f_next[170] ),
    .X(_11779_));
 sg13g2_xnor2_1 _18837_ (.Y(_11780_),
    .A(\u_inv.f_next[170] ),
    .B(\u_inv.f_reg[170] ));
 sg13g2_nor2_1 _18838_ (.A(_11776_),
    .B(_11779_),
    .Y(_11781_));
 sg13g2_nand2_1 _18839_ (.Y(_11782_),
    .A(\u_inv.f_next[168] ),
    .B(\u_inv.f_reg[168] ));
 sg13g2_xor2_1 _18840_ (.B(\u_inv.f_reg[168] ),
    .A(\u_inv.f_next[168] ),
    .X(_11783_));
 sg13g2_xnor2_1 _18841_ (.Y(_11784_),
    .A(\u_inv.f_next[168] ),
    .B(\u_inv.f_reg[168] ));
 sg13g2_xnor2_1 _18842_ (.Y(_11785_),
    .A(\u_inv.f_next[169] ),
    .B(\u_inv.f_reg[169] ));
 sg13g2_nand3_1 _18843_ (.B(_11784_),
    .C(_11785_),
    .A(_11781_),
    .Y(_11786_));
 sg13g2_nor2_1 _18844_ (.A(_11775_),
    .B(_11786_),
    .Y(_11787_));
 sg13g2_xnor2_1 _18845_ (.Y(_11788_),
    .A(\u_inv.f_next[163] ),
    .B(\u_inv.f_reg[163] ));
 sg13g2_nand2_1 _18846_ (.Y(_11789_),
    .A(\u_inv.f_next[162] ),
    .B(\u_inv.f_reg[162] ));
 sg13g2_xnor2_1 _18847_ (.Y(_11790_),
    .A(\u_inv.f_next[162] ),
    .B(\u_inv.f_reg[162] ));
 sg13g2_inv_1 _18848_ (.Y(_11791_),
    .A(_11790_));
 sg13g2_xnor2_1 _18849_ (.Y(_11792_),
    .A(\u_inv.f_next[160] ),
    .B(\u_inv.f_reg[160] ));
 sg13g2_xnor2_1 _18850_ (.Y(_11793_),
    .A(\u_inv.f_next[161] ),
    .B(\u_inv.f_reg[161] ));
 sg13g2_and4_1 _18851_ (.A(_11788_),
    .B(_11790_),
    .C(net4432),
    .D(_11793_),
    .X(_11794_));
 sg13g2_xnor2_1 _18852_ (.Y(_11795_),
    .A(\u_inv.f_next[167] ),
    .B(\u_inv.f_reg[167] ));
 sg13g2_nand2_1 _18853_ (.Y(_11796_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_xnor2_1 _18854_ (.Y(_11797_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_xor2_1 _18855_ (.B(\u_inv.f_reg[164] ),
    .A(\u_inv.f_next[164] ),
    .X(_11798_));
 sg13g2_xor2_1 _18856_ (.B(\u_inv.f_reg[165] ),
    .A(\u_inv.f_next[165] ),
    .X(_11799_));
 sg13g2_xnor2_1 _18857_ (.Y(_11800_),
    .A(\u_inv.f_next[165] ),
    .B(\u_inv.f_reg[165] ));
 sg13g2_nand3_1 _18858_ (.B(_11797_),
    .C(_11800_),
    .A(_11795_),
    .Y(_11801_));
 sg13g2_nor2_1 _18859_ (.A(_11798_),
    .B(_11801_),
    .Y(_11802_));
 sg13g2_and2_1 _18860_ (.A(_11794_),
    .B(_11802_),
    .X(_11803_));
 sg13g2_nand2_1 _18861_ (.Y(_11804_),
    .A(_11787_),
    .B(_11803_));
 sg13g2_nand4_1 _18862_ (.B(_11767_),
    .C(_11787_),
    .A(_11729_),
    .Y(_11805_),
    .D(_11803_));
 sg13g2_nor2_1 _18863_ (.A(_10427_),
    .B(\u_inv.f_reg[154] ),
    .Y(_11806_));
 sg13g2_nand2_1 _18864_ (.Y(_11807_),
    .A(\u_inv.f_next[153] ),
    .B(_10737_));
 sg13g2_nor2_1 _18865_ (.A(_10429_),
    .B(\u_inv.f_reg[152] ),
    .Y(_11808_));
 sg13g2_nand2b_1 _18866_ (.Y(_11809_),
    .B(_11808_),
    .A_N(_11652_));
 sg13g2_a21oi_1 _18867_ (.A1(_11807_),
    .A2(_11809_),
    .Y(_11810_),
    .B1(_11654_));
 sg13g2_o21ai_1 _18868_ (.B1(_11656_),
    .Y(_11811_),
    .A1(_11806_),
    .A2(_11810_));
 sg13g2_o21ai_1 _18869_ (.B1(_11811_),
    .Y(_11812_),
    .A1(_10426_),
    .A2(\u_inv.f_reg[155] ));
 sg13g2_inv_1 _18870_ (.Y(_11813_),
    .A(_11812_));
 sg13g2_nand2_1 _18871_ (.Y(_11814_),
    .A(\u_inv.f_next[151] ),
    .B(_10739_));
 sg13g2_nand2_1 _18872_ (.Y(_11815_),
    .A(\u_inv.f_next[148] ),
    .B(_10742_));
 sg13g2_nor2_1 _18873_ (.A(_10437_),
    .B(\u_inv.f_reg[144] ),
    .Y(_11816_));
 sg13g2_nand2_1 _18874_ (.Y(_11817_),
    .A(_11674_),
    .B(_11816_));
 sg13g2_o21ai_1 _18875_ (.B1(_11817_),
    .Y(_11818_),
    .A1(_10436_),
    .A2(\u_inv.f_reg[145] ));
 sg13g2_nand2_1 _18876_ (.Y(_11819_),
    .A(_11669_),
    .B(_11818_));
 sg13g2_nand2_1 _18877_ (.Y(_11820_),
    .A(\u_inv.f_next[146] ),
    .B(_10744_));
 sg13g2_a21oi_1 _18878_ (.A1(_11819_),
    .A2(_11820_),
    .Y(_11821_),
    .B1(_11672_));
 sg13g2_a21o_1 _18879_ (.A2(_10743_),
    .A1(\u_inv.f_next[147] ),
    .B1(_11821_),
    .X(_11822_));
 sg13g2_nand2_1 _18880_ (.Y(_11823_),
    .A(_11664_),
    .B(_11822_));
 sg13g2_nor2_1 _18881_ (.A(_10431_),
    .B(\u_inv.f_reg[150] ),
    .Y(_11824_));
 sg13g2_nor2_1 _18882_ (.A(_10432_),
    .B(\u_inv.f_reg[149] ),
    .Y(_11825_));
 sg13g2_a21oi_1 _18883_ (.A1(_11815_),
    .A2(_11823_),
    .Y(_11826_),
    .B1(_11659_));
 sg13g2_o21ai_1 _18884_ (.B1(_11662_),
    .Y(_11827_),
    .A1(_11825_),
    .A2(_11826_));
 sg13g2_nor2b_1 _18885_ (.A(_11824_),
    .B_N(_11827_),
    .Y(_11828_));
 sg13g2_o21ai_1 _18886_ (.B1(_11814_),
    .Y(_11829_),
    .A1(_11665_),
    .A2(_11828_));
 sg13g2_a21oi_1 _18887_ (.A1(_11657_),
    .A2(_11829_),
    .Y(_11830_),
    .B1(_11812_));
 sg13g2_nor2_1 _18888_ (.A(_11685_),
    .B(_11830_),
    .Y(_11831_));
 sg13g2_nor2_1 _18889_ (.A(_10423_),
    .B(\u_inv.f_reg[158] ),
    .Y(_11832_));
 sg13g2_nand2_1 _18890_ (.Y(_11833_),
    .A(\u_inv.f_next[157] ),
    .B(_10733_));
 sg13g2_nor2_1 _18891_ (.A(_10425_),
    .B(\u_inv.f_reg[156] ),
    .Y(_11834_));
 sg13g2_nand2_1 _18892_ (.Y(_11835_),
    .A(_11683_),
    .B(_11834_));
 sg13g2_a21oi_1 _18893_ (.A1(_11833_),
    .A2(_11835_),
    .Y(_11836_),
    .B1(_11680_));
 sg13g2_o21ai_1 _18894_ (.B1(_11678_),
    .Y(_11837_),
    .A1(_11832_),
    .A2(_11836_));
 sg13g2_o21ai_1 _18895_ (.B1(_11837_),
    .Y(_11838_),
    .A1(_10422_),
    .A2(\u_inv.f_reg[159] ));
 sg13g2_nand2_1 _18896_ (.Y(_11839_),
    .A(\u_inv.f_next[130] ),
    .B(_10760_));
 sg13g2_nor2_1 _18897_ (.A(_10452_),
    .B(\u_inv.f_reg[129] ),
    .Y(_11840_));
 sg13g2_nand2_1 _18898_ (.Y(_11841_),
    .A(\u_inv.f_next[128] ),
    .B(_10762_));
 sg13g2_nor2b_1 _18899_ (.A(_11841_),
    .B_N(_11725_),
    .Y(_11842_));
 sg13g2_o21ai_1 _18900_ (.B1(_11722_),
    .Y(_11843_),
    .A1(_11840_),
    .A2(_11842_));
 sg13g2_a21oi_1 _18901_ (.A1(_11839_),
    .A2(_11843_),
    .Y(_11844_),
    .B1(_11719_));
 sg13g2_a21oi_2 _18902_ (.B1(_11844_),
    .Y(_11845_),
    .A2(_10759_),
    .A1(\u_inv.f_next[131] ));
 sg13g2_nor2_1 _18903_ (.A(_10448_),
    .B(\u_inv.f_reg[133] ),
    .Y(_11846_));
 sg13g2_nor2_1 _18904_ (.A(_10449_),
    .B(\u_inv.f_reg[132] ),
    .Y(_11847_));
 sg13g2_a21oi_1 _18905_ (.A1(_11717_),
    .A2(_11847_),
    .Y(_11848_),
    .B1(_11846_));
 sg13g2_nor3_1 _18906_ (.A(_11710_),
    .B(_11713_),
    .C(_11848_),
    .Y(_11849_));
 sg13g2_nor3_1 _18907_ (.A(_10447_),
    .B(\u_inv.f_reg[134] ),
    .C(_11710_),
    .Y(_11850_));
 sg13g2_a21oi_1 _18908_ (.A1(\u_inv.f_next[135] ),
    .A2(_10755_),
    .Y(_11851_),
    .B1(_11850_));
 sg13g2_o21ai_1 _18909_ (.B1(_11851_),
    .Y(_11852_),
    .A1(_11718_),
    .A2(_11845_));
 sg13g2_nor2_1 _18910_ (.A(_11849_),
    .B(_11852_),
    .Y(_11853_));
 sg13g2_nor2_1 _18911_ (.A(_11708_),
    .B(_11853_),
    .Y(_11854_));
 sg13g2_nor2_1 _18912_ (.A(_10440_),
    .B(\u_inv.f_reg[141] ),
    .Y(_11855_));
 sg13g2_nand2_1 _18913_ (.Y(_11856_),
    .A(\u_inv.f_next[140] ),
    .B(_10750_));
 sg13g2_nor2_1 _18914_ (.A(_11695_),
    .B(_11856_),
    .Y(_11857_));
 sg13g2_o21ai_1 _18915_ (.B1(_11694_),
    .Y(_11858_),
    .A1(_11855_),
    .A2(_11857_));
 sg13g2_nand2_1 _18916_ (.Y(_11859_),
    .A(\u_inv.f_next[142] ),
    .B(_10748_));
 sg13g2_nand2_1 _18917_ (.Y(_11860_),
    .A(\u_inv.f_next[139] ),
    .B(_10751_));
 sg13g2_nor2_1 _18918_ (.A(_10443_),
    .B(\u_inv.f_reg[138] ),
    .Y(_11861_));
 sg13g2_nand2_1 _18919_ (.Y(_11862_),
    .A(\u_inv.f_next[137] ),
    .B(_10753_));
 sg13g2_nor2_1 _18920_ (.A(_10445_),
    .B(net2158),
    .Y(_11863_));
 sg13g2_nand2_1 _18921_ (.Y(_11864_),
    .A(_11706_),
    .B(_11863_));
 sg13g2_nand2_1 _18922_ (.Y(_11865_),
    .A(_11862_),
    .B(_11864_));
 sg13g2_a21oi_1 _18923_ (.A1(_11702_),
    .A2(_11865_),
    .Y(_11866_),
    .B1(_11861_));
 sg13g2_o21ai_1 _18924_ (.B1(_11860_),
    .Y(_11867_),
    .A1(_11700_),
    .A2(_11866_));
 sg13g2_nand2b_1 _18925_ (.Y(_11868_),
    .B(_11867_),
    .A_N(_11698_));
 sg13g2_o21ai_1 _18926_ (.B1(_11858_),
    .Y(_11869_),
    .A1(_11691_),
    .A2(_11859_));
 sg13g2_o21ai_1 _18927_ (.B1(_11868_),
    .Y(_11870_),
    .A1(_10438_),
    .A2(\u_inv.f_reg[143] ));
 sg13g2_nor3_1 _18928_ (.A(_11854_),
    .B(_11869_),
    .C(_11870_),
    .Y(_11871_));
 sg13g2_nor2_1 _18929_ (.A(_11687_),
    .B(_11871_),
    .Y(_11872_));
 sg13g2_nor3_2 _18930_ (.A(_11831_),
    .B(_11838_),
    .C(_11872_),
    .Y(_11873_));
 sg13g2_nor2_1 _18931_ (.A(_10414_),
    .B(\u_inv.f_reg[167] ),
    .Y(_11874_));
 sg13g2_nor2_1 _18932_ (.A(_10415_),
    .B(\u_inv.f_reg[166] ),
    .Y(_11875_));
 sg13g2_nand2_1 _18933_ (.Y(_11876_),
    .A(\u_inv.f_next[165] ),
    .B(_10725_));
 sg13g2_nand2_1 _18934_ (.Y(_11877_),
    .A(\u_inv.f_next[164] ),
    .B(_10726_));
 sg13g2_o21ai_1 _18935_ (.B1(_11876_),
    .Y(_11878_),
    .A1(_11799_),
    .A2(_11877_));
 sg13g2_nor2_1 _18936_ (.A(_10419_),
    .B(\u_inv.f_reg[162] ),
    .Y(_11879_));
 sg13g2_nand2_1 _18937_ (.Y(_11880_),
    .A(\u_inv.f_next[161] ),
    .B(_10729_));
 sg13g2_nor2_1 _18938_ (.A(_10421_),
    .B(\u_inv.f_reg[160] ),
    .Y(_11881_));
 sg13g2_nand2_1 _18939_ (.Y(_11882_),
    .A(_11793_),
    .B(_11881_));
 sg13g2_a21oi_1 _18940_ (.A1(_11880_),
    .A2(_11882_),
    .Y(_11883_),
    .B1(_11791_));
 sg13g2_o21ai_1 _18941_ (.B1(_11788_),
    .Y(_11884_),
    .A1(_11879_),
    .A2(_11883_));
 sg13g2_o21ai_1 _18942_ (.B1(_11884_),
    .Y(_11885_),
    .A1(_10418_),
    .A2(\u_inv.f_reg[163] ));
 sg13g2_nand3_1 _18943_ (.B(_11797_),
    .C(_11878_),
    .A(_11795_),
    .Y(_11886_));
 sg13g2_a221oi_1 _18944_ (.B2(_11802_),
    .C1(_11874_),
    .B1(_11885_),
    .A1(_11795_),
    .Y(_11887_),
    .A2(_11875_));
 sg13g2_nand2_2 _18945_ (.Y(_11888_),
    .A(_11886_),
    .B(_11887_));
 sg13g2_nor2_1 _18946_ (.A(_10410_),
    .B(\u_inv.f_reg[171] ),
    .Y(_11889_));
 sg13g2_nor2_1 _18947_ (.A(_10411_),
    .B(net2750),
    .Y(_11890_));
 sg13g2_nand3_1 _18948_ (.B(_10722_),
    .C(_11785_),
    .A(\u_inv.f_next[168] ),
    .Y(_11891_));
 sg13g2_o21ai_1 _18949_ (.B1(_11891_),
    .Y(_11892_),
    .A1(_10412_),
    .A2(\u_inv.f_reg[169] ));
 sg13g2_a221oi_1 _18950_ (.B2(_11781_),
    .C1(_11889_),
    .B1(_11892_),
    .A1(_11777_),
    .Y(_11893_),
    .A2(_11890_));
 sg13g2_nor2_1 _18951_ (.A(_10409_),
    .B(\u_inv.f_reg[172] ),
    .Y(_11894_));
 sg13g2_nand2_1 _18952_ (.Y(_11895_),
    .A(_11772_),
    .B(_11894_));
 sg13g2_o21ai_1 _18953_ (.B1(_11895_),
    .Y(_11896_),
    .A1(_10408_),
    .A2(\u_inv.f_reg[173] ));
 sg13g2_nand2_1 _18954_ (.Y(_11897_),
    .A(net2630),
    .B(_10716_));
 sg13g2_nor2_1 _18955_ (.A(_11768_),
    .B(_11897_),
    .Y(_11898_));
 sg13g2_a21oi_1 _18956_ (.A1(_11771_),
    .A2(_11896_),
    .Y(_11899_),
    .B1(_11898_));
 sg13g2_o21ai_1 _18957_ (.B1(_11899_),
    .Y(_11900_),
    .A1(_11775_),
    .A2(_11893_));
 sg13g2_a21oi_1 _18958_ (.A1(_11787_),
    .A2(_11888_),
    .Y(_11901_),
    .B1(_11900_));
 sg13g2_o21ai_1 _18959_ (.B1(_11901_),
    .Y(_11902_),
    .A1(_10406_),
    .A2(\u_inv.f_reg[175] ));
 sg13g2_nand2_1 _18960_ (.Y(_11903_),
    .A(\u_inv.f_next[187] ),
    .B(_10703_));
 sg13g2_nor2_1 _18961_ (.A(_10395_),
    .B(net1941),
    .Y(_11904_));
 sg13g2_nand2_1 _18962_ (.Y(_11905_),
    .A(\u_inv.f_next[185] ),
    .B(_10705_));
 sg13g2_nand2_1 _18963_ (.Y(_11906_),
    .A(\u_inv.f_next[184] ),
    .B(_10706_));
 sg13g2_o21ai_1 _18964_ (.B1(_11905_),
    .Y(_11907_),
    .A1(_11745_),
    .A2(_11906_));
 sg13g2_a21oi_1 _18965_ (.A1(_11743_),
    .A2(_11907_),
    .Y(_11908_),
    .B1(_11904_));
 sg13g2_o21ai_1 _18966_ (.B1(_11903_),
    .Y(_11909_),
    .A1(_11740_),
    .A2(_11908_));
 sg13g2_nor2b_1 _18967_ (.A(_11739_),
    .B_N(_11909_),
    .Y(_11910_));
 sg13g2_nor2_1 _18968_ (.A(_10390_),
    .B(\u_inv.f_reg[191] ),
    .Y(_11911_));
 sg13g2_nor2_1 _18969_ (.A(_10391_),
    .B(\u_inv.f_reg[190] ),
    .Y(_11912_));
 sg13g2_nor2_1 _18970_ (.A(_10393_),
    .B(\u_inv.f_reg[188] ),
    .Y(_11913_));
 sg13g2_and2_1 _18971_ (.A(_11734_),
    .B(_11913_),
    .X(_11914_));
 sg13g2_a21oi_1 _18972_ (.A1(\u_inv.f_next[189] ),
    .A2(_10701_),
    .Y(_11915_),
    .B1(_11914_));
 sg13g2_nor2_1 _18973_ (.A(_11732_),
    .B(_11915_),
    .Y(_11916_));
 sg13g2_nor2_1 _18974_ (.A(_11912_),
    .B(_11916_),
    .Y(_11917_));
 sg13g2_nor2_1 _18975_ (.A(_11730_),
    .B(_11917_),
    .Y(_11918_));
 sg13g2_nor2_1 _18976_ (.A(_10402_),
    .B(\u_inv.f_reg[179] ),
    .Y(_11919_));
 sg13g2_nor2_1 _18977_ (.A(_10403_),
    .B(\u_inv.f_reg[178] ),
    .Y(_11920_));
 sg13g2_nand2_1 _18978_ (.Y(_11921_),
    .A(\u_inv.f_next[177] ),
    .B(_10713_));
 sg13g2_nand2_1 _18979_ (.Y(_11922_),
    .A(\u_inv.f_next[176] ),
    .B(_10714_));
 sg13g2_o21ai_1 _18980_ (.B1(_11921_),
    .Y(_11923_),
    .A1(_11760_),
    .A2(_11922_));
 sg13g2_a21o_1 _18981_ (.A2(_11923_),
    .A1(net4433),
    .B1(_11920_),
    .X(_11924_));
 sg13g2_a21oi_1 _18982_ (.A1(_11764_),
    .A2(_11924_),
    .Y(_11925_),
    .B1(_11919_));
 sg13g2_nor2_1 _18983_ (.A(_11758_),
    .B(_11925_),
    .Y(_11926_));
 sg13g2_nand2_1 _18984_ (.Y(_11927_),
    .A(\u_inv.f_next[181] ),
    .B(_10709_));
 sg13g2_nor2_1 _18985_ (.A(_10401_),
    .B(\u_inv.f_reg[180] ),
    .Y(_11928_));
 sg13g2_nand2_1 _18986_ (.Y(_11929_),
    .A(_11757_),
    .B(_11928_));
 sg13g2_nand2_1 _18987_ (.Y(_11930_),
    .A(\u_inv.f_next[182] ),
    .B(_10708_));
 sg13g2_nor2_1 _18988_ (.A(_10398_),
    .B(\u_inv.f_reg[183] ),
    .Y(_11931_));
 sg13g2_a21o_1 _18989_ (.A2(_11929_),
    .A1(_11927_),
    .B1(_11752_),
    .X(_11932_));
 sg13g2_a21oi_1 _18990_ (.A1(_11930_),
    .A2(_11932_),
    .Y(_11933_),
    .B1(_11749_));
 sg13g2_nor3_1 _18991_ (.A(_11926_),
    .B(_11931_),
    .C(_11933_),
    .Y(_11934_));
 sg13g2_nor2_1 _18992_ (.A(_11804_),
    .B(_11873_),
    .Y(_11935_));
 sg13g2_o21ai_1 _18993_ (.B1(_11767_),
    .Y(_11936_),
    .A1(_11902_),
    .A2(_11935_));
 sg13g2_o21ai_1 _18994_ (.B1(_11936_),
    .Y(_11937_),
    .A1(_11748_),
    .A2(_11934_));
 sg13g2_nor4_2 _18995_ (.A(_11910_),
    .B(_11911_),
    .C(_11918_),
    .Y(_11938_),
    .D(_11937_));
 sg13g2_o21ai_1 _18996_ (.B1(_11938_),
    .Y(_11939_),
    .A1(_11650_),
    .A2(_11805_));
 sg13g2_xnor2_1 _18997_ (.Y(_11940_),
    .A(\u_inv.f_next[219] ),
    .B(\u_inv.f_reg[219] ));
 sg13g2_nor2_1 _18998_ (.A(_10363_),
    .B(_10672_),
    .Y(_11941_));
 sg13g2_xor2_1 _18999_ (.B(\u_inv.f_reg[218] ),
    .A(\u_inv.f_next[218] ),
    .X(_11942_));
 sg13g2_xnor2_1 _19000_ (.Y(_11943_),
    .A(\u_inv.f_next[218] ),
    .B(\u_inv.f_reg[218] ));
 sg13g2_xnor2_1 _19001_ (.Y(_11944_),
    .A(\u_inv.f_next[216] ),
    .B(\u_inv.f_reg[216] ));
 sg13g2_xor2_1 _19002_ (.B(\u_inv.f_reg[217] ),
    .A(\u_inv.f_next[217] ),
    .X(_11945_));
 sg13g2_nand3_1 _19003_ (.B(_11943_),
    .C(_11944_),
    .A(_11940_),
    .Y(_11946_));
 sg13g2_nor2_1 _19004_ (.A(_11945_),
    .B(_11946_),
    .Y(_11947_));
 sg13g2_xnor2_1 _19005_ (.Y(_11948_),
    .A(\u_inv.f_next[223] ),
    .B(\u_inv.f_reg[223] ));
 sg13g2_nand2_1 _19006_ (.Y(_11949_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_xnor2_1 _19007_ (.Y(_11950_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_and2_1 _19008_ (.A(_11948_),
    .B(_11950_),
    .X(_11951_));
 sg13g2_xor2_1 _19009_ (.B(\u_inv.f_reg[221] ),
    .A(\u_inv.f_next[221] ),
    .X(_11952_));
 sg13g2_xnor2_1 _19010_ (.Y(_11953_),
    .A(\u_inv.f_next[221] ),
    .B(\u_inv.f_reg[221] ));
 sg13g2_nor2_1 _19011_ (.A(_10361_),
    .B(_10670_),
    .Y(_11954_));
 sg13g2_xor2_1 _19012_ (.B(\u_inv.f_reg[220] ),
    .A(\u_inv.f_next[220] ),
    .X(_11955_));
 sg13g2_nor2_1 _19013_ (.A(_11952_),
    .B(_11955_),
    .Y(_11956_));
 sg13g2_nand3_1 _19014_ (.B(_11951_),
    .C(_11956_),
    .A(_11947_),
    .Y(_11957_));
 sg13g2_xnor2_1 _19015_ (.Y(_11958_),
    .A(\u_inv.f_next[211] ),
    .B(\u_inv.f_reg[211] ));
 sg13g2_nand2_1 _19016_ (.Y(_11959_),
    .A(\u_inv.f_next[210] ),
    .B(\u_inv.f_reg[210] ));
 sg13g2_xnor2_1 _19017_ (.Y(_11960_),
    .A(\u_inv.f_next[210] ),
    .B(\u_inv.f_reg[210] ));
 sg13g2_and2_1 _19018_ (.A(_11958_),
    .B(_11960_),
    .X(_11961_));
 sg13g2_nor2_1 _19019_ (.A(_10373_),
    .B(_10682_),
    .Y(_11962_));
 sg13g2_xor2_1 _19020_ (.B(\u_inv.f_reg[208] ),
    .A(\u_inv.f_next[208] ),
    .X(_11963_));
 sg13g2_xor2_1 _19021_ (.B(\u_inv.f_reg[209] ),
    .A(\u_inv.f_next[209] ),
    .X(_11964_));
 sg13g2_xnor2_1 _19022_ (.Y(_11965_),
    .A(\u_inv.f_next[209] ),
    .B(\u_inv.f_reg[209] ));
 sg13g2_nand3b_1 _19023_ (.B(_11965_),
    .C(_11961_),
    .Y(_11966_),
    .A_N(_11963_));
 sg13g2_xnor2_1 _19024_ (.Y(_11967_),
    .A(\u_inv.f_next[215] ),
    .B(\u_inv.f_reg[215] ));
 sg13g2_nand2_1 _19025_ (.Y(_11968_),
    .A(\u_inv.f_next[214] ),
    .B(\u_inv.f_reg[214] ));
 sg13g2_xnor2_1 _19026_ (.Y(_11969_),
    .A(\u_inv.f_next[214] ),
    .B(\u_inv.f_reg[214] ));
 sg13g2_nand2_1 _19027_ (.Y(_11970_),
    .A(_11967_),
    .B(_11969_));
 sg13g2_xnor2_1 _19028_ (.Y(_11971_),
    .A(\u_inv.f_next[213] ),
    .B(\u_inv.f_reg[213] ));
 sg13g2_inv_2 _19029_ (.Y(_11972_),
    .A(_11971_));
 sg13g2_nand2_1 _19030_ (.Y(_11973_),
    .A(\u_inv.f_next[212] ),
    .B(\u_inv.f_reg[212] ));
 sg13g2_xnor2_1 _19031_ (.Y(_11974_),
    .A(\u_inv.f_next[212] ),
    .B(\u_inv.f_reg[212] ));
 sg13g2_nand4_1 _19032_ (.B(_11969_),
    .C(_11971_),
    .A(_11967_),
    .Y(_11975_),
    .D(_11974_));
 sg13g2_or2_1 _19033_ (.X(_11976_),
    .B(_11975_),
    .A(_11966_));
 sg13g2_nor2_1 _19034_ (.A(_11957_),
    .B(_11976_),
    .Y(_11977_));
 sg13g2_xnor2_1 _19035_ (.Y(_11978_),
    .A(\u_inv.f_next[202] ),
    .B(\u_inv.f_reg[202] ));
 sg13g2_xnor2_1 _19036_ (.Y(_11979_),
    .A(\u_inv.f_next[201] ),
    .B(\u_inv.f_reg[201] ));
 sg13g2_xor2_1 _19037_ (.B(\u_inv.f_reg[203] ),
    .A(\u_inv.f_next[203] ),
    .X(_11980_));
 sg13g2_xnor2_1 _19038_ (.Y(_11981_),
    .A(\u_inv.f_next[203] ),
    .B(\u_inv.f_reg[203] ));
 sg13g2_xnor2_1 _19039_ (.Y(_11982_),
    .A(\u_inv.f_next[205] ),
    .B(\u_inv.f_reg[205] ));
 sg13g2_nand2_1 _19040_ (.Y(_11983_),
    .A(\u_inv.f_next[204] ),
    .B(\u_inv.f_reg[204] ));
 sg13g2_xnor2_1 _19041_ (.Y(_11984_),
    .A(\u_inv.f_next[204] ),
    .B(\u_inv.f_reg[204] ));
 sg13g2_nand2_1 _19042_ (.Y(_11985_),
    .A(_11982_),
    .B(_11984_));
 sg13g2_xor2_1 _19043_ (.B(\u_inv.f_reg[207] ),
    .A(\u_inv.f_next[207] ),
    .X(_11986_));
 sg13g2_nand2_1 _19044_ (.Y(_11987_),
    .A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ));
 sg13g2_nor2_1 _19045_ (.A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ),
    .Y(_11988_));
 sg13g2_xor2_1 _19046_ (.B(\u_inv.f_reg[206] ),
    .A(\u_inv.f_next[206] ),
    .X(_11989_));
 sg13g2_nand2_1 _19047_ (.Y(_11990_),
    .A(\u_inv.f_next[200] ),
    .B(\u_inv.f_reg[200] ));
 sg13g2_xor2_1 _19048_ (.B(\u_inv.f_reg[200] ),
    .A(\u_inv.f_next[200] ),
    .X(_11991_));
 sg13g2_inv_2 _19049_ (.Y(_11992_),
    .A(_11991_));
 sg13g2_nand4_1 _19050_ (.B(_11979_),
    .C(_11981_),
    .A(_11978_),
    .Y(_11993_),
    .D(_11992_));
 sg13g2_nor4_1 _19051_ (.A(_11985_),
    .B(_11986_),
    .C(_11989_),
    .D(_11993_),
    .Y(_11994_));
 sg13g2_xnor2_1 _19052_ (.Y(_11995_),
    .A(\u_inv.f_next[195] ),
    .B(\u_inv.f_reg[195] ));
 sg13g2_nand2_1 _19053_ (.Y(_11996_),
    .A(\u_inv.f_next[194] ),
    .B(\u_inv.f_reg[194] ));
 sg13g2_xnor2_1 _19054_ (.Y(_11997_),
    .A(\u_inv.f_next[194] ),
    .B(\u_inv.f_reg[194] ));
 sg13g2_nand2_1 _19055_ (.Y(_11998_),
    .A(_11995_),
    .B(_11997_));
 sg13g2_xor2_1 _19056_ (.B(\u_inv.f_reg[192] ),
    .A(\u_inv.f_next[192] ),
    .X(_11999_));
 sg13g2_xnor2_1 _19057_ (.Y(_12000_),
    .A(\u_inv.f_next[192] ),
    .B(\u_inv.f_reg[192] ));
 sg13g2_xor2_1 _19058_ (.B(\u_inv.f_reg[193] ),
    .A(\u_inv.f_next[193] ),
    .X(_12001_));
 sg13g2_nor3_1 _19059_ (.A(_11998_),
    .B(_11999_),
    .C(_12001_),
    .Y(_12002_));
 sg13g2_nand2_1 _19060_ (.Y(_12003_),
    .A(\u_inv.f_next[199] ),
    .B(\u_inv.f_reg[199] ));
 sg13g2_xor2_1 _19061_ (.B(\u_inv.f_reg[199] ),
    .A(\u_inv.f_next[199] ),
    .X(_12004_));
 sg13g2_xnor2_1 _19062_ (.Y(_12005_),
    .A(\u_inv.f_next[199] ),
    .B(\u_inv.f_reg[199] ));
 sg13g2_nor2_1 _19063_ (.A(_10383_),
    .B(_10692_),
    .Y(_12006_));
 sg13g2_xnor2_1 _19064_ (.Y(_12007_),
    .A(\u_inv.f_next[198] ),
    .B(\u_inv.f_reg[198] ));
 sg13g2_and2_1 _19065_ (.A(_12005_),
    .B(_12007_),
    .X(_12008_));
 sg13g2_xor2_1 _19066_ (.B(\u_inv.f_reg[197] ),
    .A(\u_inv.f_next[197] ),
    .X(_12009_));
 sg13g2_nor2_1 _19067_ (.A(_10385_),
    .B(_10694_),
    .Y(_12010_));
 sg13g2_xor2_1 _19068_ (.B(\u_inv.f_reg[196] ),
    .A(\u_inv.f_next[196] ),
    .X(_12011_));
 sg13g2_nor2_1 _19069_ (.A(_12009_),
    .B(_12011_),
    .Y(_12012_));
 sg13g2_and3_2 _19070_ (.X(_12013_),
    .A(_12002_),
    .B(_12008_),
    .C(_12012_));
 sg13g2_and2_1 _19071_ (.A(_11994_),
    .B(_12013_),
    .X(_12014_));
 sg13g2_and2_1 _19072_ (.A(_11977_),
    .B(_12014_),
    .X(_12015_));
 sg13g2_nor2_1 _19073_ (.A(_10384_),
    .B(\u_inv.f_reg[197] ),
    .Y(_12016_));
 sg13g2_nand2_1 _19074_ (.Y(_12017_),
    .A(\u_inv.f_next[196] ),
    .B(_10694_));
 sg13g2_nor2_1 _19075_ (.A(_10387_),
    .B(\u_inv.f_reg[194] ),
    .Y(_12018_));
 sg13g2_nand2_1 _19076_ (.Y(_12019_),
    .A(net2771),
    .B(_10697_));
 sg13g2_nor2_1 _19077_ (.A(_10389_),
    .B(\u_inv.f_reg[192] ),
    .Y(_12020_));
 sg13g2_nand2b_1 _19078_ (.Y(_12021_),
    .B(_12020_),
    .A_N(_12001_));
 sg13g2_nand2_1 _19079_ (.Y(_12022_),
    .A(_12019_),
    .B(_12021_));
 sg13g2_and2_1 _19080_ (.A(_11997_),
    .B(_12022_),
    .X(_12023_));
 sg13g2_o21ai_1 _19081_ (.B1(_11995_),
    .Y(_12024_),
    .A1(_12018_),
    .A2(_12023_));
 sg13g2_o21ai_1 _19082_ (.B1(_12024_),
    .Y(_12025_),
    .A1(_10386_),
    .A2(\u_inv.f_reg[195] ));
 sg13g2_nand2b_1 _19083_ (.Y(_12026_),
    .B(_12025_),
    .A_N(_12011_));
 sg13g2_a21oi_1 _19084_ (.A1(_12017_),
    .A2(_12026_),
    .Y(_12027_),
    .B1(_12009_));
 sg13g2_o21ai_1 _19085_ (.B1(_12008_),
    .Y(_12028_),
    .A1(_12016_),
    .A2(_12027_));
 sg13g2_nor2_1 _19086_ (.A(_10383_),
    .B(\u_inv.f_reg[198] ),
    .Y(_12029_));
 sg13g2_o21ai_1 _19087_ (.B1(_12028_),
    .Y(_12030_),
    .A1(_10382_),
    .A2(\u_inv.f_reg[199] ));
 sg13g2_a21o_2 _19088_ (.A2(_12029_),
    .A1(_12005_),
    .B1(_12030_),
    .X(_12031_));
 sg13g2_nor2_1 _19089_ (.A(_10379_),
    .B(\u_inv.f_reg[202] ),
    .Y(_12032_));
 sg13g2_nand2_1 _19090_ (.Y(_12033_),
    .A(\u_inv.f_next[201] ),
    .B(_10689_));
 sg13g2_nand3_1 _19091_ (.B(_10690_),
    .C(_11979_),
    .A(\u_inv.f_next[200] ),
    .Y(_12034_));
 sg13g2_nand2_1 _19092_ (.Y(_12035_),
    .A(_12033_),
    .B(_12034_));
 sg13g2_a21oi_1 _19093_ (.A1(_11978_),
    .A2(_12035_),
    .Y(_12036_),
    .B1(_12032_));
 sg13g2_nor2_1 _19094_ (.A(_11980_),
    .B(_12036_),
    .Y(_12037_));
 sg13g2_a21oi_1 _19095_ (.A1(\u_inv.f_next[203] ),
    .A2(_10687_),
    .Y(_12038_),
    .B1(_12037_));
 sg13g2_nor2_1 _19096_ (.A(_10377_),
    .B(\u_inv.f_reg[204] ),
    .Y(_12039_));
 sg13g2_nand2_1 _19097_ (.Y(_12040_),
    .A(\u_inv.f_next[205] ),
    .B(_10685_));
 sg13g2_o21ai_1 _19098_ (.B1(_12040_),
    .Y(_12041_),
    .A1(_11985_),
    .A2(_12038_));
 sg13g2_a21oi_1 _19099_ (.A1(_11982_),
    .A2(_12039_),
    .Y(_12042_),
    .B1(_12041_));
 sg13g2_nor3_1 _19100_ (.A(_11986_),
    .B(_11989_),
    .C(_12042_),
    .Y(_12043_));
 sg13g2_nand2_1 _19101_ (.Y(_12044_),
    .A(\u_inv.f_next[206] ),
    .B(_10684_));
 sg13g2_a221oi_1 _19102_ (.B2(_12031_),
    .C1(_12043_),
    .B1(_11994_),
    .A1(\u_inv.f_next[207] ),
    .Y(_12045_),
    .A2(_10683_));
 sg13g2_o21ai_1 _19103_ (.B1(_12045_),
    .Y(_12046_),
    .A1(_11986_),
    .A2(_12044_));
 sg13g2_nor2_1 _19104_ (.A(_10367_),
    .B(\u_inv.f_reg[214] ),
    .Y(_12047_));
 sg13g2_nor2_1 _19105_ (.A(_10366_),
    .B(\u_inv.f_reg[215] ),
    .Y(_12048_));
 sg13g2_a21oi_1 _19106_ (.A1(_11967_),
    .A2(_12047_),
    .Y(_12049_),
    .B1(_12048_));
 sg13g2_nor2_1 _19107_ (.A(_10368_),
    .B(\u_inv.f_reg[213] ),
    .Y(_12050_));
 sg13g2_nor2_1 _19108_ (.A(_10369_),
    .B(\u_inv.f_reg[212] ),
    .Y(_12051_));
 sg13g2_a21oi_1 _19109_ (.A1(_11971_),
    .A2(_12051_),
    .Y(_12052_),
    .B1(_12050_));
 sg13g2_nor2_1 _19110_ (.A(_10370_),
    .B(\u_inv.f_reg[211] ),
    .Y(_12053_));
 sg13g2_nor2_1 _19111_ (.A(_10371_),
    .B(\u_inv.f_reg[210] ),
    .Y(_12054_));
 sg13g2_nand2_1 _19112_ (.Y(_12055_),
    .A(\u_inv.f_next[209] ),
    .B(_10681_));
 sg13g2_nand2_1 _19113_ (.Y(_12056_),
    .A(\u_inv.f_next[208] ),
    .B(_10682_));
 sg13g2_o21ai_1 _19114_ (.B1(_12055_),
    .Y(_12057_),
    .A1(_11964_),
    .A2(_12056_));
 sg13g2_a221oi_1 _19115_ (.B2(_11961_),
    .C1(_12053_),
    .B1(_12057_),
    .A1(_11958_),
    .Y(_12058_),
    .A2(_12054_));
 sg13g2_nor2_1 _19116_ (.A(_11975_),
    .B(_12058_),
    .Y(_12059_));
 sg13g2_o21ai_1 _19117_ (.B1(_12049_),
    .Y(_12060_),
    .A1(_11970_),
    .A2(_12052_));
 sg13g2_nor2_1 _19118_ (.A(_12059_),
    .B(_12060_),
    .Y(_12061_));
 sg13g2_nor2_1 _19119_ (.A(_10363_),
    .B(\u_inv.f_reg[218] ),
    .Y(_12062_));
 sg13g2_nor2_1 _19120_ (.A(_10365_),
    .B(\u_inv.f_reg[216] ),
    .Y(_12063_));
 sg13g2_nor3_1 _19121_ (.A(_10365_),
    .B(\u_inv.f_reg[216] ),
    .C(_11945_),
    .Y(_12064_));
 sg13g2_a21oi_1 _19122_ (.A1(\u_inv.f_next[217] ),
    .A2(_10673_),
    .Y(_12065_),
    .B1(_12064_));
 sg13g2_nor2_1 _19123_ (.A(_11942_),
    .B(_12065_),
    .Y(_12066_));
 sg13g2_o21ai_1 _19124_ (.B1(_11940_),
    .Y(_12067_),
    .A1(_12062_),
    .A2(_12066_));
 sg13g2_o21ai_1 _19125_ (.B1(_12067_),
    .Y(_12068_),
    .A1(_10362_),
    .A2(\u_inv.f_reg[219] ));
 sg13g2_nand2_1 _19126_ (.Y(_12069_),
    .A(\u_inv.f_next[220] ),
    .B(_10670_));
 sg13g2_nor2_1 _19127_ (.A(_10360_),
    .B(\u_inv.f_reg[221] ),
    .Y(_12070_));
 sg13g2_a21oi_1 _19128_ (.A1(_11956_),
    .A2(_12068_),
    .Y(_12071_),
    .B1(_12070_));
 sg13g2_o21ai_1 _19129_ (.B1(_12071_),
    .Y(_12072_),
    .A1(_11952_),
    .A2(_12069_));
 sg13g2_nor2_1 _19130_ (.A(_10359_),
    .B(\u_inv.f_reg[222] ),
    .Y(_12073_));
 sg13g2_and2_1 _19131_ (.A(_11948_),
    .B(_12073_),
    .X(_12074_));
 sg13g2_a221oi_1 _19132_ (.B2(_12072_),
    .C1(_12074_),
    .B1(_11951_),
    .A1(\u_inv.f_next[223] ),
    .Y(_12075_),
    .A2(_10667_));
 sg13g2_o21ai_1 _19133_ (.B1(_12075_),
    .Y(_12076_),
    .A1(_11957_),
    .A2(_12061_));
 sg13g2_a21oi_1 _19134_ (.A1(_11977_),
    .A2(_12046_),
    .Y(_12077_),
    .B1(_12076_));
 sg13g2_inv_1 _19135_ (.Y(_12078_),
    .A(_12077_));
 sg13g2_a21o_2 _19136_ (.A2(_12015_),
    .A1(_11939_),
    .B1(_12078_),
    .X(_12079_));
 sg13g2_nand2_1 _19137_ (.Y(_12080_),
    .A(\u_inv.f_next[226] ),
    .B(\u_inv.f_reg[226] ));
 sg13g2_xor2_1 _19138_ (.B(\u_inv.f_reg[226] ),
    .A(\u_inv.f_next[226] ),
    .X(_12081_));
 sg13g2_xnor2_1 _19139_ (.Y(_12082_),
    .A(\u_inv.f_next[226] ),
    .B(\u_inv.f_reg[226] ));
 sg13g2_xor2_1 _19140_ (.B(\u_inv.f_reg[227] ),
    .A(\u_inv.f_next[227] ),
    .X(_12083_));
 sg13g2_xnor2_1 _19141_ (.Y(_12084_),
    .A(\u_inv.f_next[227] ),
    .B(\u_inv.f_reg[227] ));
 sg13g2_xor2_1 _19142_ (.B(\u_inv.f_reg[224] ),
    .A(\u_inv.f_next[224] ),
    .X(_12085_));
 sg13g2_inv_2 _19143_ (.Y(_12086_),
    .A(_12085_));
 sg13g2_xor2_1 _19144_ (.B(\u_inv.f_reg[225] ),
    .A(\u_inv.f_next[225] ),
    .X(_12087_));
 sg13g2_nor4_2 _19145_ (.A(_12081_),
    .B(_12083_),
    .C(_12085_),
    .Y(_12088_),
    .D(_12087_));
 sg13g2_xor2_1 _19146_ (.B(\u_inv.f_reg[231] ),
    .A(\u_inv.f_next[231] ),
    .X(_12089_));
 sg13g2_nand2_1 _19147_ (.Y(_12090_),
    .A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ));
 sg13g2_xor2_1 _19148_ (.B(\u_inv.f_reg[230] ),
    .A(\u_inv.f_next[230] ),
    .X(_12091_));
 sg13g2_xnor2_1 _19149_ (.Y(_12092_),
    .A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ));
 sg13g2_xor2_1 _19150_ (.B(\u_inv.f_reg[229] ),
    .A(\u_inv.f_next[229] ),
    .X(_12093_));
 sg13g2_xnor2_1 _19151_ (.Y(_12094_),
    .A(\u_inv.f_next[229] ),
    .B(\u_inv.f_reg[229] ));
 sg13g2_xor2_1 _19152_ (.B(\u_inv.f_reg[228] ),
    .A(\u_inv.f_next[228] ),
    .X(_12095_));
 sg13g2_xnor2_1 _19153_ (.Y(_12096_),
    .A(\u_inv.f_next[228] ),
    .B(\u_inv.f_reg[228] ));
 sg13g2_nor4_1 _19154_ (.A(_12089_),
    .B(_12091_),
    .C(_12093_),
    .D(_12095_),
    .Y(_12097_));
 sg13g2_xnor2_1 _19155_ (.Y(_12098_),
    .A(\u_inv.f_next[235] ),
    .B(\u_inv.f_reg[235] ));
 sg13g2_nand2_1 _19156_ (.Y(_12099_),
    .A(\u_inv.f_next[234] ),
    .B(\u_inv.f_reg[234] ));
 sg13g2_xnor2_1 _19157_ (.Y(_12100_),
    .A(\u_inv.f_next[234] ),
    .B(\u_inv.f_reg[234] ));
 sg13g2_and2_1 _19158_ (.A(_12098_),
    .B(_12100_),
    .X(_12101_));
 sg13g2_nand2_1 _19159_ (.Y(_12102_),
    .A(\u_inv.f_next[232] ),
    .B(\u_inv.f_reg[232] ));
 sg13g2_xnor2_1 _19160_ (.Y(_12103_),
    .A(\u_inv.f_next[232] ),
    .B(\u_inv.f_reg[232] ));
 sg13g2_xor2_1 _19161_ (.B(\u_inv.f_reg[233] ),
    .A(\u_inv.f_next[233] ),
    .X(_12104_));
 sg13g2_xnor2_1 _19162_ (.Y(_12105_),
    .A(\u_inv.f_next[233] ),
    .B(\u_inv.f_reg[233] ));
 sg13g2_nand3_1 _19163_ (.B(_12103_),
    .C(_12105_),
    .A(_12101_),
    .Y(_12106_));
 sg13g2_inv_1 _19164_ (.Y(_12107_),
    .A(_12106_));
 sg13g2_nand2_1 _19165_ (.Y(_12108_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_inv_1 _19166_ (.Y(_12109_),
    .A(_12108_));
 sg13g2_xnor2_1 _19167_ (.Y(_12110_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_inv_1 _19168_ (.Y(_12111_),
    .A(_12110_));
 sg13g2_xnor2_1 _19169_ (.Y(_12112_),
    .A(\u_inv.f_next[237] ),
    .B(\u_inv.f_reg[237] ));
 sg13g2_nand2_1 _19170_ (.Y(_12113_),
    .A(_12110_),
    .B(_12112_));
 sg13g2_xor2_1 _19171_ (.B(\u_inv.f_reg[239] ),
    .A(\u_inv.f_next[239] ),
    .X(_12114_));
 sg13g2_nand2_1 _19172_ (.Y(_12115_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_xnor2_1 _19173_ (.Y(_12116_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_inv_1 _19174_ (.Y(_12117_),
    .A(_12116_));
 sg13g2_or3_1 _19175_ (.A(_12113_),
    .B(_12114_),
    .C(_12117_),
    .X(_12118_));
 sg13g2_nor2_1 _19176_ (.A(_12106_),
    .B(_12118_),
    .Y(_12119_));
 sg13g2_and3_1 _19177_ (.X(_12120_),
    .A(_12088_),
    .B(_12097_),
    .C(_12119_));
 sg13g2_nor2_1 _19178_ (.A(_10352_),
    .B(\u_inv.f_reg[229] ),
    .Y(_12121_));
 sg13g2_nand2_1 _19179_ (.Y(_12122_),
    .A(\u_inv.f_next[228] ),
    .B(_10662_));
 sg13g2_nand2_1 _19180_ (.Y(_12123_),
    .A(\u_inv.f_next[227] ),
    .B(_10663_));
 sg13g2_nor2_1 _19181_ (.A(_10355_),
    .B(\u_inv.f_reg[226] ),
    .Y(_12124_));
 sg13g2_nand2_1 _19182_ (.Y(_12125_),
    .A(\u_inv.f_next[225] ),
    .B(_10665_));
 sg13g2_nand2_1 _19183_ (.Y(_12126_),
    .A(\u_inv.f_next[224] ),
    .B(_10666_));
 sg13g2_o21ai_1 _19184_ (.B1(_12125_),
    .Y(_12127_),
    .A1(_12087_),
    .A2(_12126_));
 sg13g2_a21oi_1 _19185_ (.A1(_12082_),
    .A2(_12127_),
    .Y(_12128_),
    .B1(_12124_));
 sg13g2_o21ai_1 _19186_ (.B1(_12123_),
    .Y(_12129_),
    .A1(_12083_),
    .A2(_12128_));
 sg13g2_nand2_1 _19187_ (.Y(_12130_),
    .A(_12096_),
    .B(_12129_));
 sg13g2_a21oi_1 _19188_ (.A1(_12122_),
    .A2(_12130_),
    .Y(_12131_),
    .B1(_12093_));
 sg13g2_nor2_1 _19189_ (.A(_12121_),
    .B(_12131_),
    .Y(_12132_));
 sg13g2_nor3_1 _19190_ (.A(_12089_),
    .B(_12091_),
    .C(_12132_),
    .Y(_12133_));
 sg13g2_nand2_1 _19191_ (.Y(_12134_),
    .A(\u_inv.f_next[230] ),
    .B(_10660_));
 sg13g2_a21oi_1 _19192_ (.A1(\u_inv.f_next[231] ),
    .A2(_10659_),
    .Y(_12135_),
    .B1(_12133_));
 sg13g2_o21ai_1 _19193_ (.B1(_12135_),
    .Y(_12136_),
    .A1(_12089_),
    .A2(_12134_));
 sg13g2_nor2_1 _19194_ (.A(_10345_),
    .B(\u_inv.f_reg[236] ),
    .Y(_12137_));
 sg13g2_nand2_1 _19195_ (.Y(_12138_),
    .A(_12112_),
    .B(_12137_));
 sg13g2_o21ai_1 _19196_ (.B1(_12138_),
    .Y(_12139_),
    .A1(_10344_),
    .A2(\u_inv.f_reg[237] ));
 sg13g2_nor2_1 _19197_ (.A(_10343_),
    .B(\u_inv.f_reg[238] ),
    .Y(_12140_));
 sg13g2_a21oi_1 _19198_ (.A1(_12116_),
    .A2(_12139_),
    .Y(_12141_),
    .B1(_12140_));
 sg13g2_nor2_1 _19199_ (.A(_12114_),
    .B(_12141_),
    .Y(_12142_));
 sg13g2_a21oi_1 _19200_ (.A1(\u_inv.f_next[239] ),
    .A2(_10651_),
    .Y(_12143_),
    .B1(_12142_));
 sg13g2_nor2_1 _19201_ (.A(_10346_),
    .B(\u_inv.f_reg[235] ),
    .Y(_12144_));
 sg13g2_nor2_1 _19202_ (.A(_10347_),
    .B(\u_inv.f_reg[234] ),
    .Y(_12145_));
 sg13g2_nor2_1 _19203_ (.A(_10348_),
    .B(\u_inv.f_reg[233] ),
    .Y(_12146_));
 sg13g2_nand2_1 _19204_ (.Y(_12147_),
    .A(\u_inv.f_next[232] ),
    .B(_10658_));
 sg13g2_nor2_1 _19205_ (.A(_12104_),
    .B(_12147_),
    .Y(_12148_));
 sg13g2_or2_1 _19206_ (.X(_12149_),
    .B(_12148_),
    .A(_12146_));
 sg13g2_a221oi_1 _19207_ (.B2(_12101_),
    .C1(_12144_),
    .B1(_12149_),
    .A1(_12098_),
    .Y(_12150_),
    .A2(_12145_));
 sg13g2_o21ai_1 _19208_ (.B1(_12143_),
    .Y(_12151_),
    .A1(_12118_),
    .A2(_12150_));
 sg13g2_a221oi_1 _19209_ (.B2(_12119_),
    .C1(_12151_),
    .B1(_12136_),
    .A1(_12079_),
    .Y(_12152_),
    .A2(_12120_));
 sg13g2_xor2_1 _19210_ (.B(\u_inv.f_reg[243] ),
    .A(\u_inv.f_next[243] ),
    .X(_12153_));
 sg13g2_nor2_1 _19211_ (.A(_10339_),
    .B(_10648_),
    .Y(_12154_));
 sg13g2_xor2_1 _19212_ (.B(\u_inv.f_reg[242] ),
    .A(\u_inv.f_next[242] ),
    .X(_12155_));
 sg13g2_nor2_1 _19213_ (.A(_12153_),
    .B(_12155_),
    .Y(_12156_));
 sg13g2_xor2_1 _19214_ (.B(\u_inv.f_reg[240] ),
    .A(\u_inv.f_next[240] ),
    .X(_12157_));
 sg13g2_xnor2_1 _19215_ (.Y(_12158_),
    .A(\u_inv.f_next[240] ),
    .B(\u_inv.f_reg[240] ));
 sg13g2_xor2_1 _19216_ (.B(\u_inv.f_reg[241] ),
    .A(\u_inv.f_next[241] ),
    .X(_12159_));
 sg13g2_xnor2_1 _19217_ (.Y(_12160_),
    .A(\u_inv.f_next[241] ),
    .B(\u_inv.f_reg[241] ));
 sg13g2_nand3_1 _19218_ (.B(_12158_),
    .C(_12160_),
    .A(_12156_),
    .Y(_12161_));
 sg13g2_xor2_1 _19219_ (.B(\u_inv.f_reg[245] ),
    .A(\u_inv.f_next[245] ),
    .X(_12162_));
 sg13g2_nor2_1 _19220_ (.A(_10337_),
    .B(_10646_),
    .Y(_12163_));
 sg13g2_xor2_1 _19221_ (.B(\u_inv.f_reg[244] ),
    .A(\u_inv.f_next[244] ),
    .X(_12164_));
 sg13g2_inv_1 _19222_ (.Y(_12165_),
    .A(_12164_));
 sg13g2_xnor2_1 _19223_ (.Y(_12166_),
    .A(\u_inv.f_next[247] ),
    .B(\u_inv.f_reg[247] ));
 sg13g2_nand2_1 _19224_ (.Y(_12167_),
    .A(\u_inv.f_next[246] ),
    .B(\u_inv.f_reg[246] ));
 sg13g2_xnor2_1 _19225_ (.Y(_12168_),
    .A(\u_inv.f_next[246] ),
    .B(\u_inv.f_reg[246] ));
 sg13g2_nand2_1 _19226_ (.Y(_12169_),
    .A(_12166_),
    .B(_12168_));
 sg13g2_or4_1 _19227_ (.A(_12161_),
    .B(_12162_),
    .C(_12164_),
    .D(_12169_),
    .X(_12170_));
 sg13g2_nand2_1 _19228_ (.Y(_12171_),
    .A(\u_inv.f_next[245] ),
    .B(_10645_));
 sg13g2_nor2_1 _19229_ (.A(_10337_),
    .B(\u_inv.f_reg[244] ),
    .Y(_12172_));
 sg13g2_nand2_1 _19230_ (.Y(_12173_),
    .A(\u_inv.f_next[242] ),
    .B(_10648_));
 sg13g2_nand2_1 _19231_ (.Y(_12174_),
    .A(net3309),
    .B(_10649_));
 sg13g2_nand2_1 _19232_ (.Y(_12175_),
    .A(\u_inv.f_next[240] ),
    .B(_10650_));
 sg13g2_o21ai_1 _19233_ (.B1(_12174_),
    .Y(_12176_),
    .A1(_12159_),
    .A2(_12175_));
 sg13g2_nor2_1 _19234_ (.A(_12153_),
    .B(_12173_),
    .Y(_12177_));
 sg13g2_a221oi_1 _19235_ (.B2(_12176_),
    .C1(_12177_),
    .B1(_12156_),
    .A1(\u_inv.f_next[243] ),
    .Y(_12178_),
    .A2(_10647_));
 sg13g2_nor2_1 _19236_ (.A(_12164_),
    .B(_12178_),
    .Y(_12179_));
 sg13g2_nor2_1 _19237_ (.A(_12172_),
    .B(_12179_),
    .Y(_12180_));
 sg13g2_o21ai_1 _19238_ (.B1(_12171_),
    .Y(_12181_),
    .A1(_12162_),
    .A2(_12180_));
 sg13g2_nand2b_1 _19239_ (.Y(_12182_),
    .B(_12181_),
    .A_N(_12169_));
 sg13g2_nor2_1 _19240_ (.A(_10335_),
    .B(\u_inv.f_reg[246] ),
    .Y(_12183_));
 sg13g2_o21ai_1 _19241_ (.B1(_12182_),
    .Y(_12184_),
    .A1(_10334_),
    .A2(\u_inv.f_reg[247] ));
 sg13g2_a21oi_1 _19242_ (.A1(_12166_),
    .A2(_12183_),
    .Y(_12185_),
    .B1(_12184_));
 sg13g2_o21ai_1 _19243_ (.B1(_12185_),
    .Y(_12186_),
    .A1(_12152_),
    .A2(_12170_));
 sg13g2_nand2_1 _19244_ (.Y(_12187_),
    .A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ));
 sg13g2_xnor2_1 _19245_ (.Y(_12188_),
    .A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ));
 sg13g2_xnor2_1 _19246_ (.Y(_12189_),
    .A(\u_inv.f_next[251] ),
    .B(\u_inv.f_reg[251] ));
 sg13g2_xor2_1 _19247_ (.B(\u_inv.f_reg[249] ),
    .A(\u_inv.f_next[249] ),
    .X(_12190_));
 sg13g2_xnor2_1 _19248_ (.Y(_12191_),
    .A(\u_inv.f_next[249] ),
    .B(\u_inv.f_reg[249] ));
 sg13g2_nand2_1 _19249_ (.Y(_12192_),
    .A(\u_inv.f_next[250] ),
    .B(\u_inv.f_reg[250] ));
 sg13g2_xnor2_1 _19250_ (.Y(_12193_),
    .A(\u_inv.f_next[250] ),
    .B(\u_inv.f_reg[250] ));
 sg13g2_and4_1 _19251_ (.A(_12188_),
    .B(_12189_),
    .C(_12191_),
    .D(_12193_),
    .X(_12194_));
 sg13g2_nand2_1 _19252_ (.Y(_12195_),
    .A(net3180),
    .B(_10640_));
 sg13g2_nor2_1 _19253_ (.A(_10332_),
    .B(\u_inv.f_reg[249] ),
    .Y(_12196_));
 sg13g2_nor2_1 _19254_ (.A(_10333_),
    .B(\u_inv.f_reg[248] ),
    .Y(_12197_));
 sg13g2_nor3_1 _19255_ (.A(_10333_),
    .B(\u_inv.f_reg[248] ),
    .C(_12190_),
    .Y(_12198_));
 sg13g2_o21ai_1 _19256_ (.B1(_12193_),
    .Y(_12199_),
    .A1(_12196_),
    .A2(_12198_));
 sg13g2_nand2_1 _19257_ (.Y(_12200_),
    .A(_12195_),
    .B(_12199_));
 sg13g2_and2_1 _19258_ (.A(_12189_),
    .B(_12200_),
    .X(_12201_));
 sg13g2_a221oi_1 _19259_ (.B2(_12194_),
    .C1(_12201_),
    .B1(_12186_),
    .A1(\u_inv.f_next[251] ),
    .Y(_12202_),
    .A2(_10639_));
 sg13g2_xnor2_1 _19260_ (.Y(_12203_),
    .A(\u_inv.f_next[253] ),
    .B(\u_inv.f_reg[253] ));
 sg13g2_nand2_1 _19261_ (.Y(_12204_),
    .A(\u_inv.f_next[252] ),
    .B(\u_inv.f_reg[252] ));
 sg13g2_xor2_1 _19262_ (.B(\u_inv.f_reg[252] ),
    .A(\u_inv.f_next[252] ),
    .X(_12205_));
 sg13g2_xnor2_1 _19263_ (.Y(_12206_),
    .A(\u_inv.f_next[252] ),
    .B(\u_inv.f_reg[252] ));
 sg13g2_nand2_1 _19264_ (.Y(_12207_),
    .A(_12203_),
    .B(_12206_));
 sg13g2_nor2_1 _19265_ (.A(_10328_),
    .B(\u_inv.f_reg[253] ),
    .Y(_12208_));
 sg13g2_nor2_1 _19266_ (.A(_10329_),
    .B(\u_inv.f_reg[252] ),
    .Y(_12209_));
 sg13g2_a21oi_1 _19267_ (.A1(_12203_),
    .A2(_12209_),
    .Y(_12210_),
    .B1(_12208_));
 sg13g2_o21ai_1 _19268_ (.B1(_12210_),
    .Y(_12211_),
    .A1(_12202_),
    .A2(_12207_));
 sg13g2_a21o_1 _19269_ (.A2(_12211_),
    .A1(_11078_),
    .B1(_11075_),
    .X(_12212_));
 sg13g2_nor2_1 _19270_ (.A(net4596),
    .B(\u_inv.delta_reg[9] ),
    .Y(_12213_));
 sg13g2_nand2_2 _19271_ (.Y(_12214_),
    .A(net4712),
    .B(_10631_));
 sg13g2_or3_1 _19272_ (.A(\u_inv.delta_reg[1] ),
    .B(\u_inv.delta_reg[3] ),
    .C(\u_inv.delta_reg[2] ),
    .X(_12215_));
 sg13g2_nand2b_1 _19273_ (.Y(_12216_),
    .B(_10629_),
    .A_N(_12215_));
 sg13g2_nor3_1 _19274_ (.A(\u_inv.delta_reg[5] ),
    .B(\u_inv.delta_reg[6] ),
    .C(_12216_),
    .Y(_12217_));
 sg13g2_nand2_1 _19275_ (.Y(_12218_),
    .A(_10630_),
    .B(_12217_));
 sg13g2_nor2_1 _19276_ (.A(net1873),
    .B(_12218_),
    .Y(_12219_));
 sg13g2_nor2_2 _19277_ (.A(_12214_),
    .B(_12219_),
    .Y(_12220_));
 sg13g2_a21oi_2 _19278_ (.B1(_12220_),
    .Y(_12221_),
    .A2(_12213_),
    .A1(\u_inv.delta_reg[0] ));
 sg13g2_a21o_2 _19279_ (.A2(_12213_),
    .A1(\u_inv.delta_reg[0] ),
    .B1(_12220_),
    .X(_12222_));
 sg13g2_a21oi_1 _19280_ (.A1(_11070_),
    .A2(_12212_),
    .Y(_12223_),
    .B1(net3825));
 sg13g2_o21ai_1 _19281_ (.B1(_12223_),
    .Y(_12224_),
    .A1(net4959),
    .A2(net4502));
 sg13g2_nand2_1 _19282_ (.Y(_12225_),
    .A(net4685),
    .B(net3851));
 sg13g2_nor2_1 _19283_ (.A(_12166_),
    .B(_12168_),
    .Y(_12226_));
 sg13g2_and2_1 _19284_ (.A(_12162_),
    .B(_12164_),
    .X(_12227_));
 sg13g2_nand2_1 _19285_ (.Y(_12228_),
    .A(_12226_),
    .B(_12227_));
 sg13g2_nand2_1 _19286_ (.Y(_12229_),
    .A(_12153_),
    .B(_12155_));
 sg13g2_a22oi_1 _19287_ (.Y(_12230_),
    .B1(\u_inv.f_reg[240] ),
    .B2(\u_inv.f_next[240] ),
    .A2(\u_inv.f_reg[241] ),
    .A1(\u_inv.f_next[241] ));
 sg13g2_a21o_1 _19288_ (.A2(_10649_),
    .A1(_10340_),
    .B1(_12230_),
    .X(_12231_));
 sg13g2_nor2_1 _19289_ (.A(_12229_),
    .B(_12231_),
    .Y(_12232_));
 sg13g2_o21ai_1 _19290_ (.B1(_12154_),
    .Y(_12233_),
    .A1(\u_inv.f_next[243] ),
    .A2(\u_inv.f_reg[243] ));
 sg13g2_o21ai_1 _19291_ (.B1(_12233_),
    .Y(_12234_),
    .A1(_10338_),
    .A2(_10647_));
 sg13g2_nor2_1 _19292_ (.A(_12232_),
    .B(_12234_),
    .Y(_12235_));
 sg13g2_a21oi_1 _19293_ (.A1(\u_inv.f_next[245] ),
    .A2(\u_inv.f_reg[245] ),
    .Y(_12236_),
    .B1(_12163_));
 sg13g2_a21oi_1 _19294_ (.A1(_10336_),
    .A2(_10645_),
    .Y(_12237_),
    .B1(_12236_));
 sg13g2_a21oi_1 _19295_ (.A1(_10334_),
    .A2(_10643_),
    .Y(_12238_),
    .B1(_12167_));
 sg13g2_a221oi_1 _19296_ (.B2(_12237_),
    .C1(_12238_),
    .B1(_12226_),
    .A1(\u_inv.f_next[247] ),
    .Y(_12239_),
    .A2(\u_inv.f_reg[247] ));
 sg13g2_o21ai_1 _19297_ (.B1(_12239_),
    .Y(_12240_),
    .A1(_12228_),
    .A2(_12235_));
 sg13g2_nor2_1 _19298_ (.A(_11948_),
    .B(_11950_),
    .Y(_12241_));
 sg13g2_and2_1 _19299_ (.A(_11952_),
    .B(_11955_),
    .X(_12242_));
 sg13g2_nand2_1 _19300_ (.Y(_12243_),
    .A(_12241_),
    .B(_12242_));
 sg13g2_nor2_1 _19301_ (.A(_11940_),
    .B(_11943_),
    .Y(_12244_));
 sg13g2_nand2_1 _19302_ (.Y(_12245_),
    .A(_11945_),
    .B(_12244_));
 sg13g2_nor3_2 _19303_ (.A(_11944_),
    .B(_12243_),
    .C(_12245_),
    .Y(_12246_));
 sg13g2_nor2_1 _19304_ (.A(_11967_),
    .B(_11969_),
    .Y(_12247_));
 sg13g2_nor2_1 _19305_ (.A(_11971_),
    .B(_11974_),
    .Y(_12248_));
 sg13g2_nand2_1 _19306_ (.Y(_12249_),
    .A(_12247_),
    .B(_12248_));
 sg13g2_nand2_1 _19307_ (.Y(_12250_),
    .A(_11963_),
    .B(_11964_));
 sg13g2_or2_1 _19308_ (.X(_12251_),
    .B(_11960_),
    .A(_11958_));
 sg13g2_nor3_1 _19309_ (.A(_12249_),
    .B(_12250_),
    .C(_12251_),
    .Y(_12252_));
 sg13g2_nand2_2 _19310_ (.Y(_12253_),
    .A(_12246_),
    .B(_12252_));
 sg13g2_nor2_1 _19311_ (.A(_12005_),
    .B(_12007_),
    .Y(_12254_));
 sg13g2_and2_1 _19312_ (.A(_12009_),
    .B(_12011_),
    .X(_12255_));
 sg13g2_and2_1 _19313_ (.A(_12254_),
    .B(_12255_),
    .X(_12256_));
 sg13g2_or2_1 _19314_ (.X(_12257_),
    .B(_11997_),
    .A(_11995_));
 sg13g2_a22oi_1 _19315_ (.Y(_12258_),
    .B1(\u_inv.f_reg[192] ),
    .B2(\u_inv.f_next[192] ),
    .A2(\u_inv.f_reg[193] ),
    .A1(\u_inv.f_next[193] ));
 sg13g2_a21oi_1 _19316_ (.A1(_10388_),
    .A2(_10697_),
    .Y(_12259_),
    .B1(_12258_));
 sg13g2_nor2b_1 _19317_ (.A(_12257_),
    .B_N(_12259_),
    .Y(_12260_));
 sg13g2_a22oi_1 _19318_ (.Y(_12261_),
    .B1(\u_inv.f_reg[194] ),
    .B2(\u_inv.f_next[194] ),
    .A2(\u_inv.f_reg[195] ),
    .A1(\u_inv.f_next[195] ));
 sg13g2_a21oi_1 _19319_ (.A1(_10386_),
    .A2(_10695_),
    .Y(_12262_),
    .B1(_12261_));
 sg13g2_o21ai_1 _19320_ (.B1(_12256_),
    .Y(_12263_),
    .A1(_12260_),
    .A2(_12262_));
 sg13g2_o21ai_1 _19321_ (.B1(_12006_),
    .Y(_12264_),
    .A1(\u_inv.f_next[199] ),
    .A2(\u_inv.f_reg[199] ));
 sg13g2_a21oi_1 _19322_ (.A1(\u_inv.f_next[197] ),
    .A2(\u_inv.f_reg[197] ),
    .Y(_12265_),
    .B1(_12010_));
 sg13g2_a21oi_1 _19323_ (.A1(_10384_),
    .A2(_10693_),
    .Y(_12266_),
    .B1(_12265_));
 sg13g2_nand2_1 _19324_ (.Y(_12267_),
    .A(_12254_),
    .B(_12266_));
 sg13g2_nand4_1 _19325_ (.B(_12263_),
    .C(_12264_),
    .A(_12003_),
    .Y(_12268_),
    .D(_12267_));
 sg13g2_nor2_1 _19326_ (.A(_11982_),
    .B(_11984_),
    .Y(_12269_));
 sg13g2_nand3_1 _19327_ (.B(_11989_),
    .C(_12269_),
    .A(_11986_),
    .Y(_12270_));
 sg13g2_inv_1 _19328_ (.Y(_12271_),
    .A(_12270_));
 sg13g2_nand2b_1 _19329_ (.Y(_12272_),
    .B(_11980_),
    .A_N(_11978_));
 sg13g2_nand2b_1 _19330_ (.Y(_12273_),
    .B(_11991_),
    .A_N(_11979_));
 sg13g2_nor3_1 _19331_ (.A(_12270_),
    .B(_12272_),
    .C(_12273_),
    .Y(_12274_));
 sg13g2_a22oi_1 _19332_ (.Y(_12275_),
    .B1(\u_inv.f_reg[204] ),
    .B2(\u_inv.f_next[204] ),
    .A2(\u_inv.f_reg[205] ),
    .A1(\u_inv.f_next[205] ));
 sg13g2_a21oi_1 _19333_ (.A1(_10376_),
    .A2(_10685_),
    .Y(_12276_),
    .B1(_12275_));
 sg13g2_nand3_1 _19334_ (.B(_11989_),
    .C(_12276_),
    .A(_11986_),
    .Y(_12277_));
 sg13g2_a22oi_1 _19335_ (.Y(_12278_),
    .B1(\u_inv.f_reg[206] ),
    .B2(\u_inv.f_next[206] ),
    .A2(\u_inv.f_reg[207] ),
    .A1(\u_inv.f_next[207] ));
 sg13g2_a21o_1 _19336_ (.A2(_10683_),
    .A1(_10374_),
    .B1(_12278_),
    .X(_12279_));
 sg13g2_a22oi_1 _19337_ (.Y(_12280_),
    .B1(\u_inv.f_reg[200] ),
    .B2(\u_inv.f_next[200] ),
    .A2(\u_inv.f_reg[201] ),
    .A1(\u_inv.f_next[201] ));
 sg13g2_a21o_1 _19338_ (.A2(_10689_),
    .A1(_10380_),
    .B1(_12280_),
    .X(_12281_));
 sg13g2_nor2_1 _19339_ (.A(_12272_),
    .B(_12281_),
    .Y(_12282_));
 sg13g2_a22oi_1 _19340_ (.Y(_12283_),
    .B1(\u_inv.f_reg[202] ),
    .B2(\u_inv.f_next[202] ),
    .A2(\u_inv.f_reg[203] ),
    .A1(\u_inv.f_next[203] ));
 sg13g2_a21oi_1 _19341_ (.A1(_10378_),
    .A2(_10687_),
    .Y(_12284_),
    .B1(_12283_));
 sg13g2_o21ai_1 _19342_ (.B1(_12271_),
    .Y(_12285_),
    .A1(_12282_),
    .A2(_12284_));
 sg13g2_nand3_1 _19343_ (.B(_12279_),
    .C(_12285_),
    .A(_12277_),
    .Y(_12286_));
 sg13g2_a21oi_1 _19344_ (.A1(_12268_),
    .A2(_12274_),
    .Y(_12287_),
    .B1(_12286_));
 sg13g2_a21o_1 _19345_ (.A2(_12274_),
    .A1(_12268_),
    .B1(_12286_),
    .X(_12288_));
 sg13g2_a22oi_1 _19346_ (.Y(_12289_),
    .B1(\u_inv.f_reg[216] ),
    .B2(\u_inv.f_next[216] ),
    .A2(\u_inv.f_reg[217] ),
    .A1(\u_inv.f_next[217] ));
 sg13g2_a21oi_1 _19347_ (.A1(_10364_),
    .A2(_10673_),
    .Y(_12290_),
    .B1(_12289_));
 sg13g2_o21ai_1 _19348_ (.B1(_11941_),
    .Y(_12291_),
    .A1(\u_inv.f_next[219] ),
    .A2(\u_inv.f_reg[219] ));
 sg13g2_a22oi_1 _19349_ (.Y(_12292_),
    .B1(_12244_),
    .B2(_12290_),
    .A2(\u_inv.f_reg[219] ),
    .A1(\u_inv.f_next[219] ));
 sg13g2_and2_1 _19350_ (.A(_12291_),
    .B(_12292_),
    .X(_12293_));
 sg13g2_a21oi_1 _19351_ (.A1(\u_inv.f_next[221] ),
    .A2(\u_inv.f_reg[221] ),
    .Y(_12294_),
    .B1(_11954_));
 sg13g2_a21oi_1 _19352_ (.A1(_10360_),
    .A2(_10669_),
    .Y(_12295_),
    .B1(_12294_));
 sg13g2_a21oi_1 _19353_ (.A1(_10358_),
    .A2(_10667_),
    .Y(_12296_),
    .B1(_11949_));
 sg13g2_a221oi_1 _19354_ (.B2(_12295_),
    .C1(_12296_),
    .B1(_12241_),
    .A1(\u_inv.f_next[223] ),
    .Y(_12297_),
    .A2(\u_inv.f_reg[223] ));
 sg13g2_o21ai_1 _19355_ (.B1(_12297_),
    .Y(_12298_),
    .A1(_12243_),
    .A2(_12293_));
 sg13g2_a21oi_1 _19356_ (.A1(\u_inv.f_next[209] ),
    .A2(\u_inv.f_reg[209] ),
    .Y(_12299_),
    .B1(_11962_));
 sg13g2_a21o_1 _19357_ (.A2(_10681_),
    .A1(_10372_),
    .B1(_12299_),
    .X(_12300_));
 sg13g2_nor2_1 _19358_ (.A(_12251_),
    .B(_12300_),
    .Y(_12301_));
 sg13g2_a22oi_1 _19359_ (.Y(_12302_),
    .B1(\u_inv.f_reg[210] ),
    .B2(\u_inv.f_next[210] ),
    .A2(\u_inv.f_reg[211] ),
    .A1(\u_inv.f_next[211] ));
 sg13g2_a21oi_1 _19360_ (.A1(_10370_),
    .A2(_10679_),
    .Y(_12303_),
    .B1(_12302_));
 sg13g2_nor2_1 _19361_ (.A(_12301_),
    .B(_12303_),
    .Y(_12304_));
 sg13g2_a21oi_1 _19362_ (.A1(_10366_),
    .A2(_10675_),
    .Y(_12305_),
    .B1(_11968_));
 sg13g2_a22oi_1 _19363_ (.Y(_12306_),
    .B1(\u_inv.f_reg[212] ),
    .B2(\u_inv.f_next[212] ),
    .A2(\u_inv.f_reg[213] ),
    .A1(\u_inv.f_next[213] ));
 sg13g2_a21oi_1 _19364_ (.A1(_10368_),
    .A2(_10677_),
    .Y(_12307_),
    .B1(_12306_));
 sg13g2_a221oi_1 _19365_ (.B2(_12307_),
    .C1(_12305_),
    .B1(_12247_),
    .A1(\u_inv.f_next[215] ),
    .Y(_12308_),
    .A2(\u_inv.f_reg[215] ));
 sg13g2_o21ai_1 _19366_ (.B1(_12308_),
    .Y(_12309_),
    .A1(_12249_),
    .A2(_12304_));
 sg13g2_a21oi_1 _19367_ (.A1(_12246_),
    .A2(_12309_),
    .Y(_12310_),
    .B1(_12298_));
 sg13g2_o21ai_1 _19368_ (.B1(_12310_),
    .Y(_12311_),
    .A1(_12253_),
    .A2(_12287_));
 sg13g2_nor2_1 _19369_ (.A(_11741_),
    .B(_11743_),
    .Y(_12312_));
 sg13g2_nand2_1 _19370_ (.Y(_12313_),
    .A(_11745_),
    .B(_12312_));
 sg13g2_and2_1 _19371_ (.A(_11730_),
    .B(_11732_),
    .X(_12314_));
 sg13g2_nor2_1 _19372_ (.A(_11734_),
    .B(_11737_),
    .Y(_12315_));
 sg13g2_nand2_1 _19373_ (.Y(_12316_),
    .A(_12314_),
    .B(_12315_));
 sg13g2_nor3_2 _19374_ (.A(_11744_),
    .B(_12313_),
    .C(_12316_),
    .Y(_12317_));
 sg13g2_nor2_1 _19375_ (.A(_11750_),
    .B(_11753_),
    .Y(_12318_));
 sg13g2_nor2_1 _19376_ (.A(_11756_),
    .B(_11757_),
    .Y(_12319_));
 sg13g2_nand2_1 _19377_ (.Y(_12320_),
    .A(_12318_),
    .B(_12319_));
 sg13g2_or2_1 _19378_ (.X(_12321_),
    .B(_11764_),
    .A(net4433));
 sg13g2_a22oi_1 _19379_ (.Y(_12322_),
    .B1(\u_inv.f_reg[176] ),
    .B2(\u_inv.f_next[176] ),
    .A2(\u_inv.f_reg[177] ),
    .A1(\u_inv.f_next[177] ));
 sg13g2_a21oi_1 _19380_ (.A1(_10404_),
    .A2(_10713_),
    .Y(_12323_),
    .B1(_12322_));
 sg13g2_nand2b_1 _19381_ (.Y(_12324_),
    .B(_12323_),
    .A_N(_12321_));
 sg13g2_a22oi_1 _19382_ (.Y(_12325_),
    .B1(\u_inv.f_reg[178] ),
    .B2(\u_inv.f_next[178] ),
    .A2(\u_inv.f_reg[179] ),
    .A1(\u_inv.f_next[179] ));
 sg13g2_a21o_1 _19383_ (.A2(_10711_),
    .A1(_10402_),
    .B1(_12325_),
    .X(_12326_));
 sg13g2_and2_1 _19384_ (.A(_12324_),
    .B(_12326_),
    .X(_12327_));
 sg13g2_a21oi_1 _19385_ (.A1(_10398_),
    .A2(_10707_),
    .Y(_12328_),
    .B1(_11751_));
 sg13g2_a21oi_1 _19386_ (.A1(\u_inv.f_next[183] ),
    .A2(\u_inv.f_reg[183] ),
    .Y(_12329_),
    .B1(_12328_));
 sg13g2_a21oi_1 _19387_ (.A1(\u_inv.f_next[181] ),
    .A2(\u_inv.f_reg[181] ),
    .Y(_12330_),
    .B1(_11754_));
 sg13g2_a21oi_1 _19388_ (.A1(_10400_),
    .A2(_10709_),
    .Y(_12331_),
    .B1(_12330_));
 sg13g2_o21ai_1 _19389_ (.B1(_12329_),
    .Y(_12332_),
    .A1(_12320_),
    .A2(_12327_));
 sg13g2_a21oi_1 _19390_ (.A1(_12318_),
    .A2(_12331_),
    .Y(_12333_),
    .B1(_12332_));
 sg13g2_inv_1 _19391_ (.Y(_12334_),
    .A(_12333_));
 sg13g2_a22oi_1 _19392_ (.Y(_12335_),
    .B1(\u_inv.f_reg[184] ),
    .B2(\u_inv.f_next[184] ),
    .A2(\u_inv.f_reg[185] ),
    .A1(\u_inv.f_next[185] ));
 sg13g2_a21oi_1 _19393_ (.A1(_10396_),
    .A2(_10705_),
    .Y(_12336_),
    .B1(_12335_));
 sg13g2_a21oi_1 _19394_ (.A1(_10394_),
    .A2(_10703_),
    .Y(_12337_),
    .B1(_11742_));
 sg13g2_a221oi_1 _19395_ (.B2(_12336_),
    .C1(_12337_),
    .B1(_12312_),
    .A1(\u_inv.f_next[187] ),
    .Y(_12338_),
    .A2(\u_inv.f_reg[187] ));
 sg13g2_a21oi_1 _19396_ (.A1(\u_inv.f_next[189] ),
    .A2(\u_inv.f_reg[189] ),
    .Y(_12339_),
    .B1(_11735_));
 sg13g2_a21oi_1 _19397_ (.A1(_10392_),
    .A2(_10701_),
    .Y(_12340_),
    .B1(_12339_));
 sg13g2_a21oi_1 _19398_ (.A1(_10390_),
    .A2(_10699_),
    .Y(_12341_),
    .B1(_11731_));
 sg13g2_a221oi_1 _19399_ (.B2(_12340_),
    .C1(_12341_),
    .B1(_12314_),
    .A1(\u_inv.f_next[191] ),
    .Y(_12342_),
    .A2(\u_inv.f_reg[191] ));
 sg13g2_o21ai_1 _19400_ (.B1(_12342_),
    .Y(_12343_),
    .A1(_12316_),
    .A2(_12338_));
 sg13g2_a21oi_2 _19401_ (.B1(_12343_),
    .Y(_12344_),
    .A2(_12334_),
    .A1(_12317_));
 sg13g2_nand2_1 _19402_ (.Y(_12345_),
    .A(_11759_),
    .B(_11760_));
 sg13g2_inv_1 _19403_ (.Y(_12346_),
    .A(_12345_));
 sg13g2_nor3_1 _19404_ (.A(_12320_),
    .B(_12321_),
    .C(_12345_),
    .Y(_12347_));
 sg13g2_nand2_2 _19405_ (.Y(_12348_),
    .A(_12317_),
    .B(_12347_));
 sg13g2_nand2_1 _19406_ (.Y(_12349_),
    .A(_11768_),
    .B(_11770_));
 sg13g2_or2_1 _19407_ (.X(_12350_),
    .B(_11774_),
    .A(_11772_));
 sg13g2_or2_1 _19408_ (.X(_12351_),
    .B(_12350_),
    .A(_12349_));
 sg13g2_or2_1 _19409_ (.X(_12352_),
    .B(_11785_),
    .A(_11784_));
 sg13g2_nor2_1 _19410_ (.A(_11777_),
    .B(_11780_),
    .Y(_12353_));
 sg13g2_nor4_1 _19411_ (.A(_11777_),
    .B(_11780_),
    .C(_12351_),
    .D(_12352_),
    .Y(_12354_));
 sg13g2_nor2_1 _19412_ (.A(_11795_),
    .B(_11797_),
    .Y(_12355_));
 sg13g2_and2_1 _19413_ (.A(_11798_),
    .B(_11799_),
    .X(_12356_));
 sg13g2_nand2_1 _19414_ (.Y(_12357_),
    .A(_12355_),
    .B(_12356_));
 sg13g2_nor2_1 _19415_ (.A(_11788_),
    .B(_11790_),
    .Y(_12358_));
 sg13g2_a22oi_1 _19416_ (.Y(_12359_),
    .B1(\u_inv.f_reg[160] ),
    .B2(\u_inv.f_next[160] ),
    .A2(\u_inv.f_reg[161] ),
    .A1(\u_inv.f_next[161] ));
 sg13g2_a21oi_1 _19417_ (.A1(_10420_),
    .A2(_10729_),
    .Y(_12360_),
    .B1(_12359_));
 sg13g2_a21oi_1 _19418_ (.A1(_10418_),
    .A2(_10727_),
    .Y(_12361_),
    .B1(_11789_));
 sg13g2_a221oi_1 _19419_ (.B2(_12360_),
    .C1(_12361_),
    .B1(_12358_),
    .A1(\u_inv.f_next[163] ),
    .Y(_12362_),
    .A2(\u_inv.f_reg[163] ));
 sg13g2_a21oi_1 _19420_ (.A1(_10414_),
    .A2(_10723_),
    .Y(_12363_),
    .B1(_11796_));
 sg13g2_a22oi_1 _19421_ (.Y(_12364_),
    .B1(\u_inv.f_reg[164] ),
    .B2(\u_inv.f_next[164] ),
    .A2(\u_inv.f_reg[165] ),
    .A1(\u_inv.f_next[165] ));
 sg13g2_a21oi_1 _19422_ (.A1(_10416_),
    .A2(_10725_),
    .Y(_12365_),
    .B1(_12364_));
 sg13g2_a221oi_1 _19423_ (.B2(_12365_),
    .C1(_12363_),
    .B1(_12355_),
    .A1(\u_inv.f_next[167] ),
    .Y(_12366_),
    .A2(\u_inv.f_reg[167] ));
 sg13g2_o21ai_1 _19424_ (.B1(_12366_),
    .Y(_12367_),
    .A1(_12357_),
    .A2(_12362_));
 sg13g2_a22oi_1 _19425_ (.Y(_12368_),
    .B1(\u_inv.f_reg[172] ),
    .B2(\u_inv.f_next[172] ),
    .A2(\u_inv.f_reg[173] ),
    .A1(\u_inv.f_next[173] ));
 sg13g2_a21o_1 _19426_ (.A2(_10717_),
    .A1(_10408_),
    .B1(_12368_),
    .X(_12369_));
 sg13g2_nor2_1 _19427_ (.A(_12349_),
    .B(_12369_),
    .Y(_12370_));
 sg13g2_a21oi_1 _19428_ (.A1(\u_inv.f_next[175] ),
    .A2(\u_inv.f_reg[175] ),
    .Y(_12371_),
    .B1(_11769_));
 sg13g2_a21oi_1 _19429_ (.A1(_10406_),
    .A2(_10715_),
    .Y(_12372_),
    .B1(_12371_));
 sg13g2_nor2_1 _19430_ (.A(_12370_),
    .B(_12372_),
    .Y(_12373_));
 sg13g2_a22oi_1 _19431_ (.Y(_12374_),
    .B1(\u_inv.f_reg[168] ),
    .B2(\u_inv.f_next[168] ),
    .A2(\u_inv.f_reg[169] ),
    .A1(\u_inv.f_next[169] ));
 sg13g2_a21o_1 _19432_ (.A2(_10721_),
    .A1(_10412_),
    .B1(_12374_),
    .X(_12375_));
 sg13g2_inv_1 _19433_ (.Y(_12376_),
    .A(_12375_));
 sg13g2_o21ai_1 _19434_ (.B1(_11778_),
    .Y(_12377_),
    .A1(\u_inv.f_next[171] ),
    .A2(\u_inv.f_reg[171] ));
 sg13g2_o21ai_1 _19435_ (.B1(_12377_),
    .Y(_12378_),
    .A1(_10410_),
    .A2(_10719_));
 sg13g2_a21oi_1 _19436_ (.A1(_12353_),
    .A2(_12376_),
    .Y(_12379_),
    .B1(_12378_));
 sg13g2_o21ai_1 _19437_ (.B1(_12373_),
    .Y(_12380_),
    .A1(_12351_),
    .A2(_12379_));
 sg13g2_a21oi_1 _19438_ (.A1(_12354_),
    .A2(_12367_),
    .Y(_12381_),
    .B1(_12380_));
 sg13g2_nor2_1 _19439_ (.A(_12348_),
    .B(_12381_),
    .Y(_12382_));
 sg13g2_nand2_1 _19440_ (.Y(_12383_),
    .A(_11695_),
    .B(_11696_));
 sg13g2_nor3_1 _19441_ (.A(_11688_),
    .B(_11689_),
    .C(_11693_),
    .Y(_12384_));
 sg13g2_nor2b_1 _19442_ (.A(_12383_),
    .B_N(_12384_),
    .Y(_12385_));
 sg13g2_nor2_1 _19443_ (.A(_11699_),
    .B(_11702_),
    .Y(_12386_));
 sg13g2_nand2_1 _19444_ (.Y(_12387_),
    .A(_12385_),
    .B(_12386_));
 sg13g2_a22oi_1 _19445_ (.Y(_12388_),
    .B1(\u_inv.f_reg[136] ),
    .B2(\u_inv.f_next[136] ),
    .A2(\u_inv.f_reg[137] ),
    .A1(\u_inv.f_next[137] ));
 sg13g2_nor2_1 _19446_ (.A(_11704_),
    .B(_12388_),
    .Y(_12389_));
 sg13g2_or2_1 _19447_ (.X(_12390_),
    .B(_12388_),
    .A(_11704_));
 sg13g2_a22oi_1 _19448_ (.Y(_12391_),
    .B1(\u_inv.f_reg[138] ),
    .B2(\u_inv.f_next[138] ),
    .A2(\u_inv.f_reg[139] ),
    .A1(\u_inv.f_next[139] ));
 sg13g2_a21oi_1 _19449_ (.A1(_10442_),
    .A2(_10751_),
    .Y(_12392_),
    .B1(_12391_));
 sg13g2_o21ai_1 _19450_ (.B1(_11690_),
    .Y(_12393_),
    .A1(_11688_),
    .A2(_11692_));
 sg13g2_a22oi_1 _19451_ (.Y(_12394_),
    .B1(\u_inv.f_reg[140] ),
    .B2(\u_inv.f_next[140] ),
    .A2(\u_inv.f_reg[141] ),
    .A1(\u_inv.f_next[141] ));
 sg13g2_a21oi_1 _19452_ (.A1(_10440_),
    .A2(_10749_),
    .Y(_12395_),
    .B1(_12394_));
 sg13g2_a221oi_1 _19453_ (.B2(_12384_),
    .C1(_12393_),
    .B1(_12395_),
    .A1(_12385_),
    .Y(_12396_),
    .A2(_12392_));
 sg13g2_o21ai_1 _19454_ (.B1(_12396_),
    .Y(_12397_),
    .A1(_12387_),
    .A2(_12390_));
 sg13g2_nor2_1 _19455_ (.A(_11711_),
    .B(_11714_),
    .Y(_12398_));
 sg13g2_a22oi_1 _19456_ (.Y(_12399_),
    .B1(\u_inv.f_reg[132] ),
    .B2(\u_inv.f_next[132] ),
    .A2(\u_inv.f_reg[133] ),
    .A1(\u_inv.f_next[133] ));
 sg13g2_a21oi_1 _19457_ (.A1(_10448_),
    .A2(_10757_),
    .Y(_12400_),
    .B1(_12399_));
 sg13g2_a22oi_1 _19458_ (.Y(_12401_),
    .B1(_12398_),
    .B2(_12400_),
    .A2(\u_inv.f_reg[135] ),
    .A1(\u_inv.f_next[135] ));
 sg13g2_o21ai_1 _19459_ (.B1(_12401_),
    .Y(_12402_),
    .A1(_11709_),
    .A2(_11712_));
 sg13g2_nor2_1 _19460_ (.A(_11715_),
    .B(_11717_),
    .Y(_12403_));
 sg13g2_and2_1 _19461_ (.A(_12398_),
    .B(_12403_),
    .X(_12404_));
 sg13g2_nand2_2 _19462_ (.Y(_12405_),
    .A(_12398_),
    .B(_12403_));
 sg13g2_nor2_1 _19463_ (.A(_11720_),
    .B(_11722_),
    .Y(_12406_));
 sg13g2_a22oi_1 _19464_ (.Y(_12407_),
    .B1(\u_inv.f_reg[128] ),
    .B2(\u_inv.f_next[128] ),
    .A2(\u_inv.f_reg[129] ),
    .A1(\u_inv.f_next[129] ));
 sg13g2_a21oi_1 _19465_ (.A1(_10452_),
    .A2(_10761_),
    .Y(_12408_),
    .B1(_12407_));
 sg13g2_a21oi_1 _19466_ (.A1(_10450_),
    .A2(_10759_),
    .Y(_12409_),
    .B1(_11721_));
 sg13g2_a221oi_1 _19467_ (.B2(_12408_),
    .C1(_12409_),
    .B1(_12406_),
    .A1(\u_inv.f_next[131] ),
    .Y(_12410_),
    .A2(\u_inv.f_reg[131] ));
 sg13g2_nor2_1 _19468_ (.A(_12405_),
    .B(_12410_),
    .Y(_12411_));
 sg13g2_nor2_1 _19469_ (.A(_12402_),
    .B(_12411_),
    .Y(_12412_));
 sg13g2_nor2_1 _19470_ (.A(_11703_),
    .B(_11706_),
    .Y(_12413_));
 sg13g2_nor2b_2 _19471_ (.A(_12387_),
    .B_N(_12413_),
    .Y(_12414_));
 sg13g2_nor2b_1 _19472_ (.A(_12412_),
    .B_N(_12414_),
    .Y(_12415_));
 sg13g2_nand2b_1 _19473_ (.Y(_12416_),
    .B(_11680_),
    .A_N(_11678_));
 sg13g2_nor2_1 _19474_ (.A(_11683_),
    .B(_11684_),
    .Y(_12417_));
 sg13g2_nor2b_1 _19475_ (.A(_12416_),
    .B_N(_12417_),
    .Y(_12418_));
 sg13g2_and2_1 _19476_ (.A(_11654_),
    .B(_11655_),
    .X(_12419_));
 sg13g2_nand2_1 _19477_ (.Y(_12420_),
    .A(_11651_),
    .B(_11652_));
 sg13g2_nand4_1 _19478_ (.B(_11652_),
    .C(_12418_),
    .A(_11651_),
    .Y(_12421_),
    .D(_12419_));
 sg13g2_and2_1 _19479_ (.A(_11661_),
    .B(_11665_),
    .X(_12422_));
 sg13g2_nand2_1 _19480_ (.Y(_12423_),
    .A(_11659_),
    .B(_11663_));
 sg13g2_inv_1 _19481_ (.Y(_12424_),
    .A(_12423_));
 sg13g2_nand2_1 _19482_ (.Y(_12425_),
    .A(_11668_),
    .B(_11672_));
 sg13g2_nor2_1 _19483_ (.A(_11671_),
    .B(_11674_),
    .Y(_12426_));
 sg13g2_nand2_1 _19484_ (.Y(_12427_),
    .A(_12422_),
    .B(_12426_));
 sg13g2_nor3_2 _19485_ (.A(_12423_),
    .B(_12425_),
    .C(_12427_),
    .Y(_12428_));
 sg13g2_a22oi_1 _19486_ (.Y(_12429_),
    .B1(\u_inv.f_reg[156] ),
    .B2(\u_inv.f_next[156] ),
    .A2(\u_inv.f_reg[157] ),
    .A1(\u_inv.f_next[157] ));
 sg13g2_inv_1 _19487_ (.Y(_12430_),
    .A(_12429_));
 sg13g2_nand3b_1 _19488_ (.B(_12430_),
    .C(_11682_),
    .Y(_12431_),
    .A_N(_12416_));
 sg13g2_o21ai_1 _19489_ (.B1(_11677_),
    .Y(_12432_),
    .A1(_11676_),
    .A2(_11679_));
 sg13g2_a22oi_1 _19490_ (.Y(_12433_),
    .B1(\u_inv.f_reg[152] ),
    .B2(\u_inv.f_next[152] ),
    .A2(\u_inv.f_reg[153] ),
    .A1(\u_inv.f_next[153] ));
 sg13g2_a21oi_1 _19491_ (.A1(_10428_),
    .A2(_10737_),
    .Y(_12434_),
    .B1(_12433_));
 sg13g2_o21ai_1 _19492_ (.B1(_11653_),
    .Y(_12435_),
    .A1(\u_inv.f_next[155] ),
    .A2(\u_inv.f_reg[155] ));
 sg13g2_a22oi_1 _19493_ (.Y(_12436_),
    .B1(_12419_),
    .B2(_12434_),
    .A2(\u_inv.f_reg[155] ),
    .A1(\u_inv.f_next[155] ));
 sg13g2_and2_1 _19494_ (.A(_12435_),
    .B(_12436_),
    .X(_12437_));
 sg13g2_inv_1 _19495_ (.Y(_12438_),
    .A(_12437_));
 sg13g2_a22oi_1 _19496_ (.Y(_12439_),
    .B1(\u_inv.f_reg[144] ),
    .B2(\u_inv.f_next[144] ),
    .A2(\u_inv.f_reg[145] ),
    .A1(\u_inv.f_next[145] ));
 sg13g2_a21oi_1 _19497_ (.A1(_10436_),
    .A2(_10745_),
    .Y(_12440_),
    .B1(_12439_));
 sg13g2_nand2b_1 _19498_ (.Y(_12441_),
    .B(_12440_),
    .A_N(_12425_));
 sg13g2_a22oi_1 _19499_ (.Y(_12442_),
    .B1(\u_inv.f_reg[146] ),
    .B2(\u_inv.f_next[146] ),
    .A2(\u_inv.f_reg[147] ),
    .A1(\u_inv.f_next[147] ));
 sg13g2_a21oi_1 _19500_ (.A1(_10434_),
    .A2(_10743_),
    .Y(_12443_),
    .B1(_12442_));
 sg13g2_inv_1 _19501_ (.Y(_12444_),
    .A(_12443_));
 sg13g2_a21oi_1 _19502_ (.A1(_12441_),
    .A2(_12444_),
    .Y(_12445_),
    .B1(_12423_));
 sg13g2_a22oi_1 _19503_ (.Y(_12446_),
    .B1(\u_inv.f_reg[148] ),
    .B2(\u_inv.f_next[148] ),
    .A2(\u_inv.f_reg[149] ),
    .A1(\u_inv.f_next[149] ));
 sg13g2_a21oi_1 _19504_ (.A1(_10432_),
    .A2(_10741_),
    .Y(_12447_),
    .B1(_12446_));
 sg13g2_or2_1 _19505_ (.X(_12448_),
    .B(_12447_),
    .A(_12445_));
 sg13g2_a22oi_1 _19506_ (.Y(_12449_),
    .B1(\u_inv.f_reg[150] ),
    .B2(\u_inv.f_next[150] ),
    .A2(\u_inv.f_reg[151] ),
    .A1(\u_inv.f_next[151] ));
 sg13g2_a21oi_1 _19507_ (.A1(_10430_),
    .A2(_10739_),
    .Y(_12450_),
    .B1(_12449_));
 sg13g2_a21oi_1 _19508_ (.A1(_12422_),
    .A2(_12448_),
    .Y(_12451_),
    .B1(_12450_));
 sg13g2_inv_1 _19509_ (.Y(_12452_),
    .A(_12451_));
 sg13g2_o21ai_1 _19510_ (.B1(_12428_),
    .Y(_12453_),
    .A1(_12397_),
    .A2(_12415_));
 sg13g2_nand2_1 _19511_ (.Y(_12454_),
    .A(_12414_),
    .B(_12428_));
 sg13g2_a21oi_1 _19512_ (.A1(_12451_),
    .A2(_12453_),
    .Y(_12455_),
    .B1(_12421_));
 sg13g2_a21oi_1 _19513_ (.A1(_12418_),
    .A2(_12438_),
    .Y(_12456_),
    .B1(_12455_));
 sg13g2_nand3b_1 _19514_ (.B(_12456_),
    .C(_12431_),
    .Y(_12457_),
    .A_N(_12432_));
 sg13g2_nand2b_1 _19515_ (.Y(_12458_),
    .B(_12358_),
    .A_N(_11793_));
 sg13g2_nor2_1 _19516_ (.A(_12357_),
    .B(_12458_),
    .Y(_12459_));
 sg13g2_nand2_1 _19517_ (.Y(_12460_),
    .A(_12354_),
    .B(_12459_));
 sg13g2_nor3_1 _19518_ (.A(net4432),
    .B(_12348_),
    .C(_12460_),
    .Y(_12461_));
 sg13g2_a21oi_1 _19519_ (.A1(_12457_),
    .A2(_12461_),
    .Y(_12462_),
    .B1(_12382_));
 sg13g2_and2_1 _19520_ (.A(_12344_),
    .B(_12462_),
    .X(_12463_));
 sg13g2_nor2_1 _19521_ (.A(_11578_),
    .B(_11580_),
    .Y(_12464_));
 sg13g2_nor2b_1 _19522_ (.A(_11572_),
    .B_N(_11575_),
    .Y(_12465_));
 sg13g2_nand2_1 _19523_ (.Y(_12466_),
    .A(_12464_),
    .B(_12465_));
 sg13g2_nor2_1 _19524_ (.A(_11565_),
    .B(_11566_),
    .Y(_12467_));
 sg13g2_a22oi_1 _19525_ (.Y(_12468_),
    .B1(\u_inv.f_reg[96] ),
    .B2(\u_inv.f_next[96] ),
    .A2(\u_inv.f_reg[97] ),
    .A1(\u_inv.f_next[97] ));
 sg13g2_nor2_1 _19526_ (.A(_11568_),
    .B(_12468_),
    .Y(_12469_));
 sg13g2_a22oi_1 _19527_ (.Y(_12470_),
    .B1(\u_inv.f_reg[98] ),
    .B2(\u_inv.f_next[98] ),
    .A2(\u_inv.f_reg[99] ),
    .A1(\u_inv.f_next[99] ));
 sg13g2_a21oi_1 _19528_ (.A1(_10482_),
    .A2(_10791_),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_a21oi_1 _19529_ (.A1(_12467_),
    .A2(_12469_),
    .Y(_12472_),
    .B1(_12471_));
 sg13g2_a21oi_1 _19530_ (.A1(_10478_),
    .A2(_10787_),
    .Y(_12473_),
    .B1(_11579_));
 sg13g2_a21oi_1 _19531_ (.A1(\u_inv.f_next[103] ),
    .A2(\u_inv.f_reg[103] ),
    .Y(_12474_),
    .B1(_12473_));
 sg13g2_a21oi_1 _19532_ (.A1(\u_inv.f_next[101] ),
    .A2(\u_inv.f_reg[101] ),
    .Y(_12475_),
    .B1(_11574_));
 sg13g2_a21oi_1 _19533_ (.A1(_10480_),
    .A2(_10789_),
    .Y(_12476_),
    .B1(_12475_));
 sg13g2_o21ai_1 _19534_ (.B1(_12474_),
    .Y(_12477_),
    .A1(_12466_),
    .A2(_12472_));
 sg13g2_a21oi_1 _19535_ (.A1(_12464_),
    .A2(_12476_),
    .Y(_12478_),
    .B1(_12477_));
 sg13g2_nor2_1 _19536_ (.A(_11520_),
    .B(_11522_),
    .Y(_12479_));
 sg13g2_and2_1 _19537_ (.A(_11524_),
    .B(_11526_),
    .X(_12480_));
 sg13g2_nand2_1 _19538_ (.Y(_12481_),
    .A(_12479_),
    .B(_12480_));
 sg13g2_nor2_1 _19539_ (.A(_11511_),
    .B(_11512_),
    .Y(_12482_));
 sg13g2_nand2_1 _19540_ (.Y(_12483_),
    .A(_11517_),
    .B(_12482_));
 sg13g2_nor3_1 _19541_ (.A(_11514_),
    .B(_12481_),
    .C(_12483_),
    .Y(_12484_));
 sg13g2_nor2_1 _19542_ (.A(_11537_),
    .B(_11539_),
    .Y(_12485_));
 sg13g2_nor2_1 _19543_ (.A(_11541_),
    .B(_11544_),
    .Y(_12486_));
 sg13g2_nand2_1 _19544_ (.Y(_12487_),
    .A(_11529_),
    .B(_11532_));
 sg13g2_and2_1 _19545_ (.A(_11534_),
    .B(_11535_),
    .X(_12488_));
 sg13g2_nand3_1 _19546_ (.B(_12486_),
    .C(_12488_),
    .A(_12485_),
    .Y(_12489_));
 sg13g2_nor2_1 _19547_ (.A(_12487_),
    .B(_12489_),
    .Y(_12490_));
 sg13g2_nand2_2 _19548_ (.Y(_12491_),
    .A(_12484_),
    .B(_12490_));
 sg13g2_inv_1 _19549_ (.Y(_12492_),
    .A(_12491_));
 sg13g2_and2_1 _19550_ (.A(_11550_),
    .B(_11552_),
    .X(_12493_));
 sg13g2_nor2_1 _19551_ (.A(_11554_),
    .B(_11555_),
    .Y(_12494_));
 sg13g2_nand2_1 _19552_ (.Y(_12495_),
    .A(_12493_),
    .B(_12494_));
 sg13g2_inv_1 _19553_ (.Y(_12496_),
    .A(_12495_));
 sg13g2_nor2_1 _19554_ (.A(_11560_),
    .B(_11561_),
    .Y(_12497_));
 sg13g2_nand2_1 _19555_ (.Y(_12498_),
    .A(_11557_),
    .B(_11558_));
 sg13g2_nand4_1 _19556_ (.B(_11558_),
    .C(_12496_),
    .A(_11557_),
    .Y(_12499_),
    .D(_12497_));
 sg13g2_a21oi_1 _19557_ (.A1(\u_inv.f_next[113] ),
    .A2(\u_inv.f_reg[113] ),
    .Y(_12500_),
    .B1(_11533_));
 sg13g2_a21oi_1 _19558_ (.A1(_10468_),
    .A2(_10777_),
    .Y(_12501_),
    .B1(_12500_));
 sg13g2_nand2b_1 _19559_ (.Y(_12502_),
    .B(_12501_),
    .A_N(_12487_));
 sg13g2_a22oi_1 _19560_ (.Y(_12503_),
    .B1(\u_inv.f_reg[114] ),
    .B2(\u_inv.f_next[114] ),
    .A2(\u_inv.f_reg[115] ),
    .A1(\u_inv.f_next[115] ));
 sg13g2_a21o_1 _19561_ (.A2(_10775_),
    .A1(_10466_),
    .B1(_12503_),
    .X(_12504_));
 sg13g2_nand2_1 _19562_ (.Y(_12505_),
    .A(_12502_),
    .B(_12504_));
 sg13g2_nand3_1 _19563_ (.B(_12486_),
    .C(_12505_),
    .A(_12485_),
    .Y(_12506_));
 sg13g2_a21oi_1 _19564_ (.A1(_10462_),
    .A2(_10771_),
    .Y(_12507_),
    .B1(_11538_));
 sg13g2_a21oi_1 _19565_ (.A1(\u_inv.f_next[117] ),
    .A2(\u_inv.f_reg[117] ),
    .Y(_12508_),
    .B1(_11542_));
 sg13g2_a21oi_1 _19566_ (.A1(_10464_),
    .A2(_10773_),
    .Y(_12509_),
    .B1(_12508_));
 sg13g2_a221oi_1 _19567_ (.B2(_12509_),
    .C1(_12507_),
    .B1(_12485_),
    .A1(\u_inv.f_next[119] ),
    .Y(_12510_),
    .A2(\u_inv.f_reg[119] ));
 sg13g2_nand2_1 _19568_ (.Y(_12511_),
    .A(_12506_),
    .B(_12510_));
 sg13g2_a21oi_1 _19569_ (.A1(_11513_),
    .A2(_11515_),
    .Y(_12512_),
    .B1(_11516_));
 sg13g2_a22oi_1 _19570_ (.Y(_12513_),
    .B1(\u_inv.f_reg[122] ),
    .B2(\u_inv.f_next[122] ),
    .A2(\u_inv.f_reg[123] ),
    .A1(\u_inv.f_next[123] ));
 sg13g2_a21oi_1 _19571_ (.A1(_10458_),
    .A2(_10767_),
    .Y(_12514_),
    .B1(_12513_));
 sg13g2_a21oi_2 _19572_ (.B1(_12514_),
    .Y(_12515_),
    .A2(_12512_),
    .A1(_12482_));
 sg13g2_a21oi_1 _19573_ (.A1(_10454_),
    .A2(_10763_),
    .Y(_12516_),
    .B1(_11521_));
 sg13g2_o21ai_1 _19574_ (.B1(_11525_),
    .Y(_12517_),
    .A1(\u_inv.f_next[125] ),
    .A2(\u_inv.f_reg[125] ));
 sg13g2_o21ai_1 _19575_ (.B1(_12517_),
    .Y(_12518_),
    .A1(_10456_),
    .A2(_10765_));
 sg13g2_a221oi_1 _19576_ (.B2(_12518_),
    .C1(_12516_),
    .B1(_12479_),
    .A1(\u_inv.f_next[127] ),
    .Y(_12519_),
    .A2(\u_inv.f_reg[127] ));
 sg13g2_o21ai_1 _19577_ (.B1(_12519_),
    .Y(_12520_),
    .A1(_12481_),
    .A2(_12515_));
 sg13g2_a22oi_1 _19578_ (.Y(_12521_),
    .B1(\u_inv.f_reg[104] ),
    .B2(\u_inv.f_next[104] ),
    .A2(\u_inv.f_reg[105] ),
    .A1(\u_inv.f_next[105] ));
 sg13g2_a21oi_1 _19579_ (.A1(_10476_),
    .A2(_10785_),
    .Y(_12522_),
    .B1(_12521_));
 sg13g2_inv_1 _19580_ (.Y(_12523_),
    .A(_12522_));
 sg13g2_a22oi_1 _19581_ (.Y(_12524_),
    .B1(\u_inv.f_reg[106] ),
    .B2(\u_inv.f_next[106] ),
    .A2(\u_inv.f_reg[107] ),
    .A1(\u_inv.f_next[107] ));
 sg13g2_a21o_1 _19582_ (.A2(_10783_),
    .A1(_10474_),
    .B1(_12524_),
    .X(_12525_));
 sg13g2_inv_1 _19583_ (.Y(_12526_),
    .A(_12525_));
 sg13g2_a21o_1 _19584_ (.A2(_12522_),
    .A1(_12497_),
    .B1(_12526_),
    .X(_12527_));
 sg13g2_o21ai_1 _19585_ (.B1(_11549_),
    .Y(_12528_),
    .A1(_11548_),
    .A2(_11551_));
 sg13g2_a22oi_1 _19586_ (.Y(_12529_),
    .B1(\u_inv.f_reg[108] ),
    .B2(\u_inv.f_next[108] ),
    .A2(\u_inv.f_reg[109] ),
    .A1(\u_inv.f_next[109] ));
 sg13g2_a21oi_1 _19587_ (.A1(_10472_),
    .A2(_10781_),
    .Y(_12530_),
    .B1(_12529_));
 sg13g2_a221oi_1 _19588_ (.B2(_12493_),
    .C1(_12528_),
    .B1(_12530_),
    .A1(_12496_),
    .Y(_12531_),
    .A2(_12527_));
 sg13g2_o21ai_1 _19589_ (.B1(_12531_),
    .Y(_12532_),
    .A1(_12478_),
    .A2(_12499_));
 sg13g2_a22oi_1 _19590_ (.Y(_12533_),
    .B1(_12532_),
    .B2(_12492_),
    .A2(_12511_),
    .A1(_12484_));
 sg13g2_nand2b_2 _19591_ (.Y(_12534_),
    .B(_12533_),
    .A_N(_12520_));
 sg13g2_or2_1 _19592_ (.X(_12535_),
    .B(_11438_),
    .A(_11436_));
 sg13g2_and2_1 _19593_ (.A(_11440_),
    .B(_11442_),
    .X(_12536_));
 sg13g2_nor2b_1 _19594_ (.A(_12535_),
    .B_N(_12536_),
    .Y(_12537_));
 sg13g2_and2_1 _19595_ (.A(_11448_),
    .B(_11452_),
    .X(_12538_));
 sg13g2_nand2_1 _19596_ (.Y(_12539_),
    .A(_11446_),
    .B(_11449_));
 sg13g2_nor2_1 _19597_ (.A(_11455_),
    .B(_11457_),
    .Y(_12540_));
 sg13g2_a22oi_1 _19598_ (.Y(_12541_),
    .B1(\u_inv.f_reg[84] ),
    .B2(\u_inv.f_next[84] ),
    .A2(\u_inv.f_reg[85] ),
    .A1(\u_inv.f_next[85] ));
 sg13g2_a21oi_1 _19599_ (.A1(_10496_),
    .A2(_10805_),
    .Y(_12542_),
    .B1(_12541_));
 sg13g2_a21oi_1 _19600_ (.A1(_10494_),
    .A2(_10803_),
    .Y(_12543_),
    .B1(_11456_));
 sg13g2_a221oi_1 _19601_ (.B2(_12542_),
    .C1(_12543_),
    .B1(_12540_),
    .A1(\u_inv.f_next[87] ),
    .Y(_12544_),
    .A2(\u_inv.f_reg[87] ));
 sg13g2_nor2_1 _19602_ (.A(_11459_),
    .B(_11461_),
    .Y(_12545_));
 sg13g2_nand2_1 _19603_ (.Y(_12546_),
    .A(_12540_),
    .B(_12545_));
 sg13g2_nor4_1 _19604_ (.A(_11376_),
    .B(_11378_),
    .C(_11380_),
    .D(_11382_),
    .Y(_12547_));
 sg13g2_nand2_1 _19605_ (.Y(_12548_),
    .A(_11368_),
    .B(_11370_));
 sg13g2_inv_1 _19606_ (.Y(_12549_),
    .A(_12548_));
 sg13g2_a22oi_1 _19607_ (.Y(_12550_),
    .B1(\u_inv.f_reg[72] ),
    .B2(\u_inv.f_next[72] ),
    .A2(\u_inv.f_reg[73] ),
    .A1(\u_inv.f_next[73] ));
 sg13g2_a21o_1 _19608_ (.A2(_10817_),
    .A1(_10508_),
    .B1(_12550_),
    .X(_12551_));
 sg13g2_nor2_1 _19609_ (.A(_12548_),
    .B(_12551_),
    .Y(_12552_));
 sg13g2_o21ai_1 _19610_ (.B1(_11369_),
    .Y(_12553_),
    .A1(\u_inv.f_next[75] ),
    .A2(\u_inv.f_reg[75] ));
 sg13g2_o21ai_1 _19611_ (.B1(_12553_),
    .Y(_12554_),
    .A1(_10506_),
    .A2(_10815_));
 sg13g2_o21ai_1 _19612_ (.B1(_12547_),
    .Y(_12555_),
    .A1(_12552_),
    .A2(_12554_));
 sg13g2_o21ai_1 _19613_ (.B1(_11377_),
    .Y(_12556_),
    .A1(\u_inv.f_next[79] ),
    .A2(\u_inv.f_reg[79] ));
 sg13g2_a22oi_1 _19614_ (.Y(_12557_),
    .B1(\u_inv.f_reg[76] ),
    .B2(\u_inv.f_next[76] ),
    .A2(\u_inv.f_reg[77] ),
    .A1(\u_inv.f_next[77] ));
 sg13g2_a21o_1 _19615_ (.A2(_10813_),
    .A1(_10504_),
    .B1(_12557_),
    .X(_12558_));
 sg13g2_or3_1 _19616_ (.A(_11376_),
    .B(_11378_),
    .C(_12558_),
    .X(_12559_));
 sg13g2_nand4_1 _19617_ (.B(_12555_),
    .C(_12556_),
    .A(_11375_),
    .Y(_12560_),
    .D(_12559_));
 sg13g2_inv_1 _19618_ (.Y(_12561_),
    .A(_12560_));
 sg13g2_nor2_1 _19619_ (.A(_11464_),
    .B(_11466_),
    .Y(_12562_));
 sg13g2_nand2_1 _19620_ (.Y(_12563_),
    .A(_11471_),
    .B(_12562_));
 sg13g2_inv_1 _19621_ (.Y(_12564_),
    .A(_12563_));
 sg13g2_nand3_1 _19622_ (.B(\u_inv.f_reg[80] ),
    .C(_11469_),
    .A(\u_inv.f_next[80] ),
    .Y(_12565_));
 sg13g2_nand2_1 _19623_ (.Y(_12566_),
    .A(_11470_),
    .B(_12565_));
 sg13g2_a21oi_1 _19624_ (.A1(_10498_),
    .A2(_10807_),
    .Y(_12567_),
    .B1(_11465_));
 sg13g2_a221oi_1 _19625_ (.B2(_12566_),
    .C1(_12567_),
    .B1(_12562_),
    .A1(\u_inv.f_next[83] ),
    .Y(_12568_),
    .A2(\u_inv.f_reg[83] ));
 sg13g2_inv_1 _19626_ (.Y(_12569_),
    .A(_12568_));
 sg13g2_nor2_1 _19627_ (.A(_11395_),
    .B(_11397_),
    .Y(_12570_));
 sg13g2_and2_1 _19628_ (.A(_11398_),
    .B(_11400_),
    .X(_12571_));
 sg13g2_nand2_1 _19629_ (.Y(_12572_),
    .A(_12570_),
    .B(_12571_));
 sg13g2_and2_1 _19630_ (.A(_11385_),
    .B(_11387_),
    .X(_12573_));
 sg13g2_o21ai_1 _19631_ (.B1(_11389_),
    .Y(_12574_),
    .A1(_11388_),
    .A2(_11391_));
 sg13g2_o21ai_1 _19632_ (.B1(_11386_),
    .Y(_12575_),
    .A1(\u_inv.f_next[67] ),
    .A2(\u_inv.f_reg[67] ));
 sg13g2_a22oi_1 _19633_ (.Y(_12576_),
    .B1(_12573_),
    .B2(_12574_),
    .A2(\u_inv.f_reg[67] ),
    .A1(\u_inv.f_next[67] ));
 sg13g2_and2_1 _19634_ (.A(_12575_),
    .B(_12576_),
    .X(_12577_));
 sg13g2_a21oi_1 _19635_ (.A1(_10510_),
    .A2(_10819_),
    .Y(_12578_),
    .B1(_11396_));
 sg13g2_a21oi_1 _19636_ (.A1(\u_inv.f_next[69] ),
    .A2(\u_inv.f_reg[69] ),
    .Y(_12579_),
    .B1(_11399_));
 sg13g2_a21oi_1 _19637_ (.A1(_10512_),
    .A2(_10821_),
    .Y(_12580_),
    .B1(_12579_));
 sg13g2_a221oi_1 _19638_ (.B2(_12580_),
    .C1(_12578_),
    .B1(_12570_),
    .A1(\u_inv.f_next[71] ),
    .Y(_12581_),
    .A2(\u_inv.f_reg[71] ));
 sg13g2_o21ai_1 _19639_ (.B1(_12581_),
    .Y(_12582_),
    .A1(_12572_),
    .A2(_12577_));
 sg13g2_nand2_1 _19640_ (.Y(_12583_),
    .A(_11372_),
    .B(_11373_));
 sg13g2_and4_1 _19641_ (.A(_11372_),
    .B(_11373_),
    .C(_12547_),
    .D(_12549_),
    .X(_12584_));
 sg13g2_a21oi_1 _19642_ (.A1(\u_inv.f_next[93] ),
    .A2(\u_inv.f_reg[93] ),
    .Y(_12585_),
    .B1(_11441_));
 sg13g2_a21oi_1 _19643_ (.A1(_10488_),
    .A2(_10797_),
    .Y(_12586_),
    .B1(_12585_));
 sg13g2_nor2b_2 _19644_ (.A(_12535_),
    .B_N(_12586_),
    .Y(_12587_));
 sg13g2_a21oi_1 _19645_ (.A1(_10486_),
    .A2(_10795_),
    .Y(_12588_),
    .B1(_11437_));
 sg13g2_a21oi_1 _19646_ (.A1(\u_inv.f_next[95] ),
    .A2(\u_inv.f_reg[95] ),
    .Y(_12589_),
    .B1(_12588_));
 sg13g2_a21oi_1 _19647_ (.A1(\u_inv.f_next[89] ),
    .A2(\u_inv.f_reg[89] ),
    .Y(_12590_),
    .B1(_11451_));
 sg13g2_a21oi_1 _19648_ (.A1(_10492_),
    .A2(_10801_),
    .Y(_12591_),
    .B1(_12590_));
 sg13g2_nand2b_1 _19649_ (.Y(_12592_),
    .B(_12591_),
    .A_N(_12539_));
 sg13g2_a22oi_1 _19650_ (.Y(_12593_),
    .B1(\u_inv.f_reg[90] ),
    .B2(\u_inv.f_next[90] ),
    .A2(\u_inv.f_reg[91] ),
    .A1(\u_inv.f_next[91] ));
 sg13g2_a21o_1 _19651_ (.A2(_10799_),
    .A1(_10490_),
    .B1(_12593_),
    .X(_12594_));
 sg13g2_nand2_1 _19652_ (.Y(_12595_),
    .A(_12592_),
    .B(_12594_));
 sg13g2_nand2_1 _19653_ (.Y(_12596_),
    .A(_12537_),
    .B(_12595_));
 sg13g2_o21ai_1 _19654_ (.B1(_12544_),
    .Y(_12597_),
    .A1(_12546_),
    .A2(_12568_));
 sg13g2_nand4_1 _19655_ (.B(_11449_),
    .C(_12537_),
    .A(_11446_),
    .Y(_12598_),
    .D(_12538_));
 sg13g2_nand2b_1 _19656_ (.Y(_12599_),
    .B(_12597_),
    .A_N(_12598_));
 sg13g2_nor4_1 _19657_ (.A(_11468_),
    .B(_12546_),
    .C(_12563_),
    .D(_12598_),
    .Y(_12600_));
 sg13g2_and2_1 _19658_ (.A(_12584_),
    .B(_12600_),
    .X(_12601_));
 sg13g2_a221oi_1 _19659_ (.B2(_12582_),
    .C1(_12587_),
    .B1(_12601_),
    .A1(_12560_),
    .Y(_12602_),
    .A2(_12600_));
 sg13g2_nand4_1 _19660_ (.B(_12596_),
    .C(_12599_),
    .A(_12589_),
    .Y(_12603_),
    .D(_12602_));
 sg13g2_nor2_1 _19661_ (.A(_11312_),
    .B(_11313_),
    .Y(_12604_));
 sg13g2_nand3_1 _19662_ (.B(_11310_),
    .C(_12604_),
    .A(_11309_),
    .Y(_12605_));
 sg13g2_nor2_1 _19663_ (.A(_11316_),
    .B(_11318_),
    .Y(_12606_));
 sg13g2_a22oi_1 _19664_ (.Y(_12607_),
    .B1(\u_inv.f_reg[56] ),
    .B2(\u_inv.f_next[56] ),
    .A2(\u_inv.f_reg[57] ),
    .A1(\u_inv.f_next[57] ));
 sg13g2_a21oi_1 _19665_ (.A1(_10524_),
    .A2(_10833_),
    .Y(_12608_),
    .B1(_12607_));
 sg13g2_a22oi_1 _19666_ (.Y(_12609_),
    .B1(\u_inv.f_reg[58] ),
    .B2(\u_inv.f_next[58] ),
    .A2(\u_inv.f_reg[59] ),
    .A1(\u_inv.f_next[59] ));
 sg13g2_a21oi_1 _19667_ (.A1(_10522_),
    .A2(_10831_),
    .Y(_12610_),
    .B1(_12609_));
 sg13g2_a21oi_1 _19668_ (.A1(_12606_),
    .A2(_12608_),
    .Y(_12611_),
    .B1(_12610_));
 sg13g2_nor2_1 _19669_ (.A(_11324_),
    .B(_11325_),
    .Y(_12612_));
 sg13g2_nand2_1 _19670_ (.Y(_12613_),
    .A(_11327_),
    .B(_11328_));
 sg13g2_nor3_1 _19671_ (.A(_11324_),
    .B(_11325_),
    .C(_12613_),
    .Y(_12614_));
 sg13g2_nor2_1 _19672_ (.A(_11330_),
    .B(_11331_),
    .Y(_12615_));
 sg13g2_a22oi_1 _19673_ (.Y(_12616_),
    .B1(\u_inv.f_reg[48] ),
    .B2(\u_inv.f_next[48] ),
    .A2(\u_inv.f_reg[49] ),
    .A1(\u_inv.f_next[49] ));
 sg13g2_nor4_1 _19674_ (.A(_11330_),
    .B(_11331_),
    .C(_11332_),
    .D(_12616_),
    .Y(_12617_));
 sg13g2_a22oi_1 _19675_ (.Y(_12618_),
    .B1(\u_inv.f_reg[50] ),
    .B2(\u_inv.f_next[50] ),
    .A2(\u_inv.f_reg[51] ),
    .A1(\u_inv.f_next[51] ));
 sg13g2_a21oi_1 _19676_ (.A1(_10530_),
    .A2(_10839_),
    .Y(_12619_),
    .B1(_12618_));
 sg13g2_o21ai_1 _19677_ (.B1(_12614_),
    .Y(_12620_),
    .A1(_12617_),
    .A2(_12619_));
 sg13g2_a22oi_1 _19678_ (.Y(_12621_),
    .B1(\u_inv.f_reg[52] ),
    .B2(\u_inv.f_next[52] ),
    .A2(\u_inv.f_reg[53] ),
    .A1(\u_inv.f_next[53] ));
 sg13g2_a21oi_1 _19679_ (.A1(_10528_),
    .A2(_10837_),
    .Y(_12622_),
    .B1(_12621_));
 sg13g2_a21o_1 _19680_ (.A2(_10837_),
    .A1(_10528_),
    .B1(_12621_),
    .X(_12623_));
 sg13g2_a22oi_1 _19681_ (.Y(_12624_),
    .B1(\u_inv.f_reg[54] ),
    .B2(\u_inv.f_next[54] ),
    .A2(\u_inv.f_reg[55] ),
    .A1(\u_inv.f_next[55] ));
 sg13g2_a21oi_1 _19682_ (.A1(_10526_),
    .A2(_10835_),
    .Y(_12625_),
    .B1(_12624_));
 sg13g2_a21oi_1 _19683_ (.A1(_12612_),
    .A2(_12622_),
    .Y(_12626_),
    .B1(_12625_));
 sg13g2_and2_1 _19684_ (.A(_11317_),
    .B(_11321_),
    .X(_12627_));
 sg13g2_nand2_1 _19685_ (.Y(_12628_),
    .A(_12606_),
    .B(_12627_));
 sg13g2_nor2_1 _19686_ (.A(_12605_),
    .B(_12628_),
    .Y(_12629_));
 sg13g2_inv_1 _19687_ (.Y(_12630_),
    .A(_12629_));
 sg13g2_a21oi_1 _19688_ (.A1(_12620_),
    .A2(_12626_),
    .Y(_12631_),
    .B1(_12630_));
 sg13g2_nor2_1 _19689_ (.A(_12605_),
    .B(_12611_),
    .Y(_12632_));
 sg13g2_a22oi_1 _19690_ (.Y(_12633_),
    .B1(\u_inv.f_reg[62] ),
    .B2(\u_inv.f_next[62] ),
    .A2(\u_inv.f_reg[63] ),
    .A1(\u_inv.f_next[63] ));
 sg13g2_a21oi_1 _19691_ (.A1(_10518_),
    .A2(_10827_),
    .Y(_12634_),
    .B1(_12633_));
 sg13g2_a22oi_1 _19692_ (.Y(_12635_),
    .B1(\u_inv.f_reg[60] ),
    .B2(\u_inv.f_next[60] ),
    .A2(\u_inv.f_reg[61] ),
    .A1(\u_inv.f_next[61] ));
 sg13g2_a21o_1 _19693_ (.A2(_10829_),
    .A1(_10520_),
    .B1(_12635_),
    .X(_12636_));
 sg13g2_inv_1 _19694_ (.Y(_12637_),
    .A(_12636_));
 sg13g2_and3_1 _19695_ (.X(_12638_),
    .A(_11309_),
    .B(_11310_),
    .C(_12637_));
 sg13g2_nor4_1 _19696_ (.A(_12631_),
    .B(_12632_),
    .C(_12634_),
    .D(_12638_),
    .Y(_12639_));
 sg13g2_a22oi_1 _19697_ (.Y(_12640_),
    .B1(\u_inv.f_reg[40] ),
    .B2(\u_inv.f_next[40] ),
    .A2(\u_inv.f_reg[41] ),
    .A1(\u_inv.f_next[41] ));
 sg13g2_a21oi_1 _19698_ (.A1(_10540_),
    .A2(_10849_),
    .Y(_12641_),
    .B1(_12640_));
 sg13g2_nor2_1 _19699_ (.A(_11285_),
    .B(_11288_),
    .Y(_12642_));
 sg13g2_nor2_1 _19700_ (.A(_11281_),
    .B(_11282_),
    .Y(_12643_));
 sg13g2_nand2_1 _19701_ (.Y(_12644_),
    .A(_12642_),
    .B(_12643_));
 sg13g2_nand2_1 _19702_ (.Y(_12645_),
    .A(_11274_),
    .B(_11275_));
 sg13g2_inv_1 _19703_ (.Y(_12646_),
    .A(_12645_));
 sg13g2_a22oi_1 _19704_ (.Y(_12647_),
    .B1(\u_inv.f_reg[42] ),
    .B2(\u_inv.f_next[42] ),
    .A2(\u_inv.f_reg[43] ),
    .A1(\u_inv.f_next[43] ));
 sg13g2_a21oi_1 _19705_ (.A1(_10538_),
    .A2(_10847_),
    .Y(_12648_),
    .B1(_12647_));
 sg13g2_inv_1 _19706_ (.Y(_12649_),
    .A(_12648_));
 sg13g2_a21oi_1 _19707_ (.A1(_10534_),
    .A2(_10843_),
    .Y(_12650_),
    .B1(_11286_));
 sg13g2_a21oi_1 _19708_ (.A1(\u_inv.f_next[47] ),
    .A2(\u_inv.f_reg[47] ),
    .Y(_12651_),
    .B1(_12650_));
 sg13g2_a22oi_1 _19709_ (.Y(_12652_),
    .B1(\u_inv.f_reg[44] ),
    .B2(\u_inv.f_next[44] ),
    .A2(\u_inv.f_reg[45] ),
    .A1(\u_inv.f_next[45] ));
 sg13g2_a21oi_1 _19710_ (.A1(_10536_),
    .A2(_10845_),
    .Y(_12653_),
    .B1(_12652_));
 sg13g2_a21oi_1 _19711_ (.A1(_12641_),
    .A2(_12646_),
    .Y(_12654_),
    .B1(_12648_));
 sg13g2_o21ai_1 _19712_ (.B1(_12651_),
    .Y(_12655_),
    .A1(_12644_),
    .A2(_12654_));
 sg13g2_o21ai_1 _19713_ (.B1(_11238_),
    .Y(_12656_),
    .A1(_11234_),
    .A2(_11237_));
 sg13g2_nand2_1 _19714_ (.Y(_12657_),
    .A(_11242_),
    .B(_11243_));
 sg13g2_or3_1 _19715_ (.A(_11247_),
    .B(_11250_),
    .C(_12657_),
    .X(_12658_));
 sg13g2_and2_1 _19716_ (.A(_11231_),
    .B(_11232_),
    .X(_12659_));
 sg13g2_a22oi_1 _19717_ (.Y(_12660_),
    .B1(\u_inv.f_reg[34] ),
    .B2(\u_inv.f_next[34] ),
    .A2(\u_inv.f_reg[35] ),
    .A1(\u_inv.f_next[35] ));
 sg13g2_a21oi_1 _19718_ (.A1(_10546_),
    .A2(_10855_),
    .Y(_12661_),
    .B1(_12660_));
 sg13g2_a21oi_1 _19719_ (.A1(_11245_),
    .A2(_11248_),
    .Y(_12662_),
    .B1(_11246_));
 sg13g2_a22oi_1 _19720_ (.Y(_12663_),
    .B1(\u_inv.f_reg[36] ),
    .B2(\u_inv.f_next[36] ),
    .A2(\u_inv.f_reg[37] ),
    .A1(\u_inv.f_next[37] ));
 sg13g2_a21o_1 _19721_ (.A2(_10853_),
    .A1(_10544_),
    .B1(_12663_),
    .X(_12664_));
 sg13g2_nor3_1 _19722_ (.A(_11247_),
    .B(_11250_),
    .C(_12664_),
    .Y(_12665_));
 sg13g2_a21oi_1 _19723_ (.A1(_12656_),
    .A2(_12659_),
    .Y(_12666_),
    .B1(_12661_));
 sg13g2_o21ai_1 _19724_ (.B1(_12662_),
    .Y(_12667_),
    .A1(_12658_),
    .A2(_12666_));
 sg13g2_nor2_1 _19725_ (.A(_12665_),
    .B(_12667_),
    .Y(_12668_));
 sg13g2_o21ai_1 _19726_ (.B1(_11105_),
    .Y(_12669_),
    .A1(_11104_),
    .A2(_11152_));
 sg13g2_inv_1 _19727_ (.Y(_12670_),
    .A(_12669_));
 sg13g2_nand2_1 _19728_ (.Y(_12671_),
    .A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ));
 sg13g2_nor2_1 _19729_ (.A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ),
    .Y(_12672_));
 sg13g2_and2_1 _19730_ (.A(\u_inv.f_next[6] ),
    .B(\u_inv.f_reg[6] ),
    .X(_12673_));
 sg13g2_and2_1 _19731_ (.A(\u_inv.f_next[4] ),
    .B(\u_inv.f_reg[4] ),
    .X(_12674_));
 sg13g2_nand2_1 _19732_ (.Y(_12675_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_xnor2_1 _19733_ (.Y(_12676_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_nand2_1 _19734_ (.Y(_12677_),
    .A(net4639),
    .B(\u_inv.f_reg[0] ));
 sg13g2_o21ai_1 _19735_ (.B1(_12675_),
    .Y(_12678_),
    .A1(_12676_),
    .A2(_12677_));
 sg13g2_a21oi_1 _19736_ (.A1(_11132_),
    .A2(_12678_),
    .Y(_12679_),
    .B1(_11130_));
 sg13g2_o21ai_1 _19737_ (.B1(_11126_),
    .Y(_12680_),
    .A1(_11127_),
    .A2(_12679_));
 sg13g2_a21oi_1 _19738_ (.A1(_11124_),
    .A2(_12680_),
    .Y(_12681_),
    .B1(_12674_));
 sg13g2_o21ai_1 _19739_ (.B1(_11121_),
    .Y(_12682_),
    .A1(_11122_),
    .A2(_12681_));
 sg13g2_a21oi_1 _19740_ (.A1(_11119_),
    .A2(_12682_),
    .Y(_12683_),
    .B1(_12673_));
 sg13g2_o21ai_1 _19741_ (.B1(_11116_),
    .Y(_12684_),
    .A1(_11117_),
    .A2(_12683_));
 sg13g2_a21oi_1 _19742_ (.A1(_11114_),
    .A2(_12684_),
    .Y(_12685_),
    .B1(_11113_));
 sg13g2_a221oi_1 _19743_ (.B2(_12684_),
    .C1(_11113_),
    .B1(_11114_),
    .A1(\u_inv.f_next[9] ),
    .Y(_12686_),
    .A2(\u_inv.f_reg[9] ));
 sg13g2_or3_1 _19744_ (.A(_11109_),
    .B(_11111_),
    .C(_12686_),
    .X(_12687_));
 sg13g2_nand2_1 _19745_ (.Y(_12688_),
    .A(_11107_),
    .B(_12687_));
 sg13g2_o21ai_1 _19746_ (.B1(_12671_),
    .Y(_12689_),
    .A1(_11107_),
    .A2(_12672_));
 sg13g2_xnor2_1 _19747_ (.Y(_12690_),
    .A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ));
 sg13g2_nor4_1 _19748_ (.A(_11109_),
    .B(_11111_),
    .C(_12686_),
    .D(_12690_),
    .Y(_12691_));
 sg13g2_nor2_1 _19749_ (.A(_12689_),
    .B(_12691_),
    .Y(_12692_));
 sg13g2_nand2b_1 _19750_ (.Y(_12693_),
    .B(_11153_),
    .A_N(_11106_));
 sg13g2_o21ai_1 _19751_ (.B1(_12670_),
    .Y(_12694_),
    .A1(_12692_),
    .A2(_12693_));
 sg13g2_nand3b_1 _19752_ (.B(_11102_),
    .C(_12669_),
    .Y(_12695_),
    .A_N(_11100_));
 sg13g2_nor3_1 _19753_ (.A(_11100_),
    .B(_11103_),
    .C(_12693_),
    .Y(_12696_));
 sg13g2_o21ai_1 _19754_ (.B1(_12696_),
    .Y(_12697_),
    .A1(_12689_),
    .A2(_12691_));
 sg13g2_o21ai_1 _19755_ (.B1(_11101_),
    .Y(_12698_),
    .A1(\u_inv.f_next[15] ),
    .A2(\u_inv.f_reg[15] ));
 sg13g2_nand4_1 _19756_ (.B(_12695_),
    .C(_12697_),
    .A(_11099_),
    .Y(_12699_),
    .D(_12698_));
 sg13g2_nand2_1 _19757_ (.Y(_12700_),
    .A(_11094_),
    .B(_11168_));
 sg13g2_nor2b_1 _19758_ (.A(_12700_),
    .B_N(_12699_),
    .Y(_12701_));
 sg13g2_o21ai_1 _19759_ (.B1(_11096_),
    .Y(_12702_),
    .A1(_11091_),
    .A2(_11095_));
 sg13g2_a21oi_1 _19760_ (.A1(\u_inv.f_next[17] ),
    .A2(\u_inv.f_reg[17] ),
    .Y(_12703_),
    .B1(_11167_));
 sg13g2_a21oi_1 _19761_ (.A1(_10564_),
    .A2(_10872_),
    .Y(_12704_),
    .B1(_12703_));
 sg13g2_nor2_1 _19762_ (.A(_11093_),
    .B(_11098_),
    .Y(_12705_));
 sg13g2_nor3_1 _19763_ (.A(_11093_),
    .B(_11098_),
    .C(_12700_),
    .Y(_12706_));
 sg13g2_a221oi_1 _19764_ (.B2(_12699_),
    .C1(_12702_),
    .B1(_12706_),
    .A1(_12704_),
    .Y(_12707_),
    .A2(_12705_));
 sg13g2_and2_1 _19765_ (.A(_11186_),
    .B(_11188_),
    .X(_12708_));
 sg13g2_nor2_1 _19766_ (.A(_11183_),
    .B(_11187_),
    .Y(_12709_));
 sg13g2_nand2_1 _19767_ (.Y(_12710_),
    .A(_12708_),
    .B(_12709_));
 sg13g2_a21oi_1 _19768_ (.A1(_10558_),
    .A2(_10866_),
    .Y(_12711_),
    .B1(_11185_));
 sg13g2_a22oi_1 _19769_ (.Y(_12712_),
    .B1(\u_inv.f_reg[20] ),
    .B2(\u_inv.f_next[20] ),
    .A2(\u_inv.f_reg[21] ),
    .A1(\u_inv.f_next[21] ));
 sg13g2_a21oi_1 _19770_ (.A1(_10560_),
    .A2(_10868_),
    .Y(_12713_),
    .B1(_12712_));
 sg13g2_a221oi_1 _19771_ (.B2(_12713_),
    .C1(_12711_),
    .B1(_12708_),
    .A1(\u_inv.f_next[23] ),
    .Y(_12714_),
    .A2(\u_inv.f_reg[23] ));
 sg13g2_o21ai_1 _19772_ (.B1(_12714_),
    .Y(_12715_),
    .A1(_12707_),
    .A2(_12710_));
 sg13g2_nand2_1 _19773_ (.Y(_12716_),
    .A(_11079_),
    .B(_11082_));
 sg13g2_nand2_1 _19774_ (.Y(_12717_),
    .A(_11085_),
    .B(_11088_));
 sg13g2_nor2_1 _19775_ (.A(_12716_),
    .B(_12717_),
    .Y(_12718_));
 sg13g2_nor2b_1 _19776_ (.A(_11206_),
    .B_N(_11208_),
    .Y(_12719_));
 sg13g2_nand2_1 _19777_ (.Y(_12720_),
    .A(_12718_),
    .B(_12719_));
 sg13g2_nor3_1 _19778_ (.A(_11201_),
    .B(_11204_),
    .C(_12720_),
    .Y(_12721_));
 sg13g2_a22oi_1 _19779_ (.Y(_12722_),
    .B1(\u_inv.f_reg[24] ),
    .B2(\u_inv.f_next[24] ),
    .A2(\u_inv.f_reg[25] ),
    .A1(\u_inv.f_next[25] ));
 sg13g2_a21o_1 _19780_ (.A2(_10864_),
    .A1(_10556_),
    .B1(_12722_),
    .X(_12723_));
 sg13g2_a21oi_1 _19781_ (.A1(\u_inv.f_next[27] ),
    .A2(\u_inv.f_reg[27] ),
    .Y(_12724_),
    .B1(_11205_));
 sg13g2_a21oi_1 _19782_ (.A1(_10554_),
    .A2(_10862_),
    .Y(_12725_),
    .B1(_12724_));
 sg13g2_a21oi_1 _19783_ (.A1(_10550_),
    .A2(_10858_),
    .Y(_12726_),
    .B1(_11081_));
 sg13g2_a21oi_1 _19784_ (.A1(\u_inv.f_next[31] ),
    .A2(\u_inv.f_reg[31] ),
    .Y(_12727_),
    .B1(_12726_));
 sg13g2_a22oi_1 _19785_ (.Y(_12728_),
    .B1(\u_inv.f_reg[28] ),
    .B2(\u_inv.f_next[28] ),
    .A2(\u_inv.f_reg[29] ),
    .A1(\u_inv.f_next[29] ));
 sg13g2_a21o_1 _19786_ (.A2(_10860_),
    .A1(_10552_),
    .B1(_12728_),
    .X(_12729_));
 sg13g2_o21ai_1 _19787_ (.B1(_12727_),
    .Y(_12730_),
    .A1(_12716_),
    .A2(_12729_));
 sg13g2_a21oi_1 _19788_ (.A1(_12718_),
    .A2(_12725_),
    .Y(_12731_),
    .B1(_12730_));
 sg13g2_o21ai_1 _19789_ (.B1(_12731_),
    .Y(_12732_),
    .A1(_12720_),
    .A2(_12723_));
 sg13g2_a21oi_2 _19790_ (.B1(_12732_),
    .Y(_12733_),
    .A2(_12721_),
    .A1(_12715_));
 sg13g2_nor2_1 _19791_ (.A(_11235_),
    .B(_11240_),
    .Y(_12734_));
 sg13g2_nand3b_1 _19792_ (.B(_12659_),
    .C(_12734_),
    .Y(_12735_),
    .A_N(_12658_));
 sg13g2_o21ai_1 _19793_ (.B1(_12668_),
    .Y(_12736_),
    .A1(_12733_),
    .A2(_12735_));
 sg13g2_nor4_1 _19794_ (.A(_11277_),
    .B(_11278_),
    .C(_12644_),
    .D(_12645_),
    .Y(_12737_));
 sg13g2_a221oi_1 _19795_ (.B2(_12737_),
    .C1(_12655_),
    .B1(_12736_),
    .A1(_12642_),
    .Y(_12738_),
    .A2(_12653_));
 sg13g2_nor2_1 _19796_ (.A(_11323_),
    .B(_11333_),
    .Y(_12739_));
 sg13g2_nand4_1 _19797_ (.B(_12615_),
    .C(_12629_),
    .A(_12614_),
    .Y(_12740_),
    .D(_12739_));
 sg13g2_o21ai_1 _19798_ (.B1(_12639_),
    .Y(_12741_),
    .A1(_12738_),
    .A2(_12740_));
 sg13g2_nand2_1 _19799_ (.Y(_12742_),
    .A(_11390_),
    .B(_12573_));
 sg13g2_nor2_1 _19800_ (.A(_12572_),
    .B(_12742_),
    .Y(_12743_));
 sg13g2_and3_2 _19801_ (.X(_12744_),
    .A(_11392_),
    .B(_12601_),
    .C(_12743_));
 sg13g2_a21oi_2 _19802_ (.B1(_12603_),
    .Y(_12745_),
    .A2(_12744_),
    .A1(_12741_));
 sg13g2_a21o_2 _19803_ (.A2(_12744_),
    .A1(_12741_),
    .B1(_12603_),
    .X(_12746_));
 sg13g2_nand2_1 _19804_ (.Y(_12747_),
    .A(_11569_),
    .B(_12467_));
 sg13g2_or2_1 _19805_ (.X(_12748_),
    .B(_12747_),
    .A(_12466_));
 sg13g2_nor4_2 _19806_ (.A(_11567_),
    .B(_12491_),
    .C(_12499_),
    .Y(_12749_),
    .D(_12748_));
 sg13g2_a21oi_2 _19807_ (.B1(_12534_),
    .Y(_12750_),
    .A2(_12749_),
    .A1(_12746_));
 sg13g2_a21o_1 _19808_ (.A2(_12749_),
    .A1(_12746_),
    .B1(_12534_),
    .X(_12751_));
 sg13g2_or4_1 _19809_ (.A(_11720_),
    .B(_11722_),
    .C(_11724_),
    .D(_11725_),
    .X(_12752_));
 sg13g2_nor4_2 _19810_ (.A(_12405_),
    .B(_12421_),
    .C(_12454_),
    .Y(_12753_),
    .D(_12752_));
 sg13g2_nand2_1 _19811_ (.Y(_12754_),
    .A(_12461_),
    .B(_12753_));
 sg13g2_o21ai_1 _19812_ (.B1(_12463_),
    .Y(_12755_),
    .A1(_12750_),
    .A2(_12754_));
 sg13g2_and2_1 _19813_ (.A(_11999_),
    .B(_12001_),
    .X(_12756_));
 sg13g2_nand2_1 _19814_ (.Y(_12757_),
    .A(_12256_),
    .B(_12756_));
 sg13g2_nor2_2 _19815_ (.A(_12257_),
    .B(_12757_),
    .Y(_12758_));
 sg13g2_and2_1 _19816_ (.A(_12274_),
    .B(_12758_),
    .X(_12759_));
 sg13g2_nor2b_1 _19817_ (.A(_12253_),
    .B_N(_12759_),
    .Y(_12760_));
 sg13g2_a21oi_2 _19818_ (.B1(_12311_),
    .Y(_12761_),
    .A2(_12760_),
    .A1(_12755_));
 sg13g2_and2_1 _19819_ (.A(_12089_),
    .B(_12091_),
    .X(_12762_));
 sg13g2_nor2_1 _19820_ (.A(_12094_),
    .B(_12096_),
    .Y(_12763_));
 sg13g2_nand2_1 _19821_ (.Y(_12764_),
    .A(_12762_),
    .B(_12763_));
 sg13g2_nand2_1 _19822_ (.Y(_12765_),
    .A(_12114_),
    .B(_12117_));
 sg13g2_nor2_1 _19823_ (.A(_12110_),
    .B(_12112_),
    .Y(_12766_));
 sg13g2_nor2b_1 _19824_ (.A(_12765_),
    .B_N(_12766_),
    .Y(_12767_));
 sg13g2_nor2_1 _19825_ (.A(_12098_),
    .B(_12100_),
    .Y(_12768_));
 sg13g2_nor2_1 _19826_ (.A(_12103_),
    .B(_12105_),
    .Y(_12769_));
 sg13g2_and2_1 _19827_ (.A(_12768_),
    .B(_12769_),
    .X(_12770_));
 sg13g2_inv_1 _19828_ (.Y(_12771_),
    .A(_12770_));
 sg13g2_nand2_1 _19829_ (.Y(_12772_),
    .A(_12767_),
    .B(_12770_));
 sg13g2_nor2_1 _19830_ (.A(_12082_),
    .B(_12084_),
    .Y(_12773_));
 sg13g2_nand3_1 _19831_ (.B(_12087_),
    .C(_12773_),
    .A(_12085_),
    .Y(_12774_));
 sg13g2_or3_1 _19832_ (.A(_12764_),
    .B(_12772_),
    .C(_12774_),
    .X(_12775_));
 sg13g2_a22oi_1 _19833_ (.Y(_12776_),
    .B1(\u_inv.f_reg[224] ),
    .B2(\u_inv.f_next[224] ),
    .A2(\u_inv.f_reg[225] ),
    .A1(\u_inv.f_next[225] ));
 sg13g2_a21oi_1 _19834_ (.A1(_10356_),
    .A2(_10665_),
    .Y(_12777_),
    .B1(_12776_));
 sg13g2_a21oi_1 _19835_ (.A1(_10354_),
    .A2(_10663_),
    .Y(_12778_),
    .B1(_12080_));
 sg13g2_a221oi_1 _19836_ (.B2(_12777_),
    .C1(_12778_),
    .B1(_12773_),
    .A1(\u_inv.f_next[227] ),
    .Y(_12779_),
    .A2(\u_inv.f_reg[227] ));
 sg13g2_nor3_1 _19837_ (.A(_12764_),
    .B(_12772_),
    .C(_12779_),
    .Y(_12780_));
 sg13g2_a22oi_1 _19838_ (.Y(_12781_),
    .B1(\u_inv.f_reg[232] ),
    .B2(\u_inv.f_next[232] ),
    .A2(\u_inv.f_reg[233] ),
    .A1(\u_inv.f_next[233] ));
 sg13g2_a21oi_1 _19839_ (.A1(_10348_),
    .A2(_10657_),
    .Y(_12782_),
    .B1(_12781_));
 sg13g2_a21oi_1 _19840_ (.A1(_10346_),
    .A2(_10655_),
    .Y(_12783_),
    .B1(_12099_));
 sg13g2_a221oi_1 _19841_ (.B2(_12782_),
    .C1(_12783_),
    .B1(_12768_),
    .A1(\u_inv.f_next[235] ),
    .Y(_12784_),
    .A2(\u_inv.f_reg[235] ));
 sg13g2_nand2b_1 _19842_ (.Y(_12785_),
    .B(_12767_),
    .A_N(_12784_));
 sg13g2_a22oi_1 _19843_ (.Y(_12786_),
    .B1(\u_inv.f_reg[228] ),
    .B2(\u_inv.f_next[228] ),
    .A2(\u_inv.f_reg[229] ),
    .A1(\u_inv.f_next[229] ));
 sg13g2_a21oi_1 _19844_ (.A1(_10352_),
    .A2(_10661_),
    .Y(_12787_),
    .B1(_12786_));
 sg13g2_a21oi_1 _19845_ (.A1(_10350_),
    .A2(_10659_),
    .Y(_12788_),
    .B1(_12090_));
 sg13g2_a221oi_1 _19846_ (.B2(_12787_),
    .C1(_12788_),
    .B1(_12762_),
    .A1(\u_inv.f_next[231] ),
    .Y(_12789_),
    .A2(\u_inv.f_reg[231] ));
 sg13g2_nor2_1 _19847_ (.A(_12772_),
    .B(_12789_),
    .Y(_12790_));
 sg13g2_a21oi_1 _19848_ (.A1(\u_inv.f_next[237] ),
    .A2(\u_inv.f_reg[237] ),
    .Y(_12791_),
    .B1(_12109_));
 sg13g2_a21oi_1 _19849_ (.A1(_10344_),
    .A2(_10653_),
    .Y(_12792_),
    .B1(_12791_));
 sg13g2_nor2b_1 _19850_ (.A(_12765_),
    .B_N(_12792_),
    .Y(_12793_));
 sg13g2_a21oi_1 _19851_ (.A1(_10342_),
    .A2(_10651_),
    .Y(_12794_),
    .B1(_12115_));
 sg13g2_a21oi_1 _19852_ (.A1(\u_inv.f_next[239] ),
    .A2(\u_inv.f_reg[239] ),
    .Y(_12795_),
    .B1(_12794_));
 sg13g2_nand2_1 _19853_ (.Y(_12796_),
    .A(_12785_),
    .B(_12795_));
 sg13g2_nor4_1 _19854_ (.A(_12780_),
    .B(_12790_),
    .C(_12793_),
    .D(_12796_),
    .Y(_12797_));
 sg13g2_o21ai_1 _19855_ (.B1(_12797_),
    .Y(_12798_),
    .A1(_12761_),
    .A2(_12775_));
 sg13g2_nor4_1 _19856_ (.A(_12158_),
    .B(_12160_),
    .C(_12228_),
    .D(_12229_),
    .Y(_12799_));
 sg13g2_a21oi_2 _19857_ (.B1(_12240_),
    .Y(_12800_),
    .A2(_12799_),
    .A1(_12798_));
 sg13g2_nor2_1 _19858_ (.A(_12189_),
    .B(_12193_),
    .Y(_12801_));
 sg13g2_nor2_1 _19859_ (.A(_12188_),
    .B(_12191_),
    .Y(_12802_));
 sg13g2_nand2_1 _19860_ (.Y(_12803_),
    .A(_12801_),
    .B(_12802_));
 sg13g2_a21oi_1 _19861_ (.A1(_10330_),
    .A2(_10639_),
    .Y(_12804_),
    .B1(_12192_));
 sg13g2_a22oi_1 _19862_ (.Y(_12805_),
    .B1(\u_inv.f_reg[248] ),
    .B2(\u_inv.f_next[248] ),
    .A2(\u_inv.f_reg[249] ),
    .A1(\u_inv.f_next[249] ));
 sg13g2_a21oi_1 _19863_ (.A1(_10332_),
    .A2(_10641_),
    .Y(_12806_),
    .B1(_12805_));
 sg13g2_a221oi_1 _19864_ (.B2(_12806_),
    .C1(_12804_),
    .B1(_12801_),
    .A1(\u_inv.f_next[251] ),
    .Y(_12807_),
    .A2(\u_inv.f_reg[251] ));
 sg13g2_o21ai_1 _19865_ (.B1(_12807_),
    .Y(_12808_),
    .A1(_12800_),
    .A2(_12803_));
 sg13g2_nor2_1 _19866_ (.A(_12203_),
    .B(_12206_),
    .Y(_12809_));
 sg13g2_a21oi_1 _19867_ (.A1(_10328_),
    .A2(_10637_),
    .Y(_12810_),
    .B1(_12204_));
 sg13g2_a221oi_1 _19868_ (.B2(_12809_),
    .C1(_12810_),
    .B1(_12808_),
    .A1(\u_inv.f_next[253] ),
    .Y(_12811_),
    .A2(\u_inv.f_reg[253] ));
 sg13g2_a22oi_1 _19869_ (.Y(_12812_),
    .B1(\u_inv.f_reg[254] ),
    .B2(\u_inv.f_next[254] ),
    .A2(\u_inv.f_reg[255] ),
    .A1(\u_inv.f_next[255] ));
 sg13g2_o21ai_1 _19870_ (.B1(_12812_),
    .Y(_12813_),
    .A1(_11077_),
    .A2(_12811_));
 sg13g2_a21oi_1 _19871_ (.A1(_11071_),
    .A2(_12813_),
    .Y(_12814_),
    .B1(_11070_));
 sg13g2_a21oi_1 _19872_ (.A1(net4959),
    .A2(net4725),
    .Y(_12815_),
    .B1(_12814_));
 sg13g2_o21ai_1 _19873_ (.B1(_12224_),
    .Y(_12816_),
    .A1(net3722),
    .A2(_12815_));
 sg13g2_nor2_2 _19874_ (.A(net4444),
    .B(net3950),
    .Y(_12817_));
 sg13g2_nand2_1 _19875_ (.Y(_12818_),
    .A(net4838),
    .B(net4378));
 sg13g2_nor2_1 _19876_ (.A(net4526),
    .B(net4232),
    .Y(_12819_));
 sg13g2_a21o_1 _19877_ (.A2(_12819_),
    .A1(_12816_),
    .B1(_11069_),
    .X(_00010_));
 sg13g2_nand2_1 _19878_ (.Y(_12820_),
    .A(_10626_),
    .B(net10));
 sg13g2_o21ai_1 _19879_ (.B1(\state[1] ),
    .Y(_12821_),
    .A1(rd_prev),
    .A2(_12820_));
 sg13g2_a21oi_2 _19880_ (.B1(_11050_),
    .Y(_12822_),
    .A2(_12821_),
    .A1(_11053_));
 sg13g2_a221oi_1 _19881_ (.B2(net1),
    .C1(net4058),
    .B1(net4241),
    .A1(net1427),
    .Y(_12823_),
    .A2(net4389));
 sg13g2_a21oi_1 _19882_ (.A1(_10988_),
    .A2(net4058),
    .Y(_00011_),
    .B1(_12823_));
 sg13g2_a221oi_1 _19883_ (.B2(net2),
    .C1(net4057),
    .B1(net4241),
    .A1(\inv_result[1] ),
    .Y(_12824_),
    .A2(net4390));
 sg13g2_a21oi_1 _19884_ (.A1(_10989_),
    .A2(net4058),
    .Y(_00012_),
    .B1(_12824_));
 sg13g2_a221oi_1 _19885_ (.B2(net3),
    .C1(net4057),
    .B1(net4241),
    .A1(net1172),
    .Y(_12825_),
    .A2(net4390));
 sg13g2_a21oi_1 _19886_ (.A1(_10990_),
    .A2(net4058),
    .Y(_00013_),
    .B1(_12825_));
 sg13g2_a221oi_1 _19887_ (.B2(net4),
    .C1(net4056),
    .B1(net4241),
    .A1(\inv_result[3] ),
    .Y(_12826_),
    .A2(net4390));
 sg13g2_a21oi_1 _19888_ (.A1(_10991_),
    .A2(net4060),
    .Y(_00014_),
    .B1(_12826_));
 sg13g2_a221oi_1 _19889_ (.B2(net5),
    .C1(net4060),
    .B1(net4241),
    .A1(\inv_result[4] ),
    .Y(_12827_),
    .A2(net4391));
 sg13g2_a21oi_1 _19890_ (.A1(_10992_),
    .A2(net4060),
    .Y(_00015_),
    .B1(_12827_));
 sg13g2_a221oi_1 _19891_ (.B2(net6),
    .C1(net4061),
    .B1(net4241),
    .A1(\inv_result[5] ),
    .Y(_12828_),
    .A2(net4391));
 sg13g2_a21oi_1 _19892_ (.A1(_10993_),
    .A2(net4061),
    .Y(_00016_),
    .B1(_12828_));
 sg13g2_a221oi_1 _19893_ (.B2(net7),
    .C1(net4060),
    .B1(net4241),
    .A1(net1426),
    .Y(_12829_),
    .A2(net4389));
 sg13g2_a21oi_1 _19894_ (.A1(_10994_),
    .A2(net4060),
    .Y(_00017_),
    .B1(_12829_));
 sg13g2_a221oi_1 _19895_ (.B2(net8),
    .C1(net4060),
    .B1(net4241),
    .A1(net1117),
    .Y(_12830_),
    .A2(net4391));
 sg13g2_a21oi_1 _19896_ (.A1(_10995_),
    .A2(net4061),
    .Y(_00018_),
    .B1(_12830_));
 sg13g2_nor2_1 _19897_ (.A(_10988_),
    .B(net4389),
    .Y(_12831_));
 sg13g2_a21oi_1 _19898_ (.A1(\inv_result[8] ),
    .A2(net4389),
    .Y(_12832_),
    .B1(_12831_));
 sg13g2_nand2_1 _19899_ (.Y(_12833_),
    .A(net1446),
    .B(net4058));
 sg13g2_o21ai_1 _19900_ (.B1(_12833_),
    .Y(_00019_),
    .A1(net4058),
    .A2(_12832_));
 sg13g2_nor2_1 _19901_ (.A(_10989_),
    .B(net4389),
    .Y(_12834_));
 sg13g2_a21oi_1 _19902_ (.A1(net1206),
    .A2(net4389),
    .Y(_12835_),
    .B1(_12834_));
 sg13g2_nand2_1 _19903_ (.Y(_12836_),
    .A(net1249),
    .B(net4059));
 sg13g2_o21ai_1 _19904_ (.B1(_12836_),
    .Y(_00020_),
    .A1(net4059),
    .A2(_12835_));
 sg13g2_nor2_1 _19905_ (.A(_10990_),
    .B(net4390),
    .Y(_12837_));
 sg13g2_a21oi_1 _19906_ (.A1(\inv_result[10] ),
    .A2(net4389),
    .Y(_12838_),
    .B1(_12837_));
 sg13g2_nand2_1 _19907_ (.Y(_12839_),
    .A(net1593),
    .B(net4058));
 sg13g2_o21ai_1 _19908_ (.B1(_12839_),
    .Y(_00021_),
    .A1(net4058),
    .A2(_12838_));
 sg13g2_nor2_1 _19909_ (.A(_10991_),
    .B(net4390),
    .Y(_12840_));
 sg13g2_a21oi_1 _19910_ (.A1(\inv_result[11] ),
    .A2(net4389),
    .Y(_12841_),
    .B1(_12840_));
 sg13g2_nand2_1 _19911_ (.Y(_12842_),
    .A(net1241),
    .B(net4060));
 sg13g2_o21ai_1 _19912_ (.B1(_12842_),
    .Y(_00022_),
    .A1(net4060),
    .A2(_12841_));
 sg13g2_nor2_1 _19913_ (.A(_10992_),
    .B(net4391),
    .Y(_12843_));
 sg13g2_a21oi_1 _19914_ (.A1(\inv_result[12] ),
    .A2(net4392),
    .Y(_12844_),
    .B1(_12843_));
 sg13g2_nand2_1 _19915_ (.Y(_12845_),
    .A(net1212),
    .B(net4071));
 sg13g2_o21ai_1 _19916_ (.B1(_12845_),
    .Y(_00023_),
    .A1(net4062),
    .A2(_12844_));
 sg13g2_nor2_1 _19917_ (.A(_10993_),
    .B(net4393),
    .Y(_12846_));
 sg13g2_a21oi_1 _19918_ (.A1(\inv_result[13] ),
    .A2(net4393),
    .Y(_12847_),
    .B1(_12846_));
 sg13g2_nand2_1 _19919_ (.Y(_12848_),
    .A(net1143),
    .B(net4071));
 sg13g2_o21ai_1 _19920_ (.B1(_12848_),
    .Y(_00024_),
    .A1(net4071),
    .A2(_12847_));
 sg13g2_nor2_1 _19921_ (.A(_10994_),
    .B(net4392),
    .Y(_12849_));
 sg13g2_a21oi_1 _19922_ (.A1(net1734),
    .A2(net4392),
    .Y(_12850_),
    .B1(_12849_));
 sg13g2_nand2_1 _19923_ (.Y(_12851_),
    .A(net1880),
    .B(net4062));
 sg13g2_o21ai_1 _19924_ (.B1(_12851_),
    .Y(_00025_),
    .A1(net4062),
    .A2(_12850_));
 sg13g2_nor2_1 _19925_ (.A(_10995_),
    .B(net4392),
    .Y(_12852_));
 sg13g2_a21oi_1 _19926_ (.A1(net1560),
    .A2(net4393),
    .Y(_12853_),
    .B1(_12852_));
 sg13g2_nand2_1 _19927_ (.Y(_12854_),
    .A(net2310),
    .B(net4071));
 sg13g2_o21ai_1 _19928_ (.B1(_12854_),
    .Y(_00026_),
    .A1(net4062),
    .A2(_12853_));
 sg13g2_and2_1 _19929_ (.A(net1446),
    .B(net4453),
    .X(_12855_));
 sg13g2_a21oi_1 _19930_ (.A1(net1453),
    .A2(net4392),
    .Y(_12856_),
    .B1(_12855_));
 sg13g2_nand2_1 _19931_ (.Y(_12857_),
    .A(net2283),
    .B(net4059));
 sg13g2_o21ai_1 _19932_ (.B1(_12857_),
    .Y(_00027_),
    .A1(net4059),
    .A2(_12856_));
 sg13g2_and2_1 _19933_ (.A(net1249),
    .B(net4453),
    .X(_12858_));
 sg13g2_a21oi_1 _19934_ (.A1(\inv_result[17] ),
    .A2(net4392),
    .Y(_12859_),
    .B1(_12858_));
 sg13g2_nand2_1 _19935_ (.Y(_12860_),
    .A(net2038),
    .B(net4059));
 sg13g2_o21ai_1 _19936_ (.B1(_12860_),
    .Y(_00028_),
    .A1(net4059),
    .A2(_12859_));
 sg13g2_and2_1 _19937_ (.A(net1593),
    .B(net4453),
    .X(_12861_));
 sg13g2_a21oi_1 _19938_ (.A1(net1647),
    .A2(net4392),
    .Y(_12862_),
    .B1(_12861_));
 sg13g2_nand2_1 _19939_ (.Y(_12863_),
    .A(net2138),
    .B(net4071));
 sg13g2_o21ai_1 _19940_ (.B1(_12863_),
    .Y(_00029_),
    .A1(net4059),
    .A2(_12862_));
 sg13g2_and2_1 _19941_ (.A(net1241),
    .B(net4454),
    .X(_12864_));
 sg13g2_a21oi_1 _19942_ (.A1(net1668),
    .A2(net4392),
    .Y(_12865_),
    .B1(_12864_));
 sg13g2_nand2_1 _19943_ (.Y(_12866_),
    .A(net1871),
    .B(net4071));
 sg13g2_o21ai_1 _19944_ (.B1(_12866_),
    .Y(_00030_),
    .A1(net4071),
    .A2(_12865_));
 sg13g2_and2_1 _19945_ (.A(net1212),
    .B(net4453),
    .X(_12867_));
 sg13g2_a21oi_1 _19946_ (.A1(net1342),
    .A2(net4395),
    .Y(_12868_),
    .B1(_12867_));
 sg13g2_nand2_1 _19947_ (.Y(_12869_),
    .A(net1419),
    .B(net4068));
 sg13g2_o21ai_1 _19948_ (.B1(_12869_),
    .Y(_00031_),
    .A1(net4068),
    .A2(_12868_));
 sg13g2_and2_1 _19949_ (.A(net1143),
    .B(net4453),
    .X(_12870_));
 sg13g2_a21oi_1 _19950_ (.A1(\inv_result[21] ),
    .A2(net4395),
    .Y(_12871_),
    .B1(_12870_));
 sg13g2_nand2_1 _19951_ (.Y(_12872_),
    .A(net1251),
    .B(net4068));
 sg13g2_o21ai_1 _19952_ (.B1(_12872_),
    .Y(_00032_),
    .A1(net4068),
    .A2(_12871_));
 sg13g2_and2_1 _19953_ (.A(\shift_reg[14] ),
    .B(net4460),
    .X(_12873_));
 sg13g2_a21oi_1 _19954_ (.A1(\inv_result[22] ),
    .A2(net4395),
    .Y(_12874_),
    .B1(_12873_));
 sg13g2_nand2_1 _19955_ (.Y(_12875_),
    .A(net1359),
    .B(net4068));
 sg13g2_o21ai_1 _19956_ (.B1(_12875_),
    .Y(_00033_),
    .A1(net4070),
    .A2(_12874_));
 sg13g2_and2_1 _19957_ (.A(\shift_reg[15] ),
    .B(net4460),
    .X(_12876_));
 sg13g2_a21oi_1 _19958_ (.A1(net1321),
    .A2(net4395),
    .Y(_12877_),
    .B1(_12876_));
 sg13g2_nand2_1 _19959_ (.Y(_12878_),
    .A(net1487),
    .B(net4068));
 sg13g2_o21ai_1 _19960_ (.B1(_12878_),
    .Y(_00034_),
    .A1(net4069),
    .A2(_12877_));
 sg13g2_and2_1 _19961_ (.A(\shift_reg[16] ),
    .B(net4458),
    .X(_12879_));
 sg13g2_a21oi_1 _19962_ (.A1(\inv_result[24] ),
    .A2(net4396),
    .Y(_12880_),
    .B1(_12879_));
 sg13g2_nand2_1 _19963_ (.Y(_12881_),
    .A(net1633),
    .B(net4070));
 sg13g2_o21ai_1 _19964_ (.B1(_12881_),
    .Y(_00035_),
    .A1(net4070),
    .A2(_12880_));
 sg13g2_and2_1 _19965_ (.A(\shift_reg[17] ),
    .B(net4460),
    .X(_12882_));
 sg13g2_a21oi_1 _19966_ (.A1(\inv_result[25] ),
    .A2(net4395),
    .Y(_12883_),
    .B1(_12882_));
 sg13g2_nand2_1 _19967_ (.Y(_12884_),
    .A(net1230),
    .B(net4068));
 sg13g2_o21ai_1 _19968_ (.B1(_12884_),
    .Y(_00036_),
    .A1(net4068),
    .A2(_12883_));
 sg13g2_and2_1 _19969_ (.A(\shift_reg[18] ),
    .B(net4458),
    .X(_12885_));
 sg13g2_a21oi_1 _19970_ (.A1(\inv_result[26] ),
    .A2(net4396),
    .Y(_12886_),
    .B1(_12885_));
 sg13g2_nand2_1 _19971_ (.Y(_12887_),
    .A(net1210),
    .B(net4070));
 sg13g2_o21ai_1 _19972_ (.B1(_12887_),
    .Y(_00037_),
    .A1(net4070),
    .A2(_12886_));
 sg13g2_and2_1 _19973_ (.A(\shift_reg[19] ),
    .B(net4459),
    .X(_12888_));
 sg13g2_a21oi_1 _19974_ (.A1(\inv_result[27] ),
    .A2(net4395),
    .Y(_12889_),
    .B1(_12888_));
 sg13g2_nand2_1 _19975_ (.Y(_12890_),
    .A(net1584),
    .B(net4069));
 sg13g2_o21ai_1 _19976_ (.B1(_12890_),
    .Y(_00038_),
    .A1(net4069),
    .A2(_12889_));
 sg13g2_and2_1 _19977_ (.A(\shift_reg[20] ),
    .B(net4459),
    .X(_12891_));
 sg13g2_a21oi_1 _19978_ (.A1(\inv_result[28] ),
    .A2(net4396),
    .Y(_12892_),
    .B1(_12891_));
 sg13g2_nand2_1 _19979_ (.Y(_12893_),
    .A(net1160),
    .B(net4069));
 sg13g2_o21ai_1 _19980_ (.B1(_12893_),
    .Y(_00039_),
    .A1(net4069),
    .A2(_12892_));
 sg13g2_and2_1 _19981_ (.A(net1251),
    .B(net4459),
    .X(_12894_));
 sg13g2_a21oi_1 _19982_ (.A1(\inv_result[29] ),
    .A2(net4396),
    .Y(_12895_),
    .B1(_12894_));
 sg13g2_nand2_1 _19983_ (.Y(_12896_),
    .A(net1461),
    .B(net4069));
 sg13g2_o21ai_1 _19984_ (.B1(_12896_),
    .Y(_00040_),
    .A1(net4070),
    .A2(_12895_));
 sg13g2_and2_1 _19985_ (.A(\shift_reg[22] ),
    .B(net4458),
    .X(_12897_));
 sg13g2_a21oi_1 _19986_ (.A1(\inv_result[30] ),
    .A2(net4395),
    .Y(_12898_),
    .B1(_12897_));
 sg13g2_nand2_1 _19987_ (.Y(_12899_),
    .A(net1155),
    .B(net4078));
 sg13g2_o21ai_1 _19988_ (.B1(_12899_),
    .Y(_00041_),
    .A1(net4070),
    .A2(_12898_));
 sg13g2_and2_1 _19989_ (.A(\shift_reg[23] ),
    .B(net4458),
    .X(_12900_));
 sg13g2_a21oi_1 _19990_ (.A1(\inv_result[31] ),
    .A2(net4395),
    .Y(_12901_),
    .B1(_12900_));
 sg13g2_nand2_1 _19991_ (.Y(_12902_),
    .A(net1148),
    .B(net4077));
 sg13g2_o21ai_1 _19992_ (.B1(_12902_),
    .Y(_00042_),
    .A1(net4069),
    .A2(_12901_));
 sg13g2_and2_1 _19993_ (.A(\shift_reg[24] ),
    .B(net4463),
    .X(_12903_));
 sg13g2_a21oi_1 _19994_ (.A1(net1184),
    .A2(net4400),
    .Y(_12904_),
    .B1(_12903_));
 sg13g2_nand2_1 _19995_ (.Y(_12905_),
    .A(net1384),
    .B(net4078));
 sg13g2_o21ai_1 _19996_ (.B1(_12905_),
    .Y(_00043_),
    .A1(net4078),
    .A2(_12904_));
 sg13g2_and2_1 _19997_ (.A(\shift_reg[25] ),
    .B(net4459),
    .X(_12906_));
 sg13g2_a21oi_1 _19998_ (.A1(\inv_result[33] ),
    .A2(net4400),
    .Y(_12907_),
    .B1(_12906_));
 sg13g2_nand2_1 _19999_ (.Y(_12908_),
    .A(net1132),
    .B(net4077));
 sg13g2_o21ai_1 _20000_ (.B1(_12908_),
    .Y(_00044_),
    .A1(net4078),
    .A2(_12907_));
 sg13g2_and2_1 _20001_ (.A(net1210),
    .B(net4458),
    .X(_12909_));
 sg13g2_a21oi_1 _20002_ (.A1(\inv_result[34] ),
    .A2(net4400),
    .Y(_12910_),
    .B1(_12909_));
 sg13g2_nand2_1 _20003_ (.Y(_12911_),
    .A(net1388),
    .B(net4078));
 sg13g2_o21ai_1 _20004_ (.B1(_12911_),
    .Y(_00045_),
    .A1(net4078),
    .A2(_12910_));
 sg13g2_and2_1 _20005_ (.A(\shift_reg[27] ),
    .B(net4463),
    .X(_12912_));
 sg13g2_a21oi_1 _20006_ (.A1(net1074),
    .A2(net4400),
    .Y(_12913_),
    .B1(_12912_));
 sg13g2_nand2_1 _20007_ (.Y(_12914_),
    .A(net1162),
    .B(net4077));
 sg13g2_o21ai_1 _20008_ (.B1(_12914_),
    .Y(_00046_),
    .A1(net4081),
    .A2(_12913_));
 sg13g2_and2_1 _20009_ (.A(net1160),
    .B(net4459),
    .X(_12915_));
 sg13g2_a21oi_1 _20010_ (.A1(\inv_result[36] ),
    .A2(net4400),
    .Y(_12916_),
    .B1(_12915_));
 sg13g2_nand2_1 _20011_ (.Y(_12917_),
    .A(net1429),
    .B(net4077));
 sg13g2_o21ai_1 _20012_ (.B1(_12917_),
    .Y(_00047_),
    .A1(net4077),
    .A2(_12916_));
 sg13g2_and2_1 _20013_ (.A(\shift_reg[29] ),
    .B(net4458),
    .X(_12918_));
 sg13g2_a21oi_1 _20014_ (.A1(net1072),
    .A2(net4401),
    .Y(_12919_),
    .B1(_12918_));
 sg13g2_nand2_1 _20015_ (.Y(_12920_),
    .A(net1355),
    .B(net4077));
 sg13g2_o21ai_1 _20016_ (.B1(_12920_),
    .Y(_00048_),
    .A1(net4077),
    .A2(_12919_));
 sg13g2_and2_1 _20017_ (.A(net1155),
    .B(net4458),
    .X(_12921_));
 sg13g2_a21oi_1 _20018_ (.A1(\inv_result[38] ),
    .A2(net4400),
    .Y(_12922_),
    .B1(_12921_));
 sg13g2_nand2_1 _20019_ (.Y(_12923_),
    .A(net1261),
    .B(net4078));
 sg13g2_o21ai_1 _20020_ (.B1(_12923_),
    .Y(_00049_),
    .A1(net4078),
    .A2(_12922_));
 sg13g2_and2_1 _20021_ (.A(net1148),
    .B(net4458),
    .X(_12924_));
 sg13g2_a21oi_1 _20022_ (.A1(\inv_result[39] ),
    .A2(net4401),
    .Y(_12925_),
    .B1(_12924_));
 sg13g2_nand2_1 _20023_ (.Y(_12926_),
    .A(net1479),
    .B(net4079));
 sg13g2_o21ai_1 _20024_ (.B1(_12926_),
    .Y(_00050_),
    .A1(net4077),
    .A2(_12925_));
 sg13g2_and2_1 _20025_ (.A(\shift_reg[32] ),
    .B(net4463),
    .X(_12927_));
 sg13g2_a21oi_1 _20026_ (.A1(net1223),
    .A2(net4401),
    .Y(_12928_),
    .B1(_12927_));
 sg13g2_nand2_1 _20027_ (.Y(_12929_),
    .A(net1336),
    .B(net4080));
 sg13g2_o21ai_1 _20028_ (.B1(_12929_),
    .Y(_00051_),
    .A1(net4080),
    .A2(_12928_));
 sg13g2_and2_1 _20029_ (.A(net1132),
    .B(net4463),
    .X(_12930_));
 sg13g2_a21oi_1 _20030_ (.A1(\inv_result[41] ),
    .A2(net4401),
    .Y(_12931_),
    .B1(_12930_));
 sg13g2_nand2_1 _20031_ (.Y(_12932_),
    .A(net1310),
    .B(net4079));
 sg13g2_o21ai_1 _20032_ (.B1(_12932_),
    .Y(_00052_),
    .A1(net4079),
    .A2(_12931_));
 sg13g2_and2_1 _20033_ (.A(\shift_reg[34] ),
    .B(net4463),
    .X(_12933_));
 sg13g2_a21oi_1 _20034_ (.A1(net1078),
    .A2(net4400),
    .Y(_12934_),
    .B1(_12933_));
 sg13g2_nand2_1 _20035_ (.Y(_12935_),
    .A(net1274),
    .B(net4080));
 sg13g2_o21ai_1 _20036_ (.B1(_12935_),
    .Y(_00053_),
    .A1(net4080),
    .A2(_12934_));
 sg13g2_and2_1 _20037_ (.A(net1162),
    .B(net4463),
    .X(_12936_));
 sg13g2_a21oi_1 _20038_ (.A1(net1077),
    .A2(net4400),
    .Y(_12937_),
    .B1(_12936_));
 sg13g2_nand2_1 _20039_ (.Y(_12938_),
    .A(net1483),
    .B(net4079));
 sg13g2_o21ai_1 _20040_ (.B1(_12938_),
    .Y(_00054_),
    .A1(net4079),
    .A2(_12937_));
 sg13g2_and2_1 _20041_ (.A(\shift_reg[36] ),
    .B(net4464),
    .X(_12939_));
 sg13g2_a21oi_1 _20042_ (.A1(\inv_result[44] ),
    .A2(net4402),
    .Y(_12940_),
    .B1(_12939_));
 sg13g2_nand2_1 _20043_ (.Y(_12941_),
    .A(net1151),
    .B(net4080));
 sg13g2_o21ai_1 _20044_ (.B1(_12941_),
    .Y(_00055_),
    .A1(net4081),
    .A2(_12940_));
 sg13g2_nor2_1 _20045_ (.A(_10996_),
    .B(net4464),
    .Y(_12942_));
 sg13g2_a21oi_1 _20046_ (.A1(net1355),
    .A2(net4464),
    .Y(_12943_),
    .B1(_12942_));
 sg13g2_nand2_1 _20047_ (.Y(_12944_),
    .A(net2136),
    .B(net4079));
 sg13g2_o21ai_1 _20048_ (.B1(_12944_),
    .Y(_00056_),
    .A1(net4081),
    .A2(_12943_));
 sg13g2_and2_1 _20049_ (.A(net1261),
    .B(net4463),
    .X(_12945_));
 sg13g2_a21oi_1 _20050_ (.A1(net1502),
    .A2(net4402),
    .Y(_12946_),
    .B1(_12945_));
 sg13g2_nand2_1 _20051_ (.Y(_12947_),
    .A(net1842),
    .B(net4080));
 sg13g2_o21ai_1 _20052_ (.B1(_12947_),
    .Y(_00057_),
    .A1(net4080),
    .A2(_12946_));
 sg13g2_and2_1 _20053_ (.A(net1479),
    .B(net4464),
    .X(_12948_));
 sg13g2_a21oi_1 _20054_ (.A1(\inv_result[47] ),
    .A2(net4402),
    .Y(_12949_),
    .B1(_12948_));
 sg13g2_nand2_1 _20055_ (.Y(_12950_),
    .A(net1711),
    .B(net4079));
 sg13g2_o21ai_1 _20056_ (.B1(_12950_),
    .Y(_00058_),
    .A1(net4079),
    .A2(_12949_));
 sg13g2_and2_1 _20057_ (.A(net1336),
    .B(net4464),
    .X(_12951_));
 sg13g2_a21oi_2 _20058_ (.B1(_12951_),
    .Y(_12952_),
    .A2(net4399),
    .A1(net1141));
 sg13g2_nand2_1 _20059_ (.Y(_12953_),
    .A(net1804),
    .B(net4088));
 sg13g2_o21ai_1 _20060_ (.B1(_12953_),
    .Y(_00059_),
    .A1(net4088),
    .A2(_12952_));
 sg13g2_and2_1 _20061_ (.A(net1310),
    .B(net4464),
    .X(_12954_));
 sg13g2_a21oi_1 _20062_ (.A1(\inv_result[49] ),
    .A2(net4408),
    .Y(_12955_),
    .B1(_12954_));
 sg13g2_nand2_1 _20063_ (.Y(_12956_),
    .A(net1420),
    .B(net4092));
 sg13g2_o21ai_1 _20064_ (.B1(_12956_),
    .Y(_00060_),
    .A1(net4088),
    .A2(_12955_));
 sg13g2_and2_1 _20065_ (.A(\shift_reg[42] ),
    .B(net4463),
    .X(_12957_));
 sg13g2_a21oi_1 _20066_ (.A1(\inv_result[50] ),
    .A2(net4408),
    .Y(_12958_),
    .B1(_12957_));
 sg13g2_nand2_1 _20067_ (.Y(_12959_),
    .A(net1198),
    .B(net4092));
 sg13g2_o21ai_1 _20068_ (.B1(_12959_),
    .Y(_00061_),
    .A1(net4088),
    .A2(_12958_));
 sg13g2_and2_1 _20069_ (.A(\shift_reg[43] ),
    .B(net4464),
    .X(_12960_));
 sg13g2_a21oi_1 _20070_ (.A1(\inv_result[51] ),
    .A2(net4408),
    .Y(_12961_),
    .B1(_12960_));
 sg13g2_nand2_1 _20071_ (.Y(_12962_),
    .A(net1123),
    .B(net4088));
 sg13g2_o21ai_1 _20072_ (.B1(_12962_),
    .Y(_00062_),
    .A1(net4088),
    .A2(_12961_));
 sg13g2_and2_1 _20073_ (.A(net1151),
    .B(net4464),
    .X(_12963_));
 sg13g2_a21oi_1 _20074_ (.A1(net1256),
    .A2(net4408),
    .Y(_12964_),
    .B1(_12963_));
 sg13g2_nand2_1 _20075_ (.Y(_12965_),
    .A(net1278),
    .B(net4090));
 sg13g2_o21ai_1 _20076_ (.B1(_12965_),
    .Y(_00063_),
    .A1(net4090),
    .A2(_12964_));
 sg13g2_nor2_1 _20077_ (.A(_10997_),
    .B(net4467),
    .Y(_12966_));
 sg13g2_a21oi_1 _20078_ (.A1(\shift_reg[45] ),
    .A2(net4470),
    .Y(_12967_),
    .B1(_12966_));
 sg13g2_nand2_1 _20079_ (.Y(_12968_),
    .A(net1541),
    .B(net4088));
 sg13g2_o21ai_1 _20080_ (.B1(_12968_),
    .Y(_00064_),
    .A1(net4088),
    .A2(_12967_));
 sg13g2_and2_1 _20081_ (.A(\shift_reg[46] ),
    .B(net4470),
    .X(_12969_));
 sg13g2_a21oi_1 _20082_ (.A1(net1094),
    .A2(net4407),
    .Y(_12970_),
    .B1(_12969_));
 sg13g2_nand2_1 _20083_ (.Y(_12971_),
    .A(net1284),
    .B(net4091));
 sg13g2_o21ai_1 _20084_ (.B1(_12971_),
    .Y(_00065_),
    .A1(net4091),
    .A2(_12970_));
 sg13g2_and2_1 _20085_ (.A(\shift_reg[47] ),
    .B(net4470),
    .X(_12972_));
 sg13g2_a21oi_1 _20086_ (.A1(\inv_result[55] ),
    .A2(net4407),
    .Y(_12973_),
    .B1(_12972_));
 sg13g2_nand2_1 _20087_ (.Y(_12974_),
    .A(net1232),
    .B(net4089));
 sg13g2_o21ai_1 _20088_ (.B1(_12974_),
    .Y(_00066_),
    .A1(net4089),
    .A2(_12973_));
 sg13g2_and2_1 _20089_ (.A(\shift_reg[48] ),
    .B(net4470),
    .X(_12975_));
 sg13g2_a21oi_1 _20090_ (.A1(net1080),
    .A2(net4405),
    .Y(_12976_),
    .B1(_12975_));
 sg13g2_nand2_1 _20091_ (.Y(_12977_),
    .A(net1350),
    .B(net4091));
 sg13g2_o21ai_1 _20092_ (.B1(_12977_),
    .Y(_00067_),
    .A1(net4091),
    .A2(_12976_));
 sg13g2_and2_1 _20093_ (.A(net1420),
    .B(net4470),
    .X(_12978_));
 sg13g2_a21oi_1 _20094_ (.A1(net1508),
    .A2(net4406),
    .Y(_12979_),
    .B1(_12978_));
 sg13g2_nand2_1 _20095_ (.Y(_12980_),
    .A(net1650),
    .B(net4089));
 sg13g2_o21ai_1 _20096_ (.B1(_12980_),
    .Y(_00068_),
    .A1(net4089),
    .A2(_12979_));
 sg13g2_and2_1 _20097_ (.A(net1198),
    .B(net4471),
    .X(_12981_));
 sg13g2_a21oi_1 _20098_ (.A1(\inv_result[58] ),
    .A2(net4406),
    .Y(_12982_),
    .B1(_12981_));
 sg13g2_nand2_1 _20099_ (.Y(_12983_),
    .A(net1572),
    .B(net4089));
 sg13g2_o21ai_1 _20100_ (.B1(_12983_),
    .Y(_00069_),
    .A1(net4090),
    .A2(_12982_));
 sg13g2_and2_1 _20101_ (.A(net1123),
    .B(net4470),
    .X(_12984_));
 sg13g2_a21oi_1 _20102_ (.A1(net1299),
    .A2(net4407),
    .Y(_12985_),
    .B1(_12984_));
 sg13g2_nand2_1 _20103_ (.Y(_12986_),
    .A(net1383),
    .B(net4089));
 sg13g2_o21ai_1 _20104_ (.B1(_12986_),
    .Y(_00070_),
    .A1(net4089),
    .A2(_12985_));
 sg13g2_and2_1 _20105_ (.A(net1278),
    .B(net4471),
    .X(_12987_));
 sg13g2_a21oi_1 _20106_ (.A1(\inv_result[60] ),
    .A2(net4406),
    .Y(_12988_),
    .B1(_12987_));
 sg13g2_nand2_1 _20107_ (.Y(_12989_),
    .A(net1589),
    .B(net4091));
 sg13g2_o21ai_1 _20108_ (.B1(_12989_),
    .Y(_00071_),
    .A1(net4091),
    .A2(_12988_));
 sg13g2_and2_1 _20109_ (.A(net1541),
    .B(net4471),
    .X(_12990_));
 sg13g2_a21oi_1 _20110_ (.A1(net1377),
    .A2(net4406),
    .Y(_12991_),
    .B1(_12990_));
 sg13g2_nand2_1 _20111_ (.Y(_12992_),
    .A(net2363),
    .B(net4089));
 sg13g2_o21ai_1 _20112_ (.B1(_12992_),
    .Y(_00072_),
    .A1(net4090),
    .A2(_12991_));
 sg13g2_and2_1 _20113_ (.A(net1284),
    .B(net4469),
    .X(_12993_));
 sg13g2_a21oi_1 _20114_ (.A1(net1095),
    .A2(net4406),
    .Y(_12994_),
    .B1(_12993_));
 sg13g2_nand2_1 _20115_ (.Y(_12995_),
    .A(net1332),
    .B(net4095));
 sg13g2_o21ai_1 _20116_ (.B1(_12995_),
    .Y(_00073_),
    .A1(net4095),
    .A2(_12994_));
 sg13g2_and2_1 _20117_ (.A(net1232),
    .B(net4469),
    .X(_12996_));
 sg13g2_a21oi_1 _20118_ (.A1(\inv_result[63] ),
    .A2(net4406),
    .Y(_12997_),
    .B1(_12996_));
 sg13g2_nand2_1 _20119_ (.Y(_12998_),
    .A(net1519),
    .B(net4099));
 sg13g2_o21ai_1 _20120_ (.B1(_12998_),
    .Y(_00074_),
    .A1(net4099),
    .A2(_12997_));
 sg13g2_and2_1 _20121_ (.A(net1350),
    .B(net4469),
    .X(_12999_));
 sg13g2_a21oi_1 _20122_ (.A1(net1393),
    .A2(net4406),
    .Y(_13000_),
    .B1(_12999_));
 sg13g2_nand2_1 _20123_ (.Y(_13001_),
    .A(net1579),
    .B(net4096));
 sg13g2_o21ai_1 _20124_ (.B1(_13001_),
    .Y(_00075_),
    .A1(net4096),
    .A2(_13000_));
 sg13g2_and2_1 _20125_ (.A(\shift_reg[57] ),
    .B(net4469),
    .X(_13002_));
 sg13g2_a21oi_1 _20126_ (.A1(net1236),
    .A2(net4406),
    .Y(_13003_),
    .B1(_13002_));
 sg13g2_nand2_1 _20127_ (.Y(_13004_),
    .A(net1473),
    .B(net4095));
 sg13g2_o21ai_1 _20128_ (.B1(_13004_),
    .Y(_00076_),
    .A1(net4095),
    .A2(_13003_));
 sg13g2_and2_1 _20129_ (.A(\shift_reg[58] ),
    .B(net4469),
    .X(_13005_));
 sg13g2_a21oi_1 _20130_ (.A1(\inv_result[66] ),
    .A2(net4410),
    .Y(_13006_),
    .B1(_13005_));
 sg13g2_nand2_1 _20131_ (.Y(_13007_),
    .A(net1485),
    .B(net4095));
 sg13g2_o21ai_1 _20132_ (.B1(_13007_),
    .Y(_00077_),
    .A1(net4096),
    .A2(_13006_));
 sg13g2_and2_1 _20133_ (.A(net1383),
    .B(net4469),
    .X(_13008_));
 sg13g2_a21oi_1 _20134_ (.A1(\inv_result[67] ),
    .A2(net4407),
    .Y(_13009_),
    .B1(_13008_));
 sg13g2_nand2_1 _20135_ (.Y(_13010_),
    .A(net1386),
    .B(net4099));
 sg13g2_o21ai_1 _20136_ (.B1(_13010_),
    .Y(_00078_),
    .A1(net4099),
    .A2(_13009_));
 sg13g2_and2_1 _20137_ (.A(\shift_reg[60] ),
    .B(net4469),
    .X(_13011_));
 sg13g2_a21oi_1 _20138_ (.A1(\inv_result[68] ),
    .A2(net4410),
    .Y(_13012_),
    .B1(_13011_));
 sg13g2_nand2_1 _20139_ (.Y(_13013_),
    .A(net1286),
    .B(net4096));
 sg13g2_o21ai_1 _20140_ (.B1(_13013_),
    .Y(_00079_),
    .A1(net4095),
    .A2(_13012_));
 sg13g2_and2_1 _20141_ (.A(\shift_reg[61] ),
    .B(net4473),
    .X(_13014_));
 sg13g2_a21oi_1 _20142_ (.A1(\inv_result[69] ),
    .A2(net4410),
    .Y(_13015_),
    .B1(_13014_));
 sg13g2_nand2_1 _20143_ (.Y(_13016_),
    .A(net1157),
    .B(net4095));
 sg13g2_o21ai_1 _20144_ (.B1(_13016_),
    .Y(_00080_),
    .A1(net4095),
    .A2(_13015_));
 sg13g2_and2_1 _20145_ (.A(net1332),
    .B(net4474),
    .X(_13017_));
 sg13g2_a21oi_1 _20146_ (.A1(net1185),
    .A2(net4412),
    .Y(_13018_),
    .B1(_13017_));
 sg13g2_nand2_1 _20147_ (.Y(_13019_),
    .A(net1408),
    .B(net4097));
 sg13g2_o21ai_1 _20148_ (.B1(_13019_),
    .Y(_00081_),
    .A1(net4097),
    .A2(_13018_));
 sg13g2_and2_1 _20149_ (.A(\shift_reg[63] ),
    .B(net4473),
    .X(_13020_));
 sg13g2_a21oi_1 _20150_ (.A1(\inv_result[71] ),
    .A2(net4410),
    .Y(_13021_),
    .B1(_13020_));
 sg13g2_nand2_1 _20151_ (.Y(_13022_),
    .A(net1257),
    .B(net4097));
 sg13g2_o21ai_1 _20152_ (.B1(_13022_),
    .Y(_00082_),
    .A1(net4098),
    .A2(_13021_));
 sg13g2_and2_1 _20153_ (.A(\shift_reg[64] ),
    .B(net4473),
    .X(_13023_));
 sg13g2_a21oi_1 _20154_ (.A1(\inv_result[72] ),
    .A2(net4410),
    .Y(_13024_),
    .B1(_13023_));
 sg13g2_nand2_1 _20155_ (.Y(_13025_),
    .A(net1208),
    .B(net4097));
 sg13g2_o21ai_1 _20156_ (.B1(_13025_),
    .Y(_00083_),
    .A1(net4097),
    .A2(_13024_));
 sg13g2_and2_1 _20157_ (.A(net1473),
    .B(net4473),
    .X(_13026_));
 sg13g2_a21oi_1 _20158_ (.A1(\inv_result[73] ),
    .A2(net4410),
    .Y(_13027_),
    .B1(_13026_));
 sg13g2_nand2_1 _20159_ (.Y(_13028_),
    .A(net1570),
    .B(net4098));
 sg13g2_o21ai_1 _20160_ (.B1(_13028_),
    .Y(_00084_),
    .A1(net4098),
    .A2(_13027_));
 sg13g2_and2_1 _20161_ (.A(\shift_reg[66] ),
    .B(net4474),
    .X(_13029_));
 sg13g2_a21oi_1 _20162_ (.A1(net1101),
    .A2(net4411),
    .Y(_13030_),
    .B1(_13029_));
 sg13g2_nand2_1 _20163_ (.Y(_13031_),
    .A(net1238),
    .B(net4102));
 sg13g2_o21ai_1 _20164_ (.B1(_13031_),
    .Y(_00085_),
    .A1(net4102),
    .A2(_13030_));
 sg13g2_and2_1 _20165_ (.A(net1386),
    .B(net4477),
    .X(_13032_));
 sg13g2_a21oi_1 _20166_ (.A1(\inv_result[75] ),
    .A2(net4411),
    .Y(_13033_),
    .B1(_13032_));
 sg13g2_nand2_1 _20167_ (.Y(_13034_),
    .A(net1402),
    .B(net4103));
 sg13g2_o21ai_1 _20168_ (.B1(_13034_),
    .Y(_00086_),
    .A1(net4103),
    .A2(_13033_));
 sg13g2_and2_1 _20169_ (.A(net1286),
    .B(net4473),
    .X(_13035_));
 sg13g2_a21oi_1 _20170_ (.A1(\inv_result[76] ),
    .A2(net4410),
    .Y(_13036_),
    .B1(_13035_));
 sg13g2_nand2_1 _20171_ (.Y(_13037_),
    .A(net1459),
    .B(net4103));
 sg13g2_o21ai_1 _20172_ (.B1(_13037_),
    .Y(_00087_),
    .A1(net4097),
    .A2(_13036_));
 sg13g2_and2_1 _20173_ (.A(net1157),
    .B(net4473),
    .X(_13038_));
 sg13g2_a21oi_1 _20174_ (.A1(\inv_result[77] ),
    .A2(net4411),
    .Y(_13039_),
    .B1(_13038_));
 sg13g2_nand2_1 _20175_ (.Y(_13040_),
    .A(net1477),
    .B(net4100));
 sg13g2_o21ai_1 _20176_ (.B1(_13040_),
    .Y(_00088_),
    .A1(net4100),
    .A2(_13039_));
 sg13g2_and2_1 _20177_ (.A(\shift_reg[70] ),
    .B(net4474),
    .X(_13041_));
 sg13g2_a21oi_1 _20178_ (.A1(\inv_result[78] ),
    .A2(net4410),
    .Y(_13042_),
    .B1(_13041_));
 sg13g2_nand2_1 _20179_ (.Y(_13043_),
    .A(net1380),
    .B(net4100));
 sg13g2_o21ai_1 _20180_ (.B1(_13043_),
    .Y(_00089_),
    .A1(net4100),
    .A2(_13042_));
 sg13g2_and2_1 _20181_ (.A(net1257),
    .B(net4474),
    .X(_13044_));
 sg13g2_a21oi_1 _20182_ (.A1(\inv_result[79] ),
    .A2(net4411),
    .Y(_13045_),
    .B1(_13044_));
 sg13g2_nand2_1 _20183_ (.Y(_13046_),
    .A(net1317),
    .B(net4102));
 sg13g2_o21ai_1 _20184_ (.B1(_13046_),
    .Y(_00090_),
    .A1(net4102),
    .A2(_13045_));
 sg13g2_and2_1 _20185_ (.A(net1208),
    .B(net4474),
    .X(_13047_));
 sg13g2_a21oi_1 _20186_ (.A1(net1134),
    .A2(net4411),
    .Y(_13048_),
    .B1(_13047_));
 sg13g2_nand2_1 _20187_ (.Y(_13049_),
    .A(net1339),
    .B(net4100));
 sg13g2_o21ai_1 _20188_ (.B1(_13049_),
    .Y(_00091_),
    .A1(net4100),
    .A2(_13048_));
 sg13g2_nor2_1 _20189_ (.A(_10998_),
    .B(net4476),
    .Y(_13050_));
 sg13g2_a21oi_1 _20190_ (.A1(\shift_reg[73] ),
    .A2(net4476),
    .Y(_13051_),
    .B1(_13050_));
 sg13g2_nand2_1 _20191_ (.Y(_13052_),
    .A(net1282),
    .B(net4101));
 sg13g2_o21ai_1 _20192_ (.B1(_13052_),
    .Y(_00092_),
    .A1(net4101),
    .A2(_13051_));
 sg13g2_and2_1 _20193_ (.A(net1238),
    .B(net4475),
    .X(_13053_));
 sg13g2_a21oi_1 _20194_ (.A1(\inv_result[82] ),
    .A2(net4414),
    .Y(_13054_),
    .B1(_13053_));
 sg13g2_nand2_1 _20195_ (.Y(_13055_),
    .A(net1465),
    .B(net4105));
 sg13g2_o21ai_1 _20196_ (.B1(_13055_),
    .Y(_00093_),
    .A1(net4105),
    .A2(_13054_));
 sg13g2_nor2_1 _20197_ (.A(_10999_),
    .B(net4475),
    .Y(_13056_));
 sg13g2_a21oi_1 _20198_ (.A1(\shift_reg[75] ),
    .A2(net4475),
    .Y(_13057_),
    .B1(_13056_));
 sg13g2_nand2_1 _20199_ (.Y(_13058_),
    .A(net1343),
    .B(net4102));
 sg13g2_o21ai_1 _20200_ (.B1(_13058_),
    .Y(_00094_),
    .A1(net4102),
    .A2(_13057_));
 sg13g2_and2_1 _20201_ (.A(net1459),
    .B(net4476),
    .X(_13059_));
 sg13g2_a21oi_1 _20202_ (.A1(\inv_result[84] ),
    .A2(net4411),
    .Y(_13060_),
    .B1(_13059_));
 sg13g2_nand2_1 _20203_ (.Y(_13061_),
    .A(net1471),
    .B(net4101));
 sg13g2_o21ai_1 _20204_ (.B1(_13061_),
    .Y(_00095_),
    .A1(net4101),
    .A2(_13060_));
 sg13g2_nor2_1 _20205_ (.A(_11000_),
    .B(net4476),
    .Y(_13062_));
 sg13g2_a21oi_1 _20206_ (.A1(\shift_reg[77] ),
    .A2(net4476),
    .Y(_13063_),
    .B1(_13062_));
 sg13g2_nand2_1 _20207_ (.Y(_13064_),
    .A(net1253),
    .B(net4101));
 sg13g2_o21ai_1 _20208_ (.B1(_13064_),
    .Y(_00096_),
    .A1(net4101),
    .A2(_13063_));
 sg13g2_and2_1 _20209_ (.A(net1380),
    .B(net4476),
    .X(_13065_));
 sg13g2_a21oi_1 _20210_ (.A1(net1434),
    .A2(net4412),
    .Y(_13066_),
    .B1(_13065_));
 sg13g2_nand2_1 _20211_ (.Y(_13067_),
    .A(net1444),
    .B(net4101));
 sg13g2_o21ai_1 _20212_ (.B1(_13067_),
    .Y(_00097_),
    .A1(net4101),
    .A2(_13066_));
 sg13g2_and2_1 _20213_ (.A(\shift_reg[79] ),
    .B(net4475),
    .X(_13068_));
 sg13g2_a21oi_1 _20214_ (.A1(\inv_result[87] ),
    .A2(net4412),
    .Y(_13069_),
    .B1(_13068_));
 sg13g2_nand2_1 _20215_ (.Y(_13070_),
    .A(net1247),
    .B(net4102));
 sg13g2_o21ai_1 _20216_ (.B1(_13070_),
    .Y(_00098_),
    .A1(net4102),
    .A2(_13069_));
 sg13g2_and2_1 _20217_ (.A(\shift_reg[80] ),
    .B(net4476),
    .X(_13071_));
 sg13g2_a21oi_1 _20218_ (.A1(\inv_result[88] ),
    .A2(net4414),
    .Y(_13072_),
    .B1(_13071_));
 sg13g2_nand2_1 _20219_ (.Y(_13073_),
    .A(net1291),
    .B(net4105));
 sg13g2_o21ai_1 _20220_ (.B1(_13073_),
    .Y(_00099_),
    .A1(net4106),
    .A2(_13072_));
 sg13g2_nor2_1 _20221_ (.A(_11001_),
    .B(net4479),
    .Y(_13074_));
 sg13g2_a21oi_1 _20222_ (.A1(net1282),
    .A2(net4479),
    .Y(_13075_),
    .B1(_13074_));
 sg13g2_nand2_1 _20223_ (.Y(_13076_),
    .A(net1328),
    .B(net4106));
 sg13g2_o21ai_1 _20224_ (.B1(_13076_),
    .Y(_00100_),
    .A1(net4105),
    .A2(_13075_));
 sg13g2_and2_1 _20225_ (.A(\shift_reg[82] ),
    .B(net4479),
    .X(_13077_));
 sg13g2_a21oi_1 _20226_ (.A1(\inv_result[90] ),
    .A2(net4414),
    .Y(_13078_),
    .B1(_13077_));
 sg13g2_nand2_1 _20227_ (.Y(_13079_),
    .A(net1378),
    .B(net4108));
 sg13g2_o21ai_1 _20228_ (.B1(_13079_),
    .Y(_00101_),
    .A1(net4108),
    .A2(_13078_));
 sg13g2_and2_1 _20229_ (.A(net1343),
    .B(net4475),
    .X(_13080_));
 sg13g2_a21oi_1 _20230_ (.A1(net1177),
    .A2(net4414),
    .Y(_13081_),
    .B1(_13080_));
 sg13g2_nand2_1 _20231_ (.Y(_13082_),
    .A(net1615),
    .B(net4106));
 sg13g2_o21ai_1 _20232_ (.B1(_13082_),
    .Y(_00102_),
    .A1(net4106),
    .A2(_13081_));
 sg13g2_and2_1 _20233_ (.A(net1471),
    .B(net4475),
    .X(_13083_));
 sg13g2_a21oi_1 _20234_ (.A1(\inv_result[92] ),
    .A2(net4411),
    .Y(_13084_),
    .B1(_13083_));
 sg13g2_nand2_1 _20235_ (.Y(_13085_),
    .A(net1481),
    .B(net4105));
 sg13g2_o21ai_1 _20236_ (.B1(_13085_),
    .Y(_00103_),
    .A1(net4105),
    .A2(_13084_));
 sg13g2_nor2_1 _20237_ (.A(_11002_),
    .B(net4479),
    .Y(_13086_));
 sg13g2_a21oi_1 _20238_ (.A1(\shift_reg[85] ),
    .A2(net4479),
    .Y(_13087_),
    .B1(_13086_));
 sg13g2_nand2_1 _20239_ (.Y(_13088_),
    .A(net1204),
    .B(net4105));
 sg13g2_o21ai_1 _20240_ (.B1(_13088_),
    .Y(_00104_),
    .A1(net4106),
    .A2(_13087_));
 sg13g2_and2_1 _20241_ (.A(\shift_reg[86] ),
    .B(net4479),
    .X(_13089_));
 sg13g2_a21oi_1 _20242_ (.A1(\inv_result[94] ),
    .A2(net4414),
    .Y(_13090_),
    .B1(_13089_));
 sg13g2_nand2_1 _20243_ (.Y(_13091_),
    .A(net1330),
    .B(net4107));
 sg13g2_o21ai_1 _20244_ (.B1(_13091_),
    .Y(_00105_),
    .A1(net4106),
    .A2(_13090_));
 sg13g2_and2_1 _20245_ (.A(net1247),
    .B(net4475),
    .X(_13092_));
 sg13g2_a21oi_1 _20246_ (.A1(net1551),
    .A2(net4414),
    .Y(_13093_),
    .B1(_13092_));
 sg13g2_nand2_1 _20247_ (.Y(_13094_),
    .A(net1678),
    .B(net4107));
 sg13g2_o21ai_1 _20248_ (.B1(_13094_),
    .Y(_00106_),
    .A1(net4105),
    .A2(_13093_));
 sg13g2_and2_1 _20249_ (.A(net1291),
    .B(net4478),
    .X(_13095_));
 sg13g2_a21oi_1 _20250_ (.A1(net1636),
    .A2(net4415),
    .Y(_13096_),
    .B1(_13095_));
 sg13g2_nand2_1 _20251_ (.Y(_13097_),
    .A(net1731),
    .B(net4111));
 sg13g2_o21ai_1 _20252_ (.B1(_13097_),
    .Y(_00107_),
    .A1(net4110),
    .A2(_13096_));
 sg13g2_nor2_1 _20253_ (.A(_11003_),
    .B(net4478),
    .Y(_13098_));
 sg13g2_a21oi_1 _20254_ (.A1(net1328),
    .A2(net4478),
    .Y(_13099_),
    .B1(_13098_));
 sg13g2_nand2_1 _20255_ (.Y(_13100_),
    .A(net1361),
    .B(net4110));
 sg13g2_o21ai_1 _20256_ (.B1(_13100_),
    .Y(_00108_),
    .A1(net4110),
    .A2(_13099_));
 sg13g2_and2_1 _20257_ (.A(net1378),
    .B(net4478),
    .X(_13101_));
 sg13g2_a21oi_1 _20258_ (.A1(net1757),
    .A2(net4414),
    .Y(_13102_),
    .B1(_13101_));
 sg13g2_nand2_1 _20259_ (.Y(_13103_),
    .A(net1899),
    .B(net4113));
 sg13g2_o21ai_1 _20260_ (.B1(_13103_),
    .Y(_00109_),
    .A1(net4110),
    .A2(_13102_));
 sg13g2_and2_1 _20261_ (.A(\shift_reg[91] ),
    .B(net4478),
    .X(_13104_));
 sg13g2_a21oi_1 _20262_ (.A1(\inv_result[99] ),
    .A2(net4415),
    .Y(_13105_),
    .B1(_13104_));
 sg13g2_nand2_1 _20263_ (.Y(_13106_),
    .A(net1469),
    .B(net4110));
 sg13g2_o21ai_1 _20264_ (.B1(_13106_),
    .Y(_00110_),
    .A1(net4112),
    .A2(_13105_));
 sg13g2_and2_1 _20265_ (.A(net1481),
    .B(net4480),
    .X(_13107_));
 sg13g2_a21oi_1 _20266_ (.A1(net1605),
    .A2(net4415),
    .Y(_13108_),
    .B1(_13107_));
 sg13g2_nand2_1 _20267_ (.Y(_13109_),
    .A(net1766),
    .B(net4111));
 sg13g2_o21ai_1 _20268_ (.B1(_13109_),
    .Y(_00111_),
    .A1(net4110),
    .A2(_13108_));
 sg13g2_and2_1 _20269_ (.A(net1204),
    .B(net4480),
    .X(_13110_));
 sg13g2_a21oi_1 _20270_ (.A1(net1692),
    .A2(net4414),
    .Y(_13111_),
    .B1(_13110_));
 sg13g2_nand2_1 _20271_ (.Y(_13112_),
    .A(net1907),
    .B(net4111));
 sg13g2_o21ai_1 _20272_ (.B1(_13112_),
    .Y(_00112_),
    .A1(net4110),
    .A2(_13111_));
 sg13g2_and2_1 _20273_ (.A(net1330),
    .B(net4478),
    .X(_13113_));
 sg13g2_a21oi_1 _20274_ (.A1(net1135),
    .A2(net4415),
    .Y(_13114_),
    .B1(_13113_));
 sg13g2_nand2_1 _20275_ (.Y(_13115_),
    .A(net1991),
    .B(net4110));
 sg13g2_o21ai_1 _20276_ (.B1(_13115_),
    .Y(_00113_),
    .A1(net4107),
    .A2(_13114_));
 sg13g2_and2_1 _20277_ (.A(net1678),
    .B(net4478),
    .X(_13116_));
 sg13g2_a21oi_1 _20278_ (.A1(net1921),
    .A2(net4415),
    .Y(_13117_),
    .B1(_13116_));
 sg13g2_nand2_1 _20279_ (.Y(_13118_),
    .A(net2183),
    .B(net4113));
 sg13g2_o21ai_1 _20280_ (.B1(_13118_),
    .Y(_00114_),
    .A1(net4109),
    .A2(_13117_));
 sg13g2_and2_1 _20281_ (.A(net1731),
    .B(net4481),
    .X(_13119_));
 sg13g2_a21oi_1 _20282_ (.A1(net1574),
    .A2(net4416),
    .Y(_13120_),
    .B1(_13119_));
 sg13g2_nand2_1 _20283_ (.Y(_13121_),
    .A(net1736),
    .B(net4113));
 sg13g2_o21ai_1 _20284_ (.B1(_13121_),
    .Y(_00115_),
    .A1(net4113),
    .A2(_13120_));
 sg13g2_and2_1 _20285_ (.A(\shift_reg[97] ),
    .B(net4481),
    .X(_13122_));
 sg13g2_a21oi_2 _20286_ (.B1(_13122_),
    .Y(_13123_),
    .A2(net4416),
    .A1(\inv_result[105] ));
 sg13g2_nand2_1 _20287_ (.Y(_13124_),
    .A(net1173),
    .B(net4118));
 sg13g2_o21ai_1 _20288_ (.B1(_13124_),
    .Y(_00116_),
    .A1(net4118),
    .A2(_13123_));
 sg13g2_nor2_1 _20289_ (.A(_11004_),
    .B(net4481),
    .Y(_13125_));
 sg13g2_a21oi_1 _20290_ (.A1(\shift_reg[98] ),
    .A2(net4486),
    .Y(_13126_),
    .B1(_13125_));
 sg13g2_nand2_1 _20291_ (.Y(_13127_),
    .A(net1396),
    .B(net4116));
 sg13g2_o21ai_1 _20292_ (.B1(_13127_),
    .Y(_00117_),
    .A1(net4116),
    .A2(_13126_));
 sg13g2_and2_1 _20293_ (.A(\shift_reg[99] ),
    .B(net4481),
    .X(_13128_));
 sg13g2_a21oi_2 _20294_ (.B1(_13128_),
    .Y(_13129_),
    .A2(net4416),
    .A1(\inv_result[107] ));
 sg13g2_nand2_1 _20295_ (.Y(_13130_),
    .A(net1404),
    .B(net4117));
 sg13g2_o21ai_1 _20296_ (.B1(_13130_),
    .Y(_00118_),
    .A1(net4117),
    .A2(_13129_));
 sg13g2_and2_1 _20297_ (.A(\shift_reg[100] ),
    .B(net4481),
    .X(_13131_));
 sg13g2_a21oi_2 _20298_ (.B1(_13131_),
    .Y(_13132_),
    .A2(net4416),
    .A1(\inv_result[108] ));
 sg13g2_nand2_1 _20299_ (.Y(_13133_),
    .A(net1196),
    .B(net4130));
 sg13g2_o21ai_1 _20300_ (.B1(_13133_),
    .Y(_00119_),
    .A1(net4130),
    .A2(_13132_));
 sg13g2_nor2_1 _20301_ (.A(_11005_),
    .B(net4486),
    .Y(_13134_));
 sg13g2_a21oi_1 _20302_ (.A1(\shift_reg[101] ),
    .A2(net4486),
    .Y(_13135_),
    .B1(_13134_));
 sg13g2_nand2_1 _20303_ (.Y(_13136_),
    .A(net1864),
    .B(net4119));
 sg13g2_o21ai_1 _20304_ (.B1(_13136_),
    .Y(_00120_),
    .A1(net4118),
    .A2(_13135_));
 sg13g2_and2_1 _20305_ (.A(\shift_reg[102] ),
    .B(net4481),
    .X(_13137_));
 sg13g2_a21oi_1 _20306_ (.A1(net1581),
    .A2(net4416),
    .Y(_13138_),
    .B1(_13137_));
 sg13g2_nand2_1 _20307_ (.Y(_13139_),
    .A(net1776),
    .B(net4115));
 sg13g2_o21ai_1 _20308_ (.B1(_13139_),
    .Y(_00121_),
    .A1(net4115),
    .A2(_13138_));
 sg13g2_and2_1 _20309_ (.A(\shift_reg[103] ),
    .B(net4483),
    .X(_13140_));
 sg13g2_a21oi_1 _20310_ (.A1(net1511),
    .A2(net4416),
    .Y(_13141_),
    .B1(_13140_));
 sg13g2_nand2_1 _20311_ (.Y(_13142_),
    .A(net2161),
    .B(net4115));
 sg13g2_o21ai_1 _20312_ (.B1(_13142_),
    .Y(_00122_),
    .A1(net4114),
    .A2(_13141_));
 sg13g2_and2_1 _20313_ (.A(\shift_reg[104] ),
    .B(net4485),
    .X(_13143_));
 sg13g2_a21oi_1 _20314_ (.A1(\inv_result[112] ),
    .A2(net4420),
    .Y(_13144_),
    .B1(_13143_));
 sg13g2_nand2_1 _20315_ (.Y(_13145_),
    .A(net1353),
    .B(net4119));
 sg13g2_o21ai_1 _20316_ (.B1(_13145_),
    .Y(_00123_),
    .A1(net4119),
    .A2(_13144_));
 sg13g2_and2_1 _20317_ (.A(net1173),
    .B(net4484),
    .X(_13146_));
 sg13g2_a21oi_2 _20318_ (.B1(_13146_),
    .Y(_13147_),
    .A2(net4419),
    .A1(\inv_result[113] ));
 sg13g2_nand2_1 _20319_ (.Y(_13148_),
    .A(net1629),
    .B(net4137));
 sg13g2_o21ai_1 _20320_ (.B1(_13148_),
    .Y(_00124_),
    .A1(net4133),
    .A2(_13147_));
 sg13g2_and2_1 _20321_ (.A(\shift_reg[106] ),
    .B(net4485),
    .X(_13149_));
 sg13g2_a21oi_1 _20322_ (.A1(net1082),
    .A2(net4420),
    .Y(_13150_),
    .B1(_13149_));
 sg13g2_nand2_1 _20323_ (.Y(_13151_),
    .A(net1107),
    .B(net4134));
 sg13g2_o21ai_1 _20324_ (.B1(_13151_),
    .Y(_00125_),
    .A1(net4134),
    .A2(_13150_));
 sg13g2_nor2_1 _20325_ (.A(_11006_),
    .B(net4499),
    .Y(_13152_));
 sg13g2_a21oi_1 _20326_ (.A1(net1404),
    .A2(net4485),
    .Y(_13153_),
    .B1(_13152_));
 sg13g2_nand2_1 _20327_ (.Y(_13154_),
    .A(net1922),
    .B(net4118));
 sg13g2_o21ai_1 _20328_ (.B1(_13154_),
    .Y(_00126_),
    .A1(net4118),
    .A2(_13153_));
 sg13g2_and2_1 _20329_ (.A(net1196),
    .B(net4494),
    .X(_13155_));
 sg13g2_a21oi_1 _20330_ (.A1(net1591),
    .A2(net4426),
    .Y(_13156_),
    .B1(_13155_));
 sg13g2_nand2_1 _20331_ (.Y(_13157_),
    .A(net1635),
    .B(net4137));
 sg13g2_o21ai_1 _20332_ (.B1(_13157_),
    .Y(_00127_),
    .A1(net4133),
    .A2(_13156_));
 sg13g2_nor2_1 _20333_ (.A(_11007_),
    .B(net4491),
    .Y(_13158_));
 sg13g2_a21oi_1 _20334_ (.A1(\shift_reg[109] ),
    .A2(net4495),
    .Y(_13159_),
    .B1(_13158_));
 sg13g2_nand2_1 _20335_ (.Y(_13160_),
    .A(net1259),
    .B(net4139));
 sg13g2_o21ai_1 _20336_ (.B1(_13160_),
    .Y(_00128_),
    .A1(net4140),
    .A2(_13159_));
 sg13g2_and2_1 _20337_ (.A(net1776),
    .B(net4485),
    .X(_13161_));
 sg13g2_a21oi_1 _20338_ (.A1(net1120),
    .A2(net4419),
    .Y(_13162_),
    .B1(_13161_));
 sg13g2_nand2_1 _20339_ (.Y(_13163_),
    .A(net1961),
    .B(net4130));
 sg13g2_o21ai_1 _20340_ (.B1(_13163_),
    .Y(_00129_),
    .A1(net4118),
    .A2(_13162_));
 sg13g2_and2_1 _20341_ (.A(\shift_reg[111] ),
    .B(net4494),
    .X(_13164_));
 sg13g2_a21oi_1 _20342_ (.A1(\inv_result[119] ),
    .A2(net4426),
    .Y(_13165_),
    .B1(_13164_));
 sg13g2_nand2_1 _20343_ (.Y(_13166_),
    .A(net1774),
    .B(net4134));
 sg13g2_o21ai_1 _20344_ (.B1(_13166_),
    .Y(_00130_),
    .A1(net4134),
    .A2(_13165_));
 sg13g2_and2_1 _20345_ (.A(net1353),
    .B(net4485),
    .X(_13167_));
 sg13g2_a21oi_2 _20346_ (.B1(_13167_),
    .Y(_13168_),
    .A2(net4419),
    .A1(\inv_result[120] ));
 sg13g2_nand2_1 _20347_ (.Y(_13169_),
    .A(net1889),
    .B(net4141));
 sg13g2_o21ai_1 _20348_ (.B1(_13169_),
    .Y(_00131_),
    .A1(net4134),
    .A2(_13168_));
 sg13g2_nor2_1 _20349_ (.A(_11008_),
    .B(net4490),
    .Y(_13170_));
 sg13g2_a21oi_1 _20350_ (.A1(\shift_reg[113] ),
    .A2(net4498),
    .Y(_13171_),
    .B1(_13170_));
 sg13g2_nand2_1 _20351_ (.Y(_13172_),
    .A(net1500),
    .B(net4141));
 sg13g2_o21ai_1 _20352_ (.B1(_13172_),
    .Y(_00132_),
    .A1(net4141),
    .A2(_13171_));
 sg13g2_and2_1 _20353_ (.A(net1107),
    .B(net4494),
    .X(_13173_));
 sg13g2_a21oi_2 _20354_ (.B1(_13173_),
    .Y(_13174_),
    .A2(net4426),
    .A1(\inv_result[122] ));
 sg13g2_nand2_1 _20355_ (.Y(_13175_),
    .A(net1417),
    .B(net4141));
 sg13g2_o21ai_1 _20356_ (.B1(_13175_),
    .Y(_00133_),
    .A1(net4141),
    .A2(_13174_));
 sg13g2_nor2_1 _20357_ (.A(_11009_),
    .B(net4497),
    .Y(_13176_));
 sg13g2_a21oi_1 _20358_ (.A1(\shift_reg[115] ),
    .A2(net4497),
    .Y(_13177_),
    .B1(_13176_));
 sg13g2_nand2_1 _20359_ (.Y(_13178_),
    .A(net1698),
    .B(net4137));
 sg13g2_o21ai_1 _20360_ (.B1(_13178_),
    .Y(_00134_),
    .A1(net4138),
    .A2(_13177_));
 sg13g2_and2_1 _20361_ (.A(\shift_reg[116] ),
    .B(net4496),
    .X(_13179_));
 sg13g2_a21oi_1 _20362_ (.A1(\inv_result[124] ),
    .A2(net4427),
    .Y(_13180_),
    .B1(_13179_));
 sg13g2_nand2_1 _20363_ (.Y(_13181_),
    .A(net1180),
    .B(net4140));
 sg13g2_o21ai_1 _20364_ (.B1(_13181_),
    .Y(_00135_),
    .A1(net4140),
    .A2(_13180_));
 sg13g2_nor2_1 _20365_ (.A(_11010_),
    .B(net4497),
    .Y(_13182_));
 sg13g2_a21oi_1 _20366_ (.A1(net1259),
    .A2(net4497),
    .Y(_13183_),
    .B1(_13182_));
 sg13g2_nand2_1 _20367_ (.Y(_13184_),
    .A(net1986),
    .B(net4140));
 sg13g2_o21ai_1 _20368_ (.B1(_13184_),
    .Y(_00136_),
    .A1(net4139),
    .A2(_13183_));
 sg13g2_and2_1 _20369_ (.A(\shift_reg[118] ),
    .B(net4497),
    .X(_13185_));
 sg13g2_a21oi_1 _20370_ (.A1(net1111),
    .A2(net4427),
    .Y(_13186_),
    .B1(_13185_));
 sg13g2_nand2_1 _20371_ (.Y(_13187_),
    .A(net1530),
    .B(net4137));
 sg13g2_o21ai_1 _20372_ (.B1(_13187_),
    .Y(_00137_),
    .A1(net4137),
    .A2(_13186_));
 sg13g2_and2_1 _20373_ (.A(\shift_reg[119] ),
    .B(net4496),
    .X(_13188_));
 sg13g2_a21oi_1 _20374_ (.A1(\inv_result[127] ),
    .A2(net4424),
    .Y(_13189_),
    .B1(_13188_));
 sg13g2_nand2_1 _20375_ (.Y(_13190_),
    .A(net1112),
    .B(net4139));
 sg13g2_o21ai_1 _20376_ (.B1(_13190_),
    .Y(_00138_),
    .A1(net4139),
    .A2(_13189_));
 sg13g2_and2_1 _20377_ (.A(\shift_reg[120] ),
    .B(net4498),
    .X(_13191_));
 sg13g2_a21oi_1 _20378_ (.A1(\inv_result[128] ),
    .A2(net4423),
    .Y(_13192_),
    .B1(_13191_));
 sg13g2_nand2_1 _20379_ (.Y(_13193_),
    .A(net1326),
    .B(net4129));
 sg13g2_o21ai_1 _20380_ (.B1(_13193_),
    .Y(_00139_),
    .A1(net4129),
    .A2(_13192_));
 sg13g2_and2_1 _20381_ (.A(net1500),
    .B(net4496),
    .X(_13194_));
 sg13g2_a21oi_1 _20382_ (.A1(\inv_result[129] ),
    .A2(net4423),
    .Y(_13195_),
    .B1(_13194_));
 sg13g2_nand2_1 _20383_ (.Y(_13196_),
    .A(net1555),
    .B(net4127));
 sg13g2_o21ai_1 _20384_ (.B1(_13196_),
    .Y(_00140_),
    .A1(net4126),
    .A2(_13195_));
 sg13g2_and2_1 _20385_ (.A(net1417),
    .B(net4498),
    .X(_13197_));
 sg13g2_a21oi_1 _20386_ (.A1(\inv_result[130] ),
    .A2(net4424),
    .Y(_13198_),
    .B1(_13197_));
 sg13g2_nand2_1 _20387_ (.Y(_13199_),
    .A(net1606),
    .B(net4127));
 sg13g2_o21ai_1 _20388_ (.B1(_13199_),
    .Y(_00141_),
    .A1(net4126),
    .A2(_13198_));
 sg13g2_nor2_1 _20389_ (.A(_11011_),
    .B(net4490),
    .Y(_13200_));
 sg13g2_a21oi_1 _20390_ (.A1(\shift_reg[123] ),
    .A2(net4490),
    .Y(_13201_),
    .B1(_13200_));
 sg13g2_nand2_1 _20391_ (.Y(_13202_),
    .A(net1288),
    .B(net4126));
 sg13g2_o21ai_1 _20392_ (.B1(_13202_),
    .Y(_00142_),
    .A1(net4126),
    .A2(_13201_));
 sg13g2_and2_1 _20393_ (.A(net1180),
    .B(net4496),
    .X(_13203_));
 sg13g2_a21oi_1 _20394_ (.A1(net1166),
    .A2(net4421),
    .Y(_13204_),
    .B1(_13203_));
 sg13g2_nand2_1 _20395_ (.Y(_13205_),
    .A(net1218),
    .B(net4121));
 sg13g2_o21ai_1 _20396_ (.B1(_13205_),
    .Y(_00143_),
    .A1(net4122),
    .A2(_13204_));
 sg13g2_nor2_1 _20397_ (.A(_11012_),
    .B(net4487),
    .Y(_13206_));
 sg13g2_a21oi_1 _20398_ (.A1(\shift_reg[125] ),
    .A2(net4487),
    .Y(_13207_),
    .B1(_13206_));
 sg13g2_nand2_1 _20399_ (.Y(_13208_),
    .A(net1265),
    .B(net4121));
 sg13g2_o21ai_1 _20400_ (.B1(_13208_),
    .Y(_00144_),
    .A1(net4121),
    .A2(_13207_));
 sg13g2_and2_1 _20401_ (.A(\shift_reg[126] ),
    .B(net4496),
    .X(_13209_));
 sg13g2_a21oi_1 _20402_ (.A1(net1176),
    .A2(net4421),
    .Y(_13210_),
    .B1(_13209_));
 sg13g2_nand2_1 _20403_ (.Y(_13211_),
    .A(net1414),
    .B(net4122));
 sg13g2_o21ai_1 _20404_ (.B1(_13211_),
    .Y(_00145_),
    .A1(net4122),
    .A2(_13210_));
 sg13g2_and2_1 _20405_ (.A(net1112),
    .B(net4496),
    .X(_13212_));
 sg13g2_a21oi_1 _20406_ (.A1(\inv_result[135] ),
    .A2(net4421),
    .Y(_13213_),
    .B1(_13212_));
 sg13g2_nand2_1 _20407_ (.Y(_13214_),
    .A(net1394),
    .B(net4121));
 sg13g2_o21ai_1 _20408_ (.B1(_13214_),
    .Y(_00146_),
    .A1(net4122),
    .A2(_13213_));
 sg13g2_and2_1 _20409_ (.A(\shift_reg[128] ),
    .B(net4490),
    .X(_13215_));
 sg13g2_a21oi_1 _20410_ (.A1(\inv_result[136] ),
    .A2(net4422),
    .Y(_13216_),
    .B1(_13215_));
 sg13g2_nand2_1 _20411_ (.Y(_13217_),
    .A(net1221),
    .B(net4124));
 sg13g2_o21ai_1 _20412_ (.B1(_13217_),
    .Y(_00147_),
    .A1(net4124),
    .A2(_13216_));
 sg13g2_nor2_1 _20413_ (.A(_11013_),
    .B(net4492),
    .Y(_13218_));
 sg13g2_a21oi_1 _20414_ (.A1(net1555),
    .A2(net4488),
    .Y(_13219_),
    .B1(_13218_));
 sg13g2_nand2_1 _20415_ (.Y(_13220_),
    .A(net1753),
    .B(net4123));
 sg13g2_o21ai_1 _20416_ (.B1(_13220_),
    .Y(_00148_),
    .A1(net4123),
    .A2(_13219_));
 sg13g2_and2_1 _20417_ (.A(\shift_reg[130] ),
    .B(net4488),
    .X(_13221_));
 sg13g2_a21oi_1 _20418_ (.A1(\inv_result[138] ),
    .A2(net4421),
    .Y(_13222_),
    .B1(_13221_));
 sg13g2_nand2_1 _20419_ (.Y(_13223_),
    .A(net1178),
    .B(net4122));
 sg13g2_o21ai_1 _20420_ (.B1(_13223_),
    .Y(_00149_),
    .A1(net4122),
    .A2(_13222_));
 sg13g2_and2_1 _20421_ (.A(\shift_reg[131] ),
    .B(net4488),
    .X(_13224_));
 sg13g2_a21oi_1 _20422_ (.A1(\inv_result[139] ),
    .A2(net4422),
    .Y(_13225_),
    .B1(_13224_));
 sg13g2_nand2_1 _20423_ (.Y(_13226_),
    .A(net1234),
    .B(net4123));
 sg13g2_o21ai_1 _20424_ (.B1(_13226_),
    .Y(_00150_),
    .A1(net4123),
    .A2(_13225_));
 sg13g2_and2_1 _20425_ (.A(net1218),
    .B(net4487),
    .X(_13227_));
 sg13g2_a21oi_1 _20426_ (.A1(net1263),
    .A2(net4421),
    .Y(_13228_),
    .B1(_13227_));
 sg13g2_nand2_1 _20427_ (.Y(_13229_),
    .A(net1364),
    .B(net4121));
 sg13g2_o21ai_1 _20428_ (.B1(_13229_),
    .Y(_00151_),
    .A1(net4121),
    .A2(_13228_));
 sg13g2_nor2_1 _20429_ (.A(_11014_),
    .B(net4487),
    .Y(_13230_));
 sg13g2_a21oi_1 _20430_ (.A1(net1265),
    .A2(net4487),
    .Y(_13231_),
    .B1(_13230_));
 sg13g2_nand2_1 _20431_ (.Y(_13232_),
    .A(net1517),
    .B(net4121));
 sg13g2_o21ai_1 _20432_ (.B1(_13232_),
    .Y(_00152_),
    .A1(net4121),
    .A2(_13231_));
 sg13g2_and2_1 _20433_ (.A(net1414),
    .B(net4489),
    .X(_13233_));
 sg13g2_a21oi_1 _20434_ (.A1(net1553),
    .A2(net4421),
    .Y(_13234_),
    .B1(_13233_));
 sg13g2_nand2_1 _20435_ (.Y(_13235_),
    .A(net1592),
    .B(net4124));
 sg13g2_o21ai_1 _20436_ (.B1(_13235_),
    .Y(_00153_),
    .A1(net4124),
    .A2(_13234_));
 sg13g2_and2_1 _20437_ (.A(net1394),
    .B(net4487),
    .X(_13236_));
 sg13g2_a21oi_1 _20438_ (.A1(\inv_result[143] ),
    .A2(net4421),
    .Y(_13237_),
    .B1(_13236_));
 sg13g2_nand2_1 _20439_ (.Y(_13238_),
    .A(net1648),
    .B(net4123));
 sg13g2_o21ai_1 _20440_ (.B1(_13238_),
    .Y(_00154_),
    .A1(net4123),
    .A2(_13237_));
 sg13g2_and2_1 _20441_ (.A(net1221),
    .B(net4488),
    .X(_13239_));
 sg13g2_a21oi_1 _20442_ (.A1(\inv_result[144] ),
    .A2(net4425),
    .Y(_13240_),
    .B1(_13239_));
 sg13g2_nand2_1 _20443_ (.Y(_13241_),
    .A(net1536),
    .B(net4124));
 sg13g2_o21ai_1 _20444_ (.B1(_13241_),
    .Y(_00155_),
    .A1(net4124),
    .A2(_13240_));
 sg13g2_nor2_1 _20445_ (.A(_11015_),
    .B(net4489),
    .Y(_13242_));
 sg13g2_a21oi_1 _20446_ (.A1(\shift_reg[137] ),
    .A2(net4488),
    .Y(_13243_),
    .B1(_13242_));
 sg13g2_nand2_1 _20447_ (.Y(_13244_),
    .A(net1489),
    .B(net4123));
 sg13g2_o21ai_1 _20448_ (.B1(_13244_),
    .Y(_00156_),
    .A1(net4125),
    .A2(_13243_));
 sg13g2_and2_1 _20449_ (.A(net1178),
    .B(net4487),
    .X(_13245_));
 sg13g2_a21oi_1 _20450_ (.A1(net1352),
    .A2(net4422),
    .Y(_13246_),
    .B1(_13245_));
 sg13g2_nand2_1 _20451_ (.Y(_13247_),
    .A(net1869),
    .B(net4125));
 sg13g2_o21ai_1 _20452_ (.B1(_13247_),
    .Y(_00157_),
    .A1(net4123),
    .A2(_13246_));
 sg13g2_and2_1 _20453_ (.A(net1234),
    .B(net4488),
    .X(_13248_));
 sg13g2_a21oi_1 _20454_ (.A1(net1224),
    .A2(net4422),
    .Y(_13249_),
    .B1(_13248_));
 sg13g2_nand2_1 _20455_ (.Y(_13250_),
    .A(net1612),
    .B(net4126));
 sg13g2_o21ai_1 _20456_ (.B1(_13250_),
    .Y(_00158_),
    .A1(net4124),
    .A2(_13249_));
 sg13g2_and2_1 _20457_ (.A(net1364),
    .B(net4487),
    .X(_13251_));
 sg13g2_a21oi_1 _20458_ (.A1(net1431),
    .A2(net4421),
    .Y(_13252_),
    .B1(_13251_));
 sg13g2_nand2_1 _20459_ (.Y(_13253_),
    .A(net1496),
    .B(net4127));
 sg13g2_o21ai_1 _20460_ (.B1(_13253_),
    .Y(_00159_),
    .A1(net4127),
    .A2(_13252_));
 sg13g2_and2_1 _20461_ (.A(net1517),
    .B(net4489),
    .X(_13254_));
 sg13g2_a21oi_1 _20462_ (.A1(\inv_result[149] ),
    .A2(net4422),
    .Y(_13255_),
    .B1(_13254_));
 sg13g2_nand2_1 _20463_ (.Y(_13256_),
    .A(net1524),
    .B(net4126));
 sg13g2_o21ai_1 _20464_ (.B1(_13256_),
    .Y(_00160_),
    .A1(net4127),
    .A2(_13255_));
 sg13g2_and2_1 _20465_ (.A(net1592),
    .B(net4492),
    .X(_13257_));
 sg13g2_a21oi_1 _20466_ (.A1(net1187),
    .A2(net4425),
    .Y(_13258_),
    .B1(_13257_));
 sg13g2_nand2_1 _20467_ (.Y(_13259_),
    .A(net1917),
    .B(net4129));
 sg13g2_o21ai_1 _20468_ (.B1(_13259_),
    .Y(_00161_),
    .A1(net4129),
    .A2(_13258_));
 sg13g2_and2_1 _20469_ (.A(\shift_reg[143] ),
    .B(net4488),
    .X(_13260_));
 sg13g2_a21oi_1 _20470_ (.A1(net1506),
    .A2(net4422),
    .Y(_13261_),
    .B1(_13260_));
 sg13g2_nand2_1 _20471_ (.Y(_13262_),
    .A(net1600),
    .B(net4126));
 sg13g2_o21ai_1 _20472_ (.B1(_13262_),
    .Y(_00162_),
    .A1(net4126),
    .A2(_13261_));
 sg13g2_and2_1 _20473_ (.A(net1536),
    .B(net4488),
    .X(_13263_));
 sg13g2_a21oi_1 _20474_ (.A1(net1484),
    .A2(net4422),
    .Y(_13264_),
    .B1(_13263_));
 sg13g2_nand2_1 _20475_ (.Y(_13265_),
    .A(net2439),
    .B(net4128));
 sg13g2_o21ai_1 _20476_ (.B1(_13265_),
    .Y(_00163_),
    .A1(net4128),
    .A2(_13264_));
 sg13g2_nor2_1 _20477_ (.A(_11016_),
    .B(net4490),
    .Y(_13266_));
 sg13g2_a21oi_1 _20478_ (.A1(net1489),
    .A2(net4491),
    .Y(_13267_),
    .B1(_13266_));
 sg13g2_nand2_1 _20479_ (.Y(_13268_),
    .A(net1945),
    .B(net4128));
 sg13g2_o21ai_1 _20480_ (.B1(_13268_),
    .Y(_00164_),
    .A1(net4128),
    .A2(_13267_));
 sg13g2_and2_1 _20481_ (.A(\shift_reg[146] ),
    .B(net4490),
    .X(_13269_));
 sg13g2_a21oi_1 _20482_ (.A1(net1613),
    .A2(net4423),
    .Y(_13270_),
    .B1(_13269_));
 sg13g2_nand2_1 _20483_ (.Y(_13271_),
    .A(net1657),
    .B(net4135));
 sg13g2_o21ai_1 _20484_ (.B1(_13271_),
    .Y(_00165_),
    .A1(net4129),
    .A2(_13270_));
 sg13g2_nor2_1 _20485_ (.A(_11017_),
    .B(net4490),
    .Y(_13272_));
 sg13g2_a21oi_1 _20486_ (.A1(net1612),
    .A2(net4491),
    .Y(_13273_),
    .B1(_13272_));
 sg13g2_nand2_1 _20487_ (.Y(_13274_),
    .A(net1644),
    .B(net4128));
 sg13g2_o21ai_1 _20488_ (.B1(_13274_),
    .Y(_00166_),
    .A1(net4128),
    .A2(_13273_));
 sg13g2_and2_1 _20489_ (.A(net1496),
    .B(net4492),
    .X(_13275_));
 sg13g2_a21oi_1 _20490_ (.A1(net1759),
    .A2(net4424),
    .Y(_13276_),
    .B1(_13275_));
 sg13g2_nand2_1 _20491_ (.Y(_13277_),
    .A(net2442),
    .B(net4129));
 sg13g2_o21ai_1 _20492_ (.B1(_13277_),
    .Y(_00167_),
    .A1(net4129),
    .A2(_13276_));
 sg13g2_and2_1 _20493_ (.A(net1524),
    .B(net4491),
    .X(_13278_));
 sg13g2_a21oi_1 _20494_ (.A1(\inv_result[157] ),
    .A2(net4424),
    .Y(_13279_),
    .B1(_13278_));
 sg13g2_nand2_1 _20495_ (.Y(_13280_),
    .A(net1545),
    .B(net4139));
 sg13g2_o21ai_1 _20496_ (.B1(_13280_),
    .Y(_00168_),
    .A1(net4139),
    .A2(_13279_));
 sg13g2_and2_1 _20497_ (.A(\shift_reg[150] ),
    .B(net4490),
    .X(_13281_));
 sg13g2_a21oi_1 _20498_ (.A1(net1457),
    .A2(net4423),
    .Y(_13282_),
    .B1(_13281_));
 sg13g2_nand2_1 _20499_ (.Y(_13283_),
    .A(net1673),
    .B(net4135));
 sg13g2_o21ai_1 _20500_ (.B1(_13283_),
    .Y(_00169_),
    .A1(net4136),
    .A2(_13282_));
 sg13g2_and2_1 _20501_ (.A(net1600),
    .B(net4491),
    .X(_13284_));
 sg13g2_a21oi_1 _20502_ (.A1(net1409),
    .A2(net4423),
    .Y(_13285_),
    .B1(_13284_));
 sg13g2_nand2_1 _20503_ (.Y(_13286_),
    .A(net1679),
    .B(net4139));
 sg13g2_o21ai_1 _20504_ (.B1(_13286_),
    .Y(_00170_),
    .A1(net4139),
    .A2(_13285_));
 sg13g2_and2_1 _20505_ (.A(\shift_reg[152] ),
    .B(net4491),
    .X(_13287_));
 sg13g2_a21oi_1 _20506_ (.A1(\inv_result[160] ),
    .A2(net4423),
    .Y(_13288_),
    .B1(_13287_));
 sg13g2_nand2_1 _20507_ (.Y(_13289_),
    .A(net1276),
    .B(net4136));
 sg13g2_o21ai_1 _20508_ (.B1(_13289_),
    .Y(_00171_),
    .A1(net4136),
    .A2(_13288_));
 sg13g2_and2_1 _20509_ (.A(\shift_reg[153] ),
    .B(net4496),
    .X(_13290_));
 sg13g2_a21oi_1 _20510_ (.A1(\inv_result[161] ),
    .A2(net4423),
    .Y(_13291_),
    .B1(_13290_));
 sg13g2_nand2_1 _20511_ (.Y(_13292_),
    .A(net1365),
    .B(net4137));
 sg13g2_o21ai_1 _20512_ (.B1(_13292_),
    .Y(_00172_),
    .A1(net4137),
    .A2(_13291_));
 sg13g2_and2_1 _20513_ (.A(\shift_reg[154] ),
    .B(net4495),
    .X(_13293_));
 sg13g2_a21oi_1 _20514_ (.A1(\inv_result[162] ),
    .A2(net4427),
    .Y(_13294_),
    .B1(_13293_));
 sg13g2_nand2_1 _20515_ (.Y(_13295_),
    .A(net1312),
    .B(net4135));
 sg13g2_o21ai_1 _20516_ (.B1(_13295_),
    .Y(_00173_),
    .A1(net4135),
    .A2(_13294_));
 sg13g2_nor2_1 _20517_ (.A(_11018_),
    .B(net4491),
    .Y(_13296_));
 sg13g2_a21oi_1 _20518_ (.A1(net1644),
    .A2(net4495),
    .Y(_13297_),
    .B1(_13296_));
 sg13g2_nand2_1 _20519_ (.Y(_13298_),
    .A(net1702),
    .B(net4135));
 sg13g2_o21ai_1 _20520_ (.B1(_13298_),
    .Y(_00174_),
    .A1(net4136),
    .A2(_13297_));
 sg13g2_and2_1 _20521_ (.A(\shift_reg[156] ),
    .B(net4495),
    .X(_13299_));
 sg13g2_a21oi_1 _20522_ (.A1(\inv_result[164] ),
    .A2(net4423),
    .Y(_13300_),
    .B1(_13299_));
 sg13g2_nand2_1 _20523_ (.Y(_13301_),
    .A(net1243),
    .B(net4135));
 sg13g2_o21ai_1 _20524_ (.B1(_13301_),
    .Y(_00175_),
    .A1(net4135),
    .A2(_13300_));
 sg13g2_and2_1 _20525_ (.A(net1545),
    .B(net4496),
    .X(_13302_));
 sg13g2_a21oi_1 _20526_ (.A1(\inv_result[165] ),
    .A2(net4427),
    .Y(_13303_),
    .B1(_13302_));
 sg13g2_nand2_1 _20527_ (.Y(_13304_),
    .A(net1651),
    .B(net4133));
 sg13g2_o21ai_1 _20528_ (.B1(_13304_),
    .Y(_00176_),
    .A1(net4133),
    .A2(_13303_));
 sg13g2_and2_1 _20529_ (.A(\shift_reg[158] ),
    .B(net4495),
    .X(_13305_));
 sg13g2_a21oi_1 _20530_ (.A1(net1096),
    .A2(net4427),
    .Y(_13306_),
    .B1(_13305_));
 sg13g2_nand2_1 _20531_ (.Y(_13307_),
    .A(net1269),
    .B(net4137));
 sg13g2_o21ai_1 _20532_ (.B1(_13307_),
    .Y(_00177_),
    .A1(net4135),
    .A2(_13306_));
 sg13g2_and2_1 _20533_ (.A(\shift_reg[159] ),
    .B(net4493),
    .X(_13308_));
 sg13g2_a21oi_1 _20534_ (.A1(\inv_result[167] ),
    .A2(net4426),
    .Y(_13309_),
    .B1(_13308_));
 sg13g2_nand2_1 _20535_ (.Y(_13310_),
    .A(net1435),
    .B(net4132));
 sg13g2_o21ai_1 _20536_ (.B1(_13310_),
    .Y(_00178_),
    .A1(net4132),
    .A2(_13309_));
 sg13g2_and2_1 _20537_ (.A(net1276),
    .B(net4495),
    .X(_13311_));
 sg13g2_a21oi_1 _20538_ (.A1(net1240),
    .A2(net4426),
    .Y(_13312_),
    .B1(_13311_));
 sg13g2_nand2_1 _20539_ (.Y(_13313_),
    .A(net1554),
    .B(net4132));
 sg13g2_o21ai_1 _20540_ (.B1(_13313_),
    .Y(_00179_),
    .A1(net4132),
    .A2(_13312_));
 sg13g2_and2_1 _20541_ (.A(net1365),
    .B(net4495),
    .X(_13314_));
 sg13g2_a21oi_1 _20542_ (.A1(\inv_result[169] ),
    .A2(net4426),
    .Y(_13315_),
    .B1(_13314_));
 sg13g2_nand2_1 _20543_ (.Y(_13316_),
    .A(net1441),
    .B(net4132));
 sg13g2_o21ai_1 _20544_ (.B1(_13316_),
    .Y(_00180_),
    .A1(net4132),
    .A2(_13315_));
 sg13g2_and2_1 _20545_ (.A(net1312),
    .B(net4493),
    .X(_13317_));
 sg13g2_a21oi_1 _20546_ (.A1(net1093),
    .A2(net4426),
    .Y(_13318_),
    .B1(_13317_));
 sg13g2_nand2_1 _20547_ (.Y(_13319_),
    .A(net1333),
    .B(net4131));
 sg13g2_o21ai_1 _20548_ (.B1(_13319_),
    .Y(_00181_),
    .A1(net4130),
    .A2(_13318_));
 sg13g2_nor2_1 _20549_ (.A(_11019_),
    .B(net4493),
    .Y(_13320_));
 sg13g2_a21oi_1 _20550_ (.A1(\shift_reg[163] ),
    .A2(net4493),
    .Y(_13321_),
    .B1(_13320_));
 sg13g2_nand2_1 _20551_ (.Y(_13322_),
    .A(net1406),
    .B(net4131));
 sg13g2_o21ai_1 _20552_ (.B1(_13322_),
    .Y(_00182_),
    .A1(net4131),
    .A2(_13321_));
 sg13g2_and2_1 _20553_ (.A(net1243),
    .B(net4495),
    .X(_13323_));
 sg13g2_a21oi_1 _20554_ (.A1(net1085),
    .A2(net4427),
    .Y(_13324_),
    .B1(_13323_));
 sg13g2_nand2_1 _20555_ (.Y(_13325_),
    .A(net1726),
    .B(net4132));
 sg13g2_o21ai_1 _20556_ (.B1(_13325_),
    .Y(_00183_),
    .A1(net4132),
    .A2(_13324_));
 sg13g2_nor2_1 _20557_ (.A(_11020_),
    .B(net4494),
    .Y(_13326_));
 sg13g2_a21oi_1 _20558_ (.A1(\shift_reg[165] ),
    .A2(net4493),
    .Y(_13327_),
    .B1(_13326_));
 sg13g2_nand2_1 _20559_ (.Y(_13328_),
    .A(net1498),
    .B(net4130));
 sg13g2_o21ai_1 _20560_ (.B1(_13328_),
    .Y(_00184_),
    .A1(net4130),
    .A2(_13327_));
 sg13g2_and2_1 _20561_ (.A(net1269),
    .B(net4493),
    .X(_13329_));
 sg13g2_a21oi_1 _20562_ (.A1(net1308),
    .A2(net4427),
    .Y(_13330_),
    .B1(_13329_));
 sg13g2_nand2_1 _20563_ (.Y(_13331_),
    .A(net1727),
    .B(net4130));
 sg13g2_o21ai_1 _20564_ (.B1(_13331_),
    .Y(_00185_),
    .A1(net4130),
    .A2(_13330_));
 sg13g2_and2_1 _20565_ (.A(\shift_reg[167] ),
    .B(net4493),
    .X(_13332_));
 sg13g2_a21oi_1 _20566_ (.A1(\inv_result[175] ),
    .A2(net4426),
    .Y(_13333_),
    .B1(_13332_));
 sg13g2_nand2_1 _20567_ (.Y(_13334_),
    .A(net1304),
    .B(net4117));
 sg13g2_o21ai_1 _20568_ (.B1(_13334_),
    .Y(_00186_),
    .A1(net4117),
    .A2(_13333_));
 sg13g2_and2_1 _20569_ (.A(\shift_reg[168] ),
    .B(net4493),
    .X(_13335_));
 sg13g2_a21oi_1 _20570_ (.A1(\inv_result[176] ),
    .A2(net4420),
    .Y(_13336_),
    .B1(_13335_));
 sg13g2_nand2_1 _20571_ (.Y(_13337_),
    .A(net1503),
    .B(net4119));
 sg13g2_o21ai_1 _20572_ (.B1(_13337_),
    .Y(_00187_),
    .A1(net4117),
    .A2(_13336_));
 sg13g2_and2_1 _20573_ (.A(\shift_reg[169] ),
    .B(net4485),
    .X(_13338_));
 sg13g2_a21oi_1 _20574_ (.A1(\inv_result[177] ),
    .A2(net4419),
    .Y(_13339_),
    .B1(_13338_));
 sg13g2_nand2_1 _20575_ (.Y(_13340_),
    .A(net1272),
    .B(net4119));
 sg13g2_o21ai_1 _20576_ (.B1(_13340_),
    .Y(_00188_),
    .A1(net4120),
    .A2(_13339_));
 sg13g2_and2_1 _20577_ (.A(net1333),
    .B(net4484),
    .X(_13341_));
 sg13g2_a21oi_1 _20578_ (.A1(net1543),
    .A2(net4419),
    .Y(_13342_),
    .B1(_13341_));
 sg13g2_nand2_1 _20579_ (.Y(_13343_),
    .A(net1809),
    .B(net4119));
 sg13g2_o21ai_1 _20580_ (.B1(_13343_),
    .Y(_00189_),
    .A1(net4117),
    .A2(_13342_));
 sg13g2_nor2_1 _20581_ (.A(_11021_),
    .B(net4484),
    .Y(_13344_));
 sg13g2_a21oi_1 _20582_ (.A1(net1406),
    .A2(net4484),
    .Y(_13345_),
    .B1(_13344_));
 sg13g2_nand2_1 _20583_ (.Y(_13346_),
    .A(net1675),
    .B(net4116));
 sg13g2_o21ai_1 _20584_ (.B1(_13346_),
    .Y(_00190_),
    .A1(net4116),
    .A2(_13345_));
 sg13g2_and2_1 _20585_ (.A(\shift_reg[172] ),
    .B(net4484),
    .X(_13347_));
 sg13g2_a21oi_1 _20586_ (.A1(net1410),
    .A2(net4419),
    .Y(_13348_),
    .B1(_13347_));
 sg13g2_nand2_1 _20587_ (.Y(_13349_),
    .A(net1616),
    .B(net4117));
 sg13g2_o21ai_1 _20588_ (.B1(_13349_),
    .Y(_00191_),
    .A1(net4117),
    .A2(_13348_));
 sg13g2_nor2_1 _20589_ (.A(_11022_),
    .B(net4484),
    .Y(_13350_));
 sg13g2_a21oi_1 _20590_ (.A1(\shift_reg[173] ),
    .A2(net4484),
    .Y(_13351_),
    .B1(_13350_));
 sg13g2_nand2_1 _20591_ (.Y(_13352_),
    .A(net1422),
    .B(net4115));
 sg13g2_o21ai_1 _20592_ (.B1(_13352_),
    .Y(_00192_),
    .A1(net4115),
    .A2(_13351_));
 sg13g2_and2_1 _20593_ (.A(\shift_reg[174] ),
    .B(net4485),
    .X(_13353_));
 sg13g2_a21oi_1 _20594_ (.A1(net1416),
    .A2(net4419),
    .Y(_13354_),
    .B1(_13353_));
 sg13g2_nand2_1 _20595_ (.Y(_13355_),
    .A(net1596),
    .B(net4115));
 sg13g2_o21ai_1 _20596_ (.B1(_13355_),
    .Y(_00193_),
    .A1(net4116),
    .A2(_13354_));
 sg13g2_and2_1 _20597_ (.A(\shift_reg[175] ),
    .B(net4484),
    .X(_13356_));
 sg13g2_a21oi_1 _20598_ (.A1(\inv_result[183] ),
    .A2(net4419),
    .Y(_13357_),
    .B1(_13356_));
 sg13g2_nand2_1 _20599_ (.Y(_13358_),
    .A(net1167),
    .B(net4115));
 sg13g2_o21ai_1 _20600_ (.B1(_13358_),
    .Y(_00194_),
    .A1(net4115),
    .A2(_13357_));
 sg13g2_and2_1 _20601_ (.A(net1503),
    .B(net4486),
    .X(_13359_));
 sg13g2_a21oi_1 _20602_ (.A1(net1338),
    .A2(net4428),
    .Y(_13360_),
    .B1(_13359_));
 sg13g2_nand2_1 _20603_ (.Y(_13361_),
    .A(net2367),
    .B(net4113));
 sg13g2_o21ai_1 _20604_ (.B1(_13361_),
    .Y(_00195_),
    .A1(net4113),
    .A2(_13360_));
 sg13g2_and2_1 _20605_ (.A(net1272),
    .B(net4486),
    .X(_13362_));
 sg13g2_a21oi_1 _20606_ (.A1(net1293),
    .A2(net4417),
    .Y(_13363_),
    .B1(_13362_));
 sg13g2_nand2_1 _20607_ (.Y(_13364_),
    .A(net2132),
    .B(net4112));
 sg13g2_o21ai_1 _20608_ (.B1(_13364_),
    .Y(_00196_),
    .A1(net4112),
    .A2(_13363_));
 sg13g2_and2_1 _20609_ (.A(\shift_reg[178] ),
    .B(net4483),
    .X(_13365_));
 sg13g2_a21oi_1 _20610_ (.A1(net1535),
    .A2(net4416),
    .Y(_13366_),
    .B1(_13365_));
 sg13g2_nand2_1 _20611_ (.Y(_13367_),
    .A(net1687),
    .B(net4111));
 sg13g2_o21ai_1 _20612_ (.B1(_13367_),
    .Y(_00197_),
    .A1(net4111),
    .A2(_13366_));
 sg13g2_nor2_1 _20613_ (.A(_11023_),
    .B(net4482),
    .Y(_13368_));
 sg13g2_a21oi_1 _20614_ (.A1(net1675),
    .A2(net4483),
    .Y(_13369_),
    .B1(_13368_));
 sg13g2_nand2_1 _20615_ (.Y(_13370_),
    .A(net1714),
    .B(net4113));
 sg13g2_o21ai_1 _20616_ (.B1(_13370_),
    .Y(_00198_),
    .A1(net4113),
    .A2(_13369_));
 sg13g2_and2_1 _20617_ (.A(\shift_reg[180] ),
    .B(net4481),
    .X(_13371_));
 sg13g2_a21oi_1 _20618_ (.A1(net1467),
    .A2(net4416),
    .Y(_13372_),
    .B1(_13371_));
 sg13g2_nand2_1 _20619_ (.Y(_13373_),
    .A(net1513),
    .B(net4107));
 sg13g2_o21ai_1 _20620_ (.B1(_13373_),
    .Y(_00199_),
    .A1(net4107),
    .A2(_13372_));
 sg13g2_nor2_1 _20621_ (.A(_11024_),
    .B(net4482),
    .Y(_13374_));
 sg13g2_a21oi_1 _20622_ (.A1(net1422),
    .A2(net4482),
    .Y(_13375_),
    .B1(_13374_));
 sg13g2_nand2_1 _20623_ (.Y(_13376_),
    .A(net1841),
    .B(net4108));
 sg13g2_o21ai_1 _20624_ (.B1(_13376_),
    .Y(_00200_),
    .A1(net4107),
    .A2(_13375_));
 sg13g2_and2_1 _20625_ (.A(net1596),
    .B(net4481),
    .X(_13377_));
 sg13g2_a21oi_1 _20626_ (.A1(net1290),
    .A2(net4417),
    .Y(_13378_),
    .B1(_13377_));
 sg13g2_nand2_1 _20627_ (.Y(_13379_),
    .A(net1843),
    .B(net4107));
 sg13g2_o21ai_1 _20628_ (.B1(_13379_),
    .Y(_00201_),
    .A1(net4107),
    .A2(_13378_));
 sg13g2_and2_1 _20629_ (.A(net1167),
    .B(net4482),
    .X(_13380_));
 sg13g2_a21oi_2 _20630_ (.B1(_13380_),
    .Y(_13381_),
    .A2(net4417),
    .A1(\inv_result[191] ));
 sg13g2_nand2_1 _20631_ (.Y(_13382_),
    .A(net1345),
    .B(net4108));
 sg13g2_o21ai_1 _20632_ (.B1(_13382_),
    .Y(_00202_),
    .A1(net4108),
    .A2(_13381_));
 sg13g2_nor2_1 _20633_ (.A(_11025_),
    .B(net4473),
    .Y(_13383_));
 sg13g2_a21oi_1 _20634_ (.A1(\shift_reg[184] ),
    .A2(net4473),
    .Y(_13384_),
    .B1(_13383_));
 sg13g2_nand2_1 _20635_ (.Y(_13385_),
    .A(net1659),
    .B(net4097));
 sg13g2_o21ai_1 _20636_ (.B1(_13385_),
    .Y(_00203_),
    .A1(net4097),
    .A2(_13384_));
 sg13g2_and2_1 _20637_ (.A(\shift_reg[185] ),
    .B(net4477),
    .X(_13386_));
 sg13g2_a21oi_1 _20638_ (.A1(net1084),
    .A2(net4412),
    .Y(_13387_),
    .B1(_13386_));
 sg13g2_nand2_1 _20639_ (.Y(_13388_),
    .A(net1280),
    .B(net4096));
 sg13g2_o21ai_1 _20640_ (.B1(_13388_),
    .Y(_00204_),
    .A1(net4096),
    .A2(_13387_));
 sg13g2_and2_1 _20641_ (.A(\shift_reg[186] ),
    .B(net4479),
    .X(_13389_));
 sg13g2_a21oi_1 _20642_ (.A1(\inv_result[194] ),
    .A2(net4413),
    .Y(_13390_),
    .B1(_13389_));
 sg13g2_nand2_1 _20643_ (.Y(_13391_),
    .A(net1398),
    .B(net4094));
 sg13g2_o21ai_1 _20644_ (.B1(_13391_),
    .Y(_00205_),
    .A1(net4094),
    .A2(_13390_));
 sg13g2_and2_1 _20645_ (.A(net1714),
    .B(net4480),
    .X(_13392_));
 sg13g2_a21oi_1 _20646_ (.A1(net1145),
    .A2(net4413),
    .Y(_13393_),
    .B1(_13392_));
 sg13g2_nand2_1 _20647_ (.Y(_13394_),
    .A(net1763),
    .B(net4094));
 sg13g2_o21ai_1 _20648_ (.B1(_13394_),
    .Y(_00206_),
    .A1(net4094),
    .A2(_13393_));
 sg13g2_and2_1 _20649_ (.A(net1513),
    .B(net4478),
    .X(_13395_));
 sg13g2_a21oi_1 _20650_ (.A1(net1497),
    .A2(net4413),
    .Y(_13396_),
    .B1(_13395_));
 sg13g2_nand2_1 _20651_ (.Y(_13397_),
    .A(net1854),
    .B(net4094));
 sg13g2_o21ai_1 _20652_ (.B1(_13397_),
    .Y(_00207_),
    .A1(net4094),
    .A2(_13396_));
 sg13g2_and2_1 _20653_ (.A(net1841),
    .B(net4476),
    .X(_13398_));
 sg13g2_a21oi_1 _20654_ (.A1(\inv_result[197] ),
    .A2(net4413),
    .Y(_13399_),
    .B1(_13398_));
 sg13g2_nand2_1 _20655_ (.Y(_13400_),
    .A(net2057),
    .B(net4104));
 sg13g2_o21ai_1 _20656_ (.B1(_13400_),
    .Y(_00208_),
    .A1(net4104),
    .A2(_13399_));
 sg13g2_and2_1 _20657_ (.A(net1843),
    .B(net4474),
    .X(_13401_));
 sg13g2_a21oi_1 _20658_ (.A1(net1349),
    .A2(net4413),
    .Y(_13402_),
    .B1(_13401_));
 sg13g2_nand2_1 _20659_ (.Y(_13403_),
    .A(net1859),
    .B(net4094));
 sg13g2_o21ai_1 _20660_ (.B1(_13403_),
    .Y(_00209_),
    .A1(net4094),
    .A2(_13402_));
 sg13g2_and2_1 _20661_ (.A(net1345),
    .B(net4475),
    .X(_13404_));
 sg13g2_a21oi_1 _20662_ (.A1(net1654),
    .A2(net4411),
    .Y(_13405_),
    .B1(_13404_));
 sg13g2_nand2_1 _20663_ (.Y(_13406_),
    .A(net2432),
    .B(net4100));
 sg13g2_o21ai_1 _20664_ (.B1(_13406_),
    .Y(_00210_),
    .A1(net4100),
    .A2(_13405_));
 sg13g2_and2_1 _20665_ (.A(net1659),
    .B(net4468),
    .X(_13407_));
 sg13g2_a21oi_1 _20666_ (.A1(net1374),
    .A2(net4405),
    .Y(_13408_),
    .B1(_13407_));
 sg13g2_nand2_1 _20667_ (.Y(_13409_),
    .A(net1808),
    .B(net4087));
 sg13g2_o21ai_1 _20668_ (.B1(_13409_),
    .Y(_00211_),
    .A1(net4087),
    .A2(_13408_));
 sg13g2_and2_1 _20669_ (.A(net1280),
    .B(net4469),
    .X(_13410_));
 sg13g2_a21oi_1 _20670_ (.A1(\inv_result[201] ),
    .A2(net4405),
    .Y(_13411_),
    .B1(_13410_));
 sg13g2_nand2_1 _20671_ (.Y(_13412_),
    .A(net1567),
    .B(net4086));
 sg13g2_o21ai_1 _20672_ (.B1(_13412_),
    .Y(_00212_),
    .A1(net4086),
    .A2(_13411_));
 sg13g2_and2_1 _20673_ (.A(\shift_reg[194] ),
    .B(net4468),
    .X(_13413_));
 sg13g2_a21oi_1 _20674_ (.A1(net1081),
    .A2(net4405),
    .Y(_13414_),
    .B1(_13413_));
 sg13g2_nand2_1 _20675_ (.Y(_13415_),
    .A(net1357),
    .B(net4086));
 sg13g2_o21ai_1 _20676_ (.B1(_13415_),
    .Y(_00213_),
    .A1(net4086),
    .A2(_13414_));
 sg13g2_nor2_1 _20677_ (.A(_11026_),
    .B(net4468),
    .Y(_13416_));
 sg13g2_a21oi_1 _20678_ (.A1(\shift_reg[195] ),
    .A2(net4468),
    .Y(_13417_),
    .B1(_13416_));
 sg13g2_nand2_1 _20679_ (.Y(_13418_),
    .A(net1200),
    .B(net4086));
 sg13g2_o21ai_1 _20680_ (.B1(_13418_),
    .Y(_00214_),
    .A1(net4086),
    .A2(_13417_));
 sg13g2_and2_1 _20681_ (.A(\shift_reg[196] ),
    .B(net4467),
    .X(_13419_));
 sg13g2_a21oi_1 _20682_ (.A1(\inv_result[204] ),
    .A2(net4404),
    .Y(_13420_),
    .B1(_13419_));
 sg13g2_nand2_1 _20683_ (.Y(_13421_),
    .A(net1315),
    .B(net4086));
 sg13g2_o21ai_1 _20684_ (.B1(_13421_),
    .Y(_00215_),
    .A1(net4086),
    .A2(_13420_));
 sg13g2_nor2_1 _20685_ (.A(_11027_),
    .B(net4467),
    .Y(_13422_));
 sg13g2_a21oi_1 _20686_ (.A1(\shift_reg[197] ),
    .A2(net4467),
    .Y(_13423_),
    .B1(_13422_));
 sg13g2_nand2_1 _20687_ (.Y(_13424_),
    .A(net1424),
    .B(net4084));
 sg13g2_o21ai_1 _20688_ (.B1(_13424_),
    .Y(_00216_),
    .A1(net4084),
    .A2(_13423_));
 sg13g2_and2_1 _20689_ (.A(\shift_reg[198] ),
    .B(net4466),
    .X(_13425_));
 sg13g2_a21oi_1 _20690_ (.A1(net1586),
    .A2(net4404),
    .Y(_13426_),
    .B1(_13425_));
 sg13g2_nand2_1 _20691_ (.Y(_13427_),
    .A(net1805),
    .B(net4085));
 sg13g2_o21ai_1 _20692_ (.B1(_13427_),
    .Y(_00217_),
    .A1(net4085),
    .A2(_13426_));
 sg13g2_and2_1 _20693_ (.A(\shift_reg[199] ),
    .B(net4470),
    .X(_13428_));
 sg13g2_a21oi_1 _20694_ (.A1(\inv_result[207] ),
    .A2(net4404),
    .Y(_13429_),
    .B1(_13428_));
 sg13g2_nand2_1 _20695_ (.Y(_13430_),
    .A(net1323),
    .B(net4085));
 sg13g2_o21ai_1 _20696_ (.B1(_13430_),
    .Y(_00218_),
    .A1(net4085),
    .A2(_13429_));
 sg13g2_and2_1 _20697_ (.A(\shift_reg[200] ),
    .B(net4466),
    .X(_13431_));
 sg13g2_a21oi_1 _20698_ (.A1(\inv_result[208] ),
    .A2(net4404),
    .Y(_13432_),
    .B1(_13431_));
 sg13g2_nand2_1 _20699_ (.Y(_13433_),
    .A(net1371),
    .B(net4082));
 sg13g2_o21ai_1 _20700_ (.B1(_13433_),
    .Y(_00219_),
    .A1(net4082),
    .A2(_13432_));
 sg13g2_and2_1 _20701_ (.A(\shift_reg[201] ),
    .B(net4466),
    .X(_13434_));
 sg13g2_a21oi_2 _20702_ (.B1(_13434_),
    .Y(_13435_),
    .A2(net4404),
    .A1(\inv_result[209] ));
 sg13g2_nand2_1 _20703_ (.Y(_13436_),
    .A(net1164),
    .B(net4074));
 sg13g2_o21ai_1 _20704_ (.B1(_13436_),
    .Y(_00220_),
    .A1(net4074),
    .A2(_13435_));
 sg13g2_and2_1 _20705_ (.A(net1357),
    .B(net4466),
    .X(_13437_));
 sg13g2_a21oi_1 _20706_ (.A1(net1092),
    .A2(net4404),
    .Y(_13438_),
    .B1(_13437_));
 sg13g2_nand2_1 _20707_ (.Y(_13439_),
    .A(net1557),
    .B(net4082));
 sg13g2_o21ai_1 _20708_ (.B1(_13439_),
    .Y(_00221_),
    .A1(net4082),
    .A2(_13438_));
 sg13g2_nor2_1 _20709_ (.A(_11028_),
    .B(net4467),
    .Y(_13440_));
 sg13g2_a21oi_1 _20710_ (.A1(net1200),
    .A2(net4467),
    .Y(_13441_),
    .B1(_13440_));
 sg13g2_nand2_1 _20711_ (.Y(_13442_),
    .A(net1494),
    .B(net4085));
 sg13g2_o21ai_1 _20712_ (.B1(_13442_),
    .Y(_00222_),
    .A1(net4085),
    .A2(_13441_));
 sg13g2_and2_1 _20713_ (.A(net1315),
    .B(net4466),
    .X(_13443_));
 sg13g2_a21oi_1 _20714_ (.A1(net1335),
    .A2(net4404),
    .Y(_13444_),
    .B1(_13443_));
 sg13g2_nand2_1 _20715_ (.Y(_13445_),
    .A(net1618),
    .B(net4083));
 sg13g2_o21ai_1 _20716_ (.B1(_13445_),
    .Y(_00223_),
    .A1(net4083),
    .A2(_13444_));
 sg13g2_nor2_1 _20717_ (.A(_11029_),
    .B(net4468),
    .Y(_13446_));
 sg13g2_a21oi_1 _20718_ (.A1(\shift_reg[205] ),
    .A2(net4466),
    .Y(_13447_),
    .B1(_13446_));
 sg13g2_nand2_1 _20719_ (.Y(_13448_),
    .A(net1182),
    .B(net4084));
 sg13g2_o21ai_1 _20720_ (.B1(_13448_),
    .Y(_00224_),
    .A1(net4084),
    .A2(_13447_));
 sg13g2_and2_1 _20721_ (.A(\shift_reg[206] ),
    .B(net4466),
    .X(_13449_));
 sg13g2_a21oi_1 _20722_ (.A1(\inv_result[214] ),
    .A2(net4405),
    .Y(_13450_),
    .B1(_13449_));
 sg13g2_nand2_1 _20723_ (.Y(_13451_),
    .A(net1306),
    .B(net4083));
 sg13g2_o21ai_1 _20724_ (.B1(_13451_),
    .Y(_00225_),
    .A1(net4083),
    .A2(_13450_));
 sg13g2_and2_1 _20725_ (.A(\shift_reg[207] ),
    .B(net4466),
    .X(_13452_));
 sg13g2_a21oi_1 _20726_ (.A1(\inv_result[215] ),
    .A2(net4404),
    .Y(_13453_),
    .B1(_13452_));
 sg13g2_nand2_1 _20727_ (.Y(_13454_),
    .A(net1136),
    .B(net4075));
 sg13g2_o21ai_1 _20728_ (.B1(_13454_),
    .Y(_00226_),
    .A1(net4074),
    .A2(_13453_));
 sg13g2_and2_1 _20729_ (.A(\shift_reg[208] ),
    .B(net4462),
    .X(_13455_));
 sg13g2_a21oi_2 _20730_ (.B1(_13455_),
    .Y(_13456_),
    .A2(net4403),
    .A1(\inv_result[216] ));
 sg13g2_nand2_1 _20731_ (.Y(_13457_),
    .A(net1125),
    .B(net4073));
 sg13g2_o21ai_1 _20732_ (.B1(_13457_),
    .Y(_00227_),
    .A1(net4073),
    .A2(_13456_));
 sg13g2_and2_1 _20733_ (.A(net1164),
    .B(net4461),
    .X(_13458_));
 sg13g2_a21oi_1 _20734_ (.A1(net1392),
    .A2(net4403),
    .Y(_13459_),
    .B1(_13458_));
 sg13g2_nand2_1 _20735_ (.Y(_13460_),
    .A(net1443),
    .B(net4074));
 sg13g2_o21ai_1 _20736_ (.B1(_13460_),
    .Y(_00228_),
    .A1(net4074),
    .A2(_13459_));
 sg13g2_and2_1 _20737_ (.A(net1557),
    .B(net4461),
    .X(_13461_));
 sg13g2_a21oi_1 _20738_ (.A1(net1322),
    .A2(net4399),
    .Y(_13462_),
    .B1(_13461_));
 sg13g2_nand2_1 _20739_ (.Y(_13463_),
    .A(net1642),
    .B(net4074));
 sg13g2_o21ai_1 _20740_ (.B1(_13463_),
    .Y(_00229_),
    .A1(net4074),
    .A2(_13462_));
 sg13g2_and2_1 _20741_ (.A(net1494),
    .B(net4462),
    .X(_13464_));
 sg13g2_a21oi_1 _20742_ (.A1(\inv_result[219] ),
    .A2(net4399),
    .Y(_13465_),
    .B1(_13464_));
 sg13g2_nand2_1 _20743_ (.Y(_13466_),
    .A(net1587),
    .B(net4075));
 sg13g2_o21ai_1 _20744_ (.B1(_13466_),
    .Y(_00230_),
    .A1(net4074),
    .A2(_13465_));
 sg13g2_and2_1 _20745_ (.A(net1618),
    .B(net4462),
    .X(_13467_));
 sg13g2_a21oi_1 _20746_ (.A1(net1598),
    .A2(net4399),
    .Y(_13468_),
    .B1(_13467_));
 sg13g2_nand2_1 _20747_ (.Y(_13469_),
    .A(net1730),
    .B(net4082));
 sg13g2_o21ai_1 _20748_ (.B1(_13469_),
    .Y(_00231_),
    .A1(net4082),
    .A2(_13468_));
 sg13g2_nor2_1 _20749_ (.A(_11030_),
    .B(net4462),
    .Y(_13470_));
 sg13g2_a21oi_1 _20750_ (.A1(net1182),
    .A2(net4462),
    .Y(_13471_),
    .B1(_13470_));
 sg13g2_nand2_1 _20751_ (.Y(_13472_),
    .A(net2108),
    .B(net4082));
 sg13g2_o21ai_1 _20752_ (.B1(_13472_),
    .Y(_00232_),
    .A1(net4082),
    .A2(_13471_));
 sg13g2_and2_1 _20753_ (.A(net1306),
    .B(net4462),
    .X(_13473_));
 sg13g2_a21oi_1 _20754_ (.A1(net1083),
    .A2(net4403),
    .Y(_13474_),
    .B1(_13473_));
 sg13g2_nand2_1 _20755_ (.Y(_13475_),
    .A(net1602),
    .B(net4075));
 sg13g2_o21ai_1 _20756_ (.B1(_13475_),
    .Y(_00233_),
    .A1(net4075),
    .A2(_13474_));
 sg13g2_and2_1 _20757_ (.A(\shift_reg[215] ),
    .B(net4461),
    .X(_13476_));
 sg13g2_a21oi_2 _20758_ (.B1(_13476_),
    .Y(_13477_),
    .A2(net4399),
    .A1(\inv_result[223] ));
 sg13g2_nand2_1 _20759_ (.Y(_13478_),
    .A(net1090),
    .B(net4067));
 sg13g2_o21ai_1 _20760_ (.B1(_13478_),
    .Y(_00234_),
    .A1(net4067),
    .A2(_13477_));
 sg13g2_and2_1 _20761_ (.A(net1125),
    .B(net4461),
    .X(_13479_));
 sg13g2_a21oi_1 _20762_ (.A1(net1073),
    .A2(net4399),
    .Y(_13480_),
    .B1(_13479_));
 sg13g2_nand2_1 _20763_ (.Y(_13481_),
    .A(net1910),
    .B(net4073));
 sg13g2_o21ai_1 _20764_ (.B1(_13481_),
    .Y(_00235_),
    .A1(net4073),
    .A2(_13480_));
 sg13g2_and2_1 _20765_ (.A(net1443),
    .B(net4461),
    .X(_13482_));
 sg13g2_a21oi_1 _20766_ (.A1(net1382),
    .A2(net4399),
    .Y(_13483_),
    .B1(_13482_));
 sg13g2_nand2_1 _20767_ (.Y(_13484_),
    .A(net1544),
    .B(net4073));
 sg13g2_o21ai_1 _20768_ (.B1(_13484_),
    .Y(_00236_),
    .A1(net4073),
    .A2(_13483_));
 sg13g2_and2_1 _20769_ (.A(net1642),
    .B(net4461),
    .X(_13485_));
 sg13g2_a21oi_1 _20770_ (.A1(net1532),
    .A2(net4399),
    .Y(_13486_),
    .B1(_13485_));
 sg13g2_nand2_1 _20771_ (.Y(_13487_),
    .A(net1927),
    .B(net4073));
 sg13g2_o21ai_1 _20772_ (.B1(_13487_),
    .Y(_00237_),
    .A1(net4073),
    .A2(_13486_));
 sg13g2_nor2_1 _20773_ (.A(_11032_),
    .B(net4461),
    .Y(_13488_));
 sg13g2_a21oi_2 _20774_ (.B1(_13488_),
    .Y(_13489_),
    .A2(net4461),
    .A1(\shift_reg[219] ));
 sg13g2_nand2_1 _20775_ (.Y(_13490_),
    .A(net1146),
    .B(net4064));
 sg13g2_o21ai_1 _20776_ (.B1(_13490_),
    .Y(_00238_),
    .A1(net4064),
    .A2(_13489_));
 sg13g2_and2_1 _20777_ (.A(\shift_reg[220] ),
    .B(net4457),
    .X(_13491_));
 sg13g2_a21oi_1 _20778_ (.A1(net1643),
    .A2(net4397),
    .Y(_13492_),
    .B1(_13491_));
 sg13g2_nand2_1 _20779_ (.Y(_13493_),
    .A(net1685),
    .B(net4076));
 sg13g2_o21ai_1 _20780_ (.B1(_13493_),
    .Y(_00239_),
    .A1(net4076),
    .A2(_13492_));
 sg13g2_nor2_1 _20781_ (.A(_11033_),
    .B(net4457),
    .Y(_13494_));
 sg13g2_a21oi_1 _20782_ (.A1(\shift_reg[221] ),
    .A2(net4457),
    .Y(_13495_),
    .B1(_13494_));
 sg13g2_nand2_1 _20783_ (.Y(_13496_),
    .A(net1192),
    .B(net4067));
 sg13g2_o21ai_1 _20784_ (.B1(_13496_),
    .Y(_00240_),
    .A1(net4072),
    .A2(_13495_));
 sg13g2_and2_1 _20785_ (.A(\shift_reg[222] ),
    .B(net4457),
    .X(_13497_));
 sg13g2_a21oi_1 _20786_ (.A1(net1071),
    .A2(net4397),
    .Y(_13498_),
    .B1(_13497_));
 sg13g2_nand2_1 _20787_ (.Y(_13499_),
    .A(net1202),
    .B(net4064));
 sg13g2_o21ai_1 _20788_ (.B1(_13499_),
    .Y(_00241_),
    .A1(net4064),
    .A2(_13498_));
 sg13g2_and2_1 _20789_ (.A(net1090),
    .B(net4457),
    .X(_13500_));
 sg13g2_a21oi_1 _20790_ (.A1(net1454),
    .A2(net4397),
    .Y(_13501_),
    .B1(_13500_));
 sg13g2_nand2_1 _20791_ (.Y(_13502_),
    .A(net1512),
    .B(net4067));
 sg13g2_o21ai_1 _20792_ (.B1(_13502_),
    .Y(_00242_),
    .A1(net4067),
    .A2(_13501_));
 sg13g2_and2_1 _20793_ (.A(\shift_reg[224] ),
    .B(net4456),
    .X(_13503_));
 sg13g2_a21oi_1 _20794_ (.A1(\inv_result[232] ),
    .A2(net4397),
    .Y(_13504_),
    .B1(_13503_));
 sg13g2_nand2_1 _20795_ (.Y(_13505_),
    .A(net1188),
    .B(net4066));
 sg13g2_o21ai_1 _20796_ (.B1(_13505_),
    .Y(_00243_),
    .A1(net4066),
    .A2(_13504_));
 sg13g2_nor2_1 _20797_ (.A(_11034_),
    .B(net4456),
    .Y(_13506_));
 sg13g2_a21oi_1 _20798_ (.A1(\shift_reg[225] ),
    .A2(net4456),
    .Y(_13507_),
    .B1(_13506_));
 sg13g2_nand2_1 _20799_ (.Y(_13508_),
    .A(net1319),
    .B(net4067));
 sg13g2_o21ai_1 _20800_ (.B1(_13508_),
    .Y(_00244_),
    .A1(net4067),
    .A2(_13507_));
 sg13g2_and2_1 _20801_ (.A(\shift_reg[226] ),
    .B(net4455),
    .X(_13509_));
 sg13g2_a21oi_1 _20802_ (.A1(\inv_result[234] ),
    .A2(net4397),
    .Y(_13510_),
    .B1(_13509_));
 sg13g2_nand2_1 _20803_ (.Y(_13511_),
    .A(net1129),
    .B(net4064));
 sg13g2_o21ai_1 _20804_ (.B1(_13511_),
    .Y(_00245_),
    .A1(net4064),
    .A2(_13510_));
 sg13g2_nor2_1 _20805_ (.A(_11035_),
    .B(net4455),
    .Y(_13512_));
 sg13g2_a21oi_1 _20806_ (.A1(net1146),
    .A2(net4455),
    .Y(_13513_),
    .B1(_13512_));
 sg13g2_nand2_1 _20807_ (.Y(_13514_),
    .A(net1340),
    .B(net4064));
 sg13g2_o21ai_1 _20808_ (.B1(_13514_),
    .Y(_00246_),
    .A1(net4064),
    .A2(_13513_));
 sg13g2_and2_1 _20809_ (.A(\shift_reg[228] ),
    .B(net4456),
    .X(_13515_));
 sg13g2_a21oi_1 _20810_ (.A1(\inv_result[236] ),
    .A2(net4397),
    .Y(_13516_),
    .B1(_13515_));
 sg13g2_nand2_1 _20811_ (.Y(_13517_),
    .A(net1194),
    .B(net4065));
 sg13g2_o21ai_1 _20812_ (.B1(_13517_),
    .Y(_00247_),
    .A1(net4065),
    .A2(_13516_));
 sg13g2_nor2_1 _20813_ (.A(_11036_),
    .B(net4455),
    .Y(_13518_));
 sg13g2_a21oi_1 _20814_ (.A1(\shift_reg[229] ),
    .A2(net4455),
    .Y(_13519_),
    .B1(_13518_));
 sg13g2_nand2_1 _20815_ (.Y(_13520_),
    .A(net1118),
    .B(net4065));
 sg13g2_o21ai_1 _20816_ (.B1(_13520_),
    .Y(_00248_),
    .A1(net4065),
    .A2(_13519_));
 sg13g2_and2_1 _20817_ (.A(net1202),
    .B(net4455),
    .X(_13521_));
 sg13g2_a21oi_1 _20818_ (.A1(\inv_result[238] ),
    .A2(net4397),
    .Y(_13522_),
    .B1(_13521_));
 sg13g2_nand2_1 _20819_ (.Y(_13523_),
    .A(net1302),
    .B(net4065));
 sg13g2_o21ai_1 _20820_ (.B1(_13523_),
    .Y(_00249_),
    .A1(net4065),
    .A2(_13522_));
 sg13g2_and2_1 _20821_ (.A(\shift_reg[231] ),
    .B(net4455),
    .X(_13524_));
 sg13g2_a21oi_1 _20822_ (.A1(\inv_result[239] ),
    .A2(net4397),
    .Y(_13525_),
    .B1(_13524_));
 sg13g2_nand2_1 _20823_ (.Y(_13526_),
    .A(net1105),
    .B(net4053));
 sg13g2_o21ai_1 _20824_ (.B1(_13526_),
    .Y(_00250_),
    .A1(net4053),
    .A2(_13525_));
 sg13g2_and2_1 _20825_ (.A(net1188),
    .B(net4456),
    .X(_13527_));
 sg13g2_a21oi_1 _20826_ (.A1(net2032),
    .A2(net4387),
    .Y(_13528_),
    .B1(_13527_));
 sg13g2_nand2_1 _20827_ (.Y(_13529_),
    .A(net2163),
    .B(net4066));
 sg13g2_o21ai_1 _20828_ (.B1(_13529_),
    .Y(_00251_),
    .A1(net4066),
    .A2(_13528_));
 sg13g2_nor2_1 _20829_ (.A(_11037_),
    .B(net4456),
    .Y(_13530_));
 sg13g2_a21oi_2 _20830_ (.B1(_13530_),
    .Y(_13531_),
    .A2(net4455),
    .A1(\shift_reg[233] ));
 sg13g2_nand2_1 _20831_ (.Y(_13532_),
    .A(net1138),
    .B(net4053));
 sg13g2_o21ai_1 _20832_ (.B1(_13532_),
    .Y(_00252_),
    .A1(net4053),
    .A2(_13531_));
 sg13g2_and2_1 _20833_ (.A(net1129),
    .B(net4452),
    .X(_13533_));
 sg13g2_a21oi_2 _20834_ (.B1(_13533_),
    .Y(_13534_),
    .A2(net4387),
    .A1(\inv_result[242] ));
 sg13g2_nand2_1 _20835_ (.Y(_13535_),
    .A(net1549),
    .B(net4054));
 sg13g2_o21ai_1 _20836_ (.B1(_13535_),
    .Y(_00253_),
    .A1(net4054),
    .A2(_13534_));
 sg13g2_nor2_1 _20837_ (.A(_11038_),
    .B(net4452),
    .Y(_13536_));
 sg13g2_a21oi_1 _20838_ (.A1(net1340),
    .A2(net4452),
    .Y(_13537_),
    .B1(_13536_));
 sg13g2_nand2_1 _20839_ (.Y(_13538_),
    .A(net2166),
    .B(net4065));
 sg13g2_o21ai_1 _20840_ (.B1(_13538_),
    .Y(_00254_),
    .A1(net4065),
    .A2(_13537_));
 sg13g2_and2_1 _20841_ (.A(net1194),
    .B(net4452),
    .X(_13539_));
 sg13g2_a21oi_1 _20842_ (.A1(net1375),
    .A2(net4388),
    .Y(_13540_),
    .B1(_13539_));
 sg13g2_nand2_1 _20843_ (.Y(_13541_),
    .A(net1996),
    .B(net4066));
 sg13g2_o21ai_1 _20844_ (.B1(_13541_),
    .Y(_00255_),
    .A1(net4066),
    .A2(_13540_));
 sg13g2_and2_1 _20845_ (.A(net1118),
    .B(net4452),
    .X(_13542_));
 sg13g2_a21oi_1 _20846_ (.A1(\inv_result[245] ),
    .A2(net4388),
    .Y(_13543_),
    .B1(_13542_));
 sg13g2_nand2_1 _20847_ (.Y(_13544_),
    .A(net1639),
    .B(net4054));
 sg13g2_o21ai_1 _20848_ (.B1(_13544_),
    .Y(_00256_),
    .A1(net4054),
    .A2(_13543_));
 sg13g2_and2_1 _20849_ (.A(net1302),
    .B(net4454),
    .X(_13545_));
 sg13g2_a21oi_2 _20850_ (.B1(_13545_),
    .Y(_13546_),
    .A2(net4388),
    .A1(\inv_result[246] ));
 sg13g2_nand2_1 _20851_ (.Y(_13547_),
    .A(net1564),
    .B(net4053));
 sg13g2_o21ai_1 _20852_ (.B1(_13547_),
    .Y(_00257_),
    .A1(net4053),
    .A2(_13546_));
 sg13g2_and2_1 _20853_ (.A(net1105),
    .B(net4454),
    .X(_13548_));
 sg13g2_a21oi_1 _20854_ (.A1(\inv_result[247] ),
    .A2(net4388),
    .Y(_13549_),
    .B1(_13548_));
 sg13g2_nand2_1 _20855_ (.Y(_13550_),
    .A(net1706),
    .B(net4053));
 sg13g2_o21ai_1 _20856_ (.B1(_13550_),
    .Y(_00258_),
    .A1(net4053),
    .A2(_13549_));
 sg13g2_and2_1 _20857_ (.A(\shift_reg[240] ),
    .B(net4451),
    .X(_13551_));
 sg13g2_a21oi_1 _20858_ (.A1(\inv_result[248] ),
    .A2(net4387),
    .Y(_13552_),
    .B1(_13551_));
 sg13g2_nand2_1 _20859_ (.Y(_13553_),
    .A(net1127),
    .B(net4057));
 sg13g2_o21ai_1 _20860_ (.B1(_13553_),
    .Y(_00259_),
    .A1(net4057),
    .A2(_13552_));
 sg13g2_and2_1 _20861_ (.A(\shift_reg[241] ),
    .B(net4452),
    .X(_13554_));
 sg13g2_a21oi_1 _20862_ (.A1(\inv_result[249] ),
    .A2(net4387),
    .Y(_13555_),
    .B1(_13554_));
 sg13g2_nand2_1 _20863_ (.Y(_13556_),
    .A(net1097),
    .B(net4056));
 sg13g2_o21ai_1 _20864_ (.B1(_13556_),
    .Y(_00260_),
    .A1(net4056),
    .A2(_13555_));
 sg13g2_and2_1 _20865_ (.A(\shift_reg[242] ),
    .B(net4451),
    .X(_13557_));
 sg13g2_a21oi_1 _20866_ (.A1(\inv_result[250] ),
    .A2(net4387),
    .Y(_13558_),
    .B1(_13557_));
 sg13g2_nand2_1 _20867_ (.Y(_13559_),
    .A(net1086),
    .B(net4056));
 sg13g2_o21ai_1 _20868_ (.B1(_13559_),
    .Y(_00261_),
    .A1(net4056),
    .A2(_13558_));
 sg13g2_nor2_1 _20869_ (.A(_11039_),
    .B(net4451),
    .Y(_13560_));
 sg13g2_a21oi_1 _20870_ (.A1(\shift_reg[243] ),
    .A2(net4452),
    .Y(_13561_),
    .B1(_13560_));
 sg13g2_nand2_1 _20871_ (.Y(_13562_),
    .A(net1115),
    .B(net4056));
 sg13g2_o21ai_1 _20872_ (.B1(_13562_),
    .Y(_00262_),
    .A1(net4056),
    .A2(_13561_));
 sg13g2_and2_1 _20873_ (.A(\shift_reg[244] ),
    .B(net4451),
    .X(_13563_));
 sg13g2_a21oi_2 _20874_ (.B1(_13563_),
    .Y(_13564_),
    .A2(net4387),
    .A1(\inv_result[252] ));
 sg13g2_nand2_1 _20875_ (.Y(_13565_),
    .A(net1153),
    .B(net4055));
 sg13g2_o21ai_1 _20876_ (.B1(_13565_),
    .Y(_00263_),
    .A1(net4055),
    .A2(_13564_));
 sg13g2_nor2_1 _20877_ (.A(_11040_),
    .B(net4451),
    .Y(_13566_));
 sg13g2_a21oi_2 _20878_ (.B1(_13566_),
    .Y(_13567_),
    .A2(net4451),
    .A1(\shift_reg[245] ));
 sg13g2_nand2_1 _20879_ (.Y(_13568_),
    .A(net1121),
    .B(net4055));
 sg13g2_o21ai_1 _20880_ (.B1(_13568_),
    .Y(_00264_),
    .A1(net4055),
    .A2(_13567_));
 sg13g2_and2_1 _20881_ (.A(\shift_reg[246] ),
    .B(net4451),
    .X(_13569_));
 sg13g2_a21oi_2 _20882_ (.B1(_13569_),
    .Y(_13570_),
    .A2(net4387),
    .A1(\inv_result[254] ));
 sg13g2_nand2_1 _20883_ (.Y(_13571_),
    .A(net1099),
    .B(net4055));
 sg13g2_o21ai_1 _20884_ (.B1(_13571_),
    .Y(_00265_),
    .A1(net4055),
    .A2(_13570_));
 sg13g2_and2_1 _20885_ (.A(\shift_reg[247] ),
    .B(net4451),
    .X(_13572_));
 sg13g2_a21oi_2 _20886_ (.B1(_13572_),
    .Y(_13573_),
    .A2(net4387),
    .A1(\inv_result[255] ));
 sg13g2_nand2_1 _20887_ (.Y(_13574_),
    .A(net1109),
    .B(net4055));
 sg13g2_o21ai_1 _20888_ (.B1(_13574_),
    .Y(_00266_),
    .A1(net4055),
    .A2(_13573_));
 sg13g2_nor2_1 _20889_ (.A(net1150),
    .B(net4379),
    .Y(_13575_));
 sg13g2_a21oi_1 _20890_ (.A1(net1150),
    .A2(_11065_),
    .Y(_00267_),
    .B1(_13575_));
 sg13g2_a21oi_1 _20891_ (.A1(net1150),
    .A2(_11065_),
    .Y(_13576_),
    .B1(net1562));
 sg13g2_nand3_1 _20892_ (.B(net1562),
    .C(_11065_),
    .A(net1150),
    .Y(_13577_));
 sg13g2_nand2_1 _20893_ (.Y(_13578_),
    .A(_11045_),
    .B(_13577_));
 sg13g2_nor2_1 _20894_ (.A(_13576_),
    .B(_13578_),
    .Y(_00268_));
 sg13g2_nand2_1 _20895_ (.Y(_13579_),
    .A(net1150),
    .B(net1631));
 sg13g2_nand4_1 _20896_ (.B(net1562),
    .C(net1631),
    .A(net1150),
    .Y(_13580_),
    .D(net4379));
 sg13g2_nand2_1 _20897_ (.Y(_13581_),
    .A(_11045_),
    .B(_13580_));
 sg13g2_a21oi_1 _20898_ (.A1(_10633_),
    .A2(_13577_),
    .Y(_00269_),
    .B1(_13581_));
 sg13g2_nor2b_1 _20899_ (.A(net1088),
    .B_N(_13580_),
    .Y(_13582_));
 sg13g2_a21oi_1 _20900_ (.A1(net1088),
    .A2(_13581_),
    .Y(_00270_),
    .B1(_13582_));
 sg13g2_and4_1 _20901_ (.A(net1150),
    .B(net1562),
    .C(net1088),
    .D(net1631),
    .X(_13583_));
 sg13g2_a21oi_1 _20902_ (.A1(_11065_),
    .A2(_13583_),
    .Y(_13584_),
    .B1(net1857));
 sg13g2_and3_1 _20903_ (.X(_13585_),
    .A(net1857),
    .B(net4379),
    .C(_13583_));
 sg13g2_nor3_1 _20904_ (.A(_17369_[0]),
    .B(_13584_),
    .C(_13585_),
    .Y(_00271_));
 sg13g2_and2_1 _20905_ (.A(net2119),
    .B(_13585_),
    .X(_13586_));
 sg13g2_a21oi_1 _20906_ (.A1(net2119),
    .A2(_11045_),
    .Y(_13587_),
    .B1(_13585_));
 sg13g2_nor2_1 _20907_ (.A(_13586_),
    .B(net2120),
    .Y(_00272_));
 sg13g2_nand3_1 _20908_ (.B(\u_inv.counter[5] ),
    .C(_13583_),
    .A(\u_inv.counter[4] ),
    .Y(_13588_));
 sg13g2_a21o_1 _20909_ (.A2(_13586_),
    .A1(net2240),
    .B1(_17369_[0]),
    .X(_13589_));
 sg13g2_nor2_1 _20910_ (.A(net2240),
    .B(_13586_),
    .Y(_13590_));
 sg13g2_nor2_1 _20911_ (.A(_13589_),
    .B(_13590_),
    .Y(_00273_));
 sg13g2_a21oi_1 _20912_ (.A1(\u_inv.counter[6] ),
    .A2(_13586_),
    .Y(_13591_),
    .B1(net1075));
 sg13g2_a21oi_1 _20913_ (.A1(net1075),
    .A2(_13589_),
    .Y(_00274_),
    .B1(_13591_));
 sg13g2_nand2_1 _20914_ (.Y(_13592_),
    .A(net1075),
    .B(net2240));
 sg13g2_nor2_1 _20915_ (.A(_13588_),
    .B(_13592_),
    .Y(_13593_));
 sg13g2_and4_1 _20916_ (.A(net1075),
    .B(\u_inv.counter[6] ),
    .C(net1227),
    .D(_13586_),
    .X(_13594_));
 sg13g2_or2_1 _20917_ (.X(_13595_),
    .B(_13594_),
    .A(_17369_[0]));
 sg13g2_a21oi_1 _20918_ (.A1(_11065_),
    .A2(_13593_),
    .Y(_13596_),
    .B1(net1227));
 sg13g2_nor2_1 _20919_ (.A(_13595_),
    .B(net1228),
    .Y(_00275_));
 sg13g2_nor2_1 _20920_ (.A(net1067),
    .B(_13594_),
    .Y(_13597_));
 sg13g2_a21oi_1 _20921_ (.A1(net1067),
    .A2(_13595_),
    .Y(_00276_),
    .B1(_13597_));
 sg13g2_nand2b_1 _20922_ (.Y(_13598_),
    .B(\u_inv.d_reg[256] ),
    .A_N(\u_inv.d_next[256] ));
 sg13g2_nor2_1 _20923_ (.A(\u_inv.d_next[256] ),
    .B(\u_inv.d_reg[256] ),
    .Y(_13599_));
 sg13g2_xnor2_1 _20924_ (.Y(_13600_),
    .A(\u_inv.d_next[256] ),
    .B(\u_inv.d_reg[256] ));
 sg13g2_nor2_1 _20925_ (.A(\u_inv.d_next[255] ),
    .B(\u_inv.d_reg[255] ),
    .Y(_13601_));
 sg13g2_xnor2_1 _20926_ (.Y(_13602_),
    .A(\u_inv.d_next[255] ),
    .B(\u_inv.d_reg[255] ));
 sg13g2_nand2_1 _20927_ (.Y(_13603_),
    .A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ));
 sg13g2_xor2_1 _20928_ (.B(\u_inv.d_reg[254] ),
    .A(\u_inv.d_next[254] ),
    .X(_13604_));
 sg13g2_xnor2_1 _20929_ (.Y(_13605_),
    .A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ));
 sg13g2_nand2_1 _20930_ (.Y(_13606_),
    .A(_13602_),
    .B(_13605_));
 sg13g2_nor2_1 _20931_ (.A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ),
    .Y(_13607_));
 sg13g2_nand2_1 _20932_ (.Y(_13608_),
    .A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ));
 sg13g2_nand2b_2 _20933_ (.Y(_13609_),
    .B(_13608_),
    .A_N(_13607_));
 sg13g2_nand2_1 _20934_ (.Y(_13610_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_xnor2_1 _20935_ (.Y(_13611_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_and2_1 _20936_ (.A(_13609_),
    .B(_13611_),
    .X(_13612_));
 sg13g2_nand2b_1 _20937_ (.Y(_13613_),
    .B(_13612_),
    .A_N(_13606_));
 sg13g2_nand2_1 _20938_ (.Y(_13614_),
    .A(\u_inv.d_next[251] ),
    .B(\u_inv.d_reg[251] ));
 sg13g2_nor2_1 _20939_ (.A(\u_inv.d_next[251] ),
    .B(\u_inv.d_reg[251] ),
    .Y(_13615_));
 sg13g2_xnor2_1 _20940_ (.Y(_13616_),
    .A(\u_inv.d_next[251] ),
    .B(\u_inv.d_reg[251] ));
 sg13g2_nand2_1 _20941_ (.Y(_13617_),
    .A(\u_inv.d_next[250] ),
    .B(\u_inv.d_reg[250] ));
 sg13g2_xor2_1 _20942_ (.B(\u_inv.d_reg[250] ),
    .A(\u_inv.d_next[250] ),
    .X(_13618_));
 sg13g2_xnor2_1 _20943_ (.Y(_13619_),
    .A(\u_inv.d_next[250] ),
    .B(\u_inv.d_reg[250] ));
 sg13g2_nand2_1 _20944_ (.Y(_13620_),
    .A(_13616_),
    .B(_13619_));
 sg13g2_nor2_1 _20945_ (.A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ),
    .Y(_13621_));
 sg13g2_nand2_1 _20946_ (.Y(_13622_),
    .A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ));
 sg13g2_nand2b_2 _20947_ (.Y(_13623_),
    .B(_13622_),
    .A_N(_13621_));
 sg13g2_nand2_1 _20948_ (.Y(_13624_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_xnor2_1 _20949_ (.Y(_13625_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_and2_1 _20950_ (.A(_13623_),
    .B(_13625_),
    .X(_13626_));
 sg13g2_nand2_1 _20951_ (.Y(_13627_),
    .A(_13623_),
    .B(_13625_));
 sg13g2_nor3_2 _20952_ (.A(_13613_),
    .B(_13620_),
    .C(_13627_),
    .Y(_13628_));
 sg13g2_nand2_1 _20953_ (.Y(_13629_),
    .A(\u_inv.d_next[242] ),
    .B(\u_inv.d_reg[242] ));
 sg13g2_xnor2_1 _20954_ (.Y(_13630_),
    .A(\u_inv.d_next[242] ),
    .B(\u_inv.d_reg[242] ));
 sg13g2_inv_2 _20955_ (.Y(_13631_),
    .A(_13630_));
 sg13g2_nand2b_2 _20956_ (.Y(_13632_),
    .B(\u_inv.d_reg[241] ),
    .A_N(\u_inv.d_next[241] ));
 sg13g2_nor2b_1 _20957_ (.A(\u_inv.d_reg[241] ),
    .B_N(\u_inv.d_next[241] ),
    .Y(_13633_));
 sg13g2_nand2b_1 _20958_ (.Y(_13634_),
    .B(\u_inv.d_next[241] ),
    .A_N(\u_inv.d_reg[241] ));
 sg13g2_and2_1 _20959_ (.A(_13632_),
    .B(_13634_),
    .X(_13635_));
 sg13g2_nand2_2 _20960_ (.Y(_13636_),
    .A(_13632_),
    .B(_13634_));
 sg13g2_nand2_1 _20961_ (.Y(_13637_),
    .A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ));
 sg13g2_nor2_1 _20962_ (.A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ),
    .Y(_13638_));
 sg13g2_xnor2_1 _20963_ (.Y(_13639_),
    .A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ));
 sg13g2_inv_1 _20964_ (.Y(_13640_),
    .A(_13639_));
 sg13g2_nand3_1 _20965_ (.B(_13635_),
    .C(_13639_),
    .A(_13630_),
    .Y(_13641_));
 sg13g2_xnor2_1 _20966_ (.Y(_13642_),
    .A(\u_inv.d_next[245] ),
    .B(\u_inv.d_reg[245] ));
 sg13g2_nand2_1 _20967_ (.Y(_13643_),
    .A(\u_inv.d_next[244] ),
    .B(\u_inv.d_reg[244] ));
 sg13g2_xnor2_1 _20968_ (.Y(_13644_),
    .A(\u_inv.d_next[244] ),
    .B(\u_inv.d_reg[244] ));
 sg13g2_and2_1 _20969_ (.A(_13642_),
    .B(_13644_),
    .X(_13645_));
 sg13g2_nor2_1 _20970_ (.A(\u_inv.d_next[247] ),
    .B(\u_inv.d_reg[247] ),
    .Y(_13646_));
 sg13g2_xor2_1 _20971_ (.B(\u_inv.d_reg[247] ),
    .A(\u_inv.d_next[247] ),
    .X(_13647_));
 sg13g2_xnor2_1 _20972_ (.Y(_13648_),
    .A(\u_inv.d_next[247] ),
    .B(\u_inv.d_reg[247] ));
 sg13g2_and2_1 _20973_ (.A(\u_inv.d_next[246] ),
    .B(\u_inv.d_reg[246] ),
    .X(_13649_));
 sg13g2_xor2_1 _20974_ (.B(\u_inv.d_reg[246] ),
    .A(\u_inv.d_next[246] ),
    .X(_13650_));
 sg13g2_xnor2_1 _20975_ (.Y(_13651_),
    .A(\u_inv.d_next[246] ),
    .B(\u_inv.d_reg[246] ));
 sg13g2_nand3_1 _20976_ (.B(_13648_),
    .C(_13651_),
    .A(_13645_),
    .Y(_13652_));
 sg13g2_nand2_1 _20977_ (.Y(_13653_),
    .A(\u_inv.d_next[240] ),
    .B(\u_inv.d_reg[240] ));
 sg13g2_xor2_1 _20978_ (.B(\u_inv.d_reg[240] ),
    .A(\u_inv.d_next[240] ),
    .X(_13654_));
 sg13g2_nor3_1 _20979_ (.A(_13641_),
    .B(_13652_),
    .C(_13654_),
    .Y(_13655_));
 sg13g2_nand2_2 _20980_ (.Y(_13656_),
    .A(_13628_),
    .B(_13655_));
 sg13g2_nand2_1 _20981_ (.Y(_13657_),
    .A(\u_inv.d_next[234] ),
    .B(\u_inv.d_reg[234] ));
 sg13g2_xor2_1 _20982_ (.B(\u_inv.d_reg[234] ),
    .A(\u_inv.d_next[234] ),
    .X(_13658_));
 sg13g2_xnor2_1 _20983_ (.Y(_13659_),
    .A(\u_inv.d_next[234] ),
    .B(\u_inv.d_reg[234] ));
 sg13g2_nand2_1 _20984_ (.Y(_13660_),
    .A(\u_inv.d_next[232] ),
    .B(\u_inv.d_reg[232] ));
 sg13g2_xnor2_1 _20985_ (.Y(_13661_),
    .A(\u_inv.d_next[232] ),
    .B(\u_inv.d_reg[232] ));
 sg13g2_nand2b_1 _20986_ (.Y(_13662_),
    .B(\u_inv.d_reg[233] ),
    .A_N(\u_inv.d_next[233] ));
 sg13g2_nor2b_1 _20987_ (.A(\u_inv.d_reg[233] ),
    .B_N(\u_inv.d_next[233] ),
    .Y(_13663_));
 sg13g2_xnor2_1 _20988_ (.Y(_13664_),
    .A(\u_inv.d_next[233] ),
    .B(\u_inv.d_reg[233] ));
 sg13g2_nor2_1 _20989_ (.A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ),
    .Y(_13665_));
 sg13g2_nand2_1 _20990_ (.Y(_13666_),
    .A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ));
 sg13g2_nand2b_2 _20991_ (.Y(_13667_),
    .B(_13666_),
    .A_N(_13665_));
 sg13g2_nand4_1 _20992_ (.B(_13661_),
    .C(_13664_),
    .A(_13659_),
    .Y(_13668_),
    .D(_13667_));
 sg13g2_nor2_1 _20993_ (.A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ),
    .Y(_13669_));
 sg13g2_nand2_1 _20994_ (.Y(_13670_),
    .A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ));
 sg13g2_nand2b_2 _20995_ (.Y(_13671_),
    .B(_13670_),
    .A_N(_13669_));
 sg13g2_nand2_1 _20996_ (.Y(_13672_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_xnor2_1 _20997_ (.Y(_13673_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_and2_1 _20998_ (.A(_13671_),
    .B(_13673_),
    .X(_13674_));
 sg13g2_nand2_1 _20999_ (.Y(_13675_),
    .A(_13671_),
    .B(_13673_));
 sg13g2_nand2_1 _21000_ (.Y(_13676_),
    .A(\u_inv.d_next[239] ),
    .B(\u_inv.d_reg[239] ));
 sg13g2_xor2_1 _21001_ (.B(\u_inv.d_reg[239] ),
    .A(\u_inv.d_next[239] ),
    .X(_13677_));
 sg13g2_and2_1 _21002_ (.A(\u_inv.d_next[238] ),
    .B(\u_inv.d_reg[238] ),
    .X(_13678_));
 sg13g2_xor2_1 _21003_ (.B(\u_inv.d_reg[238] ),
    .A(\u_inv.d_next[238] ),
    .X(_13679_));
 sg13g2_nor2_1 _21004_ (.A(_13677_),
    .B(_13679_),
    .Y(_13680_));
 sg13g2_nor4_1 _21005_ (.A(_13668_),
    .B(_13675_),
    .C(_13677_),
    .D(_13679_),
    .Y(_13681_));
 sg13g2_nor2_1 _21006_ (.A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ),
    .Y(_13682_));
 sg13g2_xor2_1 _21007_ (.B(\u_inv.d_reg[231] ),
    .A(\u_inv.d_next[231] ),
    .X(_13683_));
 sg13g2_nand2_1 _21008_ (.Y(_13684_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_xor2_1 _21009_ (.B(\u_inv.d_reg[230] ),
    .A(\u_inv.d_next[230] ),
    .X(_13685_));
 sg13g2_xnor2_1 _21010_ (.Y(_13686_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_nor2_1 _21011_ (.A(_13683_),
    .B(_13685_),
    .Y(_13687_));
 sg13g2_nand2b_1 _21012_ (.Y(_13688_),
    .B(\u_inv.d_next[229] ),
    .A_N(net4766));
 sg13g2_nor2b_1 _21013_ (.A(\u_inv.d_next[229] ),
    .B_N(net4766),
    .Y(_13689_));
 sg13g2_xnor2_1 _21014_ (.Y(_13690_),
    .A(\u_inv.d_next[229] ),
    .B(net4766));
 sg13g2_nand2_1 _21015_ (.Y(_13691_),
    .A(\u_inv.d_next[228] ),
    .B(net4767));
 sg13g2_xor2_1 _21016_ (.B(net4767),
    .A(\u_inv.d_next[228] ),
    .X(_13692_));
 sg13g2_xnor2_1 _21017_ (.Y(_13693_),
    .A(\u_inv.d_next[228] ),
    .B(net4767));
 sg13g2_and2_1 _21018_ (.A(_13690_),
    .B(_13693_),
    .X(_13694_));
 sg13g2_and2_1 _21019_ (.A(_13687_),
    .B(_13694_),
    .X(_13695_));
 sg13g2_nand2b_1 _21020_ (.Y(_13696_),
    .B(\u_inv.d_reg[227] ),
    .A_N(\u_inv.d_next[227] ));
 sg13g2_nor2b_1 _21021_ (.A(\u_inv.d_reg[227] ),
    .B_N(\u_inv.d_next[227] ),
    .Y(_13697_));
 sg13g2_xnor2_1 _21022_ (.Y(_13698_),
    .A(\u_inv.d_next[227] ),
    .B(\u_inv.d_reg[227] ));
 sg13g2_and2_1 _21023_ (.A(\u_inv.d_next[226] ),
    .B(net4768),
    .X(_13699_));
 sg13g2_nor2_1 _21024_ (.A(\u_inv.d_next[226] ),
    .B(net4768),
    .Y(_13700_));
 sg13g2_nor2_1 _21025_ (.A(_13699_),
    .B(_13700_),
    .Y(_13701_));
 sg13g2_xnor2_1 _21026_ (.Y(_13702_),
    .A(\u_inv.d_next[226] ),
    .B(net4768));
 sg13g2_nand2_1 _21027_ (.Y(_13703_),
    .A(_13698_),
    .B(_13702_));
 sg13g2_nor2b_1 _21028_ (.A(\u_inv.d_reg[225] ),
    .B_N(\u_inv.d_next[225] ),
    .Y(_13704_));
 sg13g2_nand2b_1 _21029_ (.Y(_13705_),
    .B(\u_inv.d_reg[225] ),
    .A_N(\u_inv.d_next[225] ));
 sg13g2_xnor2_1 _21030_ (.Y(_13706_),
    .A(\u_inv.d_next[225] ),
    .B(\u_inv.d_reg[225] ));
 sg13g2_nand2_1 _21031_ (.Y(_13707_),
    .A(\u_inv.d_next[224] ),
    .B(\u_inv.d_reg[224] ));
 sg13g2_xnor2_1 _21032_ (.Y(_13708_),
    .A(\u_inv.d_next[224] ),
    .B(\u_inv.d_reg[224] ));
 sg13g2_and2_1 _21033_ (.A(_13706_),
    .B(_13708_),
    .X(_13709_));
 sg13g2_and4_1 _21034_ (.A(_13695_),
    .B(_13698_),
    .C(_13702_),
    .D(_13709_),
    .X(_13710_));
 sg13g2_nand2_1 _21035_ (.Y(_13711_),
    .A(_13681_),
    .B(_13710_));
 sg13g2_inv_1 _21036_ (.Y(_13712_),
    .A(_13711_));
 sg13g2_nand2b_2 _21037_ (.Y(_13713_),
    .B(_13712_),
    .A_N(_13656_));
 sg13g2_nor2_1 _21038_ (.A(\u_inv.d_next[207] ),
    .B(\u_inv.d_reg[207] ),
    .Y(_13714_));
 sg13g2_xnor2_1 _21039_ (.Y(_13715_),
    .A(\u_inv.d_next[207] ),
    .B(\u_inv.d_reg[207] ));
 sg13g2_nand2_1 _21040_ (.Y(_13716_),
    .A(\u_inv.d_next[206] ),
    .B(\u_inv.d_reg[206] ));
 sg13g2_xnor2_1 _21041_ (.Y(_13717_),
    .A(\u_inv.d_next[206] ),
    .B(\u_inv.d_reg[206] ));
 sg13g2_and2_1 _21042_ (.A(_13715_),
    .B(_13717_),
    .X(_13718_));
 sg13g2_nand2b_1 _21043_ (.Y(_13719_),
    .B(\u_inv.d_next[205] ),
    .A_N(\u_inv.d_reg[205] ));
 sg13g2_nor2b_1 _21044_ (.A(\u_inv.d_next[205] ),
    .B_N(\u_inv.d_reg[205] ),
    .Y(_13720_));
 sg13g2_xnor2_1 _21045_ (.Y(_13721_),
    .A(\u_inv.d_next[205] ),
    .B(\u_inv.d_reg[205] ));
 sg13g2_xor2_1 _21046_ (.B(\u_inv.d_reg[205] ),
    .A(\u_inv.d_next[205] ),
    .X(_13722_));
 sg13g2_nand2_1 _21047_ (.Y(_13723_),
    .A(\u_inv.d_next[204] ),
    .B(\u_inv.d_reg[204] ));
 sg13g2_xor2_1 _21048_ (.B(\u_inv.d_reg[204] ),
    .A(\u_inv.d_next[204] ),
    .X(_13724_));
 sg13g2_nor2_1 _21049_ (.A(_13722_),
    .B(_13724_),
    .Y(_13725_));
 sg13g2_inv_1 _21050_ (.Y(_13726_),
    .A(_13725_));
 sg13g2_nand2_1 _21051_ (.Y(_13727_),
    .A(_13718_),
    .B(_13725_));
 sg13g2_xnor2_1 _21052_ (.Y(_13728_),
    .A(\u_inv.d_next[201] ),
    .B(\u_inv.d_reg[201] ));
 sg13g2_xor2_1 _21053_ (.B(\u_inv.d_reg[201] ),
    .A(\u_inv.d_next[201] ),
    .X(_13729_));
 sg13g2_nand2_1 _21054_ (.Y(_13730_),
    .A(\u_inv.d_next[200] ),
    .B(\u_inv.d_reg[200] ));
 sg13g2_xnor2_1 _21055_ (.Y(_13731_),
    .A(\u_inv.d_next[200] ),
    .B(\u_inv.d_reg[200] ));
 sg13g2_and2_1 _21056_ (.A(_13728_),
    .B(_13731_),
    .X(_13732_));
 sg13g2_inv_1 _21057_ (.Y(_13733_),
    .A(_13732_));
 sg13g2_nor2_1 _21058_ (.A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ),
    .Y(_13734_));
 sg13g2_and2_1 _21059_ (.A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ),
    .X(_13735_));
 sg13g2_nor2_2 _21060_ (.A(_13734_),
    .B(_13735_),
    .Y(_13736_));
 sg13g2_or2_1 _21061_ (.X(_13737_),
    .B(_13735_),
    .A(_13734_));
 sg13g2_nor2b_1 _21062_ (.A(\u_inv.d_next[203] ),
    .B_N(\u_inv.d_reg[203] ),
    .Y(_13738_));
 sg13g2_nand2b_1 _21063_ (.Y(_13739_),
    .B(\u_inv.d_next[203] ),
    .A_N(\u_inv.d_reg[203] ));
 sg13g2_nand2b_2 _21064_ (.Y(_13740_),
    .B(_13739_),
    .A_N(_13738_));
 sg13g2_nor2_1 _21065_ (.A(_13736_),
    .B(_13740_),
    .Y(_13741_));
 sg13g2_nand4_1 _21066_ (.B(_13725_),
    .C(_13732_),
    .A(_13718_),
    .Y(_13742_),
    .D(_13741_));
 sg13g2_nor2b_1 _21067_ (.A(\u_inv.d_reg[199] ),
    .B_N(\u_inv.d_next[199] ),
    .Y(_13743_));
 sg13g2_nand2b_1 _21068_ (.Y(_13744_),
    .B(\u_inv.d_reg[199] ),
    .A_N(\u_inv.d_next[199] ));
 sg13g2_xnor2_1 _21069_ (.Y(_13745_),
    .A(\u_inv.d_next[199] ),
    .B(\u_inv.d_reg[199] ));
 sg13g2_nand2b_2 _21070_ (.Y(_13746_),
    .B(_13744_),
    .A_N(_13743_));
 sg13g2_nand2_1 _21071_ (.Y(_13747_),
    .A(\u_inv.d_next[198] ),
    .B(net4771));
 sg13g2_nor2_1 _21072_ (.A(\u_inv.d_next[198] ),
    .B(net4771),
    .Y(_13748_));
 sg13g2_xor2_1 _21073_ (.B(net4771),
    .A(\u_inv.d_next[198] ),
    .X(_13749_));
 sg13g2_xnor2_1 _21074_ (.Y(_13750_),
    .A(\u_inv.d_next[198] ),
    .B(net4771));
 sg13g2_nand2_1 _21075_ (.Y(_13751_),
    .A(_13745_),
    .B(_13750_));
 sg13g2_nor2_1 _21076_ (.A(\u_inv.d_next[197] ),
    .B(net4772),
    .Y(_13752_));
 sg13g2_xor2_1 _21077_ (.B(net4772),
    .A(\u_inv.d_next[197] ),
    .X(_13753_));
 sg13g2_xnor2_1 _21078_ (.Y(_13754_),
    .A(\u_inv.d_next[197] ),
    .B(net4772));
 sg13g2_nand2_1 _21079_ (.Y(_13755_),
    .A(\u_inv.d_next[196] ),
    .B(net4773));
 sg13g2_xor2_1 _21080_ (.B(net4773),
    .A(\u_inv.d_next[196] ),
    .X(_13756_));
 sg13g2_xnor2_1 _21081_ (.Y(_13757_),
    .A(\u_inv.d_next[196] ),
    .B(net4773));
 sg13g2_nand2_1 _21082_ (.Y(_13758_),
    .A(_13754_),
    .B(_13757_));
 sg13g2_nor2_1 _21083_ (.A(_13751_),
    .B(_13758_),
    .Y(_13759_));
 sg13g2_nand2b_1 _21084_ (.Y(_13760_),
    .B(\u_inv.d_reg[195] ),
    .A_N(\u_inv.d_next[195] ));
 sg13g2_nor2b_1 _21085_ (.A(\u_inv.d_reg[195] ),
    .B_N(\u_inv.d_next[195] ),
    .Y(_13761_));
 sg13g2_xnor2_1 _21086_ (.Y(_13762_),
    .A(\u_inv.d_next[195] ),
    .B(\u_inv.d_reg[195] ));
 sg13g2_nand2_1 _21087_ (.Y(_13763_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_xnor2_1 _21088_ (.Y(_13764_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_and2_1 _21089_ (.A(_13762_),
    .B(_13764_),
    .X(_13765_));
 sg13g2_nand2_1 _21090_ (.Y(_13766_),
    .A(_13762_),
    .B(_13764_));
 sg13g2_nor2b_1 _21091_ (.A(\u_inv.d_reg[193] ),
    .B_N(\u_inv.d_next[193] ),
    .Y(_13767_));
 sg13g2_nand2b_1 _21092_ (.Y(_13768_),
    .B(\u_inv.d_reg[193] ),
    .A_N(\u_inv.d_next[193] ));
 sg13g2_xnor2_1 _21093_ (.Y(_13769_),
    .A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ));
 sg13g2_inv_1 _21094_ (.Y(_13770_),
    .A(_13769_));
 sg13g2_nand2_1 _21095_ (.Y(_13771_),
    .A(\u_inv.d_next[192] ),
    .B(\u_inv.d_reg[192] ));
 sg13g2_xnor2_1 _21096_ (.Y(_13772_),
    .A(\u_inv.d_next[192] ),
    .B(\u_inv.d_reg[192] ));
 sg13g2_nand2_1 _21097_ (.Y(_13773_),
    .A(_13769_),
    .B(_13772_));
 sg13g2_nand4_1 _21098_ (.B(_13765_),
    .C(_13769_),
    .A(_13759_),
    .Y(_13774_),
    .D(_13772_));
 sg13g2_nor2_2 _21099_ (.A(_13742_),
    .B(_13774_),
    .Y(_13775_));
 sg13g2_nor2_1 _21100_ (.A(\u_inv.d_next[221] ),
    .B(\u_inv.d_reg[221] ),
    .Y(_13776_));
 sg13g2_nand2_1 _21101_ (.Y(_13777_),
    .A(\u_inv.d_next[221] ),
    .B(\u_inv.d_reg[221] ));
 sg13g2_nand2b_2 _21102_ (.Y(_13778_),
    .B(_13777_),
    .A_N(_13776_));
 sg13g2_nand2_1 _21103_ (.Y(_13779_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_xnor2_1 _21104_ (.Y(_13780_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_and2_1 _21105_ (.A(_13778_),
    .B(_13780_),
    .X(_13781_));
 sg13g2_xor2_1 _21106_ (.B(\u_inv.d_reg[223] ),
    .A(\u_inv.d_next[223] ),
    .X(_13782_));
 sg13g2_nand2_1 _21107_ (.Y(_13783_),
    .A(\u_inv.d_next[222] ),
    .B(\u_inv.d_reg[222] ));
 sg13g2_nor2_1 _21108_ (.A(\u_inv.d_next[222] ),
    .B(\u_inv.d_reg[222] ),
    .Y(_13784_));
 sg13g2_xor2_1 _21109_ (.B(\u_inv.d_reg[222] ),
    .A(\u_inv.d_next[222] ),
    .X(_13785_));
 sg13g2_nor2_1 _21110_ (.A(_13782_),
    .B(_13785_),
    .Y(_13786_));
 sg13g2_and2_1 _21111_ (.A(_13781_),
    .B(_13786_),
    .X(_13787_));
 sg13g2_nand2_1 _21112_ (.Y(_13788_),
    .A(\u_inv.d_next[216] ),
    .B(\u_inv.d_reg[216] ));
 sg13g2_xor2_1 _21113_ (.B(\u_inv.d_reg[216] ),
    .A(\u_inv.d_next[216] ),
    .X(_13789_));
 sg13g2_inv_2 _21114_ (.Y(_13790_),
    .A(_13789_));
 sg13g2_and2_1 _21115_ (.A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ),
    .X(_13791_));
 sg13g2_xor2_1 _21116_ (.B(\u_inv.d_reg[218] ),
    .A(\u_inv.d_next[218] ),
    .X(_13792_));
 sg13g2_xnor2_1 _21117_ (.Y(_13793_),
    .A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ));
 sg13g2_nor2_1 _21118_ (.A(\u_inv.d_next[217] ),
    .B(_10891_),
    .Y(_13794_));
 sg13g2_xor2_1 _21119_ (.B(\u_inv.d_reg[217] ),
    .A(\u_inv.d_next[217] ),
    .X(_13795_));
 sg13g2_nand2_1 _21120_ (.Y(_13796_),
    .A(\u_inv.d_next[219] ),
    .B(\u_inv.d_reg[219] ));
 sg13g2_xor2_1 _21121_ (.B(\u_inv.d_reg[219] ),
    .A(\u_inv.d_next[219] ),
    .X(_13797_));
 sg13g2_nor4_1 _21122_ (.A(_13789_),
    .B(_13792_),
    .C(_13795_),
    .D(_13797_),
    .Y(_13798_));
 sg13g2_and2_1 _21123_ (.A(_13787_),
    .B(_13798_),
    .X(_13799_));
 sg13g2_nor2_1 _21124_ (.A(\u_inv.d_next[215] ),
    .B(\u_inv.d_reg[215] ),
    .Y(_13800_));
 sg13g2_xnor2_1 _21125_ (.Y(_13801_),
    .A(\u_inv.d_next[215] ),
    .B(\u_inv.d_reg[215] ));
 sg13g2_nand2_1 _21126_ (.Y(_13802_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_xnor2_1 _21127_ (.Y(_13803_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_and2_1 _21128_ (.A(_13801_),
    .B(_13803_),
    .X(_13804_));
 sg13g2_nor2b_1 _21129_ (.A(\u_inv.d_reg[213] ),
    .B_N(\u_inv.d_next[213] ),
    .Y(_13805_));
 sg13g2_nand2b_1 _21130_ (.Y(_13806_),
    .B(\u_inv.d_reg[213] ),
    .A_N(\u_inv.d_next[213] ));
 sg13g2_nor2b_2 _21131_ (.A(_13805_),
    .B_N(_13806_),
    .Y(_13807_));
 sg13g2_nand2_1 _21132_ (.Y(_13808_),
    .A(\u_inv.d_next[212] ),
    .B(\u_inv.d_reg[212] ));
 sg13g2_xor2_1 _21133_ (.B(\u_inv.d_reg[212] ),
    .A(\u_inv.d_next[212] ),
    .X(_13809_));
 sg13g2_xnor2_1 _21134_ (.Y(_13810_),
    .A(\u_inv.d_next[212] ),
    .B(\u_inv.d_reg[212] ));
 sg13g2_and2_1 _21135_ (.A(_13807_),
    .B(_13810_),
    .X(_13811_));
 sg13g2_inv_1 _21136_ (.Y(_13812_),
    .A(_13811_));
 sg13g2_nand2_1 _21137_ (.Y(_13813_),
    .A(_13804_),
    .B(_13811_));
 sg13g2_nor2_1 _21138_ (.A(\u_inv.d_next[211] ),
    .B(_10894_),
    .Y(_13814_));
 sg13g2_xnor2_1 _21139_ (.Y(_13815_),
    .A(\u_inv.d_next[211] ),
    .B(\u_inv.d_reg[211] ));
 sg13g2_nor2_1 _21140_ (.A(\u_inv.d_next[210] ),
    .B(\u_inv.d_reg[210] ),
    .Y(_13816_));
 sg13g2_nand2_1 _21141_ (.Y(_13817_),
    .A(\u_inv.d_next[210] ),
    .B(\u_inv.d_reg[210] ));
 sg13g2_nor2b_2 _21142_ (.A(_13816_),
    .B_N(_13817_),
    .Y(_13818_));
 sg13g2_nor2b_1 _21143_ (.A(_13818_),
    .B_N(_13815_),
    .Y(_13819_));
 sg13g2_nor2b_1 _21144_ (.A(net4769),
    .B_N(\u_inv.d_next[209] ),
    .Y(_13820_));
 sg13g2_nand2b_1 _21145_ (.Y(_13821_),
    .B(net4769),
    .A_N(\u_inv.d_next[209] ));
 sg13g2_nor2b_2 _21146_ (.A(_13820_),
    .B_N(_13821_),
    .Y(_13822_));
 sg13g2_xor2_1 _21147_ (.B(net4769),
    .A(\u_inv.d_next[209] ),
    .X(_13823_));
 sg13g2_and2_1 _21148_ (.A(\u_inv.d_next[208] ),
    .B(net4770),
    .X(_13824_));
 sg13g2_xnor2_1 _21149_ (.Y(_13825_),
    .A(\u_inv.d_next[208] ),
    .B(net4770));
 sg13g2_nand2_1 _21150_ (.Y(_13826_),
    .A(_13822_),
    .B(net4431));
 sg13g2_nand3_1 _21151_ (.B(_13822_),
    .C(net4431),
    .A(_13819_),
    .Y(_13827_));
 sg13g2_nor2_1 _21152_ (.A(_13813_),
    .B(_13827_),
    .Y(_13828_));
 sg13g2_inv_1 _21153_ (.Y(_13829_),
    .A(_13828_));
 sg13g2_nand3_1 _21154_ (.B(_13799_),
    .C(_13828_),
    .A(_13775_),
    .Y(_13830_));
 sg13g2_or2_1 _21155_ (.X(_13831_),
    .B(_13830_),
    .A(_13713_));
 sg13g2_nor2b_1 _21156_ (.A(\u_inv.d_reg[235] ),
    .B_N(\u_inv.d_next[235] ),
    .Y(_13832_));
 sg13g2_nand2b_1 _21157_ (.Y(_13833_),
    .B(\u_inv.d_next[234] ),
    .A_N(\u_inv.d_reg[234] ));
 sg13g2_nor2b_1 _21158_ (.A(\u_inv.d_reg[232] ),
    .B_N(\u_inv.d_next[232] ),
    .Y(_13834_));
 sg13g2_o21ai_1 _21159_ (.B1(_13662_),
    .Y(_13835_),
    .A1(_13663_),
    .A2(_13834_));
 sg13g2_inv_1 _21160_ (.Y(_13836_),
    .A(_13835_));
 sg13g2_o21ai_1 _21161_ (.B1(_13833_),
    .Y(_13837_),
    .A1(_13658_),
    .A2(_13835_));
 sg13g2_a21oi_1 _21162_ (.A1(_13667_),
    .A2(_13837_),
    .Y(_13838_),
    .B1(_13832_));
 sg13g2_nor2b_1 _21163_ (.A(\u_inv.d_reg[224] ),
    .B_N(\u_inv.d_next[224] ),
    .Y(_13839_));
 sg13g2_a21o_1 _21164_ (.A2(_13839_),
    .A1(_13705_),
    .B1(_13704_),
    .X(_13840_));
 sg13g2_nand2b_1 _21165_ (.Y(_13841_),
    .B(_13840_),
    .A_N(_13703_));
 sg13g2_nor2b_1 _21166_ (.A(net4768),
    .B_N(\u_inv.d_next[226] ),
    .Y(_13842_));
 sg13g2_o21ai_1 _21167_ (.B1(_13696_),
    .Y(_13843_),
    .A1(_13697_),
    .A2(_13842_));
 sg13g2_nand2_1 _21168_ (.Y(_13844_),
    .A(_13841_),
    .B(_13843_));
 sg13g2_nand2b_1 _21169_ (.Y(_13845_),
    .B(\u_inv.d_next[230] ),
    .A_N(\u_inv.d_reg[230] ));
 sg13g2_nor2_1 _21170_ (.A(_13683_),
    .B(_13845_),
    .Y(_13846_));
 sg13g2_nand2b_1 _21171_ (.Y(_13847_),
    .B(\u_inv.d_next[228] ),
    .A_N(net4767));
 sg13g2_o21ai_1 _21172_ (.B1(_13688_),
    .Y(_13848_),
    .A1(_13689_),
    .A2(_13847_));
 sg13g2_a221oi_1 _21173_ (.B2(_13687_),
    .C1(_13846_),
    .B1(_13848_),
    .A1(_13695_),
    .Y(_13849_),
    .A2(_13844_));
 sg13g2_o21ai_1 _21174_ (.B1(_13849_),
    .Y(_13850_),
    .A1(_10579_),
    .A2(\u_inv.d_reg[231] ));
 sg13g2_nand2_1 _21175_ (.Y(_13851_),
    .A(\u_inv.d_next[238] ),
    .B(_10886_));
 sg13g2_nor2_1 _21176_ (.A(_13677_),
    .B(_13851_),
    .Y(_13852_));
 sg13g2_nand2b_1 _21177_ (.Y(_13853_),
    .B(\u_inv.d_next[239] ),
    .A_N(\u_inv.d_reg[239] ));
 sg13g2_nor2b_1 _21178_ (.A(\u_inv.d_reg[237] ),
    .B_N(\u_inv.d_next[237] ),
    .Y(_13854_));
 sg13g2_nor2b_1 _21179_ (.A(\u_inv.d_reg[236] ),
    .B_N(\u_inv.d_next[236] ),
    .Y(_13855_));
 sg13g2_a21o_1 _21180_ (.A2(_13855_),
    .A1(_13671_),
    .B1(_13854_),
    .X(_13856_));
 sg13g2_nor2_1 _21181_ (.A(_13675_),
    .B(_13838_),
    .Y(_13857_));
 sg13g2_o21ai_1 _21182_ (.B1(_13680_),
    .Y(_13858_),
    .A1(_13856_),
    .A2(_13857_));
 sg13g2_a21oi_1 _21183_ (.A1(_13681_),
    .A2(_13850_),
    .Y(_13859_),
    .B1(_13852_));
 sg13g2_nand3_1 _21184_ (.B(_13858_),
    .C(_13859_),
    .A(_13853_),
    .Y(_13860_));
 sg13g2_nor2b_1 _21185_ (.A(_13656_),
    .B_N(_13860_),
    .Y(_13861_));
 sg13g2_nor2b_1 _21186_ (.A(\u_inv.d_reg[243] ),
    .B_N(\u_inv.d_next[243] ),
    .Y(_13862_));
 sg13g2_nor2b_1 _21187_ (.A(\u_inv.d_reg[242] ),
    .B_N(\u_inv.d_next[242] ),
    .Y(_13863_));
 sg13g2_inv_1 _21188_ (.Y(_13864_),
    .A(_13863_));
 sg13g2_nor2b_1 _21189_ (.A(\u_inv.d_reg[240] ),
    .B_N(\u_inv.d_next[240] ),
    .Y(_13865_));
 sg13g2_o21ai_1 _21190_ (.B1(_13632_),
    .Y(_13866_),
    .A1(_13633_),
    .A2(_13865_));
 sg13g2_o21ai_1 _21191_ (.B1(_13864_),
    .Y(_13867_),
    .A1(_13631_),
    .A2(_13866_));
 sg13g2_a21oi_1 _21192_ (.A1(_13639_),
    .A2(_13867_),
    .Y(_13868_),
    .B1(_13862_));
 sg13g2_nor2_1 _21193_ (.A(_13652_),
    .B(_13868_),
    .Y(_13869_));
 sg13g2_nor2b_1 _21194_ (.A(\u_inv.d_reg[247] ),
    .B_N(\u_inv.d_next[247] ),
    .Y(_13870_));
 sg13g2_nand2b_1 _21195_ (.Y(_13871_),
    .B(\u_inv.d_next[246] ),
    .A_N(\u_inv.d_reg[246] ));
 sg13g2_nor2b_1 _21196_ (.A(\u_inv.d_reg[244] ),
    .B_N(\u_inv.d_next[244] ),
    .Y(_13872_));
 sg13g2_nand2_1 _21197_ (.Y(_13873_),
    .A(_13642_),
    .B(_13872_));
 sg13g2_o21ai_1 _21198_ (.B1(_13873_),
    .Y(_13874_),
    .A1(_10578_),
    .A2(\u_inv.d_reg[245] ));
 sg13g2_nand2_1 _21199_ (.Y(_13875_),
    .A(_13651_),
    .B(_13874_));
 sg13g2_a21oi_1 _21200_ (.A1(_13871_),
    .A2(_13875_),
    .Y(_13876_),
    .B1(_13647_));
 sg13g2_nor3_1 _21201_ (.A(_13869_),
    .B(_13870_),
    .C(_13876_),
    .Y(_13877_));
 sg13g2_nor2b_1 _21202_ (.A(_13877_),
    .B_N(_13628_),
    .Y(_13878_));
 sg13g2_nor2b_1 _21203_ (.A(\u_inv.d_reg[253] ),
    .B_N(\u_inv.d_next[253] ),
    .Y(_13879_));
 sg13g2_nor2b_1 _21204_ (.A(\u_inv.d_reg[252] ),
    .B_N(\u_inv.d_next[252] ),
    .Y(_13880_));
 sg13g2_a21oi_1 _21205_ (.A1(_13609_),
    .A2(_13880_),
    .Y(_13881_),
    .B1(_13879_));
 sg13g2_nor2b_1 _21206_ (.A(\u_inv.d_reg[254] ),
    .B_N(\u_inv.d_next[254] ),
    .Y(_13882_));
 sg13g2_nor2b_1 _21207_ (.A(\u_inv.d_reg[255] ),
    .B_N(\u_inv.d_next[255] ),
    .Y(_13883_));
 sg13g2_a21oi_1 _21208_ (.A1(_13602_),
    .A2(_13882_),
    .Y(_13884_),
    .B1(_13883_));
 sg13g2_o21ai_1 _21209_ (.B1(_13884_),
    .Y(_13885_),
    .A1(_13606_),
    .A2(_13881_));
 sg13g2_nor2b_1 _21210_ (.A(\u_inv.d_reg[251] ),
    .B_N(\u_inv.d_next[251] ),
    .Y(_13886_));
 sg13g2_nor2b_1 _21211_ (.A(\u_inv.d_reg[250] ),
    .B_N(\u_inv.d_next[250] ),
    .Y(_13887_));
 sg13g2_a21oi_1 _21212_ (.A1(_13616_),
    .A2(_13887_),
    .Y(_13888_),
    .B1(_13886_));
 sg13g2_nor2b_1 _21213_ (.A(\u_inv.d_reg[249] ),
    .B_N(\u_inv.d_next[249] ),
    .Y(_13889_));
 sg13g2_nor2b_1 _21214_ (.A(\u_inv.d_reg[248] ),
    .B_N(\u_inv.d_next[248] ),
    .Y(_13890_));
 sg13g2_a21o_1 _21215_ (.A2(_13890_),
    .A1(_13623_),
    .B1(_13889_),
    .X(_13891_));
 sg13g2_nand2b_1 _21216_ (.Y(_13892_),
    .B(_13891_),
    .A_N(_13620_));
 sg13g2_a21oi_1 _21217_ (.A1(_13888_),
    .A2(_13892_),
    .Y(_13893_),
    .B1(_13613_));
 sg13g2_nor3_2 _21218_ (.A(_13878_),
    .B(_13885_),
    .C(_13893_),
    .Y(_13894_));
 sg13g2_nor2b_1 _21219_ (.A(\u_inv.d_reg[192] ),
    .B_N(\u_inv.d_next[192] ),
    .Y(_13895_));
 sg13g2_a21oi_1 _21220_ (.A1(_13768_),
    .A2(_13895_),
    .Y(_13896_),
    .B1(_13767_));
 sg13g2_inv_1 _21221_ (.Y(_13897_),
    .A(_13896_));
 sg13g2_nor2b_1 _21222_ (.A(\u_inv.d_reg[194] ),
    .B_N(\u_inv.d_next[194] ),
    .Y(_13898_));
 sg13g2_o21ai_1 _21223_ (.B1(_13760_),
    .Y(_13899_),
    .A1(_13761_),
    .A2(_13898_));
 sg13g2_o21ai_1 _21224_ (.B1(_13899_),
    .Y(_13900_),
    .A1(_13766_),
    .A2(_13896_));
 sg13g2_nor2b_1 _21225_ (.A(net4771),
    .B_N(\u_inv.d_next[198] ),
    .Y(_13901_));
 sg13g2_a21oi_1 _21226_ (.A1(_13744_),
    .A2(_13901_),
    .Y(_13902_),
    .B1(_13743_));
 sg13g2_nor2b_1 _21227_ (.A(net4772),
    .B_N(\u_inv.d_next[197] ),
    .Y(_13903_));
 sg13g2_nor2b_1 _21228_ (.A(net4773),
    .B_N(\u_inv.d_next[196] ),
    .Y(_13904_));
 sg13g2_a21oi_1 _21229_ (.A1(_13754_),
    .A2(_13904_),
    .Y(_13905_),
    .B1(_13903_));
 sg13g2_o21ai_1 _21230_ (.B1(_13902_),
    .Y(_13906_),
    .A1(_13751_),
    .A2(_13905_));
 sg13g2_a21oi_2 _21231_ (.B1(_13906_),
    .Y(_13907_),
    .A2(_13900_),
    .A1(_13759_));
 sg13g2_nor2_1 _21232_ (.A(_13742_),
    .B(_13907_),
    .Y(_13908_));
 sg13g2_nor2b_1 _21233_ (.A(\u_inv.d_reg[204] ),
    .B_N(\u_inv.d_next[204] ),
    .Y(_13909_));
 sg13g2_nand2b_1 _21234_ (.Y(_13910_),
    .B(\u_inv.d_next[204] ),
    .A_N(\u_inv.d_reg[204] ));
 sg13g2_o21ai_1 _21235_ (.B1(_13719_),
    .Y(_13911_),
    .A1(_13720_),
    .A2(_13910_));
 sg13g2_nand2_1 _21236_ (.Y(_13912_),
    .A(_13718_),
    .B(_13911_));
 sg13g2_nor2b_1 _21237_ (.A(\u_inv.d_reg[207] ),
    .B_N(\u_inv.d_next[207] ),
    .Y(_13913_));
 sg13g2_nor2b_1 _21238_ (.A(\u_inv.d_reg[206] ),
    .B_N(\u_inv.d_next[206] ),
    .Y(_13914_));
 sg13g2_nand2b_1 _21239_ (.Y(_13915_),
    .B(\u_inv.d_next[206] ),
    .A_N(\u_inv.d_reg[206] ));
 sg13g2_a21oi_1 _21240_ (.A1(_13715_),
    .A2(_13914_),
    .Y(_13916_),
    .B1(_13913_));
 sg13g2_nand2_1 _21241_ (.Y(_13917_),
    .A(_13912_),
    .B(_13916_));
 sg13g2_nor2b_1 _21242_ (.A(\u_inv.d_reg[200] ),
    .B_N(\u_inv.d_next[200] ),
    .Y(_13918_));
 sg13g2_a21oi_1 _21243_ (.A1(\u_inv.d_next[201] ),
    .A2(_10896_),
    .Y(_13919_),
    .B1(_13918_));
 sg13g2_a21oi_2 _21244_ (.B1(_13919_),
    .Y(_13920_),
    .A2(\u_inv.d_reg[201] ),
    .A1(_10585_));
 sg13g2_nand2_1 _21245_ (.Y(_13921_),
    .A(_13741_),
    .B(_13920_));
 sg13g2_nand2b_1 _21246_ (.Y(_13922_),
    .B(\u_inv.d_next[202] ),
    .A_N(\u_inv.d_reg[202] ));
 sg13g2_a21o_2 _21247_ (.A2(_13922_),
    .A1(_13739_),
    .B1(_13738_),
    .X(_13923_));
 sg13g2_a21oi_1 _21248_ (.A1(_13921_),
    .A2(_13923_),
    .Y(_13924_),
    .B1(_13727_));
 sg13g2_nor3_2 _21249_ (.A(_13908_),
    .B(_13917_),
    .C(_13924_),
    .Y(_13925_));
 sg13g2_nand2b_1 _21250_ (.Y(_13926_),
    .B(\u_inv.d_next[219] ),
    .A_N(\u_inv.d_reg[219] ));
 sg13g2_nor2b_1 _21251_ (.A(\u_inv.d_reg[218] ),
    .B_N(\u_inv.d_next[218] ),
    .Y(_13927_));
 sg13g2_a22oi_1 _21252_ (.Y(_13928_),
    .B1(_10892_),
    .B2(\u_inv.d_next[216] ),
    .A2(_10891_),
    .A1(\u_inv.d_next[217] ));
 sg13g2_nor2_1 _21253_ (.A(_13794_),
    .B(_13928_),
    .Y(_13929_));
 sg13g2_a21oi_1 _21254_ (.A1(_13793_),
    .A2(_13929_),
    .Y(_13930_),
    .B1(_13927_));
 sg13g2_o21ai_1 _21255_ (.B1(_13926_),
    .Y(_13931_),
    .A1(_13797_),
    .A2(_13930_));
 sg13g2_nand2_1 _21256_ (.Y(_13932_),
    .A(\u_inv.d_next[222] ),
    .B(_10889_));
 sg13g2_nor2b_1 _21257_ (.A(\u_inv.d_reg[220] ),
    .B_N(\u_inv.d_next[220] ),
    .Y(_13933_));
 sg13g2_nand2_1 _21258_ (.Y(_13934_),
    .A(_13778_),
    .B(_13933_));
 sg13g2_o21ai_1 _21259_ (.B1(_13934_),
    .Y(_13935_),
    .A1(_10581_),
    .A2(\u_inv.d_reg[221] ));
 sg13g2_nand2b_1 _21260_ (.Y(_13936_),
    .B(_13935_),
    .A_N(_13785_));
 sg13g2_a21oi_1 _21261_ (.A1(_13932_),
    .A2(_13936_),
    .Y(_13937_),
    .B1(_13782_));
 sg13g2_a21o_1 _21262_ (.A2(_10888_),
    .A1(\u_inv.d_next[223] ),
    .B1(_13937_),
    .X(_13938_));
 sg13g2_nor2b_1 _21263_ (.A(net4770),
    .B_N(\u_inv.d_next[208] ),
    .Y(_13939_));
 sg13g2_a21o_1 _21264_ (.A2(_13939_),
    .A1(_13821_),
    .B1(_13820_),
    .X(_13940_));
 sg13g2_inv_1 _21265_ (.Y(_13941_),
    .A(_13940_));
 sg13g2_nand2_1 _21266_ (.Y(_13942_),
    .A(\u_inv.d_next[210] ),
    .B(_10895_));
 sg13g2_a22oi_1 _21267_ (.Y(_13943_),
    .B1(_10895_),
    .B2(\u_inv.d_next[210] ),
    .A2(_10894_),
    .A1(\u_inv.d_next[211] ));
 sg13g2_nor2_1 _21268_ (.A(_13814_),
    .B(_13943_),
    .Y(_13944_));
 sg13g2_a21oi_1 _21269_ (.A1(_13819_),
    .A2(_13940_),
    .Y(_13945_),
    .B1(_13944_));
 sg13g2_nor2b_1 _21270_ (.A(\u_inv.d_reg[215] ),
    .B_N(\u_inv.d_next[215] ),
    .Y(_13946_));
 sg13g2_nor2b_1 _21271_ (.A(\u_inv.d_reg[214] ),
    .B_N(\u_inv.d_next[214] ),
    .Y(_13947_));
 sg13g2_nand2b_1 _21272_ (.Y(_13948_),
    .B(\u_inv.d_next[214] ),
    .A_N(\u_inv.d_reg[214] ));
 sg13g2_nor2b_1 _21273_ (.A(\u_inv.d_reg[212] ),
    .B_N(\u_inv.d_next[212] ),
    .Y(_13949_));
 sg13g2_a21o_1 _21274_ (.A2(_13949_),
    .A1(_13806_),
    .B1(_13805_),
    .X(_13950_));
 sg13g2_a221oi_1 _21275_ (.B2(_13804_),
    .C1(_13946_),
    .B1(_13950_),
    .A1(_13801_),
    .Y(_13951_),
    .A2(_13947_));
 sg13g2_o21ai_1 _21276_ (.B1(_13951_),
    .Y(_13952_),
    .A1(_13813_),
    .A2(_13945_));
 sg13g2_inv_1 _21277_ (.Y(_13953_),
    .A(_13952_));
 sg13g2_o21ai_1 _21278_ (.B1(_13953_),
    .Y(_13954_),
    .A1(_13829_),
    .A2(_13925_));
 sg13g2_a221oi_1 _21279_ (.B2(_13799_),
    .C1(_13938_),
    .B1(_13954_),
    .A1(_13787_),
    .Y(_13955_),
    .A2(_13931_));
 sg13g2_nand2_1 _21280_ (.Y(_13956_),
    .A(\u_inv.d_next[15] ),
    .B(_10952_));
 sg13g2_nor2_1 _21281_ (.A(\u_inv.d_next[15] ),
    .B(_10952_),
    .Y(_13957_));
 sg13g2_xnor2_1 _21282_ (.Y(_13958_),
    .A(\u_inv.d_next[15] ),
    .B(\u_inv.d_reg[15] ));
 sg13g2_xor2_1 _21283_ (.B(\u_inv.d_reg[15] ),
    .A(\u_inv.d_next[15] ),
    .X(_13959_));
 sg13g2_nand2_1 _21284_ (.Y(_13960_),
    .A(\u_inv.d_next[14] ),
    .B(\u_inv.d_reg[14] ));
 sg13g2_xor2_1 _21285_ (.B(\u_inv.d_reg[14] ),
    .A(\u_inv.d_next[14] ),
    .X(_13961_));
 sg13g2_nor2_1 _21286_ (.A(_13959_),
    .B(_13961_),
    .Y(_13962_));
 sg13g2_nor2_1 _21287_ (.A(\u_inv.d_next[13] ),
    .B(\u_inv.d_reg[13] ),
    .Y(_13963_));
 sg13g2_xor2_1 _21288_ (.B(\u_inv.d_reg[13] ),
    .A(\u_inv.d_next[13] ),
    .X(_13964_));
 sg13g2_and2_1 _21289_ (.A(\u_inv.d_next[12] ),
    .B(\u_inv.d_reg[12] ),
    .X(_13965_));
 sg13g2_xor2_1 _21290_ (.B(\u_inv.d_reg[12] ),
    .A(\u_inv.d_next[12] ),
    .X(_13966_));
 sg13g2_nor2_1 _21291_ (.A(_13964_),
    .B(_13966_),
    .Y(_13967_));
 sg13g2_nand2_1 _21292_ (.Y(_13968_),
    .A(_13962_),
    .B(_13967_));
 sg13g2_nand2b_1 _21293_ (.Y(_13969_),
    .B(net4792),
    .A_N(\u_inv.d_next[11] ));
 sg13g2_nor2b_1 _21294_ (.A(net4792),
    .B_N(\u_inv.d_next[11] ),
    .Y(_13970_));
 sg13g2_xnor2_1 _21295_ (.Y(_13971_),
    .A(\u_inv.d_next[11] ),
    .B(net4792));
 sg13g2_inv_1 _21296_ (.Y(_13972_),
    .A(_13971_));
 sg13g2_nand2_1 _21297_ (.Y(_13973_),
    .A(\u_inv.d_next[10] ),
    .B(\u_inv.d_reg[10] ));
 sg13g2_xnor2_1 _21298_ (.Y(_13974_),
    .A(\u_inv.d_next[10] ),
    .B(\u_inv.d_reg[10] ));
 sg13g2_nand2_1 _21299_ (.Y(_13975_),
    .A(_13971_),
    .B(_13974_));
 sg13g2_nor2_1 _21300_ (.A(_13968_),
    .B(_13975_),
    .Y(_13976_));
 sg13g2_nand2b_1 _21301_ (.Y(_13977_),
    .B(net4794),
    .A_N(\u_inv.d_next[7] ));
 sg13g2_nand2b_1 _21302_ (.Y(_13978_),
    .B(\u_inv.d_next[7] ),
    .A_N(net4794));
 sg13g2_nand2b_1 _21303_ (.Y(_13979_),
    .B(net4806),
    .A_N(net4795));
 sg13g2_nand2_1 _21304_ (.Y(_13980_),
    .A(_13978_),
    .B(_13979_));
 sg13g2_nor2_1 _21305_ (.A(net4806),
    .B(net4795),
    .Y(_13981_));
 sg13g2_xor2_1 _21306_ (.B(net4795),
    .A(net4806),
    .X(_13982_));
 sg13g2_xnor2_1 _21307_ (.Y(_13983_),
    .A(net4806),
    .B(net4795));
 sg13g2_nor2_1 _21308_ (.A(_13980_),
    .B(_13983_),
    .Y(_13984_));
 sg13g2_a21oi_1 _21309_ (.A1(_10622_),
    .A2(net4794),
    .Y(_13985_),
    .B1(_13984_));
 sg13g2_nand2b_1 _21310_ (.Y(_13986_),
    .B(\u_inv.d_reg[5] ),
    .A_N(\u_inv.d_next[5] ));
 sg13g2_nor2b_1 _21311_ (.A(\u_inv.d_reg[3] ),
    .B_N(\u_inv.d_next[3] ),
    .Y(_13987_));
 sg13g2_xor2_1 _21312_ (.B(\u_inv.d_reg[3] ),
    .A(\u_inv.d_next[3] ),
    .X(_13988_));
 sg13g2_inv_1 _21313_ (.Y(_13989_),
    .A(_13988_));
 sg13g2_nand2b_1 _21314_ (.Y(_13990_),
    .B(\u_inv.d_next[2] ),
    .A_N(net4796));
 sg13g2_nand2_1 _21315_ (.Y(_13991_),
    .A(\u_inv.d_next[2] ),
    .B(net4796));
 sg13g2_nor2_1 _21316_ (.A(\u_inv.d_next[2] ),
    .B(net4796),
    .Y(_13992_));
 sg13g2_xor2_1 _21317_ (.B(net4796),
    .A(\u_inv.d_next[2] ),
    .X(_13993_));
 sg13g2_nor2b_1 _21318_ (.A(net4797),
    .B_N(\u_inv.d_next[1] ),
    .Y(_13994_));
 sg13g2_and2_1 _21319_ (.A(\u_inv.d_next[1] ),
    .B(net4797),
    .X(_13995_));
 sg13g2_or2_1 _21320_ (.X(_13996_),
    .B(net4797),
    .A(\u_inv.d_next[1] ));
 sg13g2_xnor2_1 _21321_ (.Y(_13997_),
    .A(\u_inv.d_next[1] ),
    .B(net4797));
 sg13g2_nand2b_1 _21322_ (.Y(_13998_),
    .B(net4799),
    .A_N(\u_inv.d_next[0] ));
 sg13g2_a21oi_1 _21323_ (.A1(_13997_),
    .A2(_13998_),
    .Y(_13999_),
    .B1(_13994_));
 sg13g2_o21ai_1 _21324_ (.B1(_13990_),
    .Y(_14000_),
    .A1(_13993_),
    .A2(_13999_));
 sg13g2_a21oi_2 _21325_ (.B1(_13987_),
    .Y(_14001_),
    .A2(_14000_),
    .A1(_13989_));
 sg13g2_and2_1 _21326_ (.A(\u_inv.d_next[4] ),
    .B(\u_inv.d_reg[4] ),
    .X(_14002_));
 sg13g2_xor2_1 _21327_ (.B(\u_inv.d_reg[4] ),
    .A(\u_inv.d_next[4] ),
    .X(_14003_));
 sg13g2_nor2_1 _21328_ (.A(_14001_),
    .B(_14003_),
    .Y(_14004_));
 sg13g2_nor2b_1 _21329_ (.A(\u_inv.d_reg[5] ),
    .B_N(\u_inv.d_next[5] ),
    .Y(_14005_));
 sg13g2_nor2b_1 _21330_ (.A(\u_inv.d_reg[4] ),
    .B_N(\u_inv.d_next[4] ),
    .Y(_14006_));
 sg13g2_xor2_1 _21331_ (.B(\u_inv.d_reg[5] ),
    .A(\u_inv.d_next[5] ),
    .X(_14007_));
 sg13g2_nor2_1 _21332_ (.A(_14003_),
    .B(_14007_),
    .Y(_14008_));
 sg13g2_inv_1 _21333_ (.Y(_14009_),
    .A(_14008_));
 sg13g2_nor2_1 _21334_ (.A(_14001_),
    .B(_14009_),
    .Y(_14010_));
 sg13g2_a21o_1 _21335_ (.A2(_14006_),
    .A1(_13986_),
    .B1(_14005_),
    .X(_14011_));
 sg13g2_or2_1 _21336_ (.X(_14012_),
    .B(_14011_),
    .A(_14010_));
 sg13g2_a21oi_1 _21337_ (.A1(_13977_),
    .A2(_13980_),
    .Y(_14013_),
    .B1(_14011_));
 sg13g2_o21ai_1 _21338_ (.B1(_14013_),
    .Y(_14014_),
    .A1(_14001_),
    .A2(_14009_));
 sg13g2_and2_1 _21339_ (.A(_13985_),
    .B(_14014_),
    .X(_14015_));
 sg13g2_xor2_1 _21340_ (.B(\u_inv.d_reg[9] ),
    .A(\u_inv.d_next[9] ),
    .X(_14016_));
 sg13g2_and2_1 _21341_ (.A(\u_inv.d_next[8] ),
    .B(\u_inv.d_reg[8] ),
    .X(_14017_));
 sg13g2_xor2_1 _21342_ (.B(\u_inv.d_reg[8] ),
    .A(\u_inv.d_next[8] ),
    .X(_14018_));
 sg13g2_nor2_1 _21343_ (.A(_14016_),
    .B(_14018_),
    .Y(_14019_));
 sg13g2_nand4_1 _21344_ (.B(_13985_),
    .C(_14014_),
    .A(_13976_),
    .Y(_14020_),
    .D(_14019_));
 sg13g2_a22oi_1 _21345_ (.Y(_14021_),
    .B1(_10956_),
    .B2(\u_inv.d_next[8] ),
    .A2(_10955_),
    .A1(\u_inv.d_next[9] ));
 sg13g2_a21oi_2 _21346_ (.B1(_14021_),
    .Y(_14022_),
    .A2(\u_inv.d_reg[9] ),
    .A1(_10621_));
 sg13g2_nor2b_1 _21347_ (.A(\u_inv.d_reg[10] ),
    .B_N(\u_inv.d_next[10] ),
    .Y(_14023_));
 sg13g2_o21ai_1 _21348_ (.B1(_13969_),
    .Y(_14024_),
    .A1(_13970_),
    .A2(_14023_));
 sg13g2_nor2_1 _21349_ (.A(_13968_),
    .B(_14024_),
    .Y(_14025_));
 sg13g2_nand2_1 _21350_ (.Y(_14026_),
    .A(\u_inv.d_next[14] ),
    .B(_10953_));
 sg13g2_o21ai_1 _21351_ (.B1(_13956_),
    .Y(_14027_),
    .A1(_13957_),
    .A2(_14026_));
 sg13g2_nand2b_1 _21352_ (.Y(_14028_),
    .B(\u_inv.d_next[13] ),
    .A_N(\u_inv.d_reg[13] ));
 sg13g2_nand2_1 _21353_ (.Y(_14029_),
    .A(\u_inv.d_next[12] ),
    .B(_10954_));
 sg13g2_o21ai_1 _21354_ (.B1(_14028_),
    .Y(_14030_),
    .A1(_13964_),
    .A2(_14029_));
 sg13g2_a221oi_1 _21355_ (.B2(_13962_),
    .C1(_14027_),
    .B1(_14030_),
    .A1(_13976_),
    .Y(_14031_),
    .A2(_14022_));
 sg13g2_nor2b_2 _21356_ (.A(_14025_),
    .B_N(_14031_),
    .Y(_14032_));
 sg13g2_and2_1 _21357_ (.A(_14020_),
    .B(_14032_),
    .X(_14033_));
 sg13g2_xnor2_1 _21358_ (.Y(_14034_),
    .A(\u_inv.d_next[31] ),
    .B(\u_inv.d_reg[31] ));
 sg13g2_xor2_1 _21359_ (.B(\u_inv.d_reg[31] ),
    .A(\u_inv.d_next[31] ),
    .X(_14035_));
 sg13g2_nand2_1 _21360_ (.Y(_14036_),
    .A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ));
 sg13g2_xor2_1 _21361_ (.B(\u_inv.d_reg[30] ),
    .A(\u_inv.d_next[30] ),
    .X(_14037_));
 sg13g2_xnor2_1 _21362_ (.Y(_14038_),
    .A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ));
 sg13g2_nor2_1 _21363_ (.A(_14035_),
    .B(_14037_),
    .Y(_14039_));
 sg13g2_xnor2_1 _21364_ (.Y(_14040_),
    .A(\u_inv.d_next[29] ),
    .B(\u_inv.d_reg[29] ));
 sg13g2_nand2_1 _21365_ (.Y(_14041_),
    .A(\u_inv.d_next[28] ),
    .B(\u_inv.d_reg[28] ));
 sg13g2_xnor2_1 _21366_ (.Y(_14042_),
    .A(\u_inv.d_next[28] ),
    .B(\u_inv.d_reg[28] ));
 sg13g2_inv_1 _21367_ (.Y(_14043_),
    .A(_14042_));
 sg13g2_and2_1 _21368_ (.A(_14040_),
    .B(_14042_),
    .X(_14044_));
 sg13g2_nand2_1 _21369_ (.Y(_14045_),
    .A(_14039_),
    .B(_14044_));
 sg13g2_nand2b_1 _21370_ (.Y(_14046_),
    .B(\u_inv.d_reg[27] ),
    .A_N(\u_inv.d_next[27] ));
 sg13g2_nand2b_1 _21371_ (.Y(_14047_),
    .B(\u_inv.d_next[27] ),
    .A_N(\u_inv.d_reg[27] ));
 sg13g2_and2_1 _21372_ (.A(_14046_),
    .B(_14047_),
    .X(_14048_));
 sg13g2_and2_1 _21373_ (.A(\u_inv.d_next[26] ),
    .B(net4787),
    .X(_14049_));
 sg13g2_nand2_1 _21374_ (.Y(_14050_),
    .A(\u_inv.d_next[26] ),
    .B(net4787));
 sg13g2_xor2_1 _21375_ (.B(net4787),
    .A(\u_inv.d_next[26] ),
    .X(_14051_));
 sg13g2_xnor2_1 _21376_ (.Y(_14052_),
    .A(\u_inv.d_next[26] ),
    .B(net4787));
 sg13g2_nand2_1 _21377_ (.Y(_14053_),
    .A(_14048_),
    .B(_14052_));
 sg13g2_nor2_1 _21378_ (.A(\u_inv.d_next[25] ),
    .B(net4788),
    .Y(_14054_));
 sg13g2_nand2_1 _21379_ (.Y(_14055_),
    .A(\u_inv.d_next[25] ),
    .B(net4788));
 sg13g2_xnor2_1 _21380_ (.Y(_14056_),
    .A(\u_inv.d_next[25] ),
    .B(net4788));
 sg13g2_nand2_1 _21381_ (.Y(_14057_),
    .A(\u_inv.d_next[24] ),
    .B(\u_inv.d_reg[24] ));
 sg13g2_xnor2_1 _21382_ (.Y(_14058_),
    .A(\u_inv.d_next[24] ),
    .B(\u_inv.d_reg[24] ));
 sg13g2_nand2_1 _21383_ (.Y(_14059_),
    .A(_14056_),
    .B(_14058_));
 sg13g2_or2_1 _21384_ (.X(_14060_),
    .B(_14059_),
    .A(_14053_));
 sg13g2_nor2_1 _21385_ (.A(_14045_),
    .B(_14060_),
    .Y(_14061_));
 sg13g2_nor2_1 _21386_ (.A(_10619_),
    .B(\u_inv.d_reg[19] ),
    .Y(_14062_));
 sg13g2_xor2_1 _21387_ (.B(\u_inv.d_reg[19] ),
    .A(\u_inv.d_next[19] ),
    .X(_14063_));
 sg13g2_xor2_1 _21388_ (.B(net4790),
    .A(\u_inv.d_next[18] ),
    .X(_14064_));
 sg13g2_xnor2_1 _21389_ (.Y(_14065_),
    .A(\u_inv.d_next[18] ),
    .B(net4790));
 sg13g2_nor2_1 _21390_ (.A(net4805),
    .B(_10950_),
    .Y(_14066_));
 sg13g2_nand2b_1 _21391_ (.Y(_14067_),
    .B(net4791),
    .A_N(net4805));
 sg13g2_xnor2_1 _21392_ (.Y(_14068_),
    .A(net4805),
    .B(net4791));
 sg13g2_xor2_1 _21393_ (.B(net4791),
    .A(net4805),
    .X(_14069_));
 sg13g2_nand2_1 _21394_ (.Y(_14070_),
    .A(\u_inv.d_next[16] ),
    .B(\u_inv.d_reg[16] ));
 sg13g2_xor2_1 _21395_ (.B(\u_inv.d_reg[16] ),
    .A(\u_inv.d_next[16] ),
    .X(_14071_));
 sg13g2_nor4_1 _21396_ (.A(_14063_),
    .B(_14064_),
    .C(_14069_),
    .D(_14071_),
    .Y(_14072_));
 sg13g2_inv_1 _21397_ (.Y(_14073_),
    .A(_14072_));
 sg13g2_nor2b_1 _21398_ (.A(\u_inv.d_next[23] ),
    .B_N(\u_inv.d_reg[23] ),
    .Y(_14074_));
 sg13g2_nand2b_1 _21399_ (.Y(_14075_),
    .B(\u_inv.d_next[23] ),
    .A_N(\u_inv.d_reg[23] ));
 sg13g2_xnor2_1 _21400_ (.Y(_14076_),
    .A(\u_inv.d_next[23] ),
    .B(\u_inv.d_reg[23] ));
 sg13g2_nand2b_1 _21401_ (.Y(_14077_),
    .B(_14075_),
    .A_N(_14074_));
 sg13g2_nand2_1 _21402_ (.Y(_14078_),
    .A(\u_inv.d_next[22] ),
    .B(net4789));
 sg13g2_nor2_1 _21403_ (.A(\u_inv.d_next[22] ),
    .B(net4789),
    .Y(_14079_));
 sg13g2_xor2_1 _21404_ (.B(net4789),
    .A(\u_inv.d_next[22] ),
    .X(_14080_));
 sg13g2_xnor2_1 _21405_ (.Y(_14081_),
    .A(\u_inv.d_next[22] ),
    .B(net4789));
 sg13g2_nor2_1 _21406_ (.A(_14077_),
    .B(_14080_),
    .Y(_14082_));
 sg13g2_nor2_1 _21407_ (.A(\u_inv.d_next[21] ),
    .B(\u_inv.d_reg[21] ),
    .Y(_14083_));
 sg13g2_xor2_1 _21408_ (.B(\u_inv.d_reg[21] ),
    .A(\u_inv.d_next[21] ),
    .X(_14084_));
 sg13g2_and2_1 _21409_ (.A(\u_inv.d_next[20] ),
    .B(\u_inv.d_reg[20] ),
    .X(_14085_));
 sg13g2_xor2_1 _21410_ (.B(\u_inv.d_reg[20] ),
    .A(\u_inv.d_next[20] ),
    .X(_14086_));
 sg13g2_nor2_1 _21411_ (.A(_14084_),
    .B(_14086_),
    .Y(_14087_));
 sg13g2_and2_1 _21412_ (.A(_14082_),
    .B(_14087_),
    .X(_14088_));
 sg13g2_nand3_1 _21413_ (.B(_14072_),
    .C(_14088_),
    .A(_14061_),
    .Y(_14089_));
 sg13g2_a21oi_2 _21414_ (.B1(_14089_),
    .Y(_14090_),
    .A2(_14032_),
    .A1(_14020_));
 sg13g2_a21o_2 _21415_ (.A2(_14032_),
    .A1(_14020_),
    .B1(_14089_),
    .X(_14091_));
 sg13g2_nand2b_1 _21416_ (.Y(_14092_),
    .B(\u_inv.d_next[22] ),
    .A_N(net4789));
 sg13g2_a21oi_1 _21417_ (.A1(_14075_),
    .A2(_14092_),
    .Y(_14093_),
    .B1(_14074_));
 sg13g2_nand2b_1 _21418_ (.Y(_14094_),
    .B(\u_inv.d_next[21] ),
    .A_N(\u_inv.d_reg[21] ));
 sg13g2_nand2b_1 _21419_ (.Y(_14095_),
    .B(\u_inv.d_next[20] ),
    .A_N(\u_inv.d_reg[20] ));
 sg13g2_o21ai_1 _21420_ (.B1(_14094_),
    .Y(_14096_),
    .A1(_14084_),
    .A2(_14095_));
 sg13g2_nor2b_1 _21421_ (.A(\u_inv.d_reg[16] ),
    .B_N(\u_inv.d_next[16] ),
    .Y(_14097_));
 sg13g2_a21oi_1 _21422_ (.A1(net4805),
    .A2(_10950_),
    .Y(_14098_),
    .B1(_14097_));
 sg13g2_nor4_1 _21423_ (.A(_14063_),
    .B(_14064_),
    .C(_14066_),
    .D(_14098_),
    .Y(_14099_));
 sg13g2_nand2b_1 _21424_ (.Y(_14100_),
    .B(\u_inv.d_next[18] ),
    .A_N(net4790));
 sg13g2_a21oi_1 _21425_ (.A1(_10619_),
    .A2(\u_inv.d_reg[19] ),
    .Y(_14101_),
    .B1(_14100_));
 sg13g2_nor3_1 _21426_ (.A(_14062_),
    .B(_14099_),
    .C(_14101_),
    .Y(_14102_));
 sg13g2_a21o_1 _21427_ (.A2(_14096_),
    .A1(_14082_),
    .B1(_14093_),
    .X(_14103_));
 sg13g2_nor2b_1 _21428_ (.A(_14102_),
    .B_N(_14088_),
    .Y(_14104_));
 sg13g2_o21ai_1 _21429_ (.B1(_14061_),
    .Y(_14105_),
    .A1(_14103_),
    .A2(_14104_));
 sg13g2_nor2b_1 _21430_ (.A(\u_inv.d_reg[28] ),
    .B_N(\u_inv.d_next[28] ),
    .Y(_14106_));
 sg13g2_nand2_1 _21431_ (.Y(_14107_),
    .A(_14040_),
    .B(_14106_));
 sg13g2_o21ai_1 _21432_ (.B1(_14107_),
    .Y(_14108_),
    .A1(_10618_),
    .A2(\u_inv.d_reg[29] ));
 sg13g2_nand2_1 _21433_ (.Y(_14109_),
    .A(\u_inv.d_next[30] ),
    .B(_10947_));
 sg13g2_a21oi_1 _21434_ (.A1(_10617_),
    .A2(\u_inv.d_reg[31] ),
    .Y(_14110_),
    .B1(_14109_));
 sg13g2_a221oi_1 _21435_ (.B2(_14108_),
    .C1(_14110_),
    .B1(_14039_),
    .A1(\u_inv.d_next[31] ),
    .Y(_14111_),
    .A2(_10946_));
 sg13g2_nor2b_1 _21436_ (.A(net4788),
    .B_N(\u_inv.d_next[25] ),
    .Y(_14112_));
 sg13g2_nor2b_1 _21437_ (.A(\u_inv.d_reg[24] ),
    .B_N(\u_inv.d_next[24] ),
    .Y(_14113_));
 sg13g2_a21oi_1 _21438_ (.A1(_14056_),
    .A2(_14113_),
    .Y(_14114_),
    .B1(_14112_));
 sg13g2_nor2b_1 _21439_ (.A(net4787),
    .B_N(\u_inv.d_next[26] ),
    .Y(_14115_));
 sg13g2_o21ai_1 _21440_ (.B1(_14047_),
    .Y(_14116_),
    .A1(_14053_),
    .A2(_14114_));
 sg13g2_a21oi_1 _21441_ (.A1(_14046_),
    .A2(_14115_),
    .Y(_14117_),
    .B1(_14116_));
 sg13g2_or2_1 _21442_ (.X(_14118_),
    .B(_14117_),
    .A(_14045_));
 sg13g2_and3_2 _21443_ (.X(_14119_),
    .A(_14105_),
    .B(_14111_),
    .C(_14118_));
 sg13g2_nand3_1 _21444_ (.B(_14111_),
    .C(_14118_),
    .A(_14105_),
    .Y(_14120_));
 sg13g2_nand2_1 _21445_ (.Y(_14121_),
    .A(_14091_),
    .B(_14119_));
 sg13g2_nor2_1 _21446_ (.A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ),
    .Y(_14122_));
 sg13g2_xnor2_1 _21447_ (.Y(_14123_),
    .A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ));
 sg13g2_nand2_1 _21448_ (.Y(_14124_),
    .A(\u_inv.d_next[62] ),
    .B(\u_inv.d_reg[62] ));
 sg13g2_xnor2_1 _21449_ (.Y(_14125_),
    .A(\u_inv.d_next[62] ),
    .B(\u_inv.d_reg[62] ));
 sg13g2_nand2_1 _21450_ (.Y(_14126_),
    .A(_14123_),
    .B(_14125_));
 sg13g2_xnor2_1 _21451_ (.Y(_14127_),
    .A(\u_inv.d_next[61] ),
    .B(\u_inv.d_reg[61] ));
 sg13g2_nand2_1 _21452_ (.Y(_14128_),
    .A(\u_inv.d_next[60] ),
    .B(\u_inv.d_reg[60] ));
 sg13g2_xor2_1 _21453_ (.B(\u_inv.d_reg[60] ),
    .A(\u_inv.d_next[60] ),
    .X(_14129_));
 sg13g2_nand2b_1 _21454_ (.Y(_14130_),
    .B(_14127_),
    .A_N(_14129_));
 sg13g2_or2_1 _21455_ (.X(_14131_),
    .B(_14130_),
    .A(_14126_));
 sg13g2_nand2b_1 _21456_ (.Y(_14132_),
    .B(\u_inv.d_reg[59] ),
    .A_N(\u_inv.d_next[59] ));
 sg13g2_nor2b_1 _21457_ (.A(\u_inv.d_reg[59] ),
    .B_N(\u_inv.d_next[59] ),
    .Y(_14133_));
 sg13g2_xnor2_1 _21458_ (.Y(_14134_),
    .A(\u_inv.d_next[59] ),
    .B(\u_inv.d_reg[59] ));
 sg13g2_xor2_1 _21459_ (.B(\u_inv.d_reg[59] ),
    .A(\u_inv.d_next[59] ),
    .X(_14135_));
 sg13g2_nand2_1 _21460_ (.Y(_14136_),
    .A(net4804),
    .B(net4785));
 sg13g2_xor2_1 _21461_ (.B(net4785),
    .A(net4804),
    .X(_14137_));
 sg13g2_xnor2_1 _21462_ (.Y(_14138_),
    .A(net4804),
    .B(net4785));
 sg13g2_nor2_1 _21463_ (.A(_14135_),
    .B(_14137_),
    .Y(_14139_));
 sg13g2_xor2_1 _21464_ (.B(\u_inv.d_reg[57] ),
    .A(\u_inv.d_next[57] ),
    .X(_14140_));
 sg13g2_and2_1 _21465_ (.A(\u_inv.d_next[56] ),
    .B(\u_inv.d_reg[56] ),
    .X(_14141_));
 sg13g2_xor2_1 _21466_ (.B(\u_inv.d_reg[56] ),
    .A(\u_inv.d_next[56] ),
    .X(_14142_));
 sg13g2_nor2_1 _21467_ (.A(_14140_),
    .B(_14142_),
    .Y(_14143_));
 sg13g2_inv_1 _21468_ (.Y(_14144_),
    .A(_14143_));
 sg13g2_nand2_1 _21469_ (.Y(_14145_),
    .A(_14139_),
    .B(_14143_));
 sg13g2_nor2b_1 _21470_ (.A(\u_inv.d_reg[55] ),
    .B_N(\u_inv.d_next[55] ),
    .Y(_14146_));
 sg13g2_nand2b_1 _21471_ (.Y(_14147_),
    .B(\u_inv.d_reg[55] ),
    .A_N(\u_inv.d_next[55] ));
 sg13g2_nor2b_2 _21472_ (.A(_14146_),
    .B_N(_14147_),
    .Y(_14148_));
 sg13g2_nand2b_1 _21473_ (.Y(_14149_),
    .B(_14147_),
    .A_N(_14146_));
 sg13g2_nand2_1 _21474_ (.Y(_14150_),
    .A(\u_inv.d_next[54] ),
    .B(\u_inv.d_reg[54] ));
 sg13g2_xor2_1 _21475_ (.B(\u_inv.d_reg[54] ),
    .A(\u_inv.d_next[54] ),
    .X(_14151_));
 sg13g2_xnor2_1 _21476_ (.Y(_14152_),
    .A(\u_inv.d_next[54] ),
    .B(\u_inv.d_reg[54] ));
 sg13g2_nand2_1 _21477_ (.Y(_14153_),
    .A(_14148_),
    .B(_14152_));
 sg13g2_nor2_1 _21478_ (.A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ),
    .Y(_14154_));
 sg13g2_nand2_1 _21479_ (.Y(_14155_),
    .A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ));
 sg13g2_nor2b_2 _21480_ (.A(_14154_),
    .B_N(_14155_),
    .Y(_14156_));
 sg13g2_xnor2_1 _21481_ (.Y(_14157_),
    .A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ));
 sg13g2_nand2_1 _21482_ (.Y(_14158_),
    .A(\u_inv.d_next[52] ),
    .B(\u_inv.d_reg[52] ));
 sg13g2_xor2_1 _21483_ (.B(\u_inv.d_reg[52] ),
    .A(\u_inv.d_next[52] ),
    .X(_14159_));
 sg13g2_xnor2_1 _21484_ (.Y(_14160_),
    .A(\u_inv.d_next[52] ),
    .B(\u_inv.d_reg[52] ));
 sg13g2_nand2_1 _21485_ (.Y(_14161_),
    .A(_14157_),
    .B(_14160_));
 sg13g2_nor2_1 _21486_ (.A(_14153_),
    .B(_14161_),
    .Y(_14162_));
 sg13g2_xnor2_1 _21487_ (.Y(_14163_),
    .A(\u_inv.d_next[51] ),
    .B(\u_inv.d_reg[51] ));
 sg13g2_nand2_1 _21488_ (.Y(_14164_),
    .A(\u_inv.d_next[50] ),
    .B(\u_inv.d_reg[50] ));
 sg13g2_xnor2_1 _21489_ (.Y(_14165_),
    .A(\u_inv.d_next[50] ),
    .B(\u_inv.d_reg[50] ));
 sg13g2_and2_1 _21490_ (.A(_14163_),
    .B(_14165_),
    .X(_14166_));
 sg13g2_nand2_1 _21491_ (.Y(_14167_),
    .A(_14163_),
    .B(_14165_));
 sg13g2_xnor2_1 _21492_ (.Y(_14168_),
    .A(\u_inv.d_next[49] ),
    .B(\u_inv.d_reg[49] ));
 sg13g2_xor2_1 _21493_ (.B(\u_inv.d_reg[49] ),
    .A(\u_inv.d_next[49] ),
    .X(_14169_));
 sg13g2_nand2_1 _21494_ (.Y(_14170_),
    .A(\u_inv.d_next[48] ),
    .B(\u_inv.d_reg[48] ));
 sg13g2_xor2_1 _21495_ (.B(\u_inv.d_reg[48] ),
    .A(\u_inv.d_next[48] ),
    .X(_14171_));
 sg13g2_nand2b_1 _21496_ (.Y(_14172_),
    .B(_14168_),
    .A_N(_14171_));
 sg13g2_or4_1 _21497_ (.A(_14153_),
    .B(_14161_),
    .C(_14167_),
    .D(_14172_),
    .X(_14173_));
 sg13g2_nor3_2 _21498_ (.A(_14131_),
    .B(_14145_),
    .C(_14173_),
    .Y(_14174_));
 sg13g2_xor2_1 _21499_ (.B(\u_inv.d_reg[47] ),
    .A(\u_inv.d_next[47] ),
    .X(_14175_));
 sg13g2_nand2_1 _21500_ (.Y(_14176_),
    .A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ));
 sg13g2_xor2_1 _21501_ (.B(\u_inv.d_reg[46] ),
    .A(\u_inv.d_next[46] ),
    .X(_14177_));
 sg13g2_xnor2_1 _21502_ (.Y(_14178_),
    .A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ));
 sg13g2_nor2_1 _21503_ (.A(_14175_),
    .B(_14177_),
    .Y(_14179_));
 sg13g2_nor2_1 _21504_ (.A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ),
    .Y(_14180_));
 sg13g2_xnor2_1 _21505_ (.Y(_14181_),
    .A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ));
 sg13g2_nand2_1 _21506_ (.Y(_14182_),
    .A(\u_inv.d_next[44] ),
    .B(\u_inv.d_reg[44] ));
 sg13g2_xnor2_1 _21507_ (.Y(_14183_),
    .A(\u_inv.d_next[44] ),
    .B(\u_inv.d_reg[44] ));
 sg13g2_and2_1 _21508_ (.A(_14181_),
    .B(_14183_),
    .X(_14184_));
 sg13g2_nand2_1 _21509_ (.Y(_14185_),
    .A(_14179_),
    .B(_14184_));
 sg13g2_nor2b_1 _21510_ (.A(\u_inv.d_reg[43] ),
    .B_N(\u_inv.d_next[43] ),
    .Y(_14186_));
 sg13g2_nand2b_1 _21511_ (.Y(_14187_),
    .B(\u_inv.d_reg[43] ),
    .A_N(\u_inv.d_next[43] ));
 sg13g2_xnor2_1 _21512_ (.Y(_14188_),
    .A(\u_inv.d_next[43] ),
    .B(\u_inv.d_reg[43] ));
 sg13g2_xor2_1 _21513_ (.B(\u_inv.d_reg[43] ),
    .A(\u_inv.d_next[43] ),
    .X(_14189_));
 sg13g2_nand2_1 _21514_ (.Y(_14190_),
    .A(\u_inv.d_next[42] ),
    .B(net4786));
 sg13g2_xnor2_1 _21515_ (.Y(_14191_),
    .A(\u_inv.d_next[42] ),
    .B(net4786));
 sg13g2_nand2_1 _21516_ (.Y(_14192_),
    .A(_14188_),
    .B(_14191_));
 sg13g2_inv_1 _21517_ (.Y(_14193_),
    .A(_14192_));
 sg13g2_or2_1 _21518_ (.X(_14194_),
    .B(\u_inv.d_reg[41] ),
    .A(\u_inv.d_next[41] ));
 sg13g2_and2_1 _21519_ (.A(\u_inv.d_next[41] ),
    .B(\u_inv.d_reg[41] ),
    .X(_14195_));
 sg13g2_xnor2_1 _21520_ (.Y(_14196_),
    .A(\u_inv.d_next[41] ),
    .B(\u_inv.d_reg[41] ));
 sg13g2_and2_1 _21521_ (.A(\u_inv.d_next[40] ),
    .B(\u_inv.d_reg[40] ),
    .X(_14197_));
 sg13g2_xor2_1 _21522_ (.B(\u_inv.d_reg[40] ),
    .A(\u_inv.d_next[40] ),
    .X(_14198_));
 sg13g2_xnor2_1 _21523_ (.Y(_14199_),
    .A(\u_inv.d_next[40] ),
    .B(\u_inv.d_reg[40] ));
 sg13g2_nand2_1 _21524_ (.Y(_14200_),
    .A(_14196_),
    .B(_14199_));
 sg13g2_nor3_1 _21525_ (.A(_14185_),
    .B(_14192_),
    .C(_14200_),
    .Y(_14201_));
 sg13g2_nand2b_1 _21526_ (.Y(_14202_),
    .B(\u_inv.d_next[39] ),
    .A_N(\u_inv.d_reg[39] ));
 sg13g2_nor2b_1 _21527_ (.A(\u_inv.d_next[39] ),
    .B_N(\u_inv.d_reg[39] ),
    .Y(_14203_));
 sg13g2_xnor2_1 _21528_ (.Y(_14204_),
    .A(\u_inv.d_next[39] ),
    .B(\u_inv.d_reg[39] ));
 sg13g2_xor2_1 _21529_ (.B(\u_inv.d_reg[39] ),
    .A(\u_inv.d_next[39] ),
    .X(_14205_));
 sg13g2_and2_1 _21530_ (.A(\u_inv.d_next[38] ),
    .B(\u_inv.d_reg[38] ),
    .X(_14206_));
 sg13g2_xor2_1 _21531_ (.B(\u_inv.d_reg[38] ),
    .A(\u_inv.d_next[38] ),
    .X(_14207_));
 sg13g2_xnor2_1 _21532_ (.Y(_14208_),
    .A(\u_inv.d_next[38] ),
    .B(\u_inv.d_reg[38] ));
 sg13g2_nor2_1 _21533_ (.A(_14205_),
    .B(_14207_),
    .Y(_14209_));
 sg13g2_nor2_1 _21534_ (.A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ),
    .Y(_14210_));
 sg13g2_nand2_1 _21535_ (.Y(_14211_),
    .A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ));
 sg13g2_nor2b_2 _21536_ (.A(_14210_),
    .B_N(_14211_),
    .Y(_14212_));
 sg13g2_xnor2_1 _21537_ (.Y(_14213_),
    .A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ));
 sg13g2_nand2_1 _21538_ (.Y(_14214_),
    .A(\u_inv.d_next[36] ),
    .B(\u_inv.d_reg[36] ));
 sg13g2_xor2_1 _21539_ (.B(\u_inv.d_reg[36] ),
    .A(\u_inv.d_next[36] ),
    .X(_14215_));
 sg13g2_xnor2_1 _21540_ (.Y(_14216_),
    .A(\u_inv.d_next[36] ),
    .B(\u_inv.d_reg[36] ));
 sg13g2_nand2_1 _21541_ (.Y(_14217_),
    .A(_14213_),
    .B(_14216_));
 sg13g2_nor3_1 _21542_ (.A(_14205_),
    .B(_14207_),
    .C(_14217_),
    .Y(_14218_));
 sg13g2_nor2b_1 _21543_ (.A(\u_inv.d_next[35] ),
    .B_N(\u_inv.d_reg[35] ),
    .Y(_14219_));
 sg13g2_nand2b_1 _21544_ (.Y(_14220_),
    .B(\u_inv.d_next[35] ),
    .A_N(\u_inv.d_reg[35] ));
 sg13g2_xnor2_1 _21545_ (.Y(_14221_),
    .A(\u_inv.d_next[35] ),
    .B(\u_inv.d_reg[35] ));
 sg13g2_nand2_1 _21546_ (.Y(_14222_),
    .A(\u_inv.d_next[34] ),
    .B(\u_inv.d_reg[34] ));
 sg13g2_nor2_1 _21547_ (.A(\u_inv.d_next[34] ),
    .B(\u_inv.d_reg[34] ),
    .Y(_14223_));
 sg13g2_xnor2_1 _21548_ (.Y(_14224_),
    .A(\u_inv.d_next[34] ),
    .B(\u_inv.d_reg[34] ));
 sg13g2_and2_1 _21549_ (.A(_14221_),
    .B(_14224_),
    .X(_14225_));
 sg13g2_nand2b_1 _21550_ (.Y(_14226_),
    .B(\u_inv.d_next[33] ),
    .A_N(\u_inv.d_reg[33] ));
 sg13g2_nor2b_1 _21551_ (.A(\u_inv.d_next[33] ),
    .B_N(\u_inv.d_reg[33] ),
    .Y(_14227_));
 sg13g2_xnor2_1 _21552_ (.Y(_14228_),
    .A(\u_inv.d_next[33] ),
    .B(\u_inv.d_reg[33] ));
 sg13g2_xor2_1 _21553_ (.B(\u_inv.d_reg[33] ),
    .A(\u_inv.d_next[33] ),
    .X(_14229_));
 sg13g2_and2_1 _21554_ (.A(\u_inv.d_next[32] ),
    .B(\u_inv.d_reg[32] ),
    .X(_14230_));
 sg13g2_xor2_1 _21555_ (.B(\u_inv.d_reg[32] ),
    .A(\u_inv.d_next[32] ),
    .X(_14231_));
 sg13g2_xnor2_1 _21556_ (.Y(_14232_),
    .A(\u_inv.d_next[32] ),
    .B(\u_inv.d_reg[32] ));
 sg13g2_nor2_1 _21557_ (.A(_14229_),
    .B(_14231_),
    .Y(_14233_));
 sg13g2_inv_1 _21558_ (.Y(_14234_),
    .A(_14233_));
 sg13g2_and3_1 _21559_ (.X(_14235_),
    .A(_14218_),
    .B(_14225_),
    .C(_14233_));
 sg13g2_and2_1 _21560_ (.A(_14201_),
    .B(_14235_),
    .X(_14236_));
 sg13g2_nand2_1 _21561_ (.Y(_14237_),
    .A(_14174_),
    .B(_14236_));
 sg13g2_a21oi_2 _21562_ (.B1(_14237_),
    .Y(_14238_),
    .A2(_14119_),
    .A1(_14091_));
 sg13g2_a21o_2 _21563_ (.A2(_14119_),
    .A1(_14091_),
    .B1(_14237_),
    .X(_14239_));
 sg13g2_nand2b_1 _21564_ (.Y(_14240_),
    .B(\u_inv.d_next[32] ),
    .A_N(\u_inv.d_reg[32] ));
 sg13g2_o21ai_1 _21565_ (.B1(_14226_),
    .Y(_14241_),
    .A1(_14227_),
    .A2(_14240_));
 sg13g2_nand2b_2 _21566_ (.Y(_14242_),
    .B(\u_inv.d_next[34] ),
    .A_N(\u_inv.d_reg[34] ));
 sg13g2_a21o_2 _21567_ (.A2(_14242_),
    .A1(_14220_),
    .B1(_14219_),
    .X(_14243_));
 sg13g2_a21oi_1 _21568_ (.A1(_14220_),
    .A2(_14242_),
    .Y(_14244_),
    .B1(_14219_));
 sg13g2_a21o_1 _21569_ (.A2(_14241_),
    .A1(_14225_),
    .B1(_14244_),
    .X(_14245_));
 sg13g2_nand2b_1 _21570_ (.Y(_14246_),
    .B(\u_inv.d_next[38] ),
    .A_N(\u_inv.d_reg[38] ));
 sg13g2_o21ai_1 _21571_ (.B1(_14202_),
    .Y(_14247_),
    .A1(_14203_),
    .A2(_14246_));
 sg13g2_nor2b_1 _21572_ (.A(\u_inv.d_reg[37] ),
    .B_N(\u_inv.d_next[37] ),
    .Y(_14248_));
 sg13g2_nor2b_1 _21573_ (.A(\u_inv.d_reg[36] ),
    .B_N(\u_inv.d_next[36] ),
    .Y(_14249_));
 sg13g2_a21o_1 _21574_ (.A2(_14249_),
    .A1(_14213_),
    .B1(_14248_),
    .X(_14250_));
 sg13g2_a221oi_1 _21575_ (.B2(_14209_),
    .C1(_14247_),
    .B1(_14250_),
    .A1(_14218_),
    .Y(_14251_),
    .A2(_14245_));
 sg13g2_nand2b_1 _21576_ (.Y(_14252_),
    .B(_14201_),
    .A_N(_14251_));
 sg13g2_nor2b_1 _21577_ (.A(\u_inv.d_reg[45] ),
    .B_N(\u_inv.d_next[45] ),
    .Y(_14253_));
 sg13g2_nor2b_1 _21578_ (.A(\u_inv.d_reg[44] ),
    .B_N(\u_inv.d_next[44] ),
    .Y(_14254_));
 sg13g2_a21o_1 _21579_ (.A2(_14254_),
    .A1(_14181_),
    .B1(_14253_),
    .X(_14255_));
 sg13g2_nand2_1 _21580_ (.Y(_14256_),
    .A(\u_inv.d_next[46] ),
    .B(_10943_));
 sg13g2_a21oi_1 _21581_ (.A1(_10615_),
    .A2(\u_inv.d_reg[47] ),
    .Y(_14257_),
    .B1(_14256_));
 sg13g2_a221oi_1 _21582_ (.B2(_14255_),
    .C1(_14257_),
    .B1(_14179_),
    .A1(\u_inv.d_next[47] ),
    .Y(_14258_),
    .A2(_10942_));
 sg13g2_nand2b_1 _21583_ (.Y(_14259_),
    .B(\u_inv.d_next[40] ),
    .A_N(\u_inv.d_reg[40] ));
 sg13g2_nor2b_1 _21584_ (.A(_14259_),
    .B_N(_14196_),
    .Y(_14260_));
 sg13g2_a21oi_1 _21585_ (.A1(\u_inv.d_next[41] ),
    .A2(_10944_),
    .Y(_14261_),
    .B1(_14260_));
 sg13g2_nor2b_1 _21586_ (.A(net4786),
    .B_N(\u_inv.d_next[42] ),
    .Y(_14262_));
 sg13g2_a21oi_1 _21587_ (.A1(_14187_),
    .A2(_14262_),
    .Y(_14263_),
    .B1(_14186_));
 sg13g2_o21ai_1 _21588_ (.B1(_14263_),
    .Y(_14264_),
    .A1(_14192_),
    .A2(_14261_));
 sg13g2_nand2b_1 _21589_ (.Y(_14265_),
    .B(_14264_),
    .A_N(_14185_));
 sg13g2_nand3_1 _21590_ (.B(_14258_),
    .C(_14265_),
    .A(_14252_),
    .Y(_14266_));
 sg13g2_inv_1 _21591_ (.Y(_14267_),
    .A(_14266_));
 sg13g2_nand2_1 _21592_ (.Y(_14268_),
    .A(_14174_),
    .B(_14266_));
 sg13g2_nor2b_1 _21593_ (.A(\u_inv.d_reg[56] ),
    .B_N(\u_inv.d_next[56] ),
    .Y(_14269_));
 sg13g2_a21oi_1 _21594_ (.A1(\u_inv.d_next[57] ),
    .A2(_10936_),
    .Y(_14270_),
    .B1(_14269_));
 sg13g2_a21oi_1 _21595_ (.A1(_10612_),
    .A2(\u_inv.d_reg[57] ),
    .Y(_14271_),
    .B1(_14270_));
 sg13g2_nor2b_1 _21596_ (.A(net4785),
    .B_N(\u_inv.d_next[58] ),
    .Y(_14272_));
 sg13g2_nand2_1 _21597_ (.Y(_14273_),
    .A(net4804),
    .B(_10935_));
 sg13g2_a21o_1 _21598_ (.A2(_14271_),
    .A1(_14139_),
    .B1(_14133_),
    .X(_14274_));
 sg13g2_a21oi_1 _21599_ (.A1(_14132_),
    .A2(_14272_),
    .Y(_14275_),
    .B1(_14274_));
 sg13g2_nor2_1 _21600_ (.A(_14131_),
    .B(_14275_),
    .Y(_14276_));
 sg13g2_nand2b_1 _21601_ (.Y(_14277_),
    .B(\u_inv.d_next[60] ),
    .A_N(\u_inv.d_reg[60] ));
 sg13g2_o21ai_1 _21602_ (.B1(_14277_),
    .Y(_14278_),
    .A1(_10611_),
    .A2(\u_inv.d_reg[61] ));
 sg13g2_o21ai_1 _21603_ (.B1(_14278_),
    .Y(_14279_),
    .A1(\u_inv.d_next[61] ),
    .A2(_10934_));
 sg13g2_nor2b_1 _21604_ (.A(\u_inv.d_reg[63] ),
    .B_N(\u_inv.d_next[63] ),
    .Y(_14280_));
 sg13g2_nor2b_1 _21605_ (.A(\u_inv.d_reg[62] ),
    .B_N(\u_inv.d_next[62] ),
    .Y(_14281_));
 sg13g2_a21oi_1 _21606_ (.A1(_14123_),
    .A2(_14281_),
    .Y(_14282_),
    .B1(_14280_));
 sg13g2_o21ai_1 _21607_ (.B1(_14282_),
    .Y(_14283_),
    .A1(_14126_),
    .A2(_14279_));
 sg13g2_nor2_1 _21608_ (.A(_14276_),
    .B(_14283_),
    .Y(_14284_));
 sg13g2_nand2b_1 _21609_ (.Y(_14285_),
    .B(\u_inv.d_next[48] ),
    .A_N(\u_inv.d_reg[48] ));
 sg13g2_o21ai_1 _21610_ (.B1(_14285_),
    .Y(_14286_),
    .A1(_10614_),
    .A2(\u_inv.d_reg[49] ));
 sg13g2_o21ai_1 _21611_ (.B1(_14286_),
    .Y(_14287_),
    .A1(\u_inv.d_next[49] ),
    .A2(_10941_));
 sg13g2_nor2_1 _21612_ (.A(_14167_),
    .B(_14287_),
    .Y(_14288_));
 sg13g2_nor2b_1 _21613_ (.A(\u_inv.d_reg[50] ),
    .B_N(\u_inv.d_next[50] ),
    .Y(_14289_));
 sg13g2_o21ai_1 _21614_ (.B1(_14289_),
    .Y(_14290_),
    .A1(\u_inv.d_next[51] ),
    .A2(_10939_));
 sg13g2_o21ai_1 _21615_ (.B1(_14290_),
    .Y(_14291_),
    .A1(_10613_),
    .A2(\u_inv.d_reg[51] ));
 sg13g2_o21ai_1 _21616_ (.B1(_14162_),
    .Y(_14292_),
    .A1(_14288_),
    .A2(_14291_));
 sg13g2_nor2b_1 _21617_ (.A(\u_inv.d_reg[54] ),
    .B_N(\u_inv.d_next[54] ),
    .Y(_14293_));
 sg13g2_a21oi_1 _21618_ (.A1(_14147_),
    .A2(_14293_),
    .Y(_14294_),
    .B1(_14146_));
 sg13g2_nand2_1 _21619_ (.Y(_14295_),
    .A(\u_inv.d_next[52] ),
    .B(_10938_));
 sg13g2_nor2_1 _21620_ (.A(_14156_),
    .B(_14295_),
    .Y(_14296_));
 sg13g2_a21oi_1 _21621_ (.A1(\u_inv.d_next[53] ),
    .A2(_10937_),
    .Y(_14297_),
    .B1(_14296_));
 sg13g2_o21ai_1 _21622_ (.B1(_14294_),
    .Y(_14298_),
    .A1(_14153_),
    .A2(_14297_));
 sg13g2_nor2b_2 _21623_ (.A(_14298_),
    .B_N(_14292_),
    .Y(_14299_));
 sg13g2_or3_1 _21624_ (.A(_14131_),
    .B(_14145_),
    .C(_14299_),
    .X(_14300_));
 sg13g2_and3_2 _21625_ (.X(_14301_),
    .A(_14268_),
    .B(_14284_),
    .C(_14300_));
 sg13g2_nand3_1 _21626_ (.B(_14284_),
    .C(_14300_),
    .A(_14268_),
    .Y(_14302_));
 sg13g2_nor2_1 _21627_ (.A(_14238_),
    .B(_14302_),
    .Y(_14303_));
 sg13g2_xnor2_1 _21628_ (.Y(_14304_),
    .A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ));
 sg13g2_nand2_1 _21629_ (.Y(_14305_),
    .A(\u_inv.d_next[126] ),
    .B(\u_inv.d_reg[126] ));
 sg13g2_xnor2_1 _21630_ (.Y(_14306_),
    .A(\u_inv.d_next[126] ),
    .B(\u_inv.d_reg[126] ));
 sg13g2_nand2_1 _21631_ (.Y(_14307_),
    .A(_14304_),
    .B(_14306_));
 sg13g2_nand2_1 _21632_ (.Y(_14308_),
    .A(\u_inv.d_next[125] ),
    .B(\u_inv.d_reg[125] ));
 sg13g2_xnor2_1 _21633_ (.Y(_14309_),
    .A(\u_inv.d_next[125] ),
    .B(\u_inv.d_reg[125] ));
 sg13g2_inv_1 _21634_ (.Y(_14310_),
    .A(_14309_));
 sg13g2_nand2_1 _21635_ (.Y(_14311_),
    .A(\u_inv.d_next[124] ),
    .B(\u_inv.d_reg[124] ));
 sg13g2_xor2_1 _21636_ (.B(\u_inv.d_reg[124] ),
    .A(\u_inv.d_next[124] ),
    .X(_14312_));
 sg13g2_inv_1 _21637_ (.Y(_14313_),
    .A(_14312_));
 sg13g2_nand2_1 _21638_ (.Y(_14314_),
    .A(_14309_),
    .B(_14313_));
 sg13g2_nor2_1 _21639_ (.A(_14307_),
    .B(_14314_),
    .Y(_14315_));
 sg13g2_and2_1 _21640_ (.A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ),
    .X(_14316_));
 sg13g2_xor2_1 _21641_ (.B(\u_inv.d_reg[122] ),
    .A(\u_inv.d_next[122] ),
    .X(_14317_));
 sg13g2_xnor2_1 _21642_ (.Y(_14318_),
    .A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ));
 sg13g2_nand2_1 _21643_ (.Y(_14319_),
    .A(\u_inv.d_next[123] ),
    .B(\u_inv.d_reg[123] ));
 sg13g2_xor2_1 _21644_ (.B(\u_inv.d_reg[123] ),
    .A(\u_inv.d_next[123] ),
    .X(_14320_));
 sg13g2_xnor2_1 _21645_ (.Y(_14321_),
    .A(\u_inv.d_next[123] ),
    .B(\u_inv.d_reg[123] ));
 sg13g2_nor2_1 _21646_ (.A(_14317_),
    .B(_14320_),
    .Y(_14322_));
 sg13g2_xnor2_1 _21647_ (.Y(_14323_),
    .A(\u_inv.d_next[121] ),
    .B(\u_inv.d_reg[121] ));
 sg13g2_nand2_1 _21648_ (.Y(_14324_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_xnor2_1 _21649_ (.Y(_14325_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_nand2_1 _21650_ (.Y(_14326_),
    .A(_14323_),
    .B(_14325_));
 sg13g2_nand4_1 _21651_ (.B(_14322_),
    .C(_14323_),
    .A(_14315_),
    .Y(_14327_),
    .D(_14325_));
 sg13g2_nor2b_1 _21652_ (.A(\u_inv.d_next[117] ),
    .B_N(\u_inv.d_reg[117] ),
    .Y(_14328_));
 sg13g2_nand2b_1 _21653_ (.Y(_14329_),
    .B(\u_inv.d_next[117] ),
    .A_N(\u_inv.d_reg[117] ));
 sg13g2_xnor2_1 _21654_ (.Y(_14330_),
    .A(\u_inv.d_next[117] ),
    .B(\u_inv.d_reg[117] ));
 sg13g2_nand2_1 _21655_ (.Y(_14331_),
    .A(\u_inv.d_next[116] ),
    .B(\u_inv.d_reg[116] ));
 sg13g2_xnor2_1 _21656_ (.Y(_14332_),
    .A(\u_inv.d_next[116] ),
    .B(\u_inv.d_reg[116] ));
 sg13g2_and2_1 _21657_ (.A(_14330_),
    .B(_14332_),
    .X(_14333_));
 sg13g2_xor2_1 _21658_ (.B(\u_inv.d_reg[119] ),
    .A(\u_inv.d_next[119] ),
    .X(_14334_));
 sg13g2_and2_1 _21659_ (.A(\u_inv.d_next[118] ),
    .B(\u_inv.d_reg[118] ),
    .X(_14335_));
 sg13g2_xor2_1 _21660_ (.B(\u_inv.d_reg[118] ),
    .A(\u_inv.d_next[118] ),
    .X(_14336_));
 sg13g2_xnor2_1 _21661_ (.Y(_14337_),
    .A(\u_inv.d_next[118] ),
    .B(\u_inv.d_reg[118] ));
 sg13g2_nor2_1 _21662_ (.A(_14334_),
    .B(_14336_),
    .Y(_14338_));
 sg13g2_and2_1 _21663_ (.A(_14333_),
    .B(_14338_),
    .X(_14339_));
 sg13g2_nand2b_1 _21664_ (.Y(_14340_),
    .B(\u_inv.d_reg[115] ),
    .A_N(\u_inv.d_next[115] ));
 sg13g2_nand2b_1 _21665_ (.Y(_14341_),
    .B(\u_inv.d_next[115] ),
    .A_N(\u_inv.d_reg[115] ));
 sg13g2_xnor2_1 _21666_ (.Y(_14342_),
    .A(\u_inv.d_next[115] ),
    .B(\u_inv.d_reg[115] ));
 sg13g2_nand2_1 _21667_ (.Y(_14343_),
    .A(_14340_),
    .B(_14341_));
 sg13g2_nand2_1 _21668_ (.Y(_14344_),
    .A(\u_inv.d_next[114] ),
    .B(\u_inv.d_reg[114] ));
 sg13g2_xnor2_1 _21669_ (.Y(_14345_),
    .A(\u_inv.d_next[114] ),
    .B(\u_inv.d_reg[114] ));
 sg13g2_inv_1 _21670_ (.Y(_14346_),
    .A(_14345_));
 sg13g2_nand2_1 _21671_ (.Y(_14347_),
    .A(_14342_),
    .B(_14345_));
 sg13g2_nor2b_1 _21672_ (.A(\u_inv.d_reg[113] ),
    .B_N(\u_inv.d_next[113] ),
    .Y(_14348_));
 sg13g2_nand2b_1 _21673_ (.Y(_14349_),
    .B(\u_inv.d_reg[113] ),
    .A_N(\u_inv.d_next[113] ));
 sg13g2_xnor2_1 _21674_ (.Y(_14350_),
    .A(\u_inv.d_next[113] ),
    .B(\u_inv.d_reg[113] ));
 sg13g2_nand2b_1 _21675_ (.Y(_14351_),
    .B(_14349_),
    .A_N(_14348_));
 sg13g2_nand2_1 _21676_ (.Y(_14352_),
    .A(\u_inv.d_next[112] ),
    .B(\u_inv.d_reg[112] ));
 sg13g2_xor2_1 _21677_ (.B(\u_inv.d_reg[112] ),
    .A(\u_inv.d_next[112] ),
    .X(_14353_));
 sg13g2_inv_1 _21678_ (.Y(_14354_),
    .A(_14353_));
 sg13g2_nor2_1 _21679_ (.A(_14351_),
    .B(_14353_),
    .Y(_14355_));
 sg13g2_nand4_1 _21680_ (.B(_14342_),
    .C(_14345_),
    .A(_14339_),
    .Y(_14356_),
    .D(_14355_));
 sg13g2_inv_1 _21681_ (.Y(_14357_),
    .A(_14356_));
 sg13g2_nor2_2 _21682_ (.A(_14327_),
    .B(_14356_),
    .Y(_14358_));
 sg13g2_xor2_1 _21683_ (.B(\u_inv.d_reg[111] ),
    .A(\u_inv.d_next[111] ),
    .X(_14359_));
 sg13g2_and2_1 _21684_ (.A(\u_inv.d_next[110] ),
    .B(\u_inv.d_reg[110] ),
    .X(_14360_));
 sg13g2_xor2_1 _21685_ (.B(\u_inv.d_reg[110] ),
    .A(\u_inv.d_next[110] ),
    .X(_14361_));
 sg13g2_xnor2_1 _21686_ (.Y(_14362_),
    .A(\u_inv.d_next[110] ),
    .B(\u_inv.d_reg[110] ));
 sg13g2_nor2_1 _21687_ (.A(_14359_),
    .B(_14361_),
    .Y(_14363_));
 sg13g2_xnor2_1 _21688_ (.Y(_14364_),
    .A(\u_inv.d_next[109] ),
    .B(\u_inv.d_reg[109] ));
 sg13g2_nand2_1 _21689_ (.Y(_14365_),
    .A(\u_inv.d_next[108] ),
    .B(\u_inv.d_reg[108] ));
 sg13g2_xnor2_1 _21690_ (.Y(_14366_),
    .A(\u_inv.d_next[108] ),
    .B(\u_inv.d_reg[108] ));
 sg13g2_and2_1 _21691_ (.A(_14364_),
    .B(_14366_),
    .X(_14367_));
 sg13g2_nand2_1 _21692_ (.Y(_14368_),
    .A(_14363_),
    .B(_14367_));
 sg13g2_nand2b_1 _21693_ (.Y(_14369_),
    .B(\u_inv.d_reg[107] ),
    .A_N(\u_inv.d_next[107] ));
 sg13g2_nand2b_1 _21694_ (.Y(_14370_),
    .B(\u_inv.d_next[107] ),
    .A_N(\u_inv.d_reg[107] ));
 sg13g2_xor2_1 _21695_ (.B(\u_inv.d_reg[107] ),
    .A(\u_inv.d_next[107] ),
    .X(_14371_));
 sg13g2_and2_1 _21696_ (.A(\u_inv.d_next[106] ),
    .B(\u_inv.d_reg[106] ),
    .X(_14372_));
 sg13g2_nand2_1 _21697_ (.Y(_14373_),
    .A(\u_inv.d_next[106] ),
    .B(\u_inv.d_reg[106] ));
 sg13g2_xor2_1 _21698_ (.B(\u_inv.d_reg[106] ),
    .A(\u_inv.d_next[106] ),
    .X(_14374_));
 sg13g2_or2_1 _21699_ (.X(_14375_),
    .B(_14374_),
    .A(_14371_));
 sg13g2_xor2_1 _21700_ (.B(\u_inv.d_reg[105] ),
    .A(\u_inv.d_next[105] ),
    .X(_14376_));
 sg13g2_and2_1 _21701_ (.A(\u_inv.d_next[104] ),
    .B(net4780),
    .X(_14377_));
 sg13g2_xor2_1 _21702_ (.B(net4780),
    .A(\u_inv.d_next[104] ),
    .X(_14378_));
 sg13g2_xnor2_1 _21703_ (.Y(_14379_),
    .A(\u_inv.d_next[104] ),
    .B(net4780));
 sg13g2_nor2_1 _21704_ (.A(_14376_),
    .B(_14378_),
    .Y(_14380_));
 sg13g2_nor4_1 _21705_ (.A(_14368_),
    .B(_14375_),
    .C(_14376_),
    .D(_14378_),
    .Y(_14381_));
 sg13g2_xnor2_1 _21706_ (.Y(_14382_),
    .A(\u_inv.d_next[103] ),
    .B(\u_inv.d_reg[103] ));
 sg13g2_xor2_1 _21707_ (.B(\u_inv.d_reg[103] ),
    .A(\u_inv.d_next[103] ),
    .X(_14383_));
 sg13g2_nand2_1 _21708_ (.Y(_14384_),
    .A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ));
 sg13g2_xor2_1 _21709_ (.B(\u_inv.d_reg[102] ),
    .A(\u_inv.d_next[102] ),
    .X(_14385_));
 sg13g2_xnor2_1 _21710_ (.Y(_14386_),
    .A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ));
 sg13g2_nor2_1 _21711_ (.A(_14383_),
    .B(_14385_),
    .Y(_14387_));
 sg13g2_nor2_1 _21712_ (.A(\u_inv.d_next[101] ),
    .B(\u_inv.d_reg[101] ),
    .Y(_14388_));
 sg13g2_xnor2_1 _21713_ (.Y(_14389_),
    .A(\u_inv.d_next[101] ),
    .B(\u_inv.d_reg[101] ));
 sg13g2_nand2_1 _21714_ (.Y(_14390_),
    .A(\u_inv.d_next[100] ),
    .B(\u_inv.d_reg[100] ));
 sg13g2_xnor2_1 _21715_ (.Y(_14391_),
    .A(\u_inv.d_next[100] ),
    .B(\u_inv.d_reg[100] ));
 sg13g2_and2_1 _21716_ (.A(_14389_),
    .B(_14391_),
    .X(_14392_));
 sg13g2_nand2_1 _21717_ (.Y(_14393_),
    .A(_14387_),
    .B(_14392_));
 sg13g2_nand2b_1 _21718_ (.Y(_14394_),
    .B(\u_inv.d_reg[99] ),
    .A_N(\u_inv.d_next[99] ));
 sg13g2_nor2b_1 _21719_ (.A(\u_inv.d_reg[99] ),
    .B_N(\u_inv.d_next[99] ),
    .Y(_14395_));
 sg13g2_xnor2_1 _21720_ (.Y(_14396_),
    .A(\u_inv.d_next[99] ),
    .B(\u_inv.d_reg[99] ));
 sg13g2_xor2_1 _21721_ (.B(\u_inv.d_reg[99] ),
    .A(\u_inv.d_next[99] ),
    .X(_14397_));
 sg13g2_nand2_1 _21722_ (.Y(_14398_),
    .A(\u_inv.d_next[98] ),
    .B(\u_inv.d_reg[98] ));
 sg13g2_xor2_1 _21723_ (.B(\u_inv.d_reg[98] ),
    .A(\u_inv.d_next[98] ),
    .X(_14399_));
 sg13g2_nand2b_1 _21724_ (.Y(_14400_),
    .B(_14396_),
    .A_N(_14399_));
 sg13g2_nor2b_1 _21725_ (.A(\u_inv.d_reg[97] ),
    .B_N(\u_inv.d_next[97] ),
    .Y(_14401_));
 sg13g2_nand2b_1 _21726_ (.Y(_14402_),
    .B(\u_inv.d_reg[97] ),
    .A_N(\u_inv.d_next[97] ));
 sg13g2_xor2_1 _21727_ (.B(\u_inv.d_reg[97] ),
    .A(\u_inv.d_next[97] ),
    .X(_14403_));
 sg13g2_and2_1 _21728_ (.A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ),
    .X(_14404_));
 sg13g2_xnor2_1 _21729_ (.Y(_14405_),
    .A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ));
 sg13g2_nand2b_1 _21730_ (.Y(_14406_),
    .B(_14405_),
    .A_N(_14403_));
 sg13g2_nor3_1 _21731_ (.A(_14393_),
    .B(_14400_),
    .C(_14406_),
    .Y(_14407_));
 sg13g2_inv_1 _21732_ (.Y(_14408_),
    .A(_14407_));
 sg13g2_and2_1 _21733_ (.A(_14381_),
    .B(_14407_),
    .X(_14409_));
 sg13g2_inv_1 _21734_ (.Y(_14410_),
    .A(_14409_));
 sg13g2_and2_1 _21735_ (.A(_14358_),
    .B(_14409_),
    .X(_14411_));
 sg13g2_nor2_1 _21736_ (.A(\u_inv.d_next[95] ),
    .B(\u_inv.d_reg[95] ),
    .Y(_14412_));
 sg13g2_xor2_1 _21737_ (.B(\u_inv.d_reg[95] ),
    .A(\u_inv.d_next[95] ),
    .X(_14413_));
 sg13g2_xnor2_1 _21738_ (.Y(_14414_),
    .A(\u_inv.d_next[95] ),
    .B(\u_inv.d_reg[95] ));
 sg13g2_nand2_1 _21739_ (.Y(_14415_),
    .A(\u_inv.d_next[94] ),
    .B(\u_inv.d_reg[94] ));
 sg13g2_xor2_1 _21740_ (.B(\u_inv.d_reg[94] ),
    .A(\u_inv.d_next[94] ),
    .X(_14416_));
 sg13g2_inv_1 _21741_ (.Y(_14417_),
    .A(_14416_));
 sg13g2_nor2_1 _21742_ (.A(_14413_),
    .B(_14416_),
    .Y(_14418_));
 sg13g2_nor2b_1 _21743_ (.A(\u_inv.d_reg[93] ),
    .B_N(\u_inv.d_next[93] ),
    .Y(_14419_));
 sg13g2_nand2b_1 _21744_ (.Y(_14420_),
    .B(\u_inv.d_reg[93] ),
    .A_N(\u_inv.d_next[93] ));
 sg13g2_nor2b_1 _21745_ (.A(_14419_),
    .B_N(_14420_),
    .Y(_14421_));
 sg13g2_xor2_1 _21746_ (.B(\u_inv.d_reg[93] ),
    .A(\u_inv.d_next[93] ),
    .X(_14422_));
 sg13g2_and2_1 _21747_ (.A(\u_inv.d_next[92] ),
    .B(\u_inv.d_reg[92] ),
    .X(_14423_));
 sg13g2_xnor2_1 _21748_ (.Y(_14424_),
    .A(\u_inv.d_next[92] ),
    .B(\u_inv.d_reg[92] ));
 sg13g2_nor2b_1 _21749_ (.A(_14422_),
    .B_N(_14424_),
    .Y(_14425_));
 sg13g2_nand2_1 _21750_ (.Y(_14426_),
    .A(_14418_),
    .B(_14425_));
 sg13g2_nand2b_1 _21751_ (.Y(_14427_),
    .B(\u_inv.d_reg[91] ),
    .A_N(\u_inv.d_next[91] ));
 sg13g2_nand2b_1 _21752_ (.Y(_14428_),
    .B(\u_inv.d_next[91] ),
    .A_N(\u_inv.d_reg[91] ));
 sg13g2_xnor2_1 _21753_ (.Y(_14429_),
    .A(\u_inv.d_next[91] ),
    .B(\u_inv.d_reg[91] ));
 sg13g2_nand2_1 _21754_ (.Y(_14430_),
    .A(_14427_),
    .B(_14428_));
 sg13g2_nand2_1 _21755_ (.Y(_14431_),
    .A(\u_inv.d_next[90] ),
    .B(\u_inv.d_reg[90] ));
 sg13g2_xnor2_1 _21756_ (.Y(_14432_),
    .A(\u_inv.d_next[90] ),
    .B(\u_inv.d_reg[90] ));
 sg13g2_inv_1 _21757_ (.Y(_14433_),
    .A(_14432_));
 sg13g2_nand2_1 _21758_ (.Y(_14434_),
    .A(_14429_),
    .B(_14432_));
 sg13g2_nor2b_1 _21759_ (.A(\u_inv.d_reg[89] ),
    .B_N(\u_inv.d_next[89] ),
    .Y(_14435_));
 sg13g2_nand2b_1 _21760_ (.Y(_14436_),
    .B(\u_inv.d_reg[89] ),
    .A_N(\u_inv.d_next[89] ));
 sg13g2_nor2b_2 _21761_ (.A(_14435_),
    .B_N(_14436_),
    .Y(_14437_));
 sg13g2_nand2b_2 _21762_ (.Y(_14438_),
    .B(_14436_),
    .A_N(_14435_));
 sg13g2_and2_1 _21763_ (.A(\u_inv.d_next[88] ),
    .B(\u_inv.d_reg[88] ),
    .X(_14439_));
 sg13g2_xor2_1 _21764_ (.B(\u_inv.d_reg[88] ),
    .A(\u_inv.d_next[88] ),
    .X(_14440_));
 sg13g2_xnor2_1 _21765_ (.Y(_14441_),
    .A(\u_inv.d_next[88] ),
    .B(\u_inv.d_reg[88] ));
 sg13g2_nor2_1 _21766_ (.A(_14438_),
    .B(_14440_),
    .Y(_14442_));
 sg13g2_nor4_1 _21767_ (.A(_14426_),
    .B(_14434_),
    .C(_14438_),
    .D(_14440_),
    .Y(_14443_));
 sg13g2_nor2b_1 _21768_ (.A(\u_inv.d_reg[87] ),
    .B_N(\u_inv.d_next[87] ),
    .Y(_14444_));
 sg13g2_nand2b_1 _21769_ (.Y(_14445_),
    .B(\u_inv.d_reg[87] ),
    .A_N(\u_inv.d_next[87] ));
 sg13g2_xnor2_1 _21770_ (.Y(_14446_),
    .A(\u_inv.d_next[87] ),
    .B(\u_inv.d_reg[87] ));
 sg13g2_nand2_1 _21771_ (.Y(_14447_),
    .A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ));
 sg13g2_nor2_1 _21772_ (.A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ),
    .Y(_14448_));
 sg13g2_xnor2_1 _21773_ (.Y(_14449_),
    .A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ));
 sg13g2_nand2_1 _21774_ (.Y(_14450_),
    .A(_14446_),
    .B(_14449_));
 sg13g2_nor2_1 _21775_ (.A(\u_inv.d_next[85] ),
    .B(\u_inv.d_reg[85] ),
    .Y(_14451_));
 sg13g2_xor2_1 _21776_ (.B(\u_inv.d_reg[85] ),
    .A(\u_inv.d_next[85] ),
    .X(_14452_));
 sg13g2_and2_1 _21777_ (.A(\u_inv.d_next[84] ),
    .B(\u_inv.d_reg[84] ),
    .X(_14453_));
 sg13g2_xor2_1 _21778_ (.B(\u_inv.d_reg[84] ),
    .A(\u_inv.d_next[84] ),
    .X(_14454_));
 sg13g2_or2_1 _21779_ (.X(_14455_),
    .B(_14454_),
    .A(_14452_));
 sg13g2_nor2_1 _21780_ (.A(_14450_),
    .B(_14455_),
    .Y(_14456_));
 sg13g2_nor2b_1 _21781_ (.A(\u_inv.d_next[83] ),
    .B_N(\u_inv.d_reg[83] ),
    .Y(_14457_));
 sg13g2_nand2b_1 _21782_ (.Y(_14458_),
    .B(\u_inv.d_next[83] ),
    .A_N(\u_inv.d_reg[83] ));
 sg13g2_xnor2_1 _21783_ (.Y(_14459_),
    .A(\u_inv.d_next[83] ),
    .B(\u_inv.d_reg[83] ));
 sg13g2_nand2_1 _21784_ (.Y(_14460_),
    .A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ));
 sg13g2_xor2_1 _21785_ (.B(\u_inv.d_reg[82] ),
    .A(\u_inv.d_next[82] ),
    .X(_14461_));
 sg13g2_xnor2_1 _21786_ (.Y(_14462_),
    .A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ));
 sg13g2_and2_1 _21787_ (.A(_14459_),
    .B(_14462_),
    .X(_14463_));
 sg13g2_nor2b_1 _21788_ (.A(\u_inv.d_reg[81] ),
    .B_N(\u_inv.d_next[81] ),
    .Y(_14464_));
 sg13g2_nand2b_1 _21789_ (.Y(_14465_),
    .B(\u_inv.d_reg[81] ),
    .A_N(\u_inv.d_next[81] ));
 sg13g2_xnor2_1 _21790_ (.Y(_14466_),
    .A(\u_inv.d_next[81] ),
    .B(\u_inv.d_reg[81] ));
 sg13g2_nand2_1 _21791_ (.Y(_14467_),
    .A(\u_inv.d_next[80] ),
    .B(\u_inv.d_reg[80] ));
 sg13g2_xor2_1 _21792_ (.B(\u_inv.d_reg[80] ),
    .A(\u_inv.d_next[80] ),
    .X(_14468_));
 sg13g2_inv_2 _21793_ (.Y(_14469_),
    .A(_14468_));
 sg13g2_nor2b_1 _21794_ (.A(_14468_),
    .B_N(_14466_),
    .Y(_14470_));
 sg13g2_inv_1 _21795_ (.Y(_14471_),
    .A(_14470_));
 sg13g2_and3_1 _21796_ (.X(_14472_),
    .A(_14456_),
    .B(_14463_),
    .C(_14470_));
 sg13g2_inv_1 _21797_ (.Y(_14473_),
    .A(_14472_));
 sg13g2_nand2_1 _21798_ (.Y(_14474_),
    .A(_14443_),
    .B(_14472_));
 sg13g2_nor2b_1 _21799_ (.A(\u_inv.d_reg[79] ),
    .B_N(\u_inv.d_next[79] ),
    .Y(_14475_));
 sg13g2_nand2b_1 _21800_ (.Y(_14476_),
    .B(\u_inv.d_reg[79] ),
    .A_N(\u_inv.d_next[79] ));
 sg13g2_xnor2_1 _21801_ (.Y(_14477_),
    .A(\u_inv.d_next[79] ),
    .B(\u_inv.d_reg[79] ));
 sg13g2_nor2_1 _21802_ (.A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ),
    .Y(_14478_));
 sg13g2_nand2_1 _21803_ (.Y(_14479_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_xnor2_1 _21804_ (.Y(_14480_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_and2_1 _21805_ (.A(_14477_),
    .B(_14480_),
    .X(_14481_));
 sg13g2_nor2_1 _21806_ (.A(\u_inv.d_next[77] ),
    .B(net4781),
    .Y(_14482_));
 sg13g2_xor2_1 _21807_ (.B(net4781),
    .A(\u_inv.d_next[77] ),
    .X(_14483_));
 sg13g2_xnor2_1 _21808_ (.Y(_14484_),
    .A(\u_inv.d_next[77] ),
    .B(net4781));
 sg13g2_nand2_1 _21809_ (.Y(_14485_),
    .A(\u_inv.d_next[76] ),
    .B(net4782));
 sg13g2_xor2_1 _21810_ (.B(net4782),
    .A(\u_inv.d_next[76] ),
    .X(_14486_));
 sg13g2_xnor2_1 _21811_ (.Y(_14487_),
    .A(\u_inv.d_next[76] ),
    .B(net4782));
 sg13g2_nand2_1 _21812_ (.Y(_14488_),
    .A(_14484_),
    .B(_14487_));
 sg13g2_nand3_1 _21813_ (.B(_14484_),
    .C(_14487_),
    .A(_14481_),
    .Y(_14489_));
 sg13g2_xnor2_1 _21814_ (.Y(_14490_),
    .A(\u_inv.d_next[75] ),
    .B(\u_inv.d_reg[75] ));
 sg13g2_xor2_1 _21815_ (.B(\u_inv.d_reg[75] ),
    .A(\u_inv.d_next[75] ),
    .X(_14491_));
 sg13g2_nand2_1 _21816_ (.Y(_14492_),
    .A(\u_inv.d_next[74] ),
    .B(\u_inv.d_reg[74] ));
 sg13g2_nor2_1 _21817_ (.A(\u_inv.d_next[74] ),
    .B(\u_inv.d_reg[74] ),
    .Y(_14493_));
 sg13g2_xor2_1 _21818_ (.B(\u_inv.d_reg[74] ),
    .A(\u_inv.d_next[74] ),
    .X(_14494_));
 sg13g2_xnor2_1 _21819_ (.Y(_14495_),
    .A(\u_inv.d_next[74] ),
    .B(\u_inv.d_reg[74] ));
 sg13g2_nor2_1 _21820_ (.A(_14491_),
    .B(_14494_),
    .Y(_14496_));
 sg13g2_nor2_2 _21821_ (.A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ),
    .Y(_14497_));
 sg13g2_and2_1 _21822_ (.A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ),
    .X(_14498_));
 sg13g2_nor2_2 _21823_ (.A(_14497_),
    .B(_14498_),
    .Y(_14499_));
 sg13g2_xnor2_1 _21824_ (.Y(_14500_),
    .A(\u_inv.d_next[72] ),
    .B(net4783));
 sg13g2_o21ai_1 _21825_ (.B1(_14500_),
    .Y(_14501_),
    .A1(_14497_),
    .A2(_14498_));
 sg13g2_or4_1 _21826_ (.A(_14489_),
    .B(_14491_),
    .C(_14494_),
    .D(_14501_),
    .X(_14502_));
 sg13g2_inv_1 _21827_ (.Y(_14503_),
    .A(_14502_));
 sg13g2_nor2b_1 _21828_ (.A(\u_inv.d_reg[71] ),
    .B_N(\u_inv.d_next[71] ),
    .Y(_14504_));
 sg13g2_nand2b_1 _21829_ (.Y(_14505_),
    .B(\u_inv.d_reg[71] ),
    .A_N(\u_inv.d_next[71] ));
 sg13g2_xnor2_1 _21830_ (.Y(_14506_),
    .A(\u_inv.d_next[71] ),
    .B(\u_inv.d_reg[71] ));
 sg13g2_nand2_1 _21831_ (.Y(_14507_),
    .A(\u_inv.d_next[70] ),
    .B(\u_inv.d_reg[70] ));
 sg13g2_nor2_1 _21832_ (.A(\u_inv.d_next[70] ),
    .B(\u_inv.d_reg[70] ),
    .Y(_14508_));
 sg13g2_xnor2_1 _21833_ (.Y(_14509_),
    .A(\u_inv.d_next[70] ),
    .B(\u_inv.d_reg[70] ));
 sg13g2_and2_1 _21834_ (.A(_14506_),
    .B(_14509_),
    .X(_14510_));
 sg13g2_nor2_1 _21835_ (.A(net4803),
    .B(\u_inv.d_reg[69] ),
    .Y(_14511_));
 sg13g2_xor2_1 _21836_ (.B(\u_inv.d_reg[69] ),
    .A(net4803),
    .X(_14512_));
 sg13g2_xnor2_1 _21837_ (.Y(_14513_),
    .A(net4803),
    .B(\u_inv.d_reg[69] ));
 sg13g2_xor2_1 _21838_ (.B(\u_inv.d_reg[68] ),
    .A(\u_inv.d_next[68] ),
    .X(_14514_));
 sg13g2_or2_1 _21839_ (.X(_14515_),
    .B(_14514_),
    .A(_14512_));
 sg13g2_nand3b_1 _21840_ (.B(_14510_),
    .C(_14513_),
    .Y(_14516_),
    .A_N(_14514_));
 sg13g2_xnor2_1 _21841_ (.Y(_14517_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_nand2_1 _21842_ (.Y(_14518_),
    .A(\u_inv.d_next[66] ),
    .B(\u_inv.d_reg[66] ));
 sg13g2_nor2_1 _21843_ (.A(\u_inv.d_next[66] ),
    .B(\u_inv.d_reg[66] ),
    .Y(_14519_));
 sg13g2_xnor2_1 _21844_ (.Y(_14520_),
    .A(\u_inv.d_next[66] ),
    .B(\u_inv.d_reg[66] ));
 sg13g2_and2_1 _21845_ (.A(_14517_),
    .B(_14520_),
    .X(_14521_));
 sg13g2_nand2_1 _21846_ (.Y(_14522_),
    .A(_14517_),
    .B(_14520_));
 sg13g2_nor2b_1 _21847_ (.A(\u_inv.d_reg[65] ),
    .B_N(\u_inv.d_next[65] ),
    .Y(_14523_));
 sg13g2_nand2b_1 _21848_ (.Y(_14524_),
    .B(\u_inv.d_reg[65] ),
    .A_N(\u_inv.d_next[65] ));
 sg13g2_nor2b_2 _21849_ (.A(_14523_),
    .B_N(_14524_),
    .Y(_14525_));
 sg13g2_xor2_1 _21850_ (.B(\u_inv.d_reg[65] ),
    .A(\u_inv.d_next[65] ),
    .X(_14526_));
 sg13g2_and2_1 _21851_ (.A(\u_inv.d_next[64] ),
    .B(net4784),
    .X(_14527_));
 sg13g2_nand2_1 _21852_ (.Y(_14528_),
    .A(\u_inv.d_next[64] ),
    .B(net4784));
 sg13g2_xor2_1 _21853_ (.B(net4784),
    .A(\u_inv.d_next[64] ),
    .X(_14529_));
 sg13g2_xnor2_1 _21854_ (.Y(_14530_),
    .A(\u_inv.d_next[64] ),
    .B(net4784));
 sg13g2_nand2_1 _21855_ (.Y(_14531_),
    .A(_14525_),
    .B(_14530_));
 sg13g2_or3_1 _21856_ (.A(_14516_),
    .B(_14522_),
    .C(_14531_),
    .X(_14532_));
 sg13g2_or2_1 _21857_ (.X(_14533_),
    .B(_14532_),
    .A(_14502_));
 sg13g2_nor2_2 _21858_ (.A(_14474_),
    .B(_14533_),
    .Y(_14534_));
 sg13g2_nand2_1 _21859_ (.Y(_14535_),
    .A(_14411_),
    .B(_14534_));
 sg13g2_a21oi_2 _21860_ (.B1(_14535_),
    .Y(_14536_),
    .A2(_14301_),
    .A1(_14239_));
 sg13g2_a21o_2 _21861_ (.A2(_14301_),
    .A1(_14239_),
    .B1(_14535_),
    .X(_14537_));
 sg13g2_nor2b_1 _21862_ (.A(net4784),
    .B_N(\u_inv.d_next[64] ),
    .Y(_14538_));
 sg13g2_a21oi_1 _21863_ (.A1(_14524_),
    .A2(_14538_),
    .Y(_14539_),
    .B1(_14523_));
 sg13g2_nor2_1 _21864_ (.A(_14522_),
    .B(_14539_),
    .Y(_14540_));
 sg13g2_nor2b_1 _21865_ (.A(\u_inv.d_reg[66] ),
    .B_N(\u_inv.d_next[66] ),
    .Y(_14541_));
 sg13g2_o21ai_1 _21866_ (.B1(_14541_),
    .Y(_14542_),
    .A1(\u_inv.d_next[67] ),
    .A2(_10933_));
 sg13g2_o21ai_1 _21867_ (.B1(_14542_),
    .Y(_14543_),
    .A1(_10610_),
    .A2(\u_inv.d_reg[67] ));
 sg13g2_nor2_1 _21868_ (.A(_14540_),
    .B(_14543_),
    .Y(_14544_));
 sg13g2_nor2_1 _21869_ (.A(_14516_),
    .B(_14544_),
    .Y(_14545_));
 sg13g2_nor2b_1 _21870_ (.A(\u_inv.d_reg[70] ),
    .B_N(\u_inv.d_next[70] ),
    .Y(_14546_));
 sg13g2_nand2b_1 _21871_ (.Y(_14547_),
    .B(\u_inv.d_next[68] ),
    .A_N(\u_inv.d_reg[68] ));
 sg13g2_nor2_1 _21872_ (.A(_14512_),
    .B(_14547_),
    .Y(_14548_));
 sg13g2_a21oi_1 _21873_ (.A1(net4803),
    .A2(_10932_),
    .Y(_14549_),
    .B1(_14548_));
 sg13g2_a21o_1 _21874_ (.A2(_10932_),
    .A1(net4803),
    .B1(_14548_),
    .X(_14550_));
 sg13g2_a221oi_1 _21875_ (.B2(_14510_),
    .C1(_14504_),
    .B1(_14550_),
    .A1(_14505_),
    .Y(_14551_),
    .A2(_14546_));
 sg13g2_nor2b_1 _21876_ (.A(_14545_),
    .B_N(_14551_),
    .Y(_14552_));
 sg13g2_o21ai_1 _21877_ (.B1(_14551_),
    .Y(_14553_),
    .A1(_14516_),
    .A2(_14544_));
 sg13g2_nand2b_1 _21878_ (.Y(_14554_),
    .B(\u_inv.d_next[77] ),
    .A_N(net4781));
 sg13g2_nand2_1 _21879_ (.Y(_14555_),
    .A(\u_inv.d_next[76] ),
    .B(_10930_));
 sg13g2_o21ai_1 _21880_ (.B1(_14554_),
    .Y(_14556_),
    .A1(_14483_),
    .A2(_14555_));
 sg13g2_inv_1 _21881_ (.Y(_14557_),
    .A(_14556_));
 sg13g2_nor2b_1 _21882_ (.A(\u_inv.d_reg[78] ),
    .B_N(\u_inv.d_next[78] ),
    .Y(_14558_));
 sg13g2_a221oi_1 _21883_ (.B2(_14476_),
    .C1(_14475_),
    .B1(_14558_),
    .A1(_14481_),
    .Y(_14559_),
    .A2(_14556_));
 sg13g2_nand2b_1 _21884_ (.Y(_14560_),
    .B(\u_inv.d_next[73] ),
    .A_N(\u_inv.d_reg[73] ));
 sg13g2_nor2b_1 _21885_ (.A(net4783),
    .B_N(\u_inv.d_next[72] ),
    .Y(_14561_));
 sg13g2_nand2b_1 _21886_ (.Y(_14562_),
    .B(\u_inv.d_next[72] ),
    .A_N(net4783));
 sg13g2_o21ai_1 _21887_ (.B1(_14560_),
    .Y(_14563_),
    .A1(_14499_),
    .A2(_14562_));
 sg13g2_nand2b_1 _21888_ (.Y(_14564_),
    .B(\u_inv.d_next[74] ),
    .A_N(\u_inv.d_reg[74] ));
 sg13g2_a21oi_1 _21889_ (.A1(_10609_),
    .A2(\u_inv.d_reg[75] ),
    .Y(_14565_),
    .B1(_14564_));
 sg13g2_a221oi_1 _21890_ (.B2(_14563_),
    .C1(_14565_),
    .B1(_14496_),
    .A1(\u_inv.d_next[75] ),
    .Y(_14566_),
    .A2(_10931_));
 sg13g2_inv_1 _21891_ (.Y(_14567_),
    .A(_14566_));
 sg13g2_o21ai_1 _21892_ (.B1(_14559_),
    .Y(_14568_),
    .A1(_14489_),
    .A2(_14566_));
 sg13g2_a21oi_2 _21893_ (.B1(_14568_),
    .Y(_14569_),
    .A2(_14553_),
    .A1(_14503_));
 sg13g2_nor2b_1 _21894_ (.A(\u_inv.d_reg[88] ),
    .B_N(\u_inv.d_next[88] ),
    .Y(_14570_));
 sg13g2_a21oi_1 _21895_ (.A1(_14436_),
    .A2(_14570_),
    .Y(_14571_),
    .B1(_14435_));
 sg13g2_nor2b_1 _21896_ (.A(\u_inv.d_reg[90] ),
    .B_N(\u_inv.d_next[90] ),
    .Y(_14572_));
 sg13g2_o21ai_1 _21897_ (.B1(_14428_),
    .Y(_14573_),
    .A1(_14434_),
    .A2(_14571_));
 sg13g2_a21oi_1 _21898_ (.A1(_14427_),
    .A2(_14572_),
    .Y(_14574_),
    .B1(_14573_));
 sg13g2_nor2b_1 _21899_ (.A(\u_inv.d_reg[92] ),
    .B_N(\u_inv.d_next[92] ),
    .Y(_14575_));
 sg13g2_a21o_1 _21900_ (.A2(_14575_),
    .A1(_14420_),
    .B1(_14419_),
    .X(_14576_));
 sg13g2_nand2b_1 _21901_ (.Y(_14577_),
    .B(\u_inv.d_next[94] ),
    .A_N(\u_inv.d_reg[94] ));
 sg13g2_nor2_1 _21902_ (.A(_14413_),
    .B(_14577_),
    .Y(_14578_));
 sg13g2_nor2b_1 _21903_ (.A(\u_inv.d_reg[80] ),
    .B_N(\u_inv.d_next[80] ),
    .Y(_14579_));
 sg13g2_a21o_1 _21904_ (.A2(_14579_),
    .A1(_14465_),
    .B1(_14464_),
    .X(_14580_));
 sg13g2_nand2b_1 _21905_ (.Y(_14581_),
    .B(\u_inv.d_next[82] ),
    .A_N(\u_inv.d_reg[82] ));
 sg13g2_o21ai_1 _21906_ (.B1(_14458_),
    .Y(_14582_),
    .A1(_14457_),
    .A2(_14581_));
 sg13g2_a21o_1 _21907_ (.A2(_14580_),
    .A1(_14463_),
    .B1(_14582_),
    .X(_14583_));
 sg13g2_nor2b_1 _21908_ (.A(\u_inv.d_reg[86] ),
    .B_N(\u_inv.d_next[86] ),
    .Y(_14584_));
 sg13g2_nand2b_1 _21909_ (.Y(_14585_),
    .B(\u_inv.d_next[84] ),
    .A_N(\u_inv.d_reg[84] ));
 sg13g2_nor2_1 _21910_ (.A(_14452_),
    .B(_14585_),
    .Y(_14586_));
 sg13g2_a21oi_1 _21911_ (.A1(\u_inv.d_next[85] ),
    .A2(_10929_),
    .Y(_14587_),
    .B1(_14586_));
 sg13g2_a221oi_1 _21912_ (.B2(_14445_),
    .C1(_14444_),
    .B1(_14584_),
    .A1(_14456_),
    .Y(_14588_),
    .A2(_14583_));
 sg13g2_o21ai_1 _21913_ (.B1(_14588_),
    .Y(_14589_),
    .A1(_14450_),
    .A2(_14587_));
 sg13g2_a22oi_1 _21914_ (.Y(_14590_),
    .B1(_14418_),
    .B2(_14576_),
    .A2(_10927_),
    .A1(\u_inv.d_next[95] ));
 sg13g2_o21ai_1 _21915_ (.B1(_14590_),
    .Y(_14591_),
    .A1(_14426_),
    .A2(_14574_));
 sg13g2_a21oi_1 _21916_ (.A1(_14443_),
    .A2(_14589_),
    .Y(_14592_),
    .B1(_14591_));
 sg13g2_o21ai_1 _21917_ (.B1(_14592_),
    .Y(_14593_),
    .A1(_14474_),
    .A2(_14569_));
 sg13g2_nor2_2 _21918_ (.A(_14578_),
    .B(_14593_),
    .Y(_14594_));
 sg13g2_o21ai_1 _21919_ (.B1(_14411_),
    .Y(_14595_),
    .A1(_14578_),
    .A2(_14593_));
 sg13g2_nor2b_1 _21920_ (.A(\u_inv.d_reg[112] ),
    .B_N(\u_inv.d_next[112] ),
    .Y(_14596_));
 sg13g2_a21oi_1 _21921_ (.A1(_14349_),
    .A2(_14596_),
    .Y(_14597_),
    .B1(_14348_));
 sg13g2_nor2_1 _21922_ (.A(_10603_),
    .B(\u_inv.d_reg[114] ),
    .Y(_14598_));
 sg13g2_o21ai_1 _21923_ (.B1(_14341_),
    .Y(_14599_),
    .A1(_14347_),
    .A2(_14597_));
 sg13g2_a21oi_1 _21924_ (.A1(_14340_),
    .A2(_14598_),
    .Y(_14600_),
    .B1(_14599_));
 sg13g2_nor2b_1 _21925_ (.A(_14600_),
    .B_N(_14339_),
    .Y(_14601_));
 sg13g2_nand2b_1 _21926_ (.Y(_14602_),
    .B(\u_inv.d_next[116] ),
    .A_N(\u_inv.d_reg[116] ));
 sg13g2_o21ai_1 _21927_ (.B1(_14329_),
    .Y(_14603_),
    .A1(_14328_),
    .A2(_14602_));
 sg13g2_nor2b_1 _21928_ (.A(\u_inv.d_reg[119] ),
    .B_N(\u_inv.d_next[119] ),
    .Y(_14604_));
 sg13g2_nand2b_1 _21929_ (.Y(_14605_),
    .B(\u_inv.d_next[118] ),
    .A_N(\u_inv.d_reg[118] ));
 sg13g2_nand2_1 _21930_ (.Y(_14606_),
    .A(_14337_),
    .B(_14603_));
 sg13g2_a21oi_1 _21931_ (.A1(_14605_),
    .A2(_14606_),
    .Y(_14607_),
    .B1(_14334_));
 sg13g2_nor3_1 _21932_ (.A(_14601_),
    .B(_14604_),
    .C(_14607_),
    .Y(_14608_));
 sg13g2_nor2_1 _21933_ (.A(_14327_),
    .B(_14608_),
    .Y(_14609_));
 sg13g2_nor2b_1 _21934_ (.A(\u_inv.d_reg[120] ),
    .B_N(\u_inv.d_next[120] ),
    .Y(_14610_));
 sg13g2_a21oi_1 _21935_ (.A1(\u_inv.d_next[121] ),
    .A2(_10921_),
    .Y(_14611_),
    .B1(_14610_));
 sg13g2_a21oi_1 _21936_ (.A1(_10602_),
    .A2(\u_inv.d_reg[121] ),
    .Y(_14612_),
    .B1(_14611_));
 sg13g2_nand2b_1 _21937_ (.Y(_14613_),
    .B(\u_inv.d_next[123] ),
    .A_N(\u_inv.d_reg[123] ));
 sg13g2_nand2b_1 _21938_ (.Y(_14614_),
    .B(\u_inv.d_next[122] ),
    .A_N(\u_inv.d_reg[122] ));
 sg13g2_o21ai_1 _21939_ (.B1(_14613_),
    .Y(_14615_),
    .A1(_14320_),
    .A2(_14614_));
 sg13g2_a21o_1 _21940_ (.A2(_14612_),
    .A1(_14322_),
    .B1(_14615_),
    .X(_14616_));
 sg13g2_nor2b_1 _21941_ (.A(\u_inv.d_reg[125] ),
    .B_N(\u_inv.d_next[125] ),
    .Y(_14617_));
 sg13g2_nor2b_1 _21942_ (.A(\u_inv.d_reg[124] ),
    .B_N(\u_inv.d_next[124] ),
    .Y(_14618_));
 sg13g2_nand2b_1 _21943_ (.Y(_14619_),
    .B(\u_inv.d_next[124] ),
    .A_N(\u_inv.d_reg[124] ));
 sg13g2_a21oi_1 _21944_ (.A1(_14309_),
    .A2(_14618_),
    .Y(_14620_),
    .B1(_14617_));
 sg13g2_nor2b_1 _21945_ (.A(\u_inv.d_reg[126] ),
    .B_N(\u_inv.d_next[126] ),
    .Y(_14621_));
 sg13g2_nor2_1 _21946_ (.A(_10601_),
    .B(\u_inv.d_reg[127] ),
    .Y(_14622_));
 sg13g2_a21oi_1 _21947_ (.A1(_14304_),
    .A2(_14621_),
    .Y(_14623_),
    .B1(_14622_));
 sg13g2_o21ai_1 _21948_ (.B1(_14623_),
    .Y(_14624_),
    .A1(_14307_),
    .A2(_14620_));
 sg13g2_a21oi_1 _21949_ (.A1(_14315_),
    .A2(_14616_),
    .Y(_14625_),
    .B1(_14624_));
 sg13g2_nor2b_1 _21950_ (.A(_14609_),
    .B_N(_14625_),
    .Y(_14626_));
 sg13g2_nor2b_1 _21951_ (.A(\u_inv.d_reg[96] ),
    .B_N(\u_inv.d_next[96] ),
    .Y(_14627_));
 sg13g2_a21oi_1 _21952_ (.A1(_14402_),
    .A2(_14627_),
    .Y(_14628_),
    .B1(_14401_));
 sg13g2_nor2b_1 _21953_ (.A(\u_inv.d_reg[98] ),
    .B_N(\u_inv.d_next[98] ),
    .Y(_14629_));
 sg13g2_o21ai_1 _21954_ (.B1(_14394_),
    .Y(_14630_),
    .A1(_14395_),
    .A2(_14629_));
 sg13g2_o21ai_1 _21955_ (.B1(_14630_),
    .Y(_14631_),
    .A1(_14400_),
    .A2(_14628_));
 sg13g2_nand2b_1 _21956_ (.Y(_14632_),
    .B(_14631_),
    .A_N(_14393_));
 sg13g2_nand2b_1 _21957_ (.Y(_14633_),
    .B(\u_inv.d_next[102] ),
    .A_N(\u_inv.d_reg[102] ));
 sg13g2_a21oi_1 _21958_ (.A1(_10607_),
    .A2(\u_inv.d_reg[103] ),
    .Y(_14634_),
    .B1(_14633_));
 sg13g2_nor2b_1 _21959_ (.A(\u_inv.d_reg[100] ),
    .B_N(\u_inv.d_next[100] ),
    .Y(_14635_));
 sg13g2_nand2_1 _21960_ (.Y(_14636_),
    .A(_14389_),
    .B(_14635_));
 sg13g2_o21ai_1 _21961_ (.B1(_14636_),
    .Y(_14637_),
    .A1(_10608_),
    .A2(\u_inv.d_reg[101] ));
 sg13g2_a221oi_1 _21962_ (.B2(_14637_),
    .C1(_14634_),
    .B1(_14387_),
    .A1(\u_inv.d_next[103] ),
    .Y(_14638_),
    .A2(_10925_));
 sg13g2_nand2_1 _21963_ (.Y(_14639_),
    .A(_14632_),
    .B(_14638_));
 sg13g2_nand2_1 _21964_ (.Y(_14640_),
    .A(_14381_),
    .B(_14639_));
 sg13g2_nand2b_1 _21965_ (.Y(_14641_),
    .B(\u_inv.d_next[104] ),
    .A_N(net4780));
 sg13g2_o21ai_1 _21966_ (.B1(_14641_),
    .Y(_14642_),
    .A1(_10606_),
    .A2(\u_inv.d_reg[105] ));
 sg13g2_o21ai_1 _21967_ (.B1(_14642_),
    .Y(_14643_),
    .A1(\u_inv.d_next[105] ),
    .A2(_10924_));
 sg13g2_nor2b_1 _21968_ (.A(\u_inv.d_reg[106] ),
    .B_N(\u_inv.d_next[106] ),
    .Y(_14644_));
 sg13g2_o21ai_1 _21969_ (.B1(_14370_),
    .Y(_14645_),
    .A1(_14375_),
    .A2(_14643_));
 sg13g2_a21oi_1 _21970_ (.A1(_14369_),
    .A2(_14644_),
    .Y(_14646_),
    .B1(_14645_));
 sg13g2_or2_1 _21971_ (.X(_14647_),
    .B(_14646_),
    .A(_14368_));
 sg13g2_nor2b_1 _21972_ (.A(\u_inv.d_reg[108] ),
    .B_N(\u_inv.d_next[108] ),
    .Y(_14648_));
 sg13g2_a21oi_1 _21973_ (.A1(\u_inv.d_next[109] ),
    .A2(_10923_),
    .Y(_14649_),
    .B1(_14648_));
 sg13g2_a21oi_1 _21974_ (.A1(_10605_),
    .A2(\u_inv.d_reg[109] ),
    .Y(_14650_),
    .B1(_14649_));
 sg13g2_nand2b_1 _21975_ (.Y(_14651_),
    .B(\u_inv.d_next[110] ),
    .A_N(\u_inv.d_reg[110] ));
 sg13g2_or2_1 _21976_ (.X(_14652_),
    .B(_14651_),
    .A(_14359_));
 sg13g2_a22oi_1 _21977_ (.Y(_14653_),
    .B1(_14363_),
    .B2(_14650_),
    .A2(_10922_),
    .A1(\u_inv.d_next[111] ));
 sg13g2_nand4_1 _21978_ (.B(_14647_),
    .C(_14652_),
    .A(_14640_),
    .Y(_14654_),
    .D(_14653_));
 sg13g2_nand2_1 _21979_ (.Y(_14655_),
    .A(_14358_),
    .B(_14654_));
 sg13g2_and3_2 _21980_ (.X(_14656_),
    .A(_14595_),
    .B(_14626_),
    .C(_14655_));
 sg13g2_nand3_1 _21981_ (.B(_14626_),
    .C(_14655_),
    .A(_14595_),
    .Y(_14657_));
 sg13g2_nand2_1 _21982_ (.Y(_14658_),
    .A(_14537_),
    .B(_14656_));
 sg13g2_nor2_1 _21983_ (.A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ),
    .Y(_14659_));
 sg13g2_nand2_1 _21984_ (.Y(_14660_),
    .A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ));
 sg13g2_xor2_1 _21985_ (.B(\u_inv.d_reg[191] ),
    .A(\u_inv.d_next[191] ),
    .X(_14661_));
 sg13g2_nand2_1 _21986_ (.Y(_14662_),
    .A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ));
 sg13g2_nor2_1 _21987_ (.A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ),
    .Y(_14663_));
 sg13g2_xor2_1 _21988_ (.B(\u_inv.d_reg[190] ),
    .A(\u_inv.d_next[190] ),
    .X(_14664_));
 sg13g2_nor2_1 _21989_ (.A(_14661_),
    .B(_14664_),
    .Y(_14665_));
 sg13g2_xor2_1 _21990_ (.B(\u_inv.d_reg[189] ),
    .A(\u_inv.d_next[189] ),
    .X(_14666_));
 sg13g2_and2_1 _21991_ (.A(\u_inv.d_next[188] ),
    .B(\u_inv.d_reg[188] ),
    .X(_14667_));
 sg13g2_xor2_1 _21992_ (.B(\u_inv.d_reg[188] ),
    .A(\u_inv.d_next[188] ),
    .X(_14668_));
 sg13g2_nor2_1 _21993_ (.A(_14666_),
    .B(_14668_),
    .Y(_14669_));
 sg13g2_inv_1 _21994_ (.Y(_14670_),
    .A(_14669_));
 sg13g2_nand2_1 _21995_ (.Y(_14671_),
    .A(_14665_),
    .B(_14669_));
 sg13g2_nand2_1 _21996_ (.Y(_14672_),
    .A(_10591_),
    .B(\u_inv.d_reg[185] ));
 sg13g2_xnor2_1 _21997_ (.Y(_14673_),
    .A(\u_inv.d_next[185] ),
    .B(\u_inv.d_reg[185] ));
 sg13g2_nand2_1 _21998_ (.Y(_14674_),
    .A(\u_inv.d_next[184] ),
    .B(\u_inv.d_reg[184] ));
 sg13g2_xor2_1 _21999_ (.B(\u_inv.d_reg[184] ),
    .A(\u_inv.d_next[184] ),
    .X(_14675_));
 sg13g2_nor2b_1 _22000_ (.A(_14675_),
    .B_N(_14673_),
    .Y(_14676_));
 sg13g2_nand2_1 _22001_ (.Y(_14677_),
    .A(\u_inv.d_next[186] ),
    .B(\u_inv.d_reg[186] ));
 sg13g2_xor2_1 _22002_ (.B(\u_inv.d_reg[186] ),
    .A(\u_inv.d_next[186] ),
    .X(_14678_));
 sg13g2_xnor2_1 _22003_ (.Y(_14679_),
    .A(\u_inv.d_next[186] ),
    .B(\u_inv.d_reg[186] ));
 sg13g2_nor2_1 _22004_ (.A(\u_inv.d_next[187] ),
    .B(net4774),
    .Y(_14680_));
 sg13g2_xor2_1 _22005_ (.B(net4774),
    .A(\u_inv.d_next[187] ),
    .X(_14681_));
 sg13g2_xnor2_1 _22006_ (.Y(_14682_),
    .A(\u_inv.d_next[187] ),
    .B(net4774));
 sg13g2_nor2_1 _22007_ (.A(_14678_),
    .B(_14681_),
    .Y(_14683_));
 sg13g2_nand2_1 _22008_ (.Y(_14684_),
    .A(_14676_),
    .B(_14683_));
 sg13g2_inv_1 _22009_ (.Y(_14685_),
    .A(_14684_));
 sg13g2_nor2_1 _22010_ (.A(_14671_),
    .B(_14684_),
    .Y(_14686_));
 sg13g2_xnor2_1 _22011_ (.Y(_14687_),
    .A(\u_inv.d_next[181] ),
    .B(\u_inv.d_reg[181] ));
 sg13g2_nand2_1 _22012_ (.Y(_14688_),
    .A(\u_inv.d_next[180] ),
    .B(\u_inv.d_reg[180] ));
 sg13g2_xor2_1 _22013_ (.B(\u_inv.d_reg[180] ),
    .A(\u_inv.d_next[180] ),
    .X(_14689_));
 sg13g2_xnor2_1 _22014_ (.Y(_14690_),
    .A(\u_inv.d_next[180] ),
    .B(\u_inv.d_reg[180] ));
 sg13g2_nand2_1 _22015_ (.Y(_14691_),
    .A(_14687_),
    .B(_14690_));
 sg13g2_nor2_1 _22016_ (.A(\u_inv.d_next[183] ),
    .B(\u_inv.d_reg[183] ),
    .Y(_14692_));
 sg13g2_xnor2_1 _22017_ (.Y(_14693_),
    .A(\u_inv.d_next[183] ),
    .B(\u_inv.d_reg[183] ));
 sg13g2_nand2_1 _22018_ (.Y(_14694_),
    .A(\u_inv.d_next[182] ),
    .B(\u_inv.d_reg[182] ));
 sg13g2_xnor2_1 _22019_ (.Y(_14695_),
    .A(\u_inv.d_next[182] ),
    .B(\u_inv.d_reg[182] ));
 sg13g2_and4_1 _22020_ (.A(_14687_),
    .B(_14690_),
    .C(_14693_),
    .D(_14695_),
    .X(_14696_));
 sg13g2_nor2_1 _22021_ (.A(\u_inv.d_next[179] ),
    .B(_10905_),
    .Y(_14697_));
 sg13g2_xnor2_1 _22022_ (.Y(_14698_),
    .A(\u_inv.d_next[179] ),
    .B(\u_inv.d_reg[179] ));
 sg13g2_xor2_1 _22023_ (.B(\u_inv.d_reg[179] ),
    .A(\u_inv.d_next[179] ),
    .X(_14699_));
 sg13g2_nand2_1 _22024_ (.Y(_14700_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_xor2_1 _22025_ (.B(\u_inv.d_reg[178] ),
    .A(\u_inv.d_next[178] ),
    .X(_14701_));
 sg13g2_xnor2_1 _22026_ (.Y(_14702_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_nor2_1 _22027_ (.A(_14699_),
    .B(_14701_),
    .Y(_14703_));
 sg13g2_nor2b_1 _22028_ (.A(\u_inv.d_reg[177] ),
    .B_N(\u_inv.d_next[177] ),
    .Y(_14704_));
 sg13g2_nand2b_1 _22029_ (.Y(_14705_),
    .B(\u_inv.d_reg[177] ),
    .A_N(\u_inv.d_next[177] ));
 sg13g2_xnor2_1 _22030_ (.Y(_14706_),
    .A(\u_inv.d_next[177] ),
    .B(\u_inv.d_reg[177] ));
 sg13g2_nand2_1 _22031_ (.Y(_14707_),
    .A(\u_inv.d_next[176] ),
    .B(\u_inv.d_reg[176] ));
 sg13g2_xnor2_1 _22032_ (.Y(_14708_),
    .A(\u_inv.d_next[176] ),
    .B(\u_inv.d_reg[176] ));
 sg13g2_nand2_1 _22033_ (.Y(_14709_),
    .A(_14706_),
    .B(_14708_));
 sg13g2_and4_1 _22034_ (.A(_14696_),
    .B(_14703_),
    .C(_14706_),
    .D(_14708_),
    .X(_14710_));
 sg13g2_inv_1 _22035_ (.Y(_14711_),
    .A(_14710_));
 sg13g2_nand2_2 _22036_ (.Y(_14712_),
    .A(_14686_),
    .B(_14710_));
 sg13g2_nor2_1 _22037_ (.A(\u_inv.d_next[175] ),
    .B(\u_inv.d_reg[175] ),
    .Y(_14713_));
 sg13g2_xnor2_1 _22038_ (.Y(_14714_),
    .A(\u_inv.d_next[175] ),
    .B(\u_inv.d_reg[175] ));
 sg13g2_nand2_1 _22039_ (.Y(_14715_),
    .A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ));
 sg13g2_xnor2_1 _22040_ (.Y(_14716_),
    .A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ));
 sg13g2_and2_1 _22041_ (.A(_14714_),
    .B(_14716_),
    .X(_14717_));
 sg13g2_nand2_1 _22042_ (.Y(_14718_),
    .A(_10593_),
    .B(\u_inv.d_reg[173] ));
 sg13g2_xnor2_1 _22043_ (.Y(_14719_),
    .A(\u_inv.d_next[173] ),
    .B(\u_inv.d_reg[173] ));
 sg13g2_nand2_1 _22044_ (.Y(_14720_),
    .A(\u_inv.d_next[172] ),
    .B(\u_inv.d_reg[172] ));
 sg13g2_xor2_1 _22045_ (.B(\u_inv.d_reg[172] ),
    .A(\u_inv.d_next[172] ),
    .X(_14721_));
 sg13g2_xnor2_1 _22046_ (.Y(_14722_),
    .A(\u_inv.d_next[172] ),
    .B(\u_inv.d_reg[172] ));
 sg13g2_nand2_1 _22047_ (.Y(_14723_),
    .A(_14719_),
    .B(_14722_));
 sg13g2_nand3_1 _22048_ (.B(_14719_),
    .C(_14722_),
    .A(_14717_),
    .Y(_14724_));
 sg13g2_xnor2_1 _22049_ (.Y(_14725_),
    .A(\u_inv.d_next[171] ),
    .B(\u_inv.d_reg[171] ));
 sg13g2_xor2_1 _22050_ (.B(\u_inv.d_reg[171] ),
    .A(\u_inv.d_next[171] ),
    .X(_14726_));
 sg13g2_nand2_1 _22051_ (.Y(_14727_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_xnor2_1 _22052_ (.Y(_14728_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_and2_1 _22053_ (.A(_14725_),
    .B(_14728_),
    .X(_14729_));
 sg13g2_nand2_1 _22054_ (.Y(_14730_),
    .A(_14725_),
    .B(_14728_));
 sg13g2_xnor2_1 _22055_ (.Y(_14731_),
    .A(\u_inv.d_next[169] ),
    .B(\u_inv.d_reg[169] ));
 sg13g2_nand2_1 _22056_ (.Y(_14732_),
    .A(\u_inv.d_next[168] ),
    .B(\u_inv.d_reg[168] ));
 sg13g2_xnor2_1 _22057_ (.Y(_14733_),
    .A(\u_inv.d_next[168] ),
    .B(\u_inv.d_reg[168] ));
 sg13g2_nand2_1 _22058_ (.Y(_14734_),
    .A(_14731_),
    .B(_14733_));
 sg13g2_nand2b_1 _22059_ (.Y(_14735_),
    .B(\u_inv.d_next[167] ),
    .A_N(\u_inv.d_reg[167] ));
 sg13g2_nor2b_1 _22060_ (.A(\u_inv.d_next[167] ),
    .B_N(\u_inv.d_reg[167] ),
    .Y(_14736_));
 sg13g2_xor2_1 _22061_ (.B(\u_inv.d_reg[167] ),
    .A(\u_inv.d_next[167] ),
    .X(_14737_));
 sg13g2_nand2_1 _22062_ (.Y(_14738_),
    .A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ));
 sg13g2_nor2_1 _22063_ (.A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ),
    .Y(_14739_));
 sg13g2_xor2_1 _22064_ (.B(\u_inv.d_reg[166] ),
    .A(\u_inv.d_next[166] ),
    .X(_14740_));
 sg13g2_nor2_1 _22065_ (.A(_14737_),
    .B(_14740_),
    .Y(_14741_));
 sg13g2_nand2_1 _22066_ (.Y(_14742_),
    .A(\u_inv.d_next[165] ),
    .B(\u_inv.d_reg[165] ));
 sg13g2_xnor2_1 _22067_ (.Y(_14743_),
    .A(\u_inv.d_next[165] ),
    .B(\u_inv.d_reg[165] ));
 sg13g2_and2_1 _22068_ (.A(\u_inv.d_next[164] ),
    .B(\u_inv.d_reg[164] ),
    .X(_14744_));
 sg13g2_or2_1 _22069_ (.X(_14745_),
    .B(\u_inv.d_reg[164] ),
    .A(\u_inv.d_next[164] ));
 sg13g2_xnor2_1 _22070_ (.Y(_14746_),
    .A(\u_inv.d_next[164] ),
    .B(\u_inv.d_reg[164] ));
 sg13g2_and2_1 _22071_ (.A(_14743_),
    .B(_14746_),
    .X(_14747_));
 sg13g2_and2_1 _22072_ (.A(_14741_),
    .B(_14747_),
    .X(_14748_));
 sg13g2_nand2b_1 _22073_ (.Y(_14749_),
    .B(\u_inv.d_reg[163] ),
    .A_N(\u_inv.d_next[163] ));
 sg13g2_nor2b_1 _22074_ (.A(\u_inv.d_reg[163] ),
    .B_N(\u_inv.d_next[163] ),
    .Y(_14750_));
 sg13g2_xnor2_1 _22075_ (.Y(_14751_),
    .A(\u_inv.d_next[163] ),
    .B(\u_inv.d_reg[163] ));
 sg13g2_xor2_1 _22076_ (.B(\u_inv.d_reg[163] ),
    .A(\u_inv.d_next[163] ),
    .X(_14752_));
 sg13g2_nand2_1 _22077_ (.Y(_14753_),
    .A(net4801),
    .B(net4775));
 sg13g2_nor2_1 _22078_ (.A(net4801),
    .B(net4775),
    .Y(_14754_));
 sg13g2_xor2_1 _22079_ (.B(net4775),
    .A(net4801),
    .X(_14755_));
 sg13g2_xnor2_1 _22080_ (.Y(_14756_),
    .A(net4801),
    .B(net4775));
 sg13g2_nand2_1 _22081_ (.Y(_14757_),
    .A(_14751_),
    .B(_14756_));
 sg13g2_nor2b_1 _22082_ (.A(\u_inv.d_reg[161] ),
    .B_N(\u_inv.d_next[161] ),
    .Y(_14758_));
 sg13g2_nand2b_1 _22083_ (.Y(_14759_),
    .B(\u_inv.d_reg[161] ),
    .A_N(\u_inv.d_next[161] ));
 sg13g2_nor2b_2 _22084_ (.A(_14758_),
    .B_N(_14759_),
    .Y(_14760_));
 sg13g2_nand2_1 _22085_ (.Y(_14761_),
    .A(\u_inv.d_next[160] ),
    .B(\u_inv.d_reg[160] ));
 sg13g2_xor2_1 _22086_ (.B(\u_inv.d_reg[160] ),
    .A(\u_inv.d_next[160] ),
    .X(_14762_));
 sg13g2_xnor2_1 _22087_ (.Y(_14763_),
    .A(\u_inv.d_next[160] ),
    .B(\u_inv.d_reg[160] ));
 sg13g2_and2_1 _22088_ (.A(_14760_),
    .B(_14763_),
    .X(_14764_));
 sg13g2_nand4_1 _22089_ (.B(_14751_),
    .C(_14756_),
    .A(_14748_),
    .Y(_14765_),
    .D(_14764_));
 sg13g2_inv_1 _22090_ (.Y(_14766_),
    .A(_14765_));
 sg13g2_or4_1 _22091_ (.A(_14724_),
    .B(_14730_),
    .C(_14734_),
    .D(_14765_),
    .X(_14767_));
 sg13g2_inv_1 _22092_ (.Y(_14768_),
    .A(_14767_));
 sg13g2_nor2_2 _22093_ (.A(_14712_),
    .B(_14767_),
    .Y(_14769_));
 sg13g2_xnor2_1 _22094_ (.Y(_14770_),
    .A(\u_inv.d_next[159] ),
    .B(\u_inv.d_reg[159] ));
 sg13g2_nand2_1 _22095_ (.Y(_14771_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_xor2_1 _22096_ (.B(\u_inv.d_reg[158] ),
    .A(\u_inv.d_next[158] ),
    .X(_14772_));
 sg13g2_xnor2_1 _22097_ (.Y(_14773_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_nand2_1 _22098_ (.Y(_14774_),
    .A(_14770_),
    .B(_14773_));
 sg13g2_xnor2_1 _22099_ (.Y(_14775_),
    .A(\u_inv.d_next[157] ),
    .B(\u_inv.d_reg[157] ));
 sg13g2_xor2_1 _22100_ (.B(\u_inv.d_reg[157] ),
    .A(\u_inv.d_next[157] ),
    .X(_14776_));
 sg13g2_and2_1 _22101_ (.A(\u_inv.d_next[156] ),
    .B(\u_inv.d_reg[156] ),
    .X(_14777_));
 sg13g2_nand2_1 _22102_ (.Y(_14778_),
    .A(\u_inv.d_next[156] ),
    .B(\u_inv.d_reg[156] ));
 sg13g2_xor2_1 _22103_ (.B(\u_inv.d_reg[156] ),
    .A(\u_inv.d_next[156] ),
    .X(_14779_));
 sg13g2_xnor2_1 _22104_ (.Y(_14780_),
    .A(\u_inv.d_next[156] ),
    .B(\u_inv.d_reg[156] ));
 sg13g2_nand2_1 _22105_ (.Y(_14781_),
    .A(_14775_),
    .B(_14780_));
 sg13g2_nor2_1 _22106_ (.A(_14774_),
    .B(_14781_),
    .Y(_14782_));
 sg13g2_nor2_1 _22107_ (.A(\u_inv.d_next[155] ),
    .B(_10915_),
    .Y(_14783_));
 sg13g2_xnor2_1 _22108_ (.Y(_14784_),
    .A(\u_inv.d_next[155] ),
    .B(\u_inv.d_reg[155] ));
 sg13g2_nand2_1 _22109_ (.Y(_14785_),
    .A(\u_inv.d_next[154] ),
    .B(\u_inv.d_reg[154] ));
 sg13g2_xnor2_1 _22110_ (.Y(_14786_),
    .A(\u_inv.d_next[154] ),
    .B(\u_inv.d_reg[154] ));
 sg13g2_and2_1 _22111_ (.A(_14784_),
    .B(_14786_),
    .X(_14787_));
 sg13g2_nor2b_1 _22112_ (.A(\u_inv.d_reg[153] ),
    .B_N(\u_inv.d_next[153] ),
    .Y(_14788_));
 sg13g2_nand2b_1 _22113_ (.Y(_14789_),
    .B(\u_inv.d_reg[153] ),
    .A_N(\u_inv.d_next[153] ));
 sg13g2_xor2_1 _22114_ (.B(\u_inv.d_reg[153] ),
    .A(\u_inv.d_next[153] ),
    .X(_14790_));
 sg13g2_and2_1 _22115_ (.A(\u_inv.d_next[152] ),
    .B(\u_inv.d_reg[152] ),
    .X(_14791_));
 sg13g2_xor2_1 _22116_ (.B(\u_inv.d_reg[152] ),
    .A(\u_inv.d_next[152] ),
    .X(_14792_));
 sg13g2_nor2_1 _22117_ (.A(_14790_),
    .B(_14792_),
    .Y(_14793_));
 sg13g2_inv_1 _22118_ (.Y(_14794_),
    .A(_14793_));
 sg13g2_nand3_1 _22119_ (.B(_14787_),
    .C(_14793_),
    .A(_14782_),
    .Y(_14795_));
 sg13g2_inv_1 _22120_ (.Y(_14796_),
    .A(_14795_));
 sg13g2_xor2_1 _22121_ (.B(\u_inv.d_reg[151] ),
    .A(\u_inv.d_next[151] ),
    .X(_14797_));
 sg13g2_nand2_1 _22122_ (.Y(_14798_),
    .A(\u_inv.d_next[150] ),
    .B(net4776));
 sg13g2_nor2_1 _22123_ (.A(\u_inv.d_next[150] ),
    .B(net4776),
    .Y(_14799_));
 sg13g2_or2_1 _22124_ (.X(_14800_),
    .B(net4776),
    .A(\u_inv.d_next[150] ));
 sg13g2_xor2_1 _22125_ (.B(net4776),
    .A(\u_inv.d_next[150] ),
    .X(_14801_));
 sg13g2_nor2_1 _22126_ (.A(_14797_),
    .B(_14801_),
    .Y(_14802_));
 sg13g2_nor2_1 _22127_ (.A(\u_inv.d_next[149] ),
    .B(\u_inv.d_reg[149] ),
    .Y(_14803_));
 sg13g2_xnor2_1 _22128_ (.Y(_14804_),
    .A(\u_inv.d_next[149] ),
    .B(\u_inv.d_reg[149] ));
 sg13g2_and2_1 _22129_ (.A(\u_inv.d_next[148] ),
    .B(\u_inv.d_reg[148] ),
    .X(_14805_));
 sg13g2_or2_1 _22130_ (.X(_14806_),
    .B(\u_inv.d_reg[148] ),
    .A(\u_inv.d_next[148] ));
 sg13g2_xnor2_1 _22131_ (.Y(_14807_),
    .A(\u_inv.d_next[148] ),
    .B(\u_inv.d_reg[148] ));
 sg13g2_and2_1 _22132_ (.A(_14804_),
    .B(_14807_),
    .X(_14808_));
 sg13g2_and2_1 _22133_ (.A(_14802_),
    .B(_14808_),
    .X(_14809_));
 sg13g2_nand2b_1 _22134_ (.Y(_14810_),
    .B(\u_inv.d_reg[147] ),
    .A_N(\u_inv.d_next[147] ));
 sg13g2_nor2b_1 _22135_ (.A(\u_inv.d_reg[147] ),
    .B_N(\u_inv.d_next[147] ),
    .Y(_14811_));
 sg13g2_xnor2_1 _22136_ (.Y(_14812_),
    .A(\u_inv.d_next[147] ),
    .B(\u_inv.d_reg[147] ));
 sg13g2_xor2_1 _22137_ (.B(\u_inv.d_reg[147] ),
    .A(\u_inv.d_next[147] ),
    .X(_14813_));
 sg13g2_and2_1 _22138_ (.A(\u_inv.d_next[146] ),
    .B(\u_inv.d_reg[146] ),
    .X(_14814_));
 sg13g2_nand2_1 _22139_ (.Y(_14815_),
    .A(\u_inv.d_next[146] ),
    .B(\u_inv.d_reg[146] ));
 sg13g2_xnor2_1 _22140_ (.Y(_14816_),
    .A(\u_inv.d_next[146] ),
    .B(\u_inv.d_reg[146] ));
 sg13g2_inv_1 _22141_ (.Y(_14817_),
    .A(_14816_));
 sg13g2_nand2_1 _22142_ (.Y(_14818_),
    .A(_14812_),
    .B(_14816_));
 sg13g2_nor2b_1 _22143_ (.A(\u_inv.d_reg[145] ),
    .B_N(\u_inv.d_next[145] ),
    .Y(_14819_));
 sg13g2_nand2b_1 _22144_ (.Y(_14820_),
    .B(\u_inv.d_reg[145] ),
    .A_N(\u_inv.d_next[145] ));
 sg13g2_xnor2_1 _22145_ (.Y(_14821_),
    .A(\u_inv.d_next[145] ),
    .B(\u_inv.d_reg[145] ));
 sg13g2_nand2_1 _22146_ (.Y(_14822_),
    .A(\u_inv.d_next[144] ),
    .B(\u_inv.d_reg[144] ));
 sg13g2_xnor2_1 _22147_ (.Y(_14823_),
    .A(\u_inv.d_next[144] ),
    .B(\u_inv.d_reg[144] ));
 sg13g2_inv_1 _22148_ (.Y(_14824_),
    .A(_14823_));
 sg13g2_and2_1 _22149_ (.A(_14821_),
    .B(_14823_),
    .X(_14825_));
 sg13g2_nand4_1 _22150_ (.B(_14812_),
    .C(_14816_),
    .A(_14809_),
    .Y(_14826_),
    .D(_14825_));
 sg13g2_inv_1 _22151_ (.Y(_14827_),
    .A(_14826_));
 sg13g2_nor2_2 _22152_ (.A(_14795_),
    .B(_14826_),
    .Y(_14828_));
 sg13g2_nor2b_1 _22153_ (.A(\u_inv.d_reg[143] ),
    .B_N(\u_inv.d_next[143] ),
    .Y(_14829_));
 sg13g2_nand2b_1 _22154_ (.Y(_14830_),
    .B(\u_inv.d_reg[143] ),
    .A_N(\u_inv.d_next[143] ));
 sg13g2_xnor2_1 _22155_ (.Y(_14831_),
    .A(\u_inv.d_next[143] ),
    .B(\u_inv.d_reg[143] ));
 sg13g2_nand2b_2 _22156_ (.Y(_14832_),
    .B(_14830_),
    .A_N(_14829_));
 sg13g2_nand2_1 _22157_ (.Y(_14833_),
    .A(\u_inv.d_next[142] ),
    .B(\u_inv.d_reg[142] ));
 sg13g2_xnor2_1 _22158_ (.Y(_14834_),
    .A(\u_inv.d_next[142] ),
    .B(\u_inv.d_reg[142] ));
 sg13g2_inv_1 _22159_ (.Y(_14835_),
    .A(_14834_));
 sg13g2_nand2_1 _22160_ (.Y(_14836_),
    .A(_14831_),
    .B(_14834_));
 sg13g2_nor2_1 _22161_ (.A(\u_inv.d_next[141] ),
    .B(\u_inv.d_reg[141] ),
    .Y(_14837_));
 sg13g2_xnor2_1 _22162_ (.Y(_14838_),
    .A(\u_inv.d_next[141] ),
    .B(\u_inv.d_reg[141] ));
 sg13g2_nand2_1 _22163_ (.Y(_14839_),
    .A(\u_inv.d_next[140] ),
    .B(\u_inv.d_reg[140] ));
 sg13g2_xnor2_1 _22164_ (.Y(_14840_),
    .A(\u_inv.d_next[140] ),
    .B(\u_inv.d_reg[140] ));
 sg13g2_and2_1 _22165_ (.A(net4430),
    .B(net4429),
    .X(_14841_));
 sg13g2_nand4_1 _22166_ (.B(_14834_),
    .C(net4430),
    .A(_14831_),
    .Y(_14842_),
    .D(net4429));
 sg13g2_inv_1 _22167_ (.Y(_14843_),
    .A(_14842_));
 sg13g2_nand2b_1 _22168_ (.Y(_14844_),
    .B(\u_inv.d_reg[139] ),
    .A_N(\u_inv.d_next[139] ));
 sg13g2_nor2b_1 _22169_ (.A(\u_inv.d_reg[139] ),
    .B_N(\u_inv.d_next[139] ),
    .Y(_14845_));
 sg13g2_xnor2_1 _22170_ (.Y(_14846_),
    .A(\u_inv.d_next[139] ),
    .B(\u_inv.d_reg[139] ));
 sg13g2_xor2_1 _22171_ (.B(\u_inv.d_reg[139] ),
    .A(\u_inv.d_next[139] ),
    .X(_14847_));
 sg13g2_nand2_1 _22172_ (.Y(_14848_),
    .A(\u_inv.d_next[138] ),
    .B(net4777));
 sg13g2_xnor2_1 _22173_ (.Y(_14849_),
    .A(\u_inv.d_next[138] ),
    .B(net4777));
 sg13g2_inv_1 _22174_ (.Y(_14850_),
    .A(_14849_));
 sg13g2_nor2_1 _22175_ (.A(_14847_),
    .B(_14850_),
    .Y(_14851_));
 sg13g2_nand2_1 _22176_ (.Y(_14852_),
    .A(_14846_),
    .B(_14849_));
 sg13g2_or2_1 _22177_ (.X(_14853_),
    .B(\u_inv.d_reg[137] ),
    .A(\u_inv.d_next[137] ));
 sg13g2_and2_1 _22178_ (.A(\u_inv.d_next[137] ),
    .B(\u_inv.d_reg[137] ),
    .X(_14854_));
 sg13g2_xor2_1 _22179_ (.B(\u_inv.d_reg[137] ),
    .A(\u_inv.d_next[137] ),
    .X(_14855_));
 sg13g2_xnor2_1 _22180_ (.Y(_14856_),
    .A(\u_inv.d_next[137] ),
    .B(\u_inv.d_reg[137] ));
 sg13g2_and2_1 _22181_ (.A(\u_inv.d_next[136] ),
    .B(\u_inv.d_reg[136] ),
    .X(_14857_));
 sg13g2_xor2_1 _22182_ (.B(\u_inv.d_reg[136] ),
    .A(\u_inv.d_next[136] ),
    .X(_14858_));
 sg13g2_xnor2_1 _22183_ (.Y(_14859_),
    .A(\u_inv.d_next[136] ),
    .B(\u_inv.d_reg[136] ));
 sg13g2_nand2_1 _22184_ (.Y(_14860_),
    .A(_14856_),
    .B(_14859_));
 sg13g2_nand4_1 _22185_ (.B(_14851_),
    .C(_14856_),
    .A(_14843_),
    .Y(_14861_),
    .D(_14859_));
 sg13g2_nand2_1 _22186_ (.Y(_14862_),
    .A(\u_inv.d_next[135] ),
    .B(_10918_));
 sg13g2_nor2_1 _22187_ (.A(\u_inv.d_next[135] ),
    .B(_10918_),
    .Y(_14863_));
 sg13g2_xnor2_1 _22188_ (.Y(_14864_),
    .A(\u_inv.d_next[135] ),
    .B(\u_inv.d_reg[135] ));
 sg13g2_xor2_1 _22189_ (.B(\u_inv.d_reg[135] ),
    .A(\u_inv.d_next[135] ),
    .X(_14865_));
 sg13g2_and2_1 _22190_ (.A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ),
    .X(_14866_));
 sg13g2_xor2_1 _22191_ (.B(\u_inv.d_reg[134] ),
    .A(\u_inv.d_next[134] ),
    .X(_14867_));
 sg13g2_xnor2_1 _22192_ (.Y(_14868_),
    .A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ));
 sg13g2_nor2_1 _22193_ (.A(_14865_),
    .B(_14867_),
    .Y(_14869_));
 sg13g2_nor2_1 _22194_ (.A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ),
    .Y(_14870_));
 sg13g2_nand2_1 _22195_ (.Y(_14871_),
    .A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ));
 sg13g2_nor2b_1 _22196_ (.A(_14870_),
    .B_N(_14871_),
    .Y(_14872_));
 sg13g2_xnor2_1 _22197_ (.Y(_14873_),
    .A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ));
 sg13g2_nand2_1 _22198_ (.Y(_14874_),
    .A(\u_inv.d_next[132] ),
    .B(\u_inv.d_reg[132] ));
 sg13g2_xnor2_1 _22199_ (.Y(_14875_),
    .A(\u_inv.d_next[132] ),
    .B(\u_inv.d_reg[132] ));
 sg13g2_and2_1 _22200_ (.A(_14873_),
    .B(_14875_),
    .X(_14876_));
 sg13g2_inv_1 _22201_ (.Y(_14877_),
    .A(_14876_));
 sg13g2_and2_1 _22202_ (.A(_14869_),
    .B(_14876_),
    .X(_14878_));
 sg13g2_nor2b_1 _22203_ (.A(\u_inv.d_next[131] ),
    .B_N(\u_inv.d_reg[131] ),
    .Y(_14879_));
 sg13g2_nand2b_1 _22204_ (.Y(_14880_),
    .B(\u_inv.d_next[131] ),
    .A_N(\u_inv.d_reg[131] ));
 sg13g2_xnor2_1 _22205_ (.Y(_14881_),
    .A(\u_inv.d_next[131] ),
    .B(\u_inv.d_reg[131] ));
 sg13g2_xor2_1 _22206_ (.B(\u_inv.d_reg[131] ),
    .A(\u_inv.d_next[131] ),
    .X(_14882_));
 sg13g2_nand2_1 _22207_ (.Y(_14883_),
    .A(net4802),
    .B(net4778));
 sg13g2_xor2_1 _22208_ (.B(net4778),
    .A(net4802),
    .X(_14884_));
 sg13g2_xnor2_1 _22209_ (.Y(_14885_),
    .A(net4802),
    .B(net4778));
 sg13g2_nand2_2 _22210_ (.Y(_14886_),
    .A(_14881_),
    .B(_14885_));
 sg13g2_nor2b_1 _22211_ (.A(net4779),
    .B_N(\u_inv.d_next[129] ),
    .Y(_14887_));
 sg13g2_nand2b_1 _22212_ (.Y(_14888_),
    .B(net4779),
    .A_N(\u_inv.d_next[129] ));
 sg13g2_nor2b_2 _22213_ (.A(_14887_),
    .B_N(_14888_),
    .Y(_14889_));
 sg13g2_xor2_1 _22214_ (.B(net4779),
    .A(\u_inv.d_next[129] ),
    .X(_14890_));
 sg13g2_and2_1 _22215_ (.A(\u_inv.d_next[128] ),
    .B(\u_inv.d_reg[128] ),
    .X(_14891_));
 sg13g2_xnor2_1 _22216_ (.Y(_14892_),
    .A(\u_inv.d_next[128] ),
    .B(\u_inv.d_reg[128] ));
 sg13g2_nor2b_1 _22217_ (.A(_14890_),
    .B_N(_14892_),
    .Y(_14893_));
 sg13g2_nand2_1 _22218_ (.Y(_14894_),
    .A(_14878_),
    .B(_14893_));
 sg13g2_nor2_1 _22219_ (.A(_14886_),
    .B(_14894_),
    .Y(_14895_));
 sg13g2_nor3_1 _22220_ (.A(_14861_),
    .B(_14886_),
    .C(_14894_),
    .Y(_14896_));
 sg13g2_inv_1 _22221_ (.Y(_14897_),
    .A(_14896_));
 sg13g2_and2_1 _22222_ (.A(_14828_),
    .B(_14896_),
    .X(_14898_));
 sg13g2_inv_1 _22223_ (.Y(_14899_),
    .A(_14898_));
 sg13g2_nand2_2 _22224_ (.Y(_14900_),
    .A(_14769_),
    .B(_14898_));
 sg13g2_a21oi_1 _22225_ (.A1(_14537_),
    .A2(_14656_),
    .Y(_14901_),
    .B1(_14900_));
 sg13g2_a21o_1 _22226_ (.A2(_14656_),
    .A1(_14537_),
    .B1(_14900_),
    .X(_14902_));
 sg13g2_nor2b_1 _22227_ (.A(\u_inv.d_reg[128] ),
    .B_N(\u_inv.d_next[128] ),
    .Y(_14903_));
 sg13g2_a21oi_2 _22228_ (.B1(_14887_),
    .Y(_14904_),
    .A2(_14903_),
    .A1(_14888_));
 sg13g2_nand2b_1 _22229_ (.Y(_14905_),
    .B(net4802),
    .A_N(net4778));
 sg13g2_a21o_2 _22230_ (.A2(_14905_),
    .A1(_14880_),
    .B1(_14879_),
    .X(_14906_));
 sg13g2_inv_1 _22231_ (.Y(_14907_),
    .A(_14906_));
 sg13g2_o21ai_1 _22232_ (.B1(_14906_),
    .Y(_14908_),
    .A1(_14886_),
    .A2(_14904_));
 sg13g2_nand2b_1 _22233_ (.Y(_14909_),
    .B(\u_inv.d_next[134] ),
    .A_N(\u_inv.d_reg[134] ));
 sg13g2_o21ai_1 _22234_ (.B1(_14862_),
    .Y(_14910_),
    .A1(_14863_),
    .A2(_14909_));
 sg13g2_nand2b_1 _22235_ (.Y(_14911_),
    .B(\u_inv.d_next[133] ),
    .A_N(\u_inv.d_reg[133] ));
 sg13g2_nand2b_1 _22236_ (.Y(_14912_),
    .B(\u_inv.d_next[132] ),
    .A_N(\u_inv.d_reg[132] ));
 sg13g2_o21ai_1 _22237_ (.B1(_14911_),
    .Y(_14913_),
    .A1(_14872_),
    .A2(_14912_));
 sg13g2_a221oi_1 _22238_ (.B2(_14869_),
    .C1(_14910_),
    .B1(_14913_),
    .A1(_14878_),
    .Y(_14914_),
    .A2(_14908_));
 sg13g2_nor2b_1 _22239_ (.A(\u_inv.d_reg[141] ),
    .B_N(\u_inv.d_next[141] ),
    .Y(_14915_));
 sg13g2_nor2b_1 _22240_ (.A(\u_inv.d_reg[140] ),
    .B_N(\u_inv.d_next[140] ),
    .Y(_14916_));
 sg13g2_a21oi_1 _22241_ (.A1(net4430),
    .A2(_14916_),
    .Y(_14917_),
    .B1(_14915_));
 sg13g2_nor2b_1 _22242_ (.A(\u_inv.d_reg[142] ),
    .B_N(\u_inv.d_next[142] ),
    .Y(_14918_));
 sg13g2_nand2_1 _22243_ (.Y(_14919_),
    .A(\u_inv.d_next[142] ),
    .B(_10917_));
 sg13g2_a21oi_1 _22244_ (.A1(_14830_),
    .A2(_14918_),
    .Y(_14920_),
    .B1(_14829_));
 sg13g2_o21ai_1 _22245_ (.B1(_14920_),
    .Y(_14921_),
    .A1(_14836_),
    .A2(_14917_));
 sg13g2_nor2b_1 _22246_ (.A(\u_inv.d_reg[137] ),
    .B_N(\u_inv.d_next[137] ),
    .Y(_14922_));
 sg13g2_nor2b_1 _22247_ (.A(\u_inv.d_reg[136] ),
    .B_N(\u_inv.d_next[136] ),
    .Y(_14923_));
 sg13g2_a21oi_1 _22248_ (.A1(_14856_),
    .A2(_14923_),
    .Y(_14924_),
    .B1(_14922_));
 sg13g2_nor2b_1 _22249_ (.A(net4777),
    .B_N(\u_inv.d_next[138] ),
    .Y(_14925_));
 sg13g2_a21oi_1 _22250_ (.A1(_14844_),
    .A2(_14925_),
    .Y(_14926_),
    .B1(_14845_));
 sg13g2_o21ai_1 _22251_ (.B1(_14926_),
    .Y(_14927_),
    .A1(_14852_),
    .A2(_14924_));
 sg13g2_a21oi_1 _22252_ (.A1(_14843_),
    .A2(_14927_),
    .Y(_14928_),
    .B1(_14921_));
 sg13g2_o21ai_1 _22253_ (.B1(_14928_),
    .Y(_14929_),
    .A1(_14861_),
    .A2(_14914_));
 sg13g2_nand2_1 _22254_ (.Y(_14930_),
    .A(_14828_),
    .B(_14929_));
 sg13g2_nor2b_1 _22255_ (.A(\u_inv.d_reg[144] ),
    .B_N(\u_inv.d_next[144] ),
    .Y(_14931_));
 sg13g2_a21oi_1 _22256_ (.A1(_14820_),
    .A2(_14931_),
    .Y(_14932_),
    .B1(_14819_));
 sg13g2_nor2b_1 _22257_ (.A(\u_inv.d_reg[146] ),
    .B_N(\u_inv.d_next[146] ),
    .Y(_14933_));
 sg13g2_a21oi_1 _22258_ (.A1(_14810_),
    .A2(_14933_),
    .Y(_14934_),
    .B1(_14811_));
 sg13g2_o21ai_1 _22259_ (.B1(_14934_),
    .Y(_14935_),
    .A1(_14818_),
    .A2(_14932_));
 sg13g2_inv_1 _22260_ (.Y(_14936_),
    .A(_14935_));
 sg13g2_nand2_1 _22261_ (.Y(_14937_),
    .A(_14809_),
    .B(_14935_));
 sg13g2_nand2b_1 _22262_ (.Y(_14938_),
    .B(\u_inv.d_next[150] ),
    .A_N(net4776));
 sg13g2_a21oi_1 _22263_ (.A1(_10599_),
    .A2(\u_inv.d_reg[151] ),
    .Y(_14939_),
    .B1(_14938_));
 sg13g2_a21oi_1 _22264_ (.A1(\u_inv.d_next[151] ),
    .A2(_10916_),
    .Y(_14940_),
    .B1(_14939_));
 sg13g2_nor2b_1 _22265_ (.A(\u_inv.d_reg[149] ),
    .B_N(\u_inv.d_next[149] ),
    .Y(_14941_));
 sg13g2_nor2b_1 _22266_ (.A(\u_inv.d_reg[148] ),
    .B_N(\u_inv.d_next[148] ),
    .Y(_14942_));
 sg13g2_a21o_1 _22267_ (.A2(_14942_),
    .A1(_14804_),
    .B1(_14941_),
    .X(_14943_));
 sg13g2_nand2_1 _22268_ (.Y(_14944_),
    .A(_14802_),
    .B(_14943_));
 sg13g2_and3_2 _22269_ (.X(_14945_),
    .A(_14937_),
    .B(_14940_),
    .C(_14944_));
 sg13g2_nand3_1 _22270_ (.B(_14940_),
    .C(_14944_),
    .A(_14937_),
    .Y(_14946_));
 sg13g2_nand2_1 _22271_ (.Y(_14947_),
    .A(_14796_),
    .B(_14946_));
 sg13g2_nor2b_1 _22272_ (.A(\u_inv.d_reg[152] ),
    .B_N(\u_inv.d_next[152] ),
    .Y(_14948_));
 sg13g2_a21o_1 _22273_ (.A2(_14948_),
    .A1(_14789_),
    .B1(_14788_),
    .X(_14949_));
 sg13g2_nand2b_1 _22274_ (.Y(_14950_),
    .B(\u_inv.d_next[154] ),
    .A_N(\u_inv.d_reg[154] ));
 sg13g2_a22oi_1 _22275_ (.Y(_14951_),
    .B1(_14787_),
    .B2(_14949_),
    .A2(_10915_),
    .A1(\u_inv.d_next[155] ));
 sg13g2_o21ai_1 _22276_ (.B1(_14951_),
    .Y(_14952_),
    .A1(_14783_),
    .A2(_14950_));
 sg13g2_nand2b_1 _22277_ (.Y(_14953_),
    .B(\u_inv.d_next[156] ),
    .A_N(\u_inv.d_reg[156] ));
 sg13g2_o21ai_1 _22278_ (.B1(_14953_),
    .Y(_14954_),
    .A1(_10598_),
    .A2(\u_inv.d_reg[157] ));
 sg13g2_o21ai_1 _22279_ (.B1(_14954_),
    .Y(_14955_),
    .A1(\u_inv.d_next[157] ),
    .A2(_10914_));
 sg13g2_nor2b_1 _22280_ (.A(\u_inv.d_reg[158] ),
    .B_N(\u_inv.d_next[158] ),
    .Y(_14956_));
 sg13g2_nor2_1 _22281_ (.A(_10597_),
    .B(\u_inv.d_reg[159] ),
    .Y(_14957_));
 sg13g2_a21oi_1 _22282_ (.A1(_14770_),
    .A2(_14956_),
    .Y(_14958_),
    .B1(_14957_));
 sg13g2_o21ai_1 _22283_ (.B1(_14958_),
    .Y(_14959_),
    .A1(_14774_),
    .A2(_14955_));
 sg13g2_a21o_1 _22284_ (.A2(_14952_),
    .A1(_14782_),
    .B1(_14959_),
    .X(_14960_));
 sg13g2_a221oi_1 _22285_ (.B2(_14796_),
    .C1(_14960_),
    .B1(_14946_),
    .A1(_14828_),
    .Y(_14961_),
    .A2(_14929_));
 sg13g2_nand3b_1 _22286_ (.B(_14947_),
    .C(_14930_),
    .Y(_14962_),
    .A_N(_14960_));
 sg13g2_nor2b_2 _22287_ (.A(_14961_),
    .B_N(_14769_),
    .Y(_14963_));
 sg13g2_nor2b_1 _22288_ (.A(\u_inv.d_reg[176] ),
    .B_N(\u_inv.d_next[176] ),
    .Y(_14964_));
 sg13g2_a21o_1 _22289_ (.A2(_14964_),
    .A1(_14705_),
    .B1(_14704_),
    .X(_14965_));
 sg13g2_nand2b_1 _22290_ (.Y(_14966_),
    .B(\u_inv.d_next[178] ),
    .A_N(\u_inv.d_reg[178] ));
 sg13g2_a22oi_1 _22291_ (.Y(_14967_),
    .B1(_14703_),
    .B2(_14965_),
    .A2(_10905_),
    .A1(\u_inv.d_next[179] ));
 sg13g2_o21ai_1 _22292_ (.B1(_14967_),
    .Y(_14968_),
    .A1(_14697_),
    .A2(_14966_));
 sg13g2_nand2b_1 _22293_ (.Y(_14969_),
    .B(\u_inv.d_next[180] ),
    .A_N(\u_inv.d_reg[180] ));
 sg13g2_o21ai_1 _22294_ (.B1(_14969_),
    .Y(_14970_),
    .A1(_10592_),
    .A2(\u_inv.d_reg[181] ));
 sg13g2_o21ai_1 _22295_ (.B1(_14970_),
    .Y(_14971_),
    .A1(\u_inv.d_next[181] ),
    .A2(_10904_));
 sg13g2_nor2b_1 _22296_ (.A(\u_inv.d_reg[182] ),
    .B_N(\u_inv.d_next[182] ),
    .Y(_14972_));
 sg13g2_nor2b_1 _22297_ (.A(_14971_),
    .B_N(_14695_),
    .Y(_14973_));
 sg13g2_o21ai_1 _22298_ (.B1(_14693_),
    .Y(_14974_),
    .A1(_14972_),
    .A2(_14973_));
 sg13g2_a22oi_1 _22299_ (.Y(_14975_),
    .B1(_14696_),
    .B2(_14968_),
    .A2(_10902_),
    .A1(\u_inv.d_next[183] ));
 sg13g2_nand2_2 _22300_ (.Y(_14976_),
    .A(_14974_),
    .B(_14975_));
 sg13g2_and2_1 _22301_ (.A(_14686_),
    .B(_14976_),
    .X(_14977_));
 sg13g2_nor2b_1 _22302_ (.A(\u_inv.d_reg[188] ),
    .B_N(\u_inv.d_next[188] ),
    .Y(_14978_));
 sg13g2_nand2b_1 _22303_ (.Y(_14979_),
    .B(_14978_),
    .A_N(_14666_));
 sg13g2_o21ai_1 _22304_ (.B1(_14979_),
    .Y(_14980_),
    .A1(_10589_),
    .A2(\u_inv.d_reg[189] ));
 sg13g2_inv_1 _22305_ (.Y(_14981_),
    .A(_14980_));
 sg13g2_nor2b_1 _22306_ (.A(\u_inv.d_reg[190] ),
    .B_N(\u_inv.d_next[190] ),
    .Y(_14982_));
 sg13g2_nand2b_1 _22307_ (.Y(_14983_),
    .B(_14982_),
    .A_N(_14661_));
 sg13g2_o21ai_1 _22308_ (.B1(_14983_),
    .Y(_14984_),
    .A1(_10588_),
    .A2(\u_inv.d_reg[191] ));
 sg13g2_a21oi_1 _22309_ (.A1(_14665_),
    .A2(_14980_),
    .Y(_14985_),
    .B1(_14984_));
 sg13g2_nand2b_1 _22310_ (.Y(_14986_),
    .B(\u_inv.d_next[184] ),
    .A_N(\u_inv.d_reg[184] ));
 sg13g2_o21ai_1 _22311_ (.B1(_14986_),
    .Y(_14987_),
    .A1(_10591_),
    .A2(\u_inv.d_reg[185] ));
 sg13g2_and2_1 _22312_ (.A(_14672_),
    .B(_14987_),
    .X(_14988_));
 sg13g2_nand2_1 _22313_ (.Y(_14989_),
    .A(_14672_),
    .B(_14987_));
 sg13g2_nor2_1 _22314_ (.A(_10590_),
    .B(\u_inv.d_reg[186] ),
    .Y(_14990_));
 sg13g2_nor2b_1 _22315_ (.A(net4774),
    .B_N(\u_inv.d_next[187] ),
    .Y(_14991_));
 sg13g2_a221oi_1 _22316_ (.B2(_14682_),
    .C1(_14991_),
    .B1(_14990_),
    .A1(_14683_),
    .Y(_14992_),
    .A2(_14988_));
 sg13g2_o21ai_1 _22317_ (.B1(_14985_),
    .Y(_14993_),
    .A1(_14671_),
    .A2(_14992_));
 sg13g2_nor2b_1 _22318_ (.A(\u_inv.d_reg[160] ),
    .B_N(\u_inv.d_next[160] ),
    .Y(_14994_));
 sg13g2_a21oi_1 _22319_ (.A1(_14759_),
    .A2(_14994_),
    .Y(_14995_),
    .B1(_14758_));
 sg13g2_nor2b_1 _22320_ (.A(net4775),
    .B_N(net4801),
    .Y(_14996_));
 sg13g2_a21oi_1 _22321_ (.A1(_14749_),
    .A2(_14996_),
    .Y(_14997_),
    .B1(_14750_));
 sg13g2_o21ai_1 _22322_ (.B1(_14997_),
    .Y(_14998_),
    .A1(_14757_),
    .A2(_14995_));
 sg13g2_inv_1 _22323_ (.Y(_14999_),
    .A(_14998_));
 sg13g2_nand2_1 _22324_ (.Y(_15000_),
    .A(\u_inv.d_next[166] ),
    .B(_10911_));
 sg13g2_o21ai_1 _22325_ (.B1(_14735_),
    .Y(_15001_),
    .A1(_14736_),
    .A2(_15000_));
 sg13g2_nor2b_1 _22326_ (.A(\u_inv.d_reg[165] ),
    .B_N(\u_inv.d_next[165] ),
    .Y(_15002_));
 sg13g2_nor2_1 _22327_ (.A(_10596_),
    .B(\u_inv.d_reg[164] ),
    .Y(_15003_));
 sg13g2_a21o_1 _22328_ (.A2(_15003_),
    .A1(_14743_),
    .B1(_15002_),
    .X(_15004_));
 sg13g2_a221oi_1 _22329_ (.B2(_14741_),
    .C1(_15001_),
    .B1(_15004_),
    .A1(_14748_),
    .Y(_15005_),
    .A2(_14998_));
 sg13g2_nor4_1 _22330_ (.A(_14724_),
    .B(_14730_),
    .C(_14734_),
    .D(_15005_),
    .Y(_15006_));
 sg13g2_nor2b_1 _22331_ (.A(\u_inv.d_reg[168] ),
    .B_N(\u_inv.d_next[168] ),
    .Y(_15007_));
 sg13g2_a21oi_1 _22332_ (.A1(\u_inv.d_next[169] ),
    .A2(_10909_),
    .Y(_15008_),
    .B1(_15007_));
 sg13g2_a21oi_2 _22333_ (.B1(_15008_),
    .Y(_15009_),
    .A2(\u_inv.d_reg[169] ),
    .A1(_10595_));
 sg13g2_nand2b_1 _22334_ (.Y(_15010_),
    .B(\u_inv.d_next[170] ),
    .A_N(\u_inv.d_reg[170] ));
 sg13g2_a21oi_1 _22335_ (.A1(_10594_),
    .A2(\u_inv.d_reg[171] ),
    .Y(_15011_),
    .B1(_15010_));
 sg13g2_a22oi_1 _22336_ (.Y(_15012_),
    .B1(_14729_),
    .B2(_15009_),
    .A2(_10908_),
    .A1(\u_inv.d_next[171] ));
 sg13g2_a221oi_1 _22337_ (.B2(_15009_),
    .C1(_15011_),
    .B1(_14729_),
    .A1(\u_inv.d_next[171] ),
    .Y(_15013_),
    .A2(_10908_));
 sg13g2_nand2b_1 _22338_ (.Y(_15014_),
    .B(_15012_),
    .A_N(_15011_));
 sg13g2_nand2b_1 _22339_ (.Y(_15015_),
    .B(\u_inv.d_next[172] ),
    .A_N(\u_inv.d_reg[172] ));
 sg13g2_o21ai_1 _22340_ (.B1(_15015_),
    .Y(_15016_),
    .A1(_10593_),
    .A2(\u_inv.d_reg[173] ));
 sg13g2_and2_1 _22341_ (.A(_14718_),
    .B(_15016_),
    .X(_15017_));
 sg13g2_nand2_1 _22342_ (.Y(_15018_),
    .A(_14718_),
    .B(_15016_));
 sg13g2_nor2b_1 _22343_ (.A(\u_inv.d_reg[175] ),
    .B_N(\u_inv.d_next[175] ),
    .Y(_15019_));
 sg13g2_nor2b_1 _22344_ (.A(\u_inv.d_reg[174] ),
    .B_N(\u_inv.d_next[174] ),
    .Y(_15020_));
 sg13g2_a22oi_1 _22345_ (.Y(_15021_),
    .B1(_15020_),
    .B2(_14714_),
    .A2(_15017_),
    .A1(_14717_));
 sg13g2_o21ai_1 _22346_ (.B1(_15021_),
    .Y(_15022_),
    .A1(_14724_),
    .A2(_15013_));
 sg13g2_nor3_2 _22347_ (.A(_15006_),
    .B(_15019_),
    .C(_15022_),
    .Y(_15023_));
 sg13g2_nor2_1 _22348_ (.A(_14712_),
    .B(_15023_),
    .Y(_15024_));
 sg13g2_nor4_2 _22349_ (.A(_14963_),
    .B(_14977_),
    .C(_14993_),
    .Y(_15025_),
    .D(_15024_));
 sg13g2_inv_1 _22350_ (.Y(_15026_),
    .A(_15025_));
 sg13g2_or2_1 _22351_ (.X(_15027_),
    .B(_14900_),
    .A(_13831_));
 sg13g2_a21oi_2 _22352_ (.B1(_15027_),
    .Y(_15028_),
    .A2(_14656_),
    .A1(_14537_));
 sg13g2_nor2_2 _22353_ (.A(_13831_),
    .B(_15025_),
    .Y(_15029_));
 sg13g2_o21ai_1 _22354_ (.B1(_13894_),
    .Y(_15030_),
    .A1(_13713_),
    .A2(_13955_));
 sg13g2_or3_1 _22355_ (.A(_13861_),
    .B(_15029_),
    .C(_15030_),
    .X(_15031_));
 sg13g2_o21ai_1 _22356_ (.B1(_13600_),
    .Y(_15032_),
    .A1(_15028_),
    .A2(_15031_));
 sg13g2_and2_1 _22357_ (.A(net3755),
    .B(_15032_),
    .X(_15033_));
 sg13g2_nand3_1 _22358_ (.B(_13598_),
    .C(_15032_),
    .A(net3755),
    .Y(_15034_));
 sg13g2_nand2b_1 _22359_ (.Y(_15035_),
    .B(_13604_),
    .A_N(_13602_));
 sg13g2_inv_1 _22360_ (.Y(_15036_),
    .A(_15035_));
 sg13g2_nor2_1 _22361_ (.A(_13609_),
    .B(_13611_),
    .Y(_15037_));
 sg13g2_nand2_1 _22362_ (.Y(_15038_),
    .A(_15036_),
    .B(_15037_));
 sg13g2_nor2_1 _22363_ (.A(_13616_),
    .B(_13619_),
    .Y(_15039_));
 sg13g2_or2_1 _22364_ (.X(_15040_),
    .B(_13625_),
    .A(_13623_));
 sg13g2_nor4_2 _22365_ (.A(_13616_),
    .B(_13619_),
    .C(_15038_),
    .Y(_15041_),
    .D(_15040_));
 sg13g2_or2_1 _22366_ (.X(_15042_),
    .B(_13644_),
    .A(_13642_));
 sg13g2_nor2_1 _22367_ (.A(_13630_),
    .B(_13639_),
    .Y(_15043_));
 sg13g2_nor2_1 _22368_ (.A(_13648_),
    .B(_13651_),
    .Y(_15044_));
 sg13g2_nand3_1 _22369_ (.B(_13654_),
    .C(_15044_),
    .A(_13636_),
    .Y(_15045_));
 sg13g2_nor4_1 _22370_ (.A(_13630_),
    .B(_13639_),
    .C(_15042_),
    .D(_15045_),
    .Y(_15046_));
 sg13g2_nand2_2 _22371_ (.Y(_15047_),
    .A(_15041_),
    .B(_15046_));
 sg13g2_nand2_1 _22372_ (.Y(_15048_),
    .A(_13677_),
    .B(_13679_));
 sg13g2_or2_1 _22373_ (.X(_15049_),
    .B(_13673_),
    .A(_13671_));
 sg13g2_nor2_1 _22374_ (.A(_15048_),
    .B(_15049_),
    .Y(_15050_));
 sg13g2_nor2_1 _22375_ (.A(_13659_),
    .B(_13667_),
    .Y(_15051_));
 sg13g2_nor2_1 _22376_ (.A(_13661_),
    .B(_13664_),
    .Y(_15052_));
 sg13g2_nand3_1 _22377_ (.B(_15051_),
    .C(_15052_),
    .A(_15050_),
    .Y(_15053_));
 sg13g2_nand2_1 _22378_ (.Y(_15054_),
    .A(_13683_),
    .B(_13685_));
 sg13g2_nor2_1 _22379_ (.A(_13690_),
    .B(_13693_),
    .Y(_15055_));
 sg13g2_nand2b_1 _22380_ (.Y(_15056_),
    .B(_15055_),
    .A_N(_15054_));
 sg13g2_or4_1 _22381_ (.A(_13698_),
    .B(_13702_),
    .C(_13706_),
    .D(_13708_),
    .X(_15057_));
 sg13g2_or2_1 _22382_ (.X(_15058_),
    .B(_15057_),
    .A(_15056_));
 sg13g2_or2_1 _22383_ (.X(_15059_),
    .B(_15058_),
    .A(_15053_));
 sg13g2_nor2_2 _22384_ (.A(_15047_),
    .B(_15059_),
    .Y(_15060_));
 sg13g2_nor2_1 _22385_ (.A(_13778_),
    .B(_13780_),
    .Y(_15061_));
 sg13g2_nand3_1 _22386_ (.B(_13785_),
    .C(_15061_),
    .A(_13782_),
    .Y(_15062_));
 sg13g2_and2_1 _22387_ (.A(_13792_),
    .B(_13797_),
    .X(_15063_));
 sg13g2_inv_1 _22388_ (.Y(_15064_),
    .A(_15063_));
 sg13g2_nand2_1 _22389_ (.Y(_15065_),
    .A(_13789_),
    .B(_13795_));
 sg13g2_nor3_1 _22390_ (.A(_15062_),
    .B(_15064_),
    .C(_15065_),
    .Y(_15066_));
 sg13g2_nor2_1 _22391_ (.A(_13801_),
    .B(_13803_),
    .Y(_15067_));
 sg13g2_nor2_1 _22392_ (.A(_13807_),
    .B(_13810_),
    .Y(_15068_));
 sg13g2_nand2_1 _22393_ (.Y(_15069_),
    .A(_15067_),
    .B(_15068_));
 sg13g2_nand2_1 _22394_ (.Y(_15070_),
    .A(\u_inv.d_next[211] ),
    .B(\u_inv.d_reg[211] ));
 sg13g2_and2_1 _22395_ (.A(\u_inv.d_next[209] ),
    .B(net4769),
    .X(_15071_));
 sg13g2_a21oi_1 _22396_ (.A1(_13823_),
    .A2(_13824_),
    .Y(_15072_),
    .B1(_15071_));
 sg13g2_inv_1 _22397_ (.Y(_15073_),
    .A(_15072_));
 sg13g2_a21o_1 _22398_ (.A2(_15072_),
    .A1(_13817_),
    .B1(_13816_),
    .X(_15074_));
 sg13g2_o21ai_1 _22399_ (.B1(_15070_),
    .Y(_15075_),
    .A1(_13815_),
    .A2(_15074_));
 sg13g2_nand2b_1 _22400_ (.Y(_15076_),
    .B(_15075_),
    .A_N(_15069_));
 sg13g2_nor2_1 _22401_ (.A(_13807_),
    .B(_13808_),
    .Y(_15077_));
 sg13g2_a21oi_1 _22402_ (.A1(\u_inv.d_next[213] ),
    .A2(\u_inv.d_reg[213] ),
    .Y(_15078_),
    .B1(_15077_));
 sg13g2_nand2b_1 _22403_ (.Y(_15079_),
    .B(_15067_),
    .A_N(_15078_));
 sg13g2_nor2_1 _22404_ (.A(_13800_),
    .B(_13802_),
    .Y(_15080_));
 sg13g2_a21oi_1 _22405_ (.A1(\u_inv.d_next[215] ),
    .A2(\u_inv.d_reg[215] ),
    .Y(_15081_),
    .B1(_15080_));
 sg13g2_nand3_1 _22406_ (.B(_15079_),
    .C(_15081_),
    .A(_15076_),
    .Y(_15082_));
 sg13g2_nor2b_1 _22407_ (.A(_13788_),
    .B_N(_13795_),
    .Y(_15083_));
 sg13g2_a21oi_1 _22408_ (.A1(\u_inv.d_next[217] ),
    .A2(\u_inv.d_reg[217] ),
    .Y(_15084_),
    .B1(_15083_));
 sg13g2_a21o_1 _22409_ (.A2(\u_inv.d_reg[217] ),
    .A1(\u_inv.d_next[217] ),
    .B1(_15083_),
    .X(_15085_));
 sg13g2_o21ai_1 _22410_ (.B1(_13791_),
    .Y(_15086_),
    .A1(\u_inv.d_next[219] ),
    .A2(\u_inv.d_reg[219] ));
 sg13g2_nand2_1 _22411_ (.Y(_15087_),
    .A(_13796_),
    .B(_15086_));
 sg13g2_a21oi_1 _22412_ (.A1(_15063_),
    .A2(_15085_),
    .Y(_15088_),
    .B1(_15087_));
 sg13g2_or2_1 _22413_ (.X(_15089_),
    .B(_15088_),
    .A(_15062_));
 sg13g2_o21ai_1 _22414_ (.B1(_13777_),
    .Y(_15090_),
    .A1(_13776_),
    .A2(_13779_));
 sg13g2_nand3_1 _22415_ (.B(_13785_),
    .C(_15090_),
    .A(_13782_),
    .Y(_15091_));
 sg13g2_a21oi_1 _22416_ (.A1(_10580_),
    .A2(_10888_),
    .Y(_15092_),
    .B1(_13783_));
 sg13g2_a21oi_1 _22417_ (.A1(\u_inv.d_next[223] ),
    .A2(\u_inv.d_reg[223] ),
    .Y(_15093_),
    .B1(_15092_));
 sg13g2_nand2b_1 _22418_ (.Y(_15094_),
    .B(_13818_),
    .A_N(_13815_));
 sg13g2_nor4_1 _22419_ (.A(_13822_),
    .B(net4431),
    .C(_15069_),
    .D(_15094_),
    .Y(_15095_));
 sg13g2_and2_1 _22420_ (.A(_15066_),
    .B(_15095_),
    .X(_15096_));
 sg13g2_or2_1 _22421_ (.X(_15097_),
    .B(_13717_),
    .A(_13715_));
 sg13g2_nand2_1 _22422_ (.Y(_15098_),
    .A(_13722_),
    .B(_13724_));
 sg13g2_inv_1 _22423_ (.Y(_15099_),
    .A(_15098_));
 sg13g2_nor2_1 _22424_ (.A(_15097_),
    .B(_15098_),
    .Y(_15100_));
 sg13g2_nand2_1 _22425_ (.Y(_15101_),
    .A(_13736_),
    .B(_13740_));
 sg13g2_nand2b_1 _22426_ (.Y(_15102_),
    .B(_13729_),
    .A_N(_13731_));
 sg13g2_nor4_1 _22427_ (.A(_15097_),
    .B(_15098_),
    .C(_15101_),
    .D(_15102_),
    .Y(_15103_));
 sg13g2_nor2_1 _22428_ (.A(_13754_),
    .B(_13757_),
    .Y(_15104_));
 sg13g2_nand3_1 _22429_ (.B(_13749_),
    .C(_15104_),
    .A(_13746_),
    .Y(_15105_));
 sg13g2_and2_1 _22430_ (.A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ),
    .X(_15106_));
 sg13g2_a22oi_1 _22431_ (.Y(_15107_),
    .B1(\u_inv.d_reg[193] ),
    .B2(\u_inv.d_next[193] ),
    .A2(\u_inv.d_reg[194] ),
    .A1(\u_inv.d_next[194] ));
 sg13g2_o21ai_1 _22432_ (.B1(_15107_),
    .Y(_15108_),
    .A1(_13769_),
    .A2(_13771_));
 sg13g2_a21oi_1 _22433_ (.A1(_10587_),
    .A2(_10898_),
    .Y(_15109_),
    .B1(_13762_));
 sg13g2_a22oi_1 _22434_ (.Y(_15110_),
    .B1(_15108_),
    .B2(_15109_),
    .A2(\u_inv.d_reg[195] ),
    .A1(\u_inv.d_next[195] ));
 sg13g2_inv_1 _22435_ (.Y(_15111_),
    .A(_15110_));
 sg13g2_a22oi_1 _22436_ (.Y(_15112_),
    .B1(net4773),
    .B2(\u_inv.d_next[196] ),
    .A2(net4772),
    .A1(\u_inv.d_next[197] ));
 sg13g2_nor2_1 _22437_ (.A(_13752_),
    .B(_15112_),
    .Y(_15113_));
 sg13g2_o21ai_1 _22438_ (.B1(_13747_),
    .Y(_15114_),
    .A1(_13752_),
    .A2(_15112_));
 sg13g2_nor2_1 _22439_ (.A(_13745_),
    .B(_13748_),
    .Y(_15115_));
 sg13g2_a22oi_1 _22440_ (.Y(_15116_),
    .B1(_15114_),
    .B2(_15115_),
    .A2(\u_inv.d_reg[199] ),
    .A1(\u_inv.d_next[199] ));
 sg13g2_o21ai_1 _22441_ (.B1(_15116_),
    .Y(_15117_),
    .A1(_15105_),
    .A2(_15110_));
 sg13g2_nand2_1 _22442_ (.Y(_15118_),
    .A(\u_inv.d_next[203] ),
    .B(\u_inv.d_reg[203] ));
 sg13g2_nand2b_1 _22443_ (.Y(_15119_),
    .B(_13729_),
    .A_N(_13730_));
 sg13g2_nand2_1 _22444_ (.Y(_15120_),
    .A(\u_inv.d_next[201] ),
    .B(\u_inv.d_reg[201] ));
 sg13g2_and2_1 _22445_ (.A(_15119_),
    .B(_15120_),
    .X(_15121_));
 sg13g2_o21ai_1 _22446_ (.B1(_15120_),
    .Y(_15122_),
    .A1(_13728_),
    .A2(_13730_));
 sg13g2_o21ai_1 _22447_ (.B1(_13740_),
    .Y(_15123_),
    .A1(_13735_),
    .A2(_15122_));
 sg13g2_o21ai_1 _22448_ (.B1(_15118_),
    .Y(_15124_),
    .A1(_13734_),
    .A2(_15123_));
 sg13g2_nor2_1 _22449_ (.A(_13714_),
    .B(_13716_),
    .Y(_15125_));
 sg13g2_a21oi_1 _22450_ (.A1(\u_inv.d_next[207] ),
    .A2(\u_inv.d_reg[207] ),
    .Y(_15126_),
    .B1(_15125_));
 sg13g2_nor2_1 _22451_ (.A(_13721_),
    .B(_13723_),
    .Y(_15127_));
 sg13g2_a21oi_1 _22452_ (.A1(\u_inv.d_next[205] ),
    .A2(\u_inv.d_reg[205] ),
    .Y(_15128_),
    .B1(_15127_));
 sg13g2_nor2_1 _22453_ (.A(_15097_),
    .B(_15128_),
    .Y(_15129_));
 sg13g2_a221oi_1 _22454_ (.B2(_15100_),
    .C1(_15129_),
    .B1(_15124_),
    .A1(_15103_),
    .Y(_15130_),
    .A2(_15117_));
 sg13g2_nand2_2 _22455_ (.Y(_15131_),
    .A(_15126_),
    .B(_15130_));
 sg13g2_a22oi_1 _22456_ (.Y(_15132_),
    .B1(_15096_),
    .B2(_15131_),
    .A2(_15082_),
    .A1(_15066_));
 sg13g2_nand4_1 _22457_ (.B(_15091_),
    .C(_15093_),
    .A(_15089_),
    .Y(_15133_),
    .D(_15132_));
 sg13g2_nand2_1 _22458_ (.Y(_15134_),
    .A(_15060_),
    .B(_15133_));
 sg13g2_a21oi_1 _22459_ (.A1(_10578_),
    .A2(_10885_),
    .Y(_15135_),
    .B1(_13643_));
 sg13g2_a21oi_1 _22460_ (.A1(\u_inv.d_next[245] ),
    .A2(\u_inv.d_reg[245] ),
    .Y(_15136_),
    .B1(_15135_));
 sg13g2_a21oi_1 _22461_ (.A1(_13629_),
    .A2(_13637_),
    .Y(_15137_),
    .B1(_13638_));
 sg13g2_nand2_1 _22462_ (.Y(_15138_),
    .A(\u_inv.d_next[241] ),
    .B(\u_inv.d_reg[241] ));
 sg13g2_nand2b_1 _22463_ (.Y(_15139_),
    .B(_13636_),
    .A_N(_13653_));
 sg13g2_and2_1 _22464_ (.A(_15138_),
    .B(_15139_),
    .X(_15140_));
 sg13g2_nand2_1 _22465_ (.Y(_15141_),
    .A(_15138_),
    .B(_15139_));
 sg13g2_a21oi_1 _22466_ (.A1(_15043_),
    .A2(_15141_),
    .Y(_15142_),
    .B1(_15137_));
 sg13g2_o21ai_1 _22467_ (.B1(_15136_),
    .Y(_15143_),
    .A1(_15042_),
    .A2(_15142_));
 sg13g2_a21oi_1 _22468_ (.A1(\u_inv.d_next[247] ),
    .A2(\u_inv.d_reg[247] ),
    .Y(_15144_),
    .B1(_13649_));
 sg13g2_nor2_1 _22469_ (.A(_13646_),
    .B(_15144_),
    .Y(_15145_));
 sg13g2_a21oi_1 _22470_ (.A1(_15044_),
    .A2(_15143_),
    .Y(_15146_),
    .B1(_15145_));
 sg13g2_inv_1 _22471_ (.Y(_15147_),
    .A(_15146_));
 sg13g2_nand2_2 _22472_ (.Y(_15148_),
    .A(_15041_),
    .B(_15147_));
 sg13g2_nand2_1 _22473_ (.Y(_15149_),
    .A(\u_inv.d_next[225] ),
    .B(\u_inv.d_reg[225] ));
 sg13g2_a22oi_1 _22474_ (.Y(_15150_),
    .B1(\u_inv.d_reg[225] ),
    .B2(\u_inv.d_next[225] ),
    .A2(net4768),
    .A1(\u_inv.d_next[226] ));
 sg13g2_o21ai_1 _22475_ (.B1(_15150_),
    .Y(_15151_),
    .A1(_13706_),
    .A2(_13707_));
 sg13g2_nor2_1 _22476_ (.A(_13698_),
    .B(_13700_),
    .Y(_15152_));
 sg13g2_a22oi_1 _22477_ (.Y(_15153_),
    .B1(_15151_),
    .B2(_15152_),
    .A2(\u_inv.d_reg[227] ),
    .A1(\u_inv.d_next[227] ));
 sg13g2_or2_1 _22478_ (.X(_15154_),
    .B(_13691_),
    .A(_13690_));
 sg13g2_nand2_1 _22479_ (.Y(_15155_),
    .A(\u_inv.d_next[229] ),
    .B(net4766));
 sg13g2_and2_1 _22480_ (.A(_15154_),
    .B(_15155_),
    .X(_15156_));
 sg13g2_nor2_1 _22481_ (.A(_15054_),
    .B(_15156_),
    .Y(_15157_));
 sg13g2_nor2_1 _22482_ (.A(_13682_),
    .B(_13684_),
    .Y(_15158_));
 sg13g2_a21oi_1 _22483_ (.A1(\u_inv.d_next[231] ),
    .A2(\u_inv.d_reg[231] ),
    .Y(_15159_),
    .B1(_15158_));
 sg13g2_o21ai_1 _22484_ (.B1(_15159_),
    .Y(_15160_),
    .A1(_15056_),
    .A2(_15153_));
 sg13g2_nor2_1 _22485_ (.A(_15157_),
    .B(_15160_),
    .Y(_15161_));
 sg13g2_o21ai_1 _22486_ (.B1(_13670_),
    .Y(_15162_),
    .A1(_13669_),
    .A2(_13672_));
 sg13g2_inv_1 _22487_ (.Y(_15163_),
    .A(_15162_));
 sg13g2_nand2b_1 _22488_ (.Y(_15164_),
    .B(_15162_),
    .A_N(_15048_));
 sg13g2_o21ai_1 _22489_ (.B1(_13678_),
    .Y(_15165_),
    .A1(\u_inv.d_next[239] ),
    .A2(\u_inv.d_reg[239] ));
 sg13g2_nand3_1 _22490_ (.B(_15164_),
    .C(_15165_),
    .A(_13676_),
    .Y(_15166_));
 sg13g2_nor2_1 _22491_ (.A(_13660_),
    .B(_13664_),
    .Y(_15167_));
 sg13g2_a21oi_1 _22492_ (.A1(\u_inv.d_next[233] ),
    .A2(\u_inv.d_reg[233] ),
    .Y(_15168_),
    .B1(_15167_));
 sg13g2_nor2b_1 _22493_ (.A(_15168_),
    .B_N(_15051_),
    .Y(_15169_));
 sg13g2_o21ai_1 _22494_ (.B1(_13666_),
    .Y(_15170_),
    .A1(_13657_),
    .A2(_13665_));
 sg13g2_o21ai_1 _22495_ (.B1(_15050_),
    .Y(_15171_),
    .A1(_15169_),
    .A2(_15170_));
 sg13g2_o21ai_1 _22496_ (.B1(_15171_),
    .Y(_15172_),
    .A1(_15053_),
    .A2(_15161_));
 sg13g2_nor2_1 _22497_ (.A(_15166_),
    .B(_15172_),
    .Y(_15173_));
 sg13g2_nor2_1 _22498_ (.A(_15047_),
    .B(_15173_),
    .Y(_15174_));
 sg13g2_o21ai_1 _22499_ (.B1(_13608_),
    .Y(_15175_),
    .A1(_13607_),
    .A2(_13610_));
 sg13g2_nor2_1 _22500_ (.A(_13601_),
    .B(_13603_),
    .Y(_15176_));
 sg13g2_a221oi_1 _22501_ (.B2(_15175_),
    .C1(_15176_),
    .B1(_15036_),
    .A1(\u_inv.d_next[255] ),
    .Y(_15177_),
    .A2(\u_inv.d_reg[255] ));
 sg13g2_o21ai_1 _22502_ (.B1(_13622_),
    .Y(_15178_),
    .A1(_13621_),
    .A2(_13624_));
 sg13g2_a21oi_1 _22503_ (.A1(_13614_),
    .A2(_13617_),
    .Y(_15179_),
    .B1(_13615_));
 sg13g2_a21oi_1 _22504_ (.A1(_15039_),
    .A2(_15178_),
    .Y(_15180_),
    .B1(_15179_));
 sg13g2_o21ai_1 _22505_ (.B1(_15177_),
    .Y(_15181_),
    .A1(_15038_),
    .A2(_15180_));
 sg13g2_nor2_1 _22506_ (.A(_15174_),
    .B(_15181_),
    .Y(_15182_));
 sg13g2_nand3_1 _22507_ (.B(_15148_),
    .C(_15182_),
    .A(_15134_),
    .Y(_15183_));
 sg13g2_nor4_1 _22508_ (.A(_13762_),
    .B(_13764_),
    .C(_13769_),
    .D(_13772_),
    .Y(_15184_));
 sg13g2_nor2b_2 _22509_ (.A(_15105_),
    .B_N(_15184_),
    .Y(_15185_));
 sg13g2_and2_1 _22510_ (.A(_15103_),
    .B(_15185_),
    .X(_15186_));
 sg13g2_and2_1 _22511_ (.A(_15096_),
    .B(_15186_),
    .X(_15187_));
 sg13g2_and2_1 _22512_ (.A(_15060_),
    .B(_15187_),
    .X(_15188_));
 sg13g2_and2_1 _22513_ (.A(_14666_),
    .B(_14668_),
    .X(_15189_));
 sg13g2_nand3_1 _22514_ (.B(_14664_),
    .C(_15189_),
    .A(_14661_),
    .Y(_15190_));
 sg13g2_nor2_1 _22515_ (.A(_14679_),
    .B(_14682_),
    .Y(_15191_));
 sg13g2_nor2b_1 _22516_ (.A(_14673_),
    .B_N(_14675_),
    .Y(_15192_));
 sg13g2_nand2_1 _22517_ (.Y(_15193_),
    .A(_15191_),
    .B(_15192_));
 sg13g2_or2_1 _22518_ (.X(_15194_),
    .B(_15193_),
    .A(_15190_));
 sg13g2_nor2_1 _22519_ (.A(_14687_),
    .B(_14690_),
    .Y(_15195_));
 sg13g2_nor4_1 _22520_ (.A(_14687_),
    .B(_14690_),
    .C(_14693_),
    .D(_14695_),
    .Y(_15196_));
 sg13g2_nor2_2 _22521_ (.A(_14706_),
    .B(_14708_),
    .Y(_15197_));
 sg13g2_nand4_1 _22522_ (.B(_14701_),
    .C(_15196_),
    .A(_14699_),
    .Y(_15198_),
    .D(_15197_));
 sg13g2_or2_1 _22523_ (.X(_15199_),
    .B(_15198_),
    .A(_15194_));
 sg13g2_nor2_1 _22524_ (.A(_14743_),
    .B(_14746_),
    .Y(_15200_));
 sg13g2_nand3_1 _22525_ (.B(_14740_),
    .C(_15200_),
    .A(_14737_),
    .Y(_15201_));
 sg13g2_nor2_1 _22526_ (.A(_14760_),
    .B(_14761_),
    .Y(_15202_));
 sg13g2_a22oi_1 _22527_ (.Y(_15203_),
    .B1(\u_inv.d_reg[161] ),
    .B2(\u_inv.d_next[161] ),
    .A2(net4775),
    .A1(net4801));
 sg13g2_o21ai_1 _22528_ (.B1(_15203_),
    .Y(_15204_),
    .A1(_14760_),
    .A2(_14761_));
 sg13g2_nor2_1 _22529_ (.A(_14751_),
    .B(_14754_),
    .Y(_15205_));
 sg13g2_a22oi_1 _22530_ (.Y(_15206_),
    .B1(_15204_),
    .B2(_15205_),
    .A2(\u_inv.d_reg[163] ),
    .A1(\u_inv.d_next[163] ));
 sg13g2_o21ai_1 _22531_ (.B1(_14744_),
    .Y(_15207_),
    .A1(\u_inv.d_next[165] ),
    .A2(\u_inv.d_reg[165] ));
 sg13g2_nand2_1 _22532_ (.Y(_15208_),
    .A(_14742_),
    .B(_15207_));
 sg13g2_nand2_1 _22533_ (.Y(_15209_),
    .A(_14740_),
    .B(_15208_));
 sg13g2_nand2_1 _22534_ (.Y(_15210_),
    .A(_14738_),
    .B(_15209_));
 sg13g2_nand2_1 _22535_ (.Y(_15211_),
    .A(\u_inv.d_next[167] ),
    .B(\u_inv.d_reg[167] ));
 sg13g2_o21ai_1 _22536_ (.B1(_15211_),
    .Y(_15212_),
    .A1(_15201_),
    .A2(_15206_));
 sg13g2_a21oi_1 _22537_ (.A1(_14737_),
    .A2(_15210_),
    .Y(_15213_),
    .B1(_15212_));
 sg13g2_or2_1 _22538_ (.X(_15214_),
    .B(_14716_),
    .A(_14714_));
 sg13g2_nor2_1 _22539_ (.A(_14719_),
    .B(_14722_),
    .Y(_15215_));
 sg13g2_nor2b_1 _22540_ (.A(_15214_),
    .B_N(_15215_),
    .Y(_15216_));
 sg13g2_o21ai_1 _22541_ (.B1(_14726_),
    .Y(_15217_),
    .A1(\u_inv.d_next[170] ),
    .A2(\u_inv.d_reg[170] ));
 sg13g2_nor2_1 _22542_ (.A(_14725_),
    .B(_14728_),
    .Y(_15218_));
 sg13g2_nor2_2 _22543_ (.A(_14731_),
    .B(_14733_),
    .Y(_15219_));
 sg13g2_nand3_1 _22544_ (.B(_15218_),
    .C(_15219_),
    .A(_15216_),
    .Y(_15220_));
 sg13g2_nor2_1 _22545_ (.A(_14731_),
    .B(_14732_),
    .Y(_15221_));
 sg13g2_a21oi_1 _22546_ (.A1(\u_inv.d_next[169] ),
    .A2(\u_inv.d_reg[169] ),
    .Y(_15222_),
    .B1(_15221_));
 sg13g2_a21oi_1 _22547_ (.A1(_14727_),
    .A2(_15222_),
    .Y(_15223_),
    .B1(_15217_));
 sg13g2_a21o_2 _22548_ (.A2(\u_inv.d_reg[171] ),
    .A1(\u_inv.d_next[171] ),
    .B1(_15223_),
    .X(_15224_));
 sg13g2_nor2_1 _22549_ (.A(_14719_),
    .B(_14720_),
    .Y(_15225_));
 sg13g2_a21oi_1 _22550_ (.A1(\u_inv.d_next[173] ),
    .A2(\u_inv.d_reg[173] ),
    .Y(_15226_),
    .B1(_15225_));
 sg13g2_nor2_1 _22551_ (.A(_14713_),
    .B(_14715_),
    .Y(_15227_));
 sg13g2_a21oi_1 _22552_ (.A1(\u_inv.d_next[175] ),
    .A2(\u_inv.d_reg[175] ),
    .Y(_15228_),
    .B1(_15227_));
 sg13g2_o21ai_1 _22553_ (.B1(_15228_),
    .Y(_15229_),
    .A1(_15214_),
    .A2(_15226_));
 sg13g2_a21oi_1 _22554_ (.A1(_15216_),
    .A2(_15224_),
    .Y(_15230_),
    .B1(_15229_));
 sg13g2_o21ai_1 _22555_ (.B1(_15230_),
    .Y(_15231_),
    .A1(_15213_),
    .A2(_15220_));
 sg13g2_nor2_1 _22556_ (.A(_14760_),
    .B(_14763_),
    .Y(_15232_));
 sg13g2_nand3_1 _22557_ (.B(_14755_),
    .C(_15232_),
    .A(_14752_),
    .Y(_15233_));
 sg13g2_or2_1 _22558_ (.X(_15234_),
    .B(_15233_),
    .A(_15201_));
 sg13g2_nor2_1 _22559_ (.A(_15220_),
    .B(_15234_),
    .Y(_15235_));
 sg13g2_nor2_1 _22560_ (.A(_14770_),
    .B(_14773_),
    .Y(_15236_));
 sg13g2_nand2_1 _22561_ (.Y(_15237_),
    .A(_14776_),
    .B(_14779_));
 sg13g2_nand3_1 _22562_ (.B(_14779_),
    .C(_15236_),
    .A(_14776_),
    .Y(_15238_));
 sg13g2_and2_1 _22563_ (.A(_14790_),
    .B(_14792_),
    .X(_15239_));
 sg13g2_nor2_1 _22564_ (.A(_14784_),
    .B(_14786_),
    .Y(_15240_));
 sg13g2_nand3b_1 _22565_ (.B(_15239_),
    .C(_15240_),
    .Y(_15241_),
    .A_N(_15238_));
 sg13g2_nor2_1 _22566_ (.A(_14804_),
    .B(_14807_),
    .Y(_15242_));
 sg13g2_nand3_1 _22567_ (.B(_14801_),
    .C(_15242_),
    .A(_14797_),
    .Y(_15243_));
 sg13g2_nor2_1 _22568_ (.A(_14821_),
    .B(_14822_),
    .Y(_15244_));
 sg13g2_a21oi_1 _22569_ (.A1(\u_inv.d_next[145] ),
    .A2(\u_inv.d_reg[145] ),
    .Y(_15245_),
    .B1(_15244_));
 sg13g2_a21o_1 _22570_ (.A2(\u_inv.d_reg[145] ),
    .A1(\u_inv.d_next[145] ),
    .B1(_15244_),
    .X(_15246_));
 sg13g2_nor2_1 _22571_ (.A(_14812_),
    .B(_14815_),
    .Y(_15247_));
 sg13g2_nor2_1 _22572_ (.A(_14812_),
    .B(_14816_),
    .Y(_15248_));
 sg13g2_a221oi_1 _22573_ (.B2(_15248_),
    .C1(_15247_),
    .B1(_15246_),
    .A1(\u_inv.d_next[147] ),
    .Y(_15249_),
    .A2(\u_inv.d_reg[147] ));
 sg13g2_nor2_1 _22574_ (.A(_15243_),
    .B(_15249_),
    .Y(_15250_));
 sg13g2_a21oi_1 _22575_ (.A1(\u_inv.d_next[149] ),
    .A2(\u_inv.d_reg[149] ),
    .Y(_15251_),
    .B1(_14805_));
 sg13g2_nor2_1 _22576_ (.A(_14803_),
    .B(_15251_),
    .Y(_15252_));
 sg13g2_o21ai_1 _22577_ (.B1(_14798_),
    .Y(_15253_),
    .A1(_14803_),
    .A2(_15251_));
 sg13g2_and2_1 _22578_ (.A(_14797_),
    .B(_14800_),
    .X(_15254_));
 sg13g2_a221oi_1 _22579_ (.B2(_15254_),
    .C1(_15250_),
    .B1(_15253_),
    .A1(\u_inv.d_next[151] ),
    .Y(_15255_),
    .A2(\u_inv.d_reg[151] ));
 sg13g2_nor2_1 _22580_ (.A(_14821_),
    .B(_14823_),
    .Y(_15256_));
 sg13g2_nand2_1 _22581_ (.Y(_15257_),
    .A(_15248_),
    .B(_15256_));
 sg13g2_nor2_1 _22582_ (.A(_15243_),
    .B(_15257_),
    .Y(_15258_));
 sg13g2_inv_1 _22583_ (.Y(_15259_),
    .A(_15258_));
 sg13g2_nor2b_1 _22584_ (.A(_15241_),
    .B_N(_15258_),
    .Y(_15260_));
 sg13g2_nor2_1 _22585_ (.A(net4430),
    .B(_14840_),
    .Y(_15261_));
 sg13g2_nor4_1 _22586_ (.A(_14831_),
    .B(_14834_),
    .C(_14838_),
    .D(net4429),
    .Y(_15262_));
 sg13g2_o21ai_1 _22587_ (.B1(_14847_),
    .Y(_15263_),
    .A1(\u_inv.d_next[138] ),
    .A2(net4777));
 sg13g2_nor2_1 _22588_ (.A(_14856_),
    .B(_14859_),
    .Y(_15264_));
 sg13g2_nor4_1 _22589_ (.A(_14846_),
    .B(_14849_),
    .C(_14856_),
    .D(_14859_),
    .Y(_15265_));
 sg13g2_nand2_1 _22590_ (.Y(_15266_),
    .A(_15262_),
    .B(_15265_));
 sg13g2_nor2_1 _22591_ (.A(_14873_),
    .B(_14875_),
    .Y(_15267_));
 sg13g2_nor4_1 _22592_ (.A(_14864_),
    .B(_14868_),
    .C(_14873_),
    .D(_14875_),
    .Y(_15268_));
 sg13g2_nand2_1 _22593_ (.Y(_15269_),
    .A(\u_inv.d_next[131] ),
    .B(\u_inv.d_reg[131] ));
 sg13g2_and2_1 _22594_ (.A(\u_inv.d_next[129] ),
    .B(net4779),
    .X(_15270_));
 sg13g2_a221oi_1 _22595_ (.B2(_14891_),
    .C1(_15270_),
    .B1(_14890_),
    .A1(net4802),
    .Y(_15271_),
    .A2(net4778));
 sg13g2_o21ai_1 _22596_ (.B1(_14882_),
    .Y(_15272_),
    .A1(\u_inv.d_next[130] ),
    .A2(net4778));
 sg13g2_o21ai_1 _22597_ (.B1(_15269_),
    .Y(_15273_),
    .A1(_15271_),
    .A2(_15272_));
 sg13g2_o21ai_1 _22598_ (.B1(_14871_),
    .Y(_15274_),
    .A1(_14870_),
    .A2(_14874_));
 sg13g2_a21o_1 _22599_ (.A2(_15274_),
    .A1(_14867_),
    .B1(_14866_),
    .X(_15275_));
 sg13g2_and2_1 _22600_ (.A(\u_inv.d_next[135] ),
    .B(\u_inv.d_reg[135] ),
    .X(_15276_));
 sg13g2_a221oi_1 _22601_ (.B2(_14865_),
    .C1(_15276_),
    .B1(_15275_),
    .A1(_15268_),
    .Y(_15277_),
    .A2(_15273_));
 sg13g2_nand2_1 _22602_ (.Y(_15278_),
    .A(\u_inv.d_next[139] ),
    .B(\u_inv.d_reg[139] ));
 sg13g2_a221oi_1 _22603_ (.B2(_14857_),
    .C1(_14854_),
    .B1(_14853_),
    .A1(\u_inv.d_next[138] ),
    .Y(_15279_),
    .A2(net4777));
 sg13g2_o21ai_1 _22604_ (.B1(_15278_),
    .Y(_15280_),
    .A1(_15263_),
    .A2(_15279_));
 sg13g2_a22oi_1 _22605_ (.Y(_15281_),
    .B1(\u_inv.d_reg[140] ),
    .B2(\u_inv.d_next[140] ),
    .A2(\u_inv.d_reg[141] ),
    .A1(\u_inv.d_next[141] ));
 sg13g2_nor2_1 _22606_ (.A(_14837_),
    .B(_15281_),
    .Y(_15282_));
 sg13g2_or3_1 _22607_ (.A(_14834_),
    .B(_14837_),
    .C(_15281_),
    .X(_15283_));
 sg13g2_a21oi_1 _22608_ (.A1(_14833_),
    .A2(_15283_),
    .Y(_15284_),
    .B1(_14831_));
 sg13g2_a221oi_1 _22609_ (.B2(_15280_),
    .C1(_15284_),
    .B1(_15262_),
    .A1(\u_inv.d_next[143] ),
    .Y(_15285_),
    .A2(\u_inv.d_reg[143] ));
 sg13g2_o21ai_1 _22610_ (.B1(_15285_),
    .Y(_15286_),
    .A1(_15266_),
    .A2(_15277_));
 sg13g2_and2_1 _22611_ (.A(\u_inv.d_next[153] ),
    .B(\u_inv.d_reg[153] ),
    .X(_15287_));
 sg13g2_a21oi_1 _22612_ (.A1(_14790_),
    .A2(_14791_),
    .Y(_15288_),
    .B1(_15287_));
 sg13g2_inv_1 _22613_ (.Y(_15289_),
    .A(_15288_));
 sg13g2_nor2_1 _22614_ (.A(_14784_),
    .B(_14785_),
    .Y(_15290_));
 sg13g2_a221oi_1 _22615_ (.B2(_15289_),
    .C1(_15290_),
    .B1(_15240_),
    .A1(\u_inv.d_next[155] ),
    .Y(_15291_),
    .A2(\u_inv.d_reg[155] ));
 sg13g2_a21oi_1 _22616_ (.A1(_10597_),
    .A2(_10913_),
    .Y(_15292_),
    .B1(_14771_));
 sg13g2_nand2_1 _22617_ (.Y(_15293_),
    .A(\u_inv.d_next[157] ),
    .B(\u_inv.d_reg[157] ));
 sg13g2_o21ai_1 _22618_ (.B1(_15293_),
    .Y(_15294_),
    .A1(_14775_),
    .A2(_14778_));
 sg13g2_a221oi_1 _22619_ (.B2(_15294_),
    .C1(_15292_),
    .B1(_15236_),
    .A1(\u_inv.d_next[159] ),
    .Y(_15295_),
    .A2(\u_inv.d_reg[159] ));
 sg13g2_o21ai_1 _22620_ (.B1(_15295_),
    .Y(_15296_),
    .A1(_15238_),
    .A2(_15291_));
 sg13g2_a21oi_1 _22621_ (.A1(_15260_),
    .A2(_15286_),
    .Y(_15297_),
    .B1(_15296_));
 sg13g2_o21ai_1 _22622_ (.B1(_15297_),
    .Y(_15298_),
    .A1(_15241_),
    .A2(_15255_));
 sg13g2_a21oi_1 _22623_ (.A1(_15235_),
    .A2(_15298_),
    .Y(_15299_),
    .B1(_15231_));
 sg13g2_or2_1 _22624_ (.X(_15300_),
    .B(_14674_),
    .A(_14673_));
 sg13g2_o21ai_1 _22625_ (.B1(_15300_),
    .Y(_15301_),
    .A1(_10591_),
    .A2(_10901_));
 sg13g2_nor2_1 _22626_ (.A(_14677_),
    .B(_14680_),
    .Y(_15302_));
 sg13g2_a221oi_1 _22627_ (.B2(_15301_),
    .C1(_15302_),
    .B1(_15191_),
    .A1(\u_inv.d_next[187] ),
    .Y(_15303_),
    .A2(\u_inv.d_reg[187] ));
 sg13g2_nor2_1 _22628_ (.A(_15190_),
    .B(_15303_),
    .Y(_15304_));
 sg13g2_a21oi_1 _22629_ (.A1(\u_inv.d_next[189] ),
    .A2(\u_inv.d_reg[189] ),
    .Y(_15305_),
    .B1(_14667_));
 sg13g2_a21oi_1 _22630_ (.A1(_10589_),
    .A2(_10899_),
    .Y(_15306_),
    .B1(_15305_));
 sg13g2_and3_1 _22631_ (.X(_15307_),
    .A(_14661_),
    .B(_14664_),
    .C(_15306_));
 sg13g2_o21ai_1 _22632_ (.B1(_14660_),
    .Y(_15308_),
    .A1(_14659_),
    .A2(_14662_));
 sg13g2_nand2_1 _22633_ (.Y(_15309_),
    .A(\u_inv.d_next[179] ),
    .B(\u_inv.d_reg[179] ));
 sg13g2_nand2_1 _22634_ (.Y(_15310_),
    .A(\u_inv.d_next[177] ),
    .B(\u_inv.d_reg[177] ));
 sg13g2_o21ai_1 _22635_ (.B1(_15310_),
    .Y(_15311_),
    .A1(_14706_),
    .A2(_14707_));
 sg13g2_nand2_1 _22636_ (.Y(_15312_),
    .A(_14701_),
    .B(_15311_));
 sg13g2_and2_1 _22637_ (.A(_14700_),
    .B(_15312_),
    .X(_15313_));
 sg13g2_o21ai_1 _22638_ (.B1(_15309_),
    .Y(_15314_),
    .A1(_14698_),
    .A2(_15313_));
 sg13g2_nor2_1 _22639_ (.A(_14687_),
    .B(_14688_),
    .Y(_15315_));
 sg13g2_a21oi_1 _22640_ (.A1(\u_inv.d_next[181] ),
    .A2(\u_inv.d_reg[181] ),
    .Y(_15316_),
    .B1(_15315_));
 sg13g2_or3_1 _22641_ (.A(_14693_),
    .B(_14695_),
    .C(_15316_),
    .X(_15317_));
 sg13g2_o21ai_1 _22642_ (.B1(_15317_),
    .Y(_15318_),
    .A1(_14692_),
    .A2(_14694_));
 sg13g2_a221oi_1 _22643_ (.B2(_15314_),
    .C1(_15318_),
    .B1(_15196_),
    .A1(\u_inv.d_next[183] ),
    .Y(_15319_),
    .A2(\u_inv.d_reg[183] ));
 sg13g2_inv_1 _22644_ (.Y(_15320_),
    .A(_15319_));
 sg13g2_nor2_1 _22645_ (.A(_15194_),
    .B(_15319_),
    .Y(_15321_));
 sg13g2_nor4_1 _22646_ (.A(_15304_),
    .B(_15307_),
    .C(_15308_),
    .D(_15321_),
    .Y(_15322_));
 sg13g2_and4_1 _22647_ (.A(_14699_),
    .B(_14701_),
    .C(_15196_),
    .D(_15197_),
    .X(_15323_));
 sg13g2_nor3_1 _22648_ (.A(_15199_),
    .B(_15220_),
    .C(_15234_),
    .Y(_15324_));
 sg13g2_o21ai_1 _22649_ (.B1(_15322_),
    .Y(_15325_),
    .A1(_15199_),
    .A2(_15299_));
 sg13g2_nor2_1 _22650_ (.A(_14309_),
    .B(_14313_),
    .Y(_15326_));
 sg13g2_nor4_1 _22651_ (.A(_14304_),
    .B(_14306_),
    .C(_14309_),
    .D(_14313_),
    .Y(_15327_));
 sg13g2_nor2_1 _22652_ (.A(_14318_),
    .B(_14321_),
    .Y(_15328_));
 sg13g2_nand2_1 _22653_ (.Y(_15329_),
    .A(_14317_),
    .B(_14320_));
 sg13g2_nor2_1 _22654_ (.A(_14323_),
    .B(_14325_),
    .Y(_15330_));
 sg13g2_inv_1 _22655_ (.Y(_15331_),
    .A(_15330_));
 sg13g2_nand2_1 _22656_ (.Y(_15332_),
    .A(_14334_),
    .B(_14336_));
 sg13g2_nor3_1 _22657_ (.A(_14330_),
    .B(_14332_),
    .C(_15332_),
    .Y(_15333_));
 sg13g2_nor4_1 _22658_ (.A(_14342_),
    .B(_14345_),
    .C(_14350_),
    .D(_14354_),
    .Y(_15334_));
 sg13g2_and2_1 _22659_ (.A(_15333_),
    .B(_15334_),
    .X(_15335_));
 sg13g2_nand4_1 _22660_ (.B(_15328_),
    .C(_15330_),
    .A(_15327_),
    .Y(_15336_),
    .D(_15335_));
 sg13g2_and2_1 _22661_ (.A(_14376_),
    .B(_14378_),
    .X(_15337_));
 sg13g2_inv_1 _22662_ (.Y(_15338_),
    .A(_15337_));
 sg13g2_nand3_1 _22663_ (.B(_14374_),
    .C(_15337_),
    .A(_14371_),
    .Y(_15339_));
 sg13g2_nor2_1 _22664_ (.A(_14364_),
    .B(_14366_),
    .Y(_15340_));
 sg13g2_nand2_1 _22665_ (.Y(_15341_),
    .A(_14359_),
    .B(_14361_));
 sg13g2_or4_1 _22666_ (.A(_14364_),
    .B(_14366_),
    .C(_15339_),
    .D(_15341_),
    .X(_15342_));
 sg13g2_nor2b_1 _22667_ (.A(_14405_),
    .B_N(_14403_),
    .Y(_15343_));
 sg13g2_nand2b_1 _22668_ (.Y(_15344_),
    .B(_14403_),
    .A_N(_14405_));
 sg13g2_nor2_1 _22669_ (.A(_14389_),
    .B(_14391_),
    .Y(_15345_));
 sg13g2_nor4_1 _22670_ (.A(_14382_),
    .B(_14386_),
    .C(_14389_),
    .D(_14391_),
    .Y(_15346_));
 sg13g2_and2_1 _22671_ (.A(_14397_),
    .B(_14399_),
    .X(_15347_));
 sg13g2_nand2_1 _22672_ (.Y(_15348_),
    .A(_14397_),
    .B(_14399_));
 sg13g2_nand3_1 _22673_ (.B(_15346_),
    .C(_15347_),
    .A(_15343_),
    .Y(_15349_));
 sg13g2_inv_1 _22674_ (.Y(_15350_),
    .A(_15349_));
 sg13g2_nand2b_2 _22675_ (.Y(_15351_),
    .B(_15350_),
    .A_N(_15342_));
 sg13g2_nor2_1 _22676_ (.A(_15336_),
    .B(_15351_),
    .Y(_15352_));
 sg13g2_nor2_1 _22677_ (.A(_14484_),
    .B(_14487_),
    .Y(_15353_));
 sg13g2_or4_1 _22678_ (.A(_14477_),
    .B(_14480_),
    .C(_14484_),
    .D(_14487_),
    .X(_15354_));
 sg13g2_nor2_1 _22679_ (.A(_14490_),
    .B(_14493_),
    .Y(_15355_));
 sg13g2_nor3_1 _22680_ (.A(_14497_),
    .B(_14498_),
    .C(_14500_),
    .Y(_15356_));
 sg13g2_nand3_1 _22681_ (.B(_14494_),
    .C(_15356_),
    .A(_14491_),
    .Y(_15357_));
 sg13g2_inv_1 _22682_ (.Y(_15358_),
    .A(_15357_));
 sg13g2_nor2_1 _22683_ (.A(_15354_),
    .B(_15357_),
    .Y(_15359_));
 sg13g2_nand2_1 _22684_ (.Y(_15360_),
    .A(_14512_),
    .B(_14514_));
 sg13g2_nor3_1 _22685_ (.A(_14506_),
    .B(_14509_),
    .C(_15360_),
    .Y(_15361_));
 sg13g2_nand2_1 _22686_ (.Y(_15362_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_and2_1 _22687_ (.A(\u_inv.d_next[65] ),
    .B(\u_inv.d_reg[65] ),
    .X(_15363_));
 sg13g2_nor2_1 _22688_ (.A(_14525_),
    .B(_14528_),
    .Y(_15364_));
 sg13g2_nor2_1 _22689_ (.A(_15363_),
    .B(_15364_),
    .Y(_15365_));
 sg13g2_a221oi_1 _22690_ (.B2(_14527_),
    .C1(_15363_),
    .B1(_14526_),
    .A1(\u_inv.d_next[66] ),
    .Y(_15366_),
    .A2(\u_inv.d_reg[66] ));
 sg13g2_or2_1 _22691_ (.X(_15367_),
    .B(_14519_),
    .A(_14517_));
 sg13g2_o21ai_1 _22692_ (.B1(_15362_),
    .Y(_15368_),
    .A1(_15366_),
    .A2(_15367_));
 sg13g2_a22oi_1 _22693_ (.Y(_15369_),
    .B1(\u_inv.d_reg[68] ),
    .B2(\u_inv.d_next[68] ),
    .A2(\u_inv.d_reg[69] ),
    .A1(net4803));
 sg13g2_nor2_1 _22694_ (.A(_14511_),
    .B(_15369_),
    .Y(_15370_));
 sg13g2_o21ai_1 _22695_ (.B1(_14507_),
    .Y(_15371_),
    .A1(_14511_),
    .A2(_15369_));
 sg13g2_nor2_1 _22696_ (.A(_14506_),
    .B(_14508_),
    .Y(_15372_));
 sg13g2_and2_1 _22697_ (.A(\u_inv.d_next[71] ),
    .B(\u_inv.d_reg[71] ),
    .X(_15373_));
 sg13g2_a21o_1 _22698_ (.A2(_15372_),
    .A1(_15371_),
    .B1(_15373_),
    .X(_15374_));
 sg13g2_a21o_2 _22699_ (.A2(_15368_),
    .A1(_15361_),
    .B1(_15374_),
    .X(_15375_));
 sg13g2_a22oi_1 _22700_ (.Y(_15376_),
    .B1(net4782),
    .B2(\u_inv.d_next[76] ),
    .A2(net4781),
    .A1(\u_inv.d_next[77] ));
 sg13g2_nor2_1 _22701_ (.A(_14482_),
    .B(_15376_),
    .Y(_15377_));
 sg13g2_o21ai_1 _22702_ (.B1(_14479_),
    .Y(_15378_),
    .A1(_14482_),
    .A2(_15376_));
 sg13g2_nor2_1 _22703_ (.A(_14477_),
    .B(_14478_),
    .Y(_15379_));
 sg13g2_a22oi_1 _22704_ (.Y(_15380_),
    .B1(_15378_),
    .B2(_15379_),
    .A2(\u_inv.d_reg[79] ),
    .A1(\u_inv.d_next[79] ));
 sg13g2_a22oi_1 _22705_ (.Y(_15381_),
    .B1(net4783),
    .B2(\u_inv.d_next[72] ),
    .A2(\u_inv.d_reg[73] ),
    .A1(\u_inv.d_next[73] ));
 sg13g2_nor2_1 _22706_ (.A(_14497_),
    .B(_15381_),
    .Y(_15382_));
 sg13g2_o21ai_1 _22707_ (.B1(_14492_),
    .Y(_15383_),
    .A1(_14497_),
    .A2(_15381_));
 sg13g2_a22oi_1 _22708_ (.Y(_15384_),
    .B1(_15355_),
    .B2(_15383_),
    .A2(\u_inv.d_reg[75] ),
    .A1(\u_inv.d_next[75] ));
 sg13g2_inv_1 _22709_ (.Y(_15385_),
    .A(_15384_));
 sg13g2_o21ai_1 _22710_ (.B1(_15380_),
    .Y(_15386_),
    .A1(_15354_),
    .A2(_15384_));
 sg13g2_a21oi_1 _22711_ (.A1(_15359_),
    .A2(_15375_),
    .Y(_15387_),
    .B1(_15386_));
 sg13g2_nand2_1 _22712_ (.Y(_15388_),
    .A(_14452_),
    .B(_14454_));
 sg13g2_or3_1 _22713_ (.A(_14446_),
    .B(_14449_),
    .C(_15388_),
    .X(_15389_));
 sg13g2_nor2_1 _22714_ (.A(_14459_),
    .B(_14462_),
    .Y(_15390_));
 sg13g2_nand2b_1 _22715_ (.Y(_15391_),
    .B(_14461_),
    .A_N(_14459_));
 sg13g2_nor2_1 _22716_ (.A(_15389_),
    .B(_15391_),
    .Y(_15392_));
 sg13g2_nand2_1 _22717_ (.Y(_15393_),
    .A(_14413_),
    .B(_14416_));
 sg13g2_nor3_1 _22718_ (.A(_14421_),
    .B(_14424_),
    .C(_15393_),
    .Y(_15394_));
 sg13g2_nor2_1 _22719_ (.A(_14437_),
    .B(_14441_),
    .Y(_15395_));
 sg13g2_nor4_1 _22720_ (.A(_14429_),
    .B(_14432_),
    .C(_14437_),
    .D(_14441_),
    .Y(_15396_));
 sg13g2_and2_1 _22721_ (.A(_15394_),
    .B(_15396_),
    .X(_15397_));
 sg13g2_nor2_2 _22722_ (.A(_14466_),
    .B(_14469_),
    .Y(_15398_));
 sg13g2_nand3_1 _22723_ (.B(_15397_),
    .C(_15398_),
    .A(_15392_),
    .Y(_15399_));
 sg13g2_nand2_1 _22724_ (.Y(_15400_),
    .A(\u_inv.d_next[91] ),
    .B(\u_inv.d_reg[91] ));
 sg13g2_and2_1 _22725_ (.A(\u_inv.d_next[89] ),
    .B(\u_inv.d_reg[89] ),
    .X(_15401_));
 sg13g2_a221oi_1 _22726_ (.B2(_14439_),
    .C1(_15401_),
    .B1(_14438_),
    .A1(\u_inv.d_next[90] ),
    .Y(_15402_),
    .A2(\u_inv.d_reg[90] ));
 sg13g2_o21ai_1 _22727_ (.B1(_14430_),
    .Y(_15403_),
    .A1(\u_inv.d_next[90] ),
    .A2(\u_inv.d_reg[90] ));
 sg13g2_o21ai_1 _22728_ (.B1(_15400_),
    .Y(_15404_),
    .A1(_15402_),
    .A2(_15403_));
 sg13g2_and2_1 _22729_ (.A(\u_inv.d_next[93] ),
    .B(\u_inv.d_reg[93] ),
    .X(_15405_));
 sg13g2_a21oi_1 _22730_ (.A1(_14422_),
    .A2(_14423_),
    .Y(_15406_),
    .B1(_15405_));
 sg13g2_or2_1 _22731_ (.X(_15407_),
    .B(_14415_),
    .A(_14412_));
 sg13g2_o21ai_1 _22732_ (.B1(_15407_),
    .Y(_15408_),
    .A1(_15393_),
    .A2(_15406_));
 sg13g2_a21o_1 _22733_ (.A2(\u_inv.d_reg[95] ),
    .A1(\u_inv.d_next[95] ),
    .B1(_15408_),
    .X(_15409_));
 sg13g2_or2_1 _22734_ (.X(_15410_),
    .B(_14467_),
    .A(_14466_));
 sg13g2_nand2_1 _22735_ (.Y(_15411_),
    .A(\u_inv.d_next[81] ),
    .B(\u_inv.d_reg[81] ));
 sg13g2_o21ai_1 _22736_ (.B1(_15411_),
    .Y(_15412_),
    .A1(_14466_),
    .A2(_14467_));
 sg13g2_nor2_1 _22737_ (.A(_14459_),
    .B(_14460_),
    .Y(_15413_));
 sg13g2_a221oi_1 _22738_ (.B2(_15412_),
    .C1(_15413_),
    .B1(_15390_),
    .A1(\u_inv.d_next[83] ),
    .Y(_15414_),
    .A2(\u_inv.d_reg[83] ));
 sg13g2_a22oi_1 _22739_ (.Y(_15415_),
    .B1(\u_inv.d_reg[84] ),
    .B2(\u_inv.d_next[84] ),
    .A2(\u_inv.d_reg[85] ),
    .A1(\u_inv.d_next[85] ));
 sg13g2_or2_1 _22740_ (.X(_15416_),
    .B(_15415_),
    .A(_14451_));
 sg13g2_o21ai_1 _22741_ (.B1(_14447_),
    .Y(_15417_),
    .A1(_14451_),
    .A2(_15415_));
 sg13g2_nor2_1 _22742_ (.A(_14446_),
    .B(_14448_),
    .Y(_15418_));
 sg13g2_a22oi_1 _22743_ (.Y(_15419_),
    .B1(_15417_),
    .B2(_15418_),
    .A2(\u_inv.d_reg[87] ),
    .A1(\u_inv.d_next[87] ));
 sg13g2_o21ai_1 _22744_ (.B1(_15419_),
    .Y(_15420_),
    .A1(_15389_),
    .A2(_15414_));
 sg13g2_a221oi_1 _22745_ (.B2(_15397_),
    .C1(_15409_),
    .B1(_15420_),
    .A1(_15394_),
    .Y(_15421_),
    .A2(_15404_));
 sg13g2_nor4_1 _22746_ (.A(_14466_),
    .B(_14469_),
    .C(_15389_),
    .D(_15391_),
    .Y(_15422_));
 sg13g2_o21ai_1 _22747_ (.B1(_15421_),
    .Y(_15423_),
    .A1(_15387_),
    .A2(_15399_));
 sg13g2_and2_1 _22748_ (.A(_15352_),
    .B(_15423_),
    .X(_15424_));
 sg13g2_nand2_1 _22749_ (.Y(_15425_),
    .A(\u_inv.d_next[115] ),
    .B(\u_inv.d_reg[115] ));
 sg13g2_nor2_1 _22750_ (.A(_14350_),
    .B(_14352_),
    .Y(_15426_));
 sg13g2_a21oi_1 _22751_ (.A1(\u_inv.d_next[113] ),
    .A2(\u_inv.d_reg[113] ),
    .Y(_15427_),
    .B1(_15426_));
 sg13g2_a221oi_1 _22752_ (.B2(\u_inv.d_next[113] ),
    .C1(_15426_),
    .B1(\u_inv.d_reg[113] ),
    .A1(\u_inv.d_next[114] ),
    .Y(_15428_),
    .A2(\u_inv.d_reg[114] ));
 sg13g2_o21ai_1 _22753_ (.B1(_14343_),
    .Y(_15429_),
    .A1(\u_inv.d_next[114] ),
    .A2(\u_inv.d_reg[114] ));
 sg13g2_o21ai_1 _22754_ (.B1(_15425_),
    .Y(_15430_),
    .A1(_15428_),
    .A2(_15429_));
 sg13g2_nor2_1 _22755_ (.A(_14330_),
    .B(_14331_),
    .Y(_15431_));
 sg13g2_inv_1 _22756_ (.Y(_15432_),
    .A(_15431_));
 sg13g2_a21oi_1 _22757_ (.A1(\u_inv.d_next[117] ),
    .A2(\u_inv.d_reg[117] ),
    .Y(_15433_),
    .B1(_15431_));
 sg13g2_o21ai_1 _22758_ (.B1(_14335_),
    .Y(_15434_),
    .A1(\u_inv.d_next[119] ),
    .A2(\u_inv.d_reg[119] ));
 sg13g2_o21ai_1 _22759_ (.B1(_15434_),
    .Y(_15435_),
    .A1(_15332_),
    .A2(_15433_));
 sg13g2_a221oi_1 _22760_ (.B2(_15430_),
    .C1(_15435_),
    .B1(_15333_),
    .A1(\u_inv.d_next[119] ),
    .Y(_15436_),
    .A2(\u_inv.d_reg[119] ));
 sg13g2_inv_1 _22761_ (.Y(_15437_),
    .A(_15436_));
 sg13g2_and4_1 _22762_ (.A(_15327_),
    .B(_15328_),
    .C(_15330_),
    .D(_15437_),
    .X(_15438_));
 sg13g2_nor2_1 _22763_ (.A(_14323_),
    .B(_14324_),
    .Y(_15439_));
 sg13g2_a21oi_1 _22764_ (.A1(\u_inv.d_next[121] ),
    .A2(\u_inv.d_reg[121] ),
    .Y(_15440_),
    .B1(_15439_));
 sg13g2_o21ai_1 _22765_ (.B1(_14316_),
    .Y(_15441_),
    .A1(\u_inv.d_next[123] ),
    .A2(\u_inv.d_reg[123] ));
 sg13g2_o21ai_1 _22766_ (.B1(_14319_),
    .Y(_15442_),
    .A1(_15329_),
    .A2(_15440_));
 sg13g2_nand2b_2 _22767_ (.Y(_15443_),
    .B(_15441_),
    .A_N(_15442_));
 sg13g2_a21oi_1 _22768_ (.A1(_10601_),
    .A2(_10920_),
    .Y(_15444_),
    .B1(_14305_));
 sg13g2_a21oi_1 _22769_ (.A1(\u_inv.d_next[127] ),
    .A2(\u_inv.d_reg[127] ),
    .Y(_15445_),
    .B1(_15444_));
 sg13g2_nand2_1 _22770_ (.Y(_15446_),
    .A(_14308_),
    .B(_14311_));
 sg13g2_o21ai_1 _22771_ (.B1(_15446_),
    .Y(_15447_),
    .A1(\u_inv.d_next[125] ),
    .A2(\u_inv.d_reg[125] ));
 sg13g2_nor3_1 _22772_ (.A(_14304_),
    .B(_14306_),
    .C(_15447_),
    .Y(_15448_));
 sg13g2_a21oi_1 _22773_ (.A1(_15327_),
    .A2(_15443_),
    .Y(_15449_),
    .B1(_15448_));
 sg13g2_nand2_1 _22774_ (.Y(_15450_),
    .A(_15445_),
    .B(_15449_));
 sg13g2_and2_1 _22775_ (.A(\u_inv.d_next[97] ),
    .B(\u_inv.d_reg[97] ),
    .X(_15451_));
 sg13g2_a21oi_1 _22776_ (.A1(_14403_),
    .A2(_14404_),
    .Y(_15452_),
    .B1(_15451_));
 sg13g2_a22oi_1 _22777_ (.Y(_15453_),
    .B1(\u_inv.d_reg[100] ),
    .B2(\u_inv.d_next[100] ),
    .A2(\u_inv.d_reg[101] ),
    .A1(\u_inv.d_next[101] ));
 sg13g2_nor2_1 _22778_ (.A(_14388_),
    .B(_15453_),
    .Y(_15454_));
 sg13g2_or3_1 _22779_ (.A(_14386_),
    .B(_14388_),
    .C(_15453_),
    .X(_15455_));
 sg13g2_a21oi_1 _22780_ (.A1(_14384_),
    .A2(_15455_),
    .Y(_15456_),
    .B1(_14382_));
 sg13g2_a21oi_1 _22781_ (.A1(\u_inv.d_next[103] ),
    .A2(\u_inv.d_reg[103] ),
    .Y(_15457_),
    .B1(_15456_));
 sg13g2_nor2_1 _22782_ (.A(_14396_),
    .B(_14398_),
    .Y(_15458_));
 sg13g2_a21o_1 _22783_ (.A2(\u_inv.d_reg[99] ),
    .A1(\u_inv.d_next[99] ),
    .B1(_15458_),
    .X(_15459_));
 sg13g2_nor2_1 _22784_ (.A(_15348_),
    .B(_15452_),
    .Y(_15460_));
 sg13g2_o21ai_1 _22785_ (.B1(_15346_),
    .Y(_15461_),
    .A1(_15459_),
    .A2(_15460_));
 sg13g2_nand2_1 _22786_ (.Y(_15462_),
    .A(_15457_),
    .B(_15461_));
 sg13g2_a21oi_1 _22787_ (.A1(_15457_),
    .A2(_15461_),
    .Y(_15463_),
    .B1(_15342_));
 sg13g2_a21oi_1 _22788_ (.A1(\u_inv.d_next[111] ),
    .A2(\u_inv.d_reg[111] ),
    .Y(_15464_),
    .B1(_14360_));
 sg13g2_a21oi_1 _22789_ (.A1(_10604_),
    .A2(_10922_),
    .Y(_15465_),
    .B1(_15464_));
 sg13g2_and2_1 _22790_ (.A(\u_inv.d_next[107] ),
    .B(\u_inv.d_reg[107] ),
    .X(_15466_));
 sg13g2_and2_1 _22791_ (.A(\u_inv.d_next[105] ),
    .B(\u_inv.d_reg[105] ),
    .X(_15467_));
 sg13g2_a21oi_1 _22792_ (.A1(_14376_),
    .A2(_14377_),
    .Y(_15468_),
    .B1(_15467_));
 sg13g2_o21ai_1 _22793_ (.B1(_14371_),
    .Y(_15469_),
    .A1(\u_inv.d_next[106] ),
    .A2(\u_inv.d_reg[106] ));
 sg13g2_a21oi_1 _22794_ (.A1(_14373_),
    .A2(_15468_),
    .Y(_15470_),
    .B1(_15469_));
 sg13g2_nor2_1 _22795_ (.A(_15466_),
    .B(_15470_),
    .Y(_15471_));
 sg13g2_o21ai_1 _22796_ (.B1(_15340_),
    .Y(_15472_),
    .A1(_15466_),
    .A2(_15470_));
 sg13g2_nor2_1 _22797_ (.A(_14364_),
    .B(_14365_),
    .Y(_15473_));
 sg13g2_a21oi_1 _22798_ (.A1(\u_inv.d_next[109] ),
    .A2(\u_inv.d_reg[109] ),
    .Y(_15474_),
    .B1(_15473_));
 sg13g2_a21oi_1 _22799_ (.A1(_15472_),
    .A2(_15474_),
    .Y(_15475_),
    .B1(_15341_));
 sg13g2_nor3_1 _22800_ (.A(_15463_),
    .B(_15465_),
    .C(_15475_),
    .Y(_15476_));
 sg13g2_nor2_1 _22801_ (.A(_15336_),
    .B(_15476_),
    .Y(_15477_));
 sg13g2_or4_1 _22802_ (.A(_15424_),
    .B(_15438_),
    .C(_15450_),
    .D(_15477_),
    .X(_15478_));
 sg13g2_nor2_1 _22803_ (.A(_14213_),
    .B(_14216_),
    .Y(_15479_));
 sg13g2_nor4_1 _22804_ (.A(_14204_),
    .B(_14208_),
    .C(_14213_),
    .D(_14216_),
    .Y(_15480_));
 sg13g2_nand2_1 _22805_ (.Y(_15481_),
    .A(\u_inv.d_next[35] ),
    .B(\u_inv.d_reg[35] ));
 sg13g2_and2_1 _22806_ (.A(\u_inv.d_next[33] ),
    .B(\u_inv.d_reg[33] ),
    .X(_15482_));
 sg13g2_a221oi_1 _22807_ (.B2(_14230_),
    .C1(_15482_),
    .B1(_14229_),
    .A1(\u_inv.d_next[34] ),
    .Y(_15483_),
    .A2(\u_inv.d_reg[34] ));
 sg13g2_or2_1 _22808_ (.X(_15484_),
    .B(_14223_),
    .A(_14221_));
 sg13g2_o21ai_1 _22809_ (.B1(_15481_),
    .Y(_15485_),
    .A1(_15483_),
    .A2(_15484_));
 sg13g2_o21ai_1 _22810_ (.B1(_14211_),
    .Y(_15486_),
    .A1(_14210_),
    .A2(_14214_));
 sg13g2_a21o_1 _22811_ (.A2(_15486_),
    .A1(_14207_),
    .B1(_14206_),
    .X(_15487_));
 sg13g2_and2_1 _22812_ (.A(\u_inv.d_next[39] ),
    .B(\u_inv.d_reg[39] ),
    .X(_15488_));
 sg13g2_a221oi_1 _22813_ (.B2(_14205_),
    .C1(_15488_),
    .B1(_15487_),
    .A1(_15480_),
    .Y(_15489_),
    .A2(_15485_));
 sg13g2_nor2_1 _22814_ (.A(_14181_),
    .B(_14183_),
    .Y(_15490_));
 sg13g2_and3_1 _22815_ (.X(_15491_),
    .A(_14175_),
    .B(_14177_),
    .C(_15490_));
 sg13g2_nor2_1 _22816_ (.A(_14188_),
    .B(_14191_),
    .Y(_15492_));
 sg13g2_nor2_1 _22817_ (.A(_14196_),
    .B(_14199_),
    .Y(_15493_));
 sg13g2_and2_1 _22818_ (.A(_15492_),
    .B(_15493_),
    .X(_15494_));
 sg13g2_nand2_1 _22819_ (.Y(_15495_),
    .A(_15491_),
    .B(_15494_));
 sg13g2_nand2_1 _22820_ (.Y(_15496_),
    .A(\u_inv.d_next[43] ),
    .B(\u_inv.d_reg[43] ));
 sg13g2_a221oi_1 _22821_ (.B2(_14197_),
    .C1(_14195_),
    .B1(_14194_),
    .A1(\u_inv.d_next[42] ),
    .Y(_15497_),
    .A2(net4786));
 sg13g2_o21ai_1 _22822_ (.B1(_14189_),
    .Y(_15498_),
    .A1(\u_inv.d_next[42] ),
    .A2(net4786));
 sg13g2_o21ai_1 _22823_ (.B1(_15496_),
    .Y(_15499_),
    .A1(_15497_),
    .A2(_15498_));
 sg13g2_a22oi_1 _22824_ (.Y(_15500_),
    .B1(\u_inv.d_reg[44] ),
    .B2(\u_inv.d_next[44] ),
    .A2(\u_inv.d_reg[45] ),
    .A1(\u_inv.d_next[45] ));
 sg13g2_nor2_1 _22825_ (.A(_14180_),
    .B(_15500_),
    .Y(_15501_));
 sg13g2_o21ai_1 _22826_ (.B1(_14176_),
    .Y(_15502_),
    .A1(_14180_),
    .A2(_15500_));
 sg13g2_o21ai_1 _22827_ (.B1(_14175_),
    .Y(_15503_),
    .A1(\u_inv.d_next[46] ),
    .A2(\u_inv.d_reg[46] ));
 sg13g2_nor2b_1 _22828_ (.A(_15503_),
    .B_N(_15502_),
    .Y(_15504_));
 sg13g2_a221oi_1 _22829_ (.B2(_15499_),
    .C1(_15504_),
    .B1(_15491_),
    .A1(\u_inv.d_next[47] ),
    .Y(_15505_),
    .A2(\u_inv.d_reg[47] ));
 sg13g2_nand3_1 _22830_ (.B(_15492_),
    .C(_15493_),
    .A(_15491_),
    .Y(_15506_));
 sg13g2_o21ai_1 _22831_ (.B1(_15505_),
    .Y(_15507_),
    .A1(_15489_),
    .A2(_15495_));
 sg13g2_nor2_1 _22832_ (.A(_14157_),
    .B(_14160_),
    .Y(_15508_));
 sg13g2_nand3_1 _22833_ (.B(_14151_),
    .C(_15508_),
    .A(_14149_),
    .Y(_15509_));
 sg13g2_nor2_1 _22834_ (.A(_14163_),
    .B(_14165_),
    .Y(_15510_));
 sg13g2_and2_1 _22835_ (.A(_14169_),
    .B(_14171_),
    .X(_15511_));
 sg13g2_nand3b_1 _22836_ (.B(_15510_),
    .C(_15511_),
    .Y(_15512_),
    .A_N(_15509_));
 sg13g2_nor2_1 _22837_ (.A(_14123_),
    .B(_14125_),
    .Y(_15513_));
 sg13g2_nor2b_1 _22838_ (.A(_14127_),
    .B_N(_14129_),
    .Y(_15514_));
 sg13g2_and2_1 _22839_ (.A(_15513_),
    .B(_15514_),
    .X(_15515_));
 sg13g2_nor2_1 _22840_ (.A(_14134_),
    .B(_14138_),
    .Y(_15516_));
 sg13g2_and2_1 _22841_ (.A(_14140_),
    .B(_14142_),
    .X(_15517_));
 sg13g2_nand2_1 _22842_ (.Y(_15518_),
    .A(\u_inv.d_next[59] ),
    .B(\u_inv.d_reg[59] ));
 sg13g2_and2_1 _22843_ (.A(_14140_),
    .B(_14141_),
    .X(_15519_));
 sg13g2_and2_1 _22844_ (.A(\u_inv.d_next[57] ),
    .B(\u_inv.d_reg[57] ),
    .X(_15520_));
 sg13g2_a221oi_1 _22845_ (.B2(_14141_),
    .C1(_15520_),
    .B1(_14140_),
    .A1(net4804),
    .Y(_15521_),
    .A2(net4785));
 sg13g2_o21ai_1 _22846_ (.B1(_14135_),
    .Y(_15522_),
    .A1(\u_inv.d_next[58] ),
    .A2(net4785));
 sg13g2_o21ai_1 _22847_ (.B1(_15518_),
    .Y(_15523_),
    .A1(_15521_),
    .A2(_15522_));
 sg13g2_nand2_1 _22848_ (.Y(_15524_),
    .A(_15515_),
    .B(_15523_));
 sg13g2_nor2_1 _22849_ (.A(_14127_),
    .B(_14128_),
    .Y(_15525_));
 sg13g2_a21oi_1 _22850_ (.A1(\u_inv.d_next[61] ),
    .A2(\u_inv.d_reg[61] ),
    .Y(_15526_),
    .B1(_15525_));
 sg13g2_nand2b_1 _22851_ (.Y(_15527_),
    .B(_15513_),
    .A_N(_15526_));
 sg13g2_nor2_1 _22852_ (.A(_14122_),
    .B(_14124_),
    .Y(_15528_));
 sg13g2_a21oi_1 _22853_ (.A1(\u_inv.d_next[63] ),
    .A2(\u_inv.d_reg[63] ),
    .Y(_15529_),
    .B1(_15528_));
 sg13g2_nand3_1 _22854_ (.B(_15527_),
    .C(_15529_),
    .A(_15524_),
    .Y(_15530_));
 sg13g2_nand2_1 _22855_ (.Y(_15531_),
    .A(\u_inv.d_next[51] ),
    .B(\u_inv.d_reg[51] ));
 sg13g2_o21ai_1 _22856_ (.B1(_15531_),
    .Y(_15532_),
    .A1(_14163_),
    .A2(_14164_));
 sg13g2_nand2b_1 _22857_ (.Y(_15533_),
    .B(_14169_),
    .A_N(_14170_));
 sg13g2_o21ai_1 _22858_ (.B1(_15533_),
    .Y(_15534_),
    .A1(_10614_),
    .A2(_10941_));
 sg13g2_a21oi_1 _22859_ (.A1(_15510_),
    .A2(_15534_),
    .Y(_15535_),
    .B1(_15532_));
 sg13g2_o21ai_1 _22860_ (.B1(_14155_),
    .Y(_15536_),
    .A1(_14154_),
    .A2(_14158_));
 sg13g2_nand2_1 _22861_ (.Y(_15537_),
    .A(_14151_),
    .B(_15536_));
 sg13g2_a21o_1 _22862_ (.A2(_15537_),
    .A1(_14150_),
    .B1(_14148_),
    .X(_15538_));
 sg13g2_o21ai_1 _22863_ (.B1(_15538_),
    .Y(_15539_),
    .A1(_15509_),
    .A2(_15535_));
 sg13g2_a21oi_1 _22864_ (.A1(\u_inv.d_next[55] ),
    .A2(\u_inv.d_reg[55] ),
    .Y(_15540_),
    .B1(_15539_));
 sg13g2_nand3_1 _22865_ (.B(_15516_),
    .C(_15517_),
    .A(_15515_),
    .Y(_15541_));
 sg13g2_nor2_1 _22866_ (.A(_15512_),
    .B(_15541_),
    .Y(_15542_));
 sg13g2_a21oi_1 _22867_ (.A1(_15507_),
    .A2(_15542_),
    .Y(_15543_),
    .B1(_15530_));
 sg13g2_o21ai_1 _22868_ (.B1(_15543_),
    .Y(_15544_),
    .A1(_15540_),
    .A2(_15541_));
 sg13g2_nand2b_1 _22869_ (.Y(_15545_),
    .B(_14069_),
    .A_N(_14070_));
 sg13g2_nand2_1 _22870_ (.Y(_15546_),
    .A(\u_inv.d_next[17] ),
    .B(\u_inv.d_reg[17] ));
 sg13g2_and2_1 _22871_ (.A(_15545_),
    .B(_15546_),
    .X(_15547_));
 sg13g2_o21ai_1 _22872_ (.B1(_15546_),
    .Y(_15548_),
    .A1(_14068_),
    .A2(_14070_));
 sg13g2_and3_1 _22873_ (.X(_15549_),
    .A(\u_inv.d_next[18] ),
    .B(net4790),
    .C(_14063_));
 sg13g2_and2_1 _22874_ (.A(_14063_),
    .B(_14064_),
    .X(_15550_));
 sg13g2_a221oi_1 _22875_ (.B2(_15550_),
    .C1(_15549_),
    .B1(_15548_),
    .A1(\u_inv.d_next[19] ),
    .Y(_15551_),
    .A2(\u_inv.d_reg[19] ));
 sg13g2_inv_1 _22876_ (.Y(_15552_),
    .A(_15551_));
 sg13g2_nor2_1 _22877_ (.A(_14040_),
    .B(_14042_),
    .Y(_15553_));
 sg13g2_nand3_1 _22878_ (.B(_14037_),
    .C(_15553_),
    .A(_14035_),
    .Y(_15554_));
 sg13g2_inv_1 _22879_ (.Y(_15555_),
    .A(_15554_));
 sg13g2_or2_1 _22880_ (.X(_15556_),
    .B(_14058_),
    .A(_14056_));
 sg13g2_or3_1 _22881_ (.A(_14048_),
    .B(_14052_),
    .C(_15556_),
    .X(_15557_));
 sg13g2_nor2_1 _22882_ (.A(_15554_),
    .B(_15557_),
    .Y(_15558_));
 sg13g2_and2_1 _22883_ (.A(_14084_),
    .B(_14086_),
    .X(_15559_));
 sg13g2_nor2_1 _22884_ (.A(_14076_),
    .B(_14081_),
    .Y(_15560_));
 sg13g2_and2_1 _22885_ (.A(_15559_),
    .B(_15560_),
    .X(_15561_));
 sg13g2_nand2_1 _22886_ (.Y(_15562_),
    .A(_15559_),
    .B(_15560_));
 sg13g2_a22oi_1 _22887_ (.Y(_15563_),
    .B1(\u_inv.d_reg[20] ),
    .B2(\u_inv.d_next[20] ),
    .A2(\u_inv.d_reg[21] ),
    .A1(\u_inv.d_next[21] ));
 sg13g2_nor2_1 _22888_ (.A(_14083_),
    .B(_15563_),
    .Y(_15564_));
 sg13g2_o21ai_1 _22889_ (.B1(_14078_),
    .Y(_15565_),
    .A1(_14083_),
    .A2(_15563_));
 sg13g2_nor2_1 _22890_ (.A(_14076_),
    .B(_14079_),
    .Y(_15566_));
 sg13g2_a22oi_1 _22891_ (.Y(_15567_),
    .B1(_15565_),
    .B2(_15566_),
    .A2(\u_inv.d_reg[23] ),
    .A1(\u_inv.d_next[23] ));
 sg13g2_a21oi_1 _22892_ (.A1(_10618_),
    .A2(_10948_),
    .Y(_15568_),
    .B1(_14041_));
 sg13g2_a21oi_1 _22893_ (.A1(\u_inv.d_next[29] ),
    .A2(\u_inv.d_reg[29] ),
    .Y(_15569_),
    .B1(_15568_));
 sg13g2_o21ai_1 _22894_ (.B1(_14035_),
    .Y(_15570_),
    .A1(\u_inv.d_next[30] ),
    .A2(\u_inv.d_reg[30] ));
 sg13g2_a21oi_1 _22895_ (.A1(_14036_),
    .A2(_15569_),
    .Y(_15571_),
    .B1(_15570_));
 sg13g2_a21oi_1 _22896_ (.A1(\u_inv.d_next[31] ),
    .A2(\u_inv.d_reg[31] ),
    .Y(_15572_),
    .B1(_15571_));
 sg13g2_nand2_1 _22897_ (.Y(_15573_),
    .A(\u_inv.d_next[27] ),
    .B(\u_inv.d_reg[27] ));
 sg13g2_o21ai_1 _22898_ (.B1(_14055_),
    .Y(_15574_),
    .A1(_14054_),
    .A2(_14057_));
 sg13g2_a21oi_1 _22899_ (.A1(_14051_),
    .A2(_15574_),
    .Y(_15575_),
    .B1(_14049_));
 sg13g2_o21ai_1 _22900_ (.B1(_15573_),
    .Y(_15576_),
    .A1(_14048_),
    .A2(_15575_));
 sg13g2_o21ai_1 _22901_ (.B1(_15567_),
    .Y(_15577_),
    .A1(_15551_),
    .A2(_15562_));
 sg13g2_a22oi_1 _22902_ (.Y(_15578_),
    .B1(_15577_),
    .B2(_15558_),
    .A2(_15576_),
    .A1(_15555_));
 sg13g2_nand2_1 _22903_ (.Y(_15579_),
    .A(_15572_),
    .B(_15578_));
 sg13g2_and2_1 _22904_ (.A(\u_inv.d_next[3] ),
    .B(\u_inv.d_reg[3] ),
    .X(_15580_));
 sg13g2_and2_1 _22905_ (.A(\u_inv.d_next[0] ),
    .B(net4799),
    .X(_15581_));
 sg13g2_a21oi_1 _22906_ (.A1(_13996_),
    .A2(_15581_),
    .Y(_15582_),
    .B1(_13995_));
 sg13g2_o21ai_1 _22907_ (.B1(_13991_),
    .Y(_15583_),
    .A1(_13992_),
    .A2(_15582_));
 sg13g2_a21oi_1 _22908_ (.A1(_13988_),
    .A2(_15583_),
    .Y(_15584_),
    .B1(_15580_));
 sg13g2_nand2b_1 _22909_ (.Y(_15585_),
    .B(_14003_),
    .A_N(_15584_));
 sg13g2_nand2b_1 _22910_ (.Y(_15586_),
    .B(_14007_),
    .A_N(_15585_));
 sg13g2_and2_1 _22911_ (.A(_13977_),
    .B(_13978_),
    .X(_15587_));
 sg13g2_nand3_1 _22912_ (.B(_14003_),
    .C(_14007_),
    .A(_13982_),
    .Y(_15588_));
 sg13g2_or2_1 _22913_ (.X(_15589_),
    .B(_15588_),
    .A(_15587_));
 sg13g2_and2_1 _22914_ (.A(\u_inv.d_next[5] ),
    .B(\u_inv.d_reg[5] ),
    .X(_15590_));
 sg13g2_and2_1 _22915_ (.A(_14002_),
    .B(_14007_),
    .X(_15591_));
 sg13g2_nor2_1 _22916_ (.A(_15590_),
    .B(_15591_),
    .Y(_15592_));
 sg13g2_a221oi_1 _22917_ (.B2(_14007_),
    .C1(_15590_),
    .B1(_14002_),
    .A1(net4806),
    .Y(_15593_),
    .A2(net4795));
 sg13g2_nor3_1 _22918_ (.A(_13981_),
    .B(_15587_),
    .C(_15593_),
    .Y(_15594_));
 sg13g2_a21oi_1 _22919_ (.A1(\u_inv.d_next[7] ),
    .A2(net4794),
    .Y(_15595_),
    .B1(_15594_));
 sg13g2_o21ai_1 _22920_ (.B1(_15595_),
    .Y(_15596_),
    .A1(_15584_),
    .A2(_15589_));
 sg13g2_nand4_1 _22921_ (.B(_13961_),
    .C(_13964_),
    .A(_13959_),
    .Y(_15597_),
    .D(_13966_));
 sg13g2_or2_1 _22922_ (.X(_15598_),
    .B(_13974_),
    .A(_13971_));
 sg13g2_nand2_1 _22923_ (.Y(_15599_),
    .A(_14016_),
    .B(_14018_));
 sg13g2_nor3_1 _22924_ (.A(_15597_),
    .B(_15598_),
    .C(_15599_),
    .Y(_15600_));
 sg13g2_and2_1 _22925_ (.A(\u_inv.d_next[11] ),
    .B(net4792),
    .X(_15601_));
 sg13g2_and2_1 _22926_ (.A(\u_inv.d_next[9] ),
    .B(\u_inv.d_reg[9] ),
    .X(_15602_));
 sg13g2_a21oi_1 _22927_ (.A1(_14016_),
    .A2(_14017_),
    .Y(_15603_),
    .B1(_15602_));
 sg13g2_o21ai_1 _22928_ (.B1(_13973_),
    .Y(_15604_),
    .A1(_13974_),
    .A2(_15603_));
 sg13g2_a21oi_1 _22929_ (.A1(_13972_),
    .A2(_15604_),
    .Y(_15605_),
    .B1(_15601_));
 sg13g2_a21oi_1 _22930_ (.A1(\u_inv.d_next[13] ),
    .A2(\u_inv.d_reg[13] ),
    .Y(_15606_),
    .B1(_13965_));
 sg13g2_nor2_1 _22931_ (.A(_13963_),
    .B(_15606_),
    .Y(_15607_));
 sg13g2_o21ai_1 _22932_ (.B1(_13960_),
    .Y(_15608_),
    .A1(_13963_),
    .A2(_15606_));
 sg13g2_a21oi_1 _22933_ (.A1(_10620_),
    .A2(_10953_),
    .Y(_15609_),
    .B1(_13958_));
 sg13g2_a22oi_1 _22934_ (.Y(_15610_),
    .B1(_15608_),
    .B2(_15609_),
    .A2(\u_inv.d_reg[15] ),
    .A1(\u_inv.d_next[15] ));
 sg13g2_o21ai_1 _22935_ (.B1(_15610_),
    .Y(_15611_),
    .A1(_15597_),
    .A2(_15605_));
 sg13g2_a21o_2 _22936_ (.A2(_15600_),
    .A1(_15596_),
    .B1(_15611_),
    .X(_15612_));
 sg13g2_and2_1 _22937_ (.A(_14069_),
    .B(_14071_),
    .X(_15613_));
 sg13g2_nand2_1 _22938_ (.Y(_15614_),
    .A(_15612_),
    .B(_15613_));
 sg13g2_and4_1 _22939_ (.A(_15550_),
    .B(_15558_),
    .C(_15561_),
    .D(_15613_),
    .X(_15615_));
 sg13g2_a21oi_2 _22940_ (.B1(_15579_),
    .Y(_15616_),
    .A2(_15615_),
    .A1(_15612_));
 sg13g2_a21o_2 _22941_ (.A2(_15615_),
    .A1(_15612_),
    .B1(_15579_),
    .X(_15617_));
 sg13g2_nor4_1 _22942_ (.A(_14221_),
    .B(_14224_),
    .C(_14228_),
    .D(_14232_),
    .Y(_15618_));
 sg13g2_nand2_2 _22943_ (.Y(_15619_),
    .A(_15480_),
    .B(_15618_));
 sg13g2_nor2_1 _22944_ (.A(_15495_),
    .B(_15619_),
    .Y(_15620_));
 sg13g2_nor4_1 _22945_ (.A(_15506_),
    .B(_15512_),
    .C(_15541_),
    .D(_15619_),
    .Y(_15621_));
 sg13g2_a21oi_2 _22946_ (.B1(_15544_),
    .Y(_15622_),
    .A2(_15621_),
    .A1(_15617_));
 sg13g2_a21o_2 _22947_ (.A2(_15621_),
    .A1(_15617_),
    .B1(_15544_),
    .X(_15623_));
 sg13g2_nor4_1 _22948_ (.A(_14517_),
    .B(_14520_),
    .C(_14525_),
    .D(_14530_),
    .Y(_15624_));
 sg13g2_and2_1 _22949_ (.A(_15361_),
    .B(_15624_),
    .X(_15625_));
 sg13g2_nand2_1 _22950_ (.Y(_15626_),
    .A(_15359_),
    .B(_15625_));
 sg13g2_and4_1 _22951_ (.A(_15359_),
    .B(_15397_),
    .C(_15422_),
    .D(_15625_),
    .X(_15627_));
 sg13g2_and2_1 _22952_ (.A(_15352_),
    .B(_15627_),
    .X(_15628_));
 sg13g2_a21oi_2 _22953_ (.B1(_15478_),
    .Y(_15629_),
    .A2(_15628_),
    .A1(_15623_));
 sg13g2_a21o_2 _22954_ (.A2(_15628_),
    .A1(_15623_),
    .B1(_15478_),
    .X(_15630_));
 sg13g2_nor2_1 _22955_ (.A(_14889_),
    .B(_14892_),
    .Y(_15631_));
 sg13g2_nor4_2 _22956_ (.A(_14881_),
    .B(_14885_),
    .C(_14889_),
    .Y(_15632_),
    .D(_14892_));
 sg13g2_nand2_1 _22957_ (.Y(_15633_),
    .A(_15268_),
    .B(_15632_));
 sg13g2_nor2_1 _22958_ (.A(_15266_),
    .B(_15633_),
    .Y(_15634_));
 sg13g2_and2_1 _22959_ (.A(_15260_),
    .B(_15634_),
    .X(_15635_));
 sg13g2_and2_1 _22960_ (.A(_15324_),
    .B(_15635_),
    .X(_15636_));
 sg13g2_a21oi_2 _22961_ (.B1(_15325_),
    .Y(_15637_),
    .A2(_15636_),
    .A1(net3586));
 sg13g2_a21o_2 _22962_ (.A2(_15636_),
    .A1(net3586),
    .B1(_15325_),
    .X(_15638_));
 sg13g2_a21oi_1 _22963_ (.A1(_15188_),
    .A2(_15638_),
    .Y(_15639_),
    .B1(_15183_));
 sg13g2_a21o_1 _22964_ (.A2(_15638_),
    .A1(_15188_),
    .B1(_15183_),
    .X(_15640_));
 sg13g2_nor2_1 _22965_ (.A(net4540),
    .B(_13600_),
    .Y(_15641_));
 sg13g2_nand2_1 _22966_ (.Y(_15642_),
    .A(_15640_),
    .B(_15641_));
 sg13g2_o21ai_1 _22967_ (.B1(net3835),
    .Y(_15643_),
    .A1(net4656),
    .A2(\u_inv.d_next[256] ));
 sg13g2_nor2_1 _22968_ (.A(_13599_),
    .B(_15643_),
    .Y(_15644_));
 sg13g2_inv_1 _22969_ (.Y(_15645_),
    .A(_15644_));
 sg13g2_a21oi_1 _22970_ (.A1(_15640_),
    .A2(_15641_),
    .Y(_15646_),
    .B1(_15645_));
 sg13g2_a21o_2 _22971_ (.A2(_15641_),
    .A1(_15640_),
    .B1(_15645_),
    .X(_15647_));
 sg13g2_and2_1 _22972_ (.A(net3491),
    .B(net3490),
    .X(_15648_));
 sg13g2_nand2_2 _22973_ (.Y(_15649_),
    .A(net3491),
    .B(net3490));
 sg13g2_nand2_1 _22974_ (.Y(_15650_),
    .A(net4799),
    .B(net3741));
 sg13g2_xnor2_1 _22975_ (.Y(_15651_),
    .A(_13997_),
    .B(_15581_));
 sg13g2_nor2_1 _22976_ (.A(net4525),
    .B(_15651_),
    .Y(_15652_));
 sg13g2_a21oi_1 _22977_ (.A1(net4525),
    .A2(_10623_),
    .Y(_15653_),
    .B1(_15652_));
 sg13g2_xor2_1 _22978_ (.B(_15653_),
    .A(_15650_),
    .X(_15654_));
 sg13g2_nor2_1 _22979_ (.A(net3467),
    .B(_15654_),
    .Y(_15655_));
 sg13g2_nand2_2 _22980_ (.Y(_15656_),
    .A(net4635),
    .B(net4799));
 sg13g2_xnor2_1 _22981_ (.Y(_15657_),
    .A(\u_inv.d_next[0] ),
    .B(_15656_));
 sg13g2_xnor2_1 _22982_ (.Y(_15658_),
    .A(_10624_),
    .B(_15656_));
 sg13g2_nand3_1 _22983_ (.B(net3490),
    .C(_15654_),
    .A(net3491),
    .Y(_15659_));
 sg13g2_nand2_1 _22984_ (.Y(_15660_),
    .A(net4305),
    .B(_15659_));
 sg13g2_nand2_1 _22985_ (.Y(_15661_),
    .A(_15654_),
    .B(net4289));
 sg13g2_o21ai_1 _22986_ (.B1(_15661_),
    .Y(_15662_),
    .A1(_15655_),
    .A2(_15660_));
 sg13g2_a22oi_1 _22987_ (.Y(_00277_),
    .B1(net3876),
    .B2(_15662_),
    .A2(net3914),
    .A1(_10624_));
 sg13g2_xnor2_1 _22988_ (.Y(_15663_),
    .A(_13993_),
    .B(_15582_));
 sg13g2_mux2_1 _22989_ (.A0(\u_inv.d_next[2] ),
    .A1(_15663_),
    .S(net4635),
    .X(_15664_));
 sg13g2_xnor2_1 _22990_ (.Y(_15665_),
    .A(_13993_),
    .B(_13999_));
 sg13g2_nor2_1 _22991_ (.A(net3823),
    .B(_15665_),
    .Y(_15666_));
 sg13g2_a21oi_2 _22992_ (.B1(_15666_),
    .Y(_15667_),
    .A2(_15664_),
    .A1(net3823));
 sg13g2_nor2_1 _22993_ (.A(net3467),
    .B(_15667_),
    .Y(_15668_));
 sg13g2_nand3_1 _22994_ (.B(net3490),
    .C(_15667_),
    .A(net3491),
    .Y(_15669_));
 sg13g2_nand3_1 _22995_ (.B(_15659_),
    .C(_15669_),
    .A(net4305),
    .Y(_15670_));
 sg13g2_a21oi_1 _22996_ (.A1(_15660_),
    .A2(_15667_),
    .Y(_15671_),
    .B1(net4232));
 sg13g2_o21ai_1 _22997_ (.B1(_15671_),
    .Y(_15672_),
    .A1(_15668_),
    .A2(_15670_));
 sg13g2_o21ai_1 _22998_ (.B1(_15672_),
    .Y(_00278_),
    .A1(_10623_),
    .A2(net4005));
 sg13g2_a21o_1 _22999_ (.A2(_15667_),
    .A1(_15654_),
    .B1(net3467),
    .X(_15673_));
 sg13g2_xnor2_1 _23000_ (.Y(_15674_),
    .A(_13988_),
    .B(_15583_));
 sg13g2_o21ai_1 _23001_ (.B1(net3823),
    .Y(_15675_),
    .A1(net4635),
    .A2(\u_inv.d_next[3] ));
 sg13g2_a21oi_1 _23002_ (.A1(net4635),
    .A2(_15674_),
    .Y(_15676_),
    .B1(_15675_));
 sg13g2_xnor2_1 _23003_ (.Y(_15677_),
    .A(_13988_),
    .B(_14000_));
 sg13g2_a21oi_1 _23004_ (.A1(net3741),
    .A2(_15677_),
    .Y(_15678_),
    .B1(_15676_));
 sg13g2_nand2_1 _23005_ (.Y(_15679_),
    .A(net3467),
    .B(_15678_));
 sg13g2_inv_1 _23006_ (.Y(_15680_),
    .A(_15679_));
 sg13g2_or2_1 _23007_ (.X(_15681_),
    .B(_15678_),
    .A(net3468));
 sg13g2_a22oi_1 _23008_ (.Y(_15682_),
    .B1(_15679_),
    .B2(_15681_),
    .A2(_15673_),
    .A1(_15670_));
 sg13g2_nand4_1 _23009_ (.B(_15673_),
    .C(_15679_),
    .A(_15670_),
    .Y(_15683_),
    .D(_15681_));
 sg13g2_nand3b_1 _23010_ (.B(_15683_),
    .C(net4305),
    .Y(_15684_),
    .A_N(_15682_));
 sg13g2_a21oi_1 _23011_ (.A1(net4289),
    .A2(_15678_),
    .Y(_15685_),
    .B1(net4232));
 sg13g2_a22oi_1 _23012_ (.Y(_15686_),
    .B1(_15684_),
    .B2(_15685_),
    .A2(net3914),
    .A1(net3030));
 sg13g2_inv_1 _23013_ (.Y(_00279_),
    .A(_15686_));
 sg13g2_xor2_1 _23014_ (.B(_14003_),
    .A(_14001_),
    .X(_15687_));
 sg13g2_nand2b_1 _23015_ (.Y(_15688_),
    .B(_15584_),
    .A_N(_14003_));
 sg13g2_nand3_1 _23016_ (.B(_15585_),
    .C(_15688_),
    .A(net4635),
    .Y(_15689_));
 sg13g2_a21oi_1 _23017_ (.A1(net4525),
    .A2(\u_inv.d_next[4] ),
    .Y(_15690_),
    .B1(net3741));
 sg13g2_nand2_1 _23018_ (.Y(_15691_),
    .A(_15689_),
    .B(_15690_));
 sg13g2_o21ai_1 _23019_ (.B1(_15691_),
    .Y(_15692_),
    .A1(net3823),
    .A2(_15687_));
 sg13g2_nand2_1 _23020_ (.Y(_15693_),
    .A(net3467),
    .B(_15692_));
 sg13g2_xnor2_1 _23021_ (.Y(_15694_),
    .A(net3467),
    .B(_15692_));
 sg13g2_inv_1 _23022_ (.Y(_15695_),
    .A(_15694_));
 sg13g2_and3_1 _23023_ (.X(_15696_),
    .A(_15670_),
    .B(_15673_),
    .C(_15681_));
 sg13g2_or3_1 _23024_ (.A(_15680_),
    .B(_15695_),
    .C(_15696_),
    .X(_15697_));
 sg13g2_o21ai_1 _23025_ (.B1(_15695_),
    .Y(_15698_),
    .A1(_15680_),
    .A2(_15696_));
 sg13g2_a21oi_1 _23026_ (.A1(_15697_),
    .A2(_15698_),
    .Y(_15699_),
    .B1(net4289));
 sg13g2_a21o_1 _23027_ (.A2(_15692_),
    .A1(net4289),
    .B1(net4232),
    .X(_15700_));
 sg13g2_nand2_1 _23028_ (.Y(_15701_),
    .A(net2797),
    .B(net3914));
 sg13g2_o21ai_1 _23029_ (.B1(_15701_),
    .Y(_00280_),
    .A1(_15699_),
    .A2(_15700_));
 sg13g2_nand2_1 _23030_ (.Y(_15702_),
    .A(net2155),
    .B(net3914));
 sg13g2_o21ai_1 _23031_ (.B1(_15697_),
    .Y(_15703_),
    .A1(net3398),
    .A2(_15692_));
 sg13g2_nor2_1 _23032_ (.A(_14002_),
    .B(_14007_),
    .Y(_15704_));
 sg13g2_a21oi_1 _23033_ (.A1(_15585_),
    .A2(_15704_),
    .Y(_15705_),
    .B1(_15591_));
 sg13g2_nand3_1 _23034_ (.B(_15586_),
    .C(_15705_),
    .A(net4635),
    .Y(_15706_));
 sg13g2_a21oi_1 _23035_ (.A1(net4525),
    .A2(\u_inv.d_next[5] ),
    .Y(_15707_),
    .B1(net3741));
 sg13g2_nor3_1 _23036_ (.A(_14004_),
    .B(_14006_),
    .C(_14007_),
    .Y(_15708_));
 sg13g2_o21ai_1 _23037_ (.B1(_14007_),
    .Y(_15709_),
    .A1(_14004_),
    .A2(_14006_));
 sg13g2_nor2_1 _23038_ (.A(net3823),
    .B(_15708_),
    .Y(_15710_));
 sg13g2_a22oi_1 _23039_ (.Y(_15711_),
    .B1(_15709_),
    .B2(_15710_),
    .A2(_15707_),
    .A1(_15706_));
 sg13g2_xnor2_1 _23040_ (.Y(_15712_),
    .A(net3393),
    .B(_15711_));
 sg13g2_o21ai_1 _23041_ (.B1(net4300),
    .Y(_15713_),
    .A1(_15703_),
    .A2(_15712_));
 sg13g2_a21oi_1 _23042_ (.A1(_15703_),
    .A2(_15712_),
    .Y(_15714_),
    .B1(_15713_));
 sg13g2_o21ai_1 _23043_ (.B1(net3874),
    .Y(_15715_),
    .A1(net4301),
    .A2(_15711_));
 sg13g2_o21ai_1 _23044_ (.B1(_15702_),
    .Y(_00281_),
    .A1(_15714_),
    .A2(_15715_));
 sg13g2_nand2_1 _23045_ (.Y(_15716_),
    .A(_13983_),
    .B(_14012_));
 sg13g2_xnor2_1 _23046_ (.Y(_15717_),
    .A(_13983_),
    .B(_14012_));
 sg13g2_nand3_1 _23047_ (.B(_15586_),
    .C(_15592_),
    .A(_13983_),
    .Y(_15718_));
 sg13g2_a21oi_1 _23048_ (.A1(_15586_),
    .A2(_15592_),
    .Y(_15719_),
    .B1(_13983_));
 sg13g2_nor2_1 _23049_ (.A(net4525),
    .B(_15719_),
    .Y(_15720_));
 sg13g2_a221oi_1 _23050_ (.B2(_15720_),
    .C1(net3741),
    .B1(_15718_),
    .A1(net4525),
    .Y(_15721_),
    .A2(net4806));
 sg13g2_a21o_2 _23051_ (.A2(_15717_),
    .A1(net3741),
    .B1(_15721_),
    .X(_15722_));
 sg13g2_or2_1 _23052_ (.X(_15723_),
    .B(_15722_),
    .A(net3393));
 sg13g2_xnor2_1 _23053_ (.Y(_15724_),
    .A(net3470),
    .B(_15722_));
 sg13g2_nand2_1 _23054_ (.Y(_15725_),
    .A(_15693_),
    .B(_15711_));
 sg13g2_o21ai_1 _23055_ (.B1(_15725_),
    .Y(_15726_),
    .A1(_15697_),
    .A2(_15712_));
 sg13g2_nand2_1 _23056_ (.Y(_15727_),
    .A(_15724_),
    .B(_15726_));
 sg13g2_xor2_1 _23057_ (.B(_15726_),
    .A(_15724_),
    .X(_15728_));
 sg13g2_o21ai_1 _23058_ (.B1(net3874),
    .Y(_15729_),
    .A1(net4289),
    .A2(_15728_));
 sg13g2_a21oi_1 _23059_ (.A1(net4289),
    .A2(_15722_),
    .Y(_15730_),
    .B1(_15729_));
 sg13g2_a21o_1 _23060_ (.A2(net3914),
    .A1(net2816),
    .B1(_15730_),
    .X(_00282_));
 sg13g2_a21oi_1 _23061_ (.A1(net4806),
    .A2(net4795),
    .Y(_15731_),
    .B1(_15719_));
 sg13g2_a21oi_1 _23062_ (.A1(_15587_),
    .A2(_15731_),
    .Y(_15732_),
    .B1(net4525));
 sg13g2_o21ai_1 _23063_ (.B1(_15732_),
    .Y(_15733_),
    .A1(_15587_),
    .A2(_15731_));
 sg13g2_a21oi_1 _23064_ (.A1(net4525),
    .A2(\u_inv.d_next[7] ),
    .Y(_15734_),
    .B1(net3741));
 sg13g2_a21oi_1 _23065_ (.A1(_13979_),
    .A2(_15716_),
    .Y(_15735_),
    .B1(_15587_));
 sg13g2_nand3_1 _23066_ (.B(_15587_),
    .C(_15716_),
    .A(_13979_),
    .Y(_15736_));
 sg13g2_nor2_1 _23067_ (.A(net3823),
    .B(_15735_),
    .Y(_15737_));
 sg13g2_a22oi_1 _23068_ (.Y(_15738_),
    .B1(_15736_),
    .B2(_15737_),
    .A2(_15734_),
    .A1(_15733_));
 sg13g2_nand2_1 _23069_ (.Y(_15739_),
    .A(net3470),
    .B(_15738_));
 sg13g2_xnor2_1 _23070_ (.Y(_15740_),
    .A(net3394),
    .B(_15738_));
 sg13g2_nand2_1 _23071_ (.Y(_15741_),
    .A(_15723_),
    .B(_15727_));
 sg13g2_xnor2_1 _23072_ (.Y(_15742_),
    .A(_15740_),
    .B(_15741_));
 sg13g2_o21ai_1 _23073_ (.B1(net3874),
    .Y(_15743_),
    .A1(net4301),
    .A2(_15738_));
 sg13g2_a21oi_1 _23074_ (.A1(net4301),
    .A2(_15742_),
    .Y(_15744_),
    .B1(_15743_));
 sg13g2_a21o_1 _23075_ (.A2(net3914),
    .A1(net4806),
    .B1(_15744_),
    .X(_00283_));
 sg13g2_nor2b_1 _23076_ (.A(_14018_),
    .B_N(_14015_),
    .Y(_15745_));
 sg13g2_xnor2_1 _23077_ (.Y(_15746_),
    .A(_14015_),
    .B(_14018_));
 sg13g2_xnor2_1 _23078_ (.Y(_15747_),
    .A(_14018_),
    .B(_15596_));
 sg13g2_o21ai_1 _23079_ (.B1(net3824),
    .Y(_15748_),
    .A1(net4634),
    .A2(\u_inv.d_next[8] ));
 sg13g2_a21oi_1 _23080_ (.A1(net4634),
    .A2(_15747_),
    .Y(_15749_),
    .B1(_15748_));
 sg13g2_a21oi_1 _23081_ (.A1(net3739),
    .A2(_15746_),
    .Y(_15750_),
    .B1(_15749_));
 sg13g2_inv_1 _23082_ (.Y(_15751_),
    .A(_15750_));
 sg13g2_xnor2_1 _23083_ (.Y(_15752_),
    .A(net3398),
    .B(_15751_));
 sg13g2_nand3b_1 _23084_ (.B(_15724_),
    .C(_15740_),
    .Y(_15753_),
    .A_N(_15712_));
 sg13g2_nor4_1 _23085_ (.A(_15680_),
    .B(_15695_),
    .C(_15696_),
    .D(_15753_),
    .Y(_15754_));
 sg13g2_nand4_1 _23086_ (.B(_15711_),
    .C(_15724_),
    .A(_15693_),
    .Y(_15755_),
    .D(_15740_));
 sg13g2_nand3_1 _23087_ (.B(_15739_),
    .C(_15755_),
    .A(_15723_),
    .Y(_15756_));
 sg13g2_or2_1 _23088_ (.X(_15757_),
    .B(_15756_),
    .A(_15754_));
 sg13g2_and2_1 _23089_ (.A(_15752_),
    .B(_15757_),
    .X(_15758_));
 sg13g2_xor2_1 _23090_ (.B(_15757_),
    .A(_15752_),
    .X(_15759_));
 sg13g2_a21oi_1 _23091_ (.A1(net4289),
    .A2(_15750_),
    .Y(_15760_),
    .B1(net4232));
 sg13g2_o21ai_1 _23092_ (.B1(_15760_),
    .Y(_15761_),
    .A1(net4289),
    .A2(_15759_));
 sg13g2_o21ai_1 _23093_ (.B1(_15761_),
    .Y(_00284_),
    .A1(_10622_),
    .A2(net4005));
 sg13g2_nand2_1 _23094_ (.Y(_15762_),
    .A(net2516),
    .B(net3913));
 sg13g2_a21oi_1 _23095_ (.A1(_14018_),
    .A2(_15596_),
    .Y(_15763_),
    .B1(_14017_));
 sg13g2_nand2b_1 _23096_ (.Y(_15764_),
    .B(_15763_),
    .A_N(_14016_));
 sg13g2_nand3_1 _23097_ (.B(_14018_),
    .C(_15596_),
    .A(_14016_),
    .Y(_15765_));
 sg13g2_a21oi_1 _23098_ (.A1(_14016_),
    .A2(_14017_),
    .Y(_15766_),
    .B1(net4524));
 sg13g2_nand3_1 _23099_ (.B(_15765_),
    .C(_15766_),
    .A(_15764_),
    .Y(_15767_));
 sg13g2_a21oi_1 _23100_ (.A1(net4524),
    .A2(\u_inv.d_next[9] ),
    .Y(_15768_),
    .B1(net3739));
 sg13g2_a21oi_1 _23101_ (.A1(\u_inv.d_next[8] ),
    .A2(_10956_),
    .Y(_15769_),
    .B1(_15745_));
 sg13g2_xnor2_1 _23102_ (.Y(_15770_),
    .A(_14016_),
    .B(_15769_));
 sg13g2_a22oi_1 _23103_ (.Y(_15771_),
    .B1(_15770_),
    .B2(net3739),
    .A2(_15768_),
    .A1(_15767_));
 sg13g2_xnor2_1 _23104_ (.Y(_15772_),
    .A(net3398),
    .B(_15771_));
 sg13g2_a21oi_1 _23105_ (.A1(net3467),
    .A2(_15751_),
    .Y(_15773_),
    .B1(_15758_));
 sg13g2_o21ai_1 _23106_ (.B1(net4305),
    .Y(_15774_),
    .A1(_15772_),
    .A2(_15773_));
 sg13g2_a21oi_1 _23107_ (.A1(_15772_),
    .A2(_15773_),
    .Y(_15775_),
    .B1(_15774_));
 sg13g2_o21ai_1 _23108_ (.B1(net3876),
    .Y(_15776_),
    .A1(net4305),
    .A2(_15771_));
 sg13g2_o21ai_1 _23109_ (.B1(_15762_),
    .Y(_00285_),
    .A1(_15775_),
    .A2(_15776_));
 sg13g2_a21oi_2 _23110_ (.B1(_14022_),
    .Y(_15777_),
    .A2(_14019_),
    .A1(_14015_));
 sg13g2_inv_1 _23111_ (.Y(_15778_),
    .A(_15777_));
 sg13g2_xor2_1 _23112_ (.B(_15777_),
    .A(_13974_),
    .X(_15779_));
 sg13g2_nand3_1 _23113_ (.B(_15603_),
    .C(_15765_),
    .A(_13974_),
    .Y(_15780_));
 sg13g2_a21o_1 _23114_ (.A2(_15765_),
    .A1(_15603_),
    .B1(_13974_),
    .X(_15781_));
 sg13g2_nand3_1 _23115_ (.B(_15780_),
    .C(_15781_),
    .A(net4634),
    .Y(_15782_));
 sg13g2_a21oi_1 _23116_ (.A1(net4524),
    .A2(\u_inv.d_next[10] ),
    .Y(_15783_),
    .B1(net3739));
 sg13g2_a22oi_1 _23117_ (.Y(_15784_),
    .B1(_15782_),
    .B2(_15783_),
    .A2(_15779_),
    .A1(net3739));
 sg13g2_nand2_1 _23118_ (.Y(_15785_),
    .A(net3398),
    .B(_15784_));
 sg13g2_xnor2_1 _23119_ (.Y(_15786_),
    .A(net3398),
    .B(_15784_));
 sg13g2_o21ai_1 _23120_ (.B1(net3467),
    .Y(_15787_),
    .A1(_15751_),
    .A2(_15771_));
 sg13g2_and2_1 _23121_ (.A(_15758_),
    .B(_15772_),
    .X(_15788_));
 sg13g2_nor2b_1 _23122_ (.A(_15788_),
    .B_N(_15787_),
    .Y(_15789_));
 sg13g2_xnor2_1 _23123_ (.Y(_15790_),
    .A(_15786_),
    .B(_15789_));
 sg13g2_o21ai_1 _23124_ (.B1(net3876),
    .Y(_15791_),
    .A1(net4305),
    .A2(_15784_));
 sg13g2_a21oi_1 _23125_ (.A1(net4305),
    .A2(_15790_),
    .Y(_15792_),
    .B1(_15791_));
 sg13g2_a21o_1 _23126_ (.A2(net3913),
    .A1(net2901),
    .B1(_15792_),
    .X(_00286_));
 sg13g2_nand2_1 _23127_ (.Y(_15793_),
    .A(net2066),
    .B(net3920));
 sg13g2_nand3_1 _23128_ (.B(_13973_),
    .C(_15781_),
    .A(_13971_),
    .Y(_15794_));
 sg13g2_a21o_1 _23129_ (.A2(_15781_),
    .A1(_13973_),
    .B1(_13971_),
    .X(_15795_));
 sg13g2_nand3_1 _23130_ (.B(_15794_),
    .C(_15795_),
    .A(net4634),
    .Y(_15796_));
 sg13g2_a21oi_1 _23131_ (.A1(net4524),
    .A2(\u_inv.d_next[11] ),
    .Y(_15797_),
    .B1(net3740));
 sg13g2_a21oi_1 _23132_ (.A1(_13974_),
    .A2(_15778_),
    .Y(_15798_),
    .B1(_14023_));
 sg13g2_xnor2_1 _23133_ (.Y(_15799_),
    .A(_13972_),
    .B(_15798_));
 sg13g2_a22oi_1 _23134_ (.Y(_15800_),
    .B1(_15799_),
    .B2(net3739),
    .A2(_15797_),
    .A1(_15796_));
 sg13g2_xnor2_1 _23135_ (.Y(_15801_),
    .A(net3398),
    .B(_15800_));
 sg13g2_o21ai_1 _23136_ (.B1(_15785_),
    .Y(_15802_),
    .A1(_15786_),
    .A2(_15789_));
 sg13g2_o21ai_1 _23137_ (.B1(net4305),
    .Y(_15803_),
    .A1(_15801_),
    .A2(_15802_));
 sg13g2_a21oi_1 _23138_ (.A1(_15801_),
    .A2(_15802_),
    .Y(_15804_),
    .B1(_15803_));
 sg13g2_o21ai_1 _23139_ (.B1(net3876),
    .Y(_15805_),
    .A1(net4306),
    .A2(_15800_));
 sg13g2_o21ai_1 _23140_ (.B1(_15793_),
    .Y(_00287_),
    .A1(_15804_),
    .A2(_15805_));
 sg13g2_o21ai_1 _23141_ (.B1(_14024_),
    .Y(_15806_),
    .A1(_13975_),
    .A2(_15777_));
 sg13g2_nand2b_1 _23142_ (.Y(_15807_),
    .B(_15806_),
    .A_N(_13966_));
 sg13g2_xor2_1 _23143_ (.B(_15806_),
    .A(_13966_),
    .X(_15808_));
 sg13g2_o21ai_1 _23144_ (.B1(_15605_),
    .Y(_15809_),
    .A1(_15598_),
    .A2(_15765_));
 sg13g2_a21oi_1 _23145_ (.A1(_13966_),
    .A2(_15809_),
    .Y(_15810_),
    .B1(net4524));
 sg13g2_o21ai_1 _23146_ (.B1(_15810_),
    .Y(_15811_),
    .A1(_13966_),
    .A2(_15809_));
 sg13g2_a21oi_1 _23147_ (.A1(net4529),
    .A2(\u_inv.d_next[12] ),
    .Y(_15812_),
    .B1(net3739));
 sg13g2_a22oi_1 _23148_ (.Y(_15813_),
    .B1(_15811_),
    .B2(_15812_),
    .A2(_15808_),
    .A1(net3739));
 sg13g2_and2_1 _23149_ (.A(net3398),
    .B(_15813_),
    .X(_15814_));
 sg13g2_xnor2_1 _23150_ (.Y(_15815_),
    .A(net3399),
    .B(_15813_));
 sg13g2_nor2_1 _23151_ (.A(_15786_),
    .B(_15801_),
    .Y(_15816_));
 sg13g2_nor3_1 _23152_ (.A(_15786_),
    .B(_15787_),
    .C(_15801_),
    .Y(_15817_));
 sg13g2_o21ai_1 _23153_ (.B1(net3398),
    .Y(_15818_),
    .A1(_15784_),
    .A2(_15800_));
 sg13g2_nand2b_1 _23154_ (.Y(_15819_),
    .B(_15818_),
    .A_N(_15817_));
 sg13g2_a21oi_1 _23155_ (.A1(_15788_),
    .A2(_15816_),
    .Y(_15820_),
    .B1(_15819_));
 sg13g2_nor2_1 _23156_ (.A(_15815_),
    .B(_15820_),
    .Y(_15821_));
 sg13g2_xnor2_1 _23157_ (.Y(_15822_),
    .A(_15815_),
    .B(_15820_));
 sg13g2_o21ai_1 _23158_ (.B1(net3876),
    .Y(_15823_),
    .A1(net4306),
    .A2(_15813_));
 sg13g2_a21oi_1 _23159_ (.A1(net4306),
    .A2(_15822_),
    .Y(_15824_),
    .B1(_15823_));
 sg13g2_a21o_1 _23160_ (.A2(net3914),
    .A1(net2492),
    .B1(_15824_),
    .X(_00288_));
 sg13g2_nand2b_1 _23161_ (.Y(_15825_),
    .B(net3824),
    .A_N(\u_inv.d_next[13] ));
 sg13g2_a21oi_1 _23162_ (.A1(_13966_),
    .A2(_15809_),
    .Y(_15826_),
    .B1(_13965_));
 sg13g2_xnor2_1 _23163_ (.Y(_15827_),
    .A(_13964_),
    .B(_15826_));
 sg13g2_a22oi_1 _23164_ (.Y(_15828_),
    .B1(_15827_),
    .B2(net4634),
    .A2(_15825_),
    .A1(net3723));
 sg13g2_and2_1 _23165_ (.A(_14029_),
    .B(_15807_),
    .X(_15829_));
 sg13g2_nor2b_1 _23166_ (.A(_15829_),
    .B_N(_13964_),
    .Y(_15830_));
 sg13g2_nor2b_1 _23167_ (.A(_13964_),
    .B_N(_15829_),
    .Y(_15831_));
 sg13g2_nor3_1 _23168_ (.A(net3824),
    .B(_15830_),
    .C(_15831_),
    .Y(_15832_));
 sg13g2_or2_1 _23169_ (.X(_15833_),
    .B(_15832_),
    .A(_15828_));
 sg13g2_nor2_1 _23170_ (.A(net3468),
    .B(_15833_),
    .Y(_15834_));
 sg13g2_nand2_1 _23171_ (.Y(_15835_),
    .A(net3468),
    .B(_15833_));
 sg13g2_xnor2_1 _23172_ (.Y(_15836_),
    .A(net3468),
    .B(_15833_));
 sg13g2_nor2_1 _23173_ (.A(_15814_),
    .B(_15821_),
    .Y(_15837_));
 sg13g2_xnor2_1 _23174_ (.Y(_15838_),
    .A(_15836_),
    .B(_15837_));
 sg13g2_nand2_1 _23175_ (.Y(_15839_),
    .A(net4306),
    .B(_15838_));
 sg13g2_a21oi_1 _23176_ (.A1(net4290),
    .A2(_15833_),
    .Y(_15840_),
    .B1(net4232));
 sg13g2_a22oi_1 _23177_ (.Y(_15841_),
    .B1(_15839_),
    .B2(_15840_),
    .A2(net3913),
    .A1(net2511));
 sg13g2_inv_1 _23178_ (.Y(_00289_),
    .A(_15841_));
 sg13g2_a21oi_1 _23179_ (.A1(_13967_),
    .A2(_15806_),
    .Y(_15842_),
    .B1(_14030_));
 sg13g2_xnor2_1 _23180_ (.Y(_15843_),
    .A(_13961_),
    .B(_15842_));
 sg13g2_nand2_1 _23181_ (.Y(_15844_),
    .A(net3740),
    .B(_15843_));
 sg13g2_and3_1 _23182_ (.X(_15845_),
    .A(_13964_),
    .B(_13966_),
    .C(_15809_));
 sg13g2_nor3_1 _23183_ (.A(_13961_),
    .B(_15607_),
    .C(_15845_),
    .Y(_15846_));
 sg13g2_o21ai_1 _23184_ (.B1(_13961_),
    .Y(_15847_),
    .A1(_15607_),
    .A2(_15845_));
 sg13g2_nand2_1 _23185_ (.Y(_15848_),
    .A(net4655),
    .B(_15847_));
 sg13g2_a21oi_1 _23186_ (.A1(net4524),
    .A2(\u_inv.d_next[14] ),
    .Y(_15849_),
    .B1(net3740));
 sg13g2_o21ai_1 _23187_ (.B1(_15849_),
    .Y(_15850_),
    .A1(_15846_),
    .A2(_15848_));
 sg13g2_nand2_2 _23188_ (.Y(_15851_),
    .A(_15844_),
    .B(_15850_));
 sg13g2_xnor2_1 _23189_ (.Y(_15852_),
    .A(net3469),
    .B(_15851_));
 sg13g2_or2_1 _23190_ (.X(_15853_),
    .B(_15834_),
    .A(_15814_));
 sg13g2_o21ai_1 _23191_ (.B1(_15835_),
    .Y(_15854_),
    .A1(_15821_),
    .A2(_15853_));
 sg13g2_or2_1 _23192_ (.X(_15855_),
    .B(_15854_),
    .A(_15852_));
 sg13g2_xor2_1 _23193_ (.B(_15854_),
    .A(_15852_),
    .X(_15856_));
 sg13g2_o21ai_1 _23194_ (.B1(net3876),
    .Y(_15857_),
    .A1(net4290),
    .A2(_15856_));
 sg13g2_a21oi_1 _23195_ (.A1(net4291),
    .A2(_15851_),
    .Y(_15858_),
    .B1(_15857_));
 sg13g2_a21o_1 _23196_ (.A2(net3913),
    .A1(net2727),
    .B1(_15858_),
    .X(_00290_));
 sg13g2_nand3_1 _23197_ (.B(_13960_),
    .C(_15847_),
    .A(_13958_),
    .Y(_15859_));
 sg13g2_a21oi_1 _23198_ (.A1(_13960_),
    .A2(_15847_),
    .Y(_15860_),
    .B1(_13958_));
 sg13g2_nand2_1 _23199_ (.Y(_15861_),
    .A(net4635),
    .B(_15859_));
 sg13g2_a21oi_1 _23200_ (.A1(net4524),
    .A2(\u_inv.d_next[15] ),
    .Y(_15862_),
    .B1(net3740));
 sg13g2_o21ai_1 _23201_ (.B1(_15862_),
    .Y(_15863_),
    .A1(_15860_),
    .A2(_15861_));
 sg13g2_o21ai_1 _23202_ (.B1(_14026_),
    .Y(_15864_),
    .A1(_13961_),
    .A2(_15842_));
 sg13g2_xnor2_1 _23203_ (.Y(_15865_),
    .A(_13959_),
    .B(_15864_));
 sg13g2_o21ai_1 _23204_ (.B1(_15863_),
    .Y(_15866_),
    .A1(net3824),
    .A2(_15865_));
 sg13g2_xnor2_1 _23205_ (.Y(_15867_),
    .A(net3469),
    .B(_15866_));
 sg13g2_o21ai_1 _23206_ (.B1(_15855_),
    .Y(_15868_),
    .A1(net3469),
    .A2(_15851_));
 sg13g2_a21oi_1 _23207_ (.A1(_15867_),
    .A2(_15868_),
    .Y(_15869_),
    .B1(net4290));
 sg13g2_o21ai_1 _23208_ (.B1(_15869_),
    .Y(_15870_),
    .A1(_15867_),
    .A2(_15868_));
 sg13g2_a21oi_1 _23209_ (.A1(net4291),
    .A2(_15866_),
    .Y(_15871_),
    .B1(net4232));
 sg13g2_a22oi_1 _23210_ (.Y(_15872_),
    .B1(_15870_),
    .B2(_15871_),
    .A2(net3913),
    .A1(net2945));
 sg13g2_inv_1 _23211_ (.Y(_00291_),
    .A(_15872_));
 sg13g2_nor2_1 _23212_ (.A(_14033_),
    .B(_14071_),
    .Y(_15873_));
 sg13g2_xnor2_1 _23213_ (.Y(_15874_),
    .A(_14033_),
    .B(_14071_));
 sg13g2_a21oi_1 _23214_ (.A1(_14071_),
    .A2(_15612_),
    .Y(_15875_),
    .B1(net4531));
 sg13g2_o21ai_1 _23215_ (.B1(_15875_),
    .Y(_15876_),
    .A1(_14071_),
    .A2(_15612_));
 sg13g2_a21oi_1 _23216_ (.A1(net4531),
    .A2(\u_inv.d_next[16] ),
    .Y(_15877_),
    .B1(net3746));
 sg13g2_a22oi_1 _23217_ (.Y(_15878_),
    .B1(_15876_),
    .B2(_15877_),
    .A2(_15874_),
    .A1(net3746));
 sg13g2_xnor2_1 _23218_ (.Y(_15879_),
    .A(net3470),
    .B(_15878_));
 sg13g2_nor2_1 _23219_ (.A(_15852_),
    .B(_15867_),
    .Y(_15880_));
 sg13g2_nor4_1 _23220_ (.A(_15815_),
    .B(_15836_),
    .C(_15852_),
    .D(_15867_),
    .Y(_15881_));
 sg13g2_a21oi_1 _23221_ (.A1(_15851_),
    .A2(_15866_),
    .Y(_15882_),
    .B1(net3469));
 sg13g2_a221oi_1 _23222_ (.B2(_15819_),
    .C1(_15882_),
    .B1(_15881_),
    .A1(_15853_),
    .Y(_15883_),
    .A2(_15880_));
 sg13g2_and4_1 _23223_ (.A(_15752_),
    .B(_15772_),
    .C(_15816_),
    .D(_15881_),
    .X(_15884_));
 sg13g2_o21ai_1 _23224_ (.B1(_15884_),
    .Y(_15885_),
    .A1(_15754_),
    .A2(_15756_));
 sg13g2_nand2_1 _23225_ (.Y(_15886_),
    .A(_15883_),
    .B(_15885_));
 sg13g2_and2_1 _23226_ (.A(_15879_),
    .B(_15886_),
    .X(_15887_));
 sg13g2_xnor2_1 _23227_ (.Y(_15888_),
    .A(_15879_),
    .B(_15886_));
 sg13g2_o21ai_1 _23228_ (.B1(net3876),
    .Y(_15889_),
    .A1(net4304),
    .A2(_15878_));
 sg13g2_a21oi_1 _23229_ (.A1(net4304),
    .A2(_15888_),
    .Y(_15890_),
    .B1(_15889_));
 sg13g2_a21o_1 _23230_ (.A2(net3913),
    .A1(net3215),
    .B1(_15890_),
    .X(_00292_));
 sg13g2_nand2_1 _23231_ (.Y(_15891_),
    .A(net2028),
    .B(net3921));
 sg13g2_a21oi_1 _23232_ (.A1(_14071_),
    .A2(_15612_),
    .Y(_15892_),
    .B1(_14069_));
 sg13g2_nand2_1 _23233_ (.Y(_15893_),
    .A(_14070_),
    .B(_15892_));
 sg13g2_nand4_1 _23234_ (.B(_15545_),
    .C(_15614_),
    .A(net4643),
    .Y(_15894_),
    .D(_15893_));
 sg13g2_a21oi_1 _23235_ (.A1(net4531),
    .A2(net4805),
    .Y(_15895_),
    .B1(net3746));
 sg13g2_nor2_1 _23236_ (.A(_14097_),
    .B(_15873_),
    .Y(_15896_));
 sg13g2_xnor2_1 _23237_ (.Y(_15897_),
    .A(_14069_),
    .B(_15896_));
 sg13g2_a22oi_1 _23238_ (.Y(_15898_),
    .B1(_15897_),
    .B2(net3746),
    .A2(_15895_),
    .A1(_15894_));
 sg13g2_xnor2_1 _23239_ (.Y(_15899_),
    .A(net3469),
    .B(_15898_));
 sg13g2_a21oi_1 _23240_ (.A1(net3399),
    .A2(_15878_),
    .Y(_15900_),
    .B1(_15887_));
 sg13g2_o21ai_1 _23241_ (.B1(net4307),
    .Y(_15901_),
    .A1(_15899_),
    .A2(_15900_));
 sg13g2_a21oi_1 _23242_ (.A1(_15899_),
    .A2(_15900_),
    .Y(_15902_),
    .B1(_15901_));
 sg13g2_o21ai_1 _23243_ (.B1(net3876),
    .Y(_15903_),
    .A1(net4307),
    .A2(_15898_));
 sg13g2_o21ai_1 _23244_ (.B1(_15891_),
    .Y(_00293_),
    .A1(_15902_),
    .A2(_15903_));
 sg13g2_a21oi_1 _23245_ (.A1(_15547_),
    .A2(_15614_),
    .Y(_15904_),
    .B1(_14065_));
 sg13g2_nand3_1 _23246_ (.B(_15547_),
    .C(_15614_),
    .A(_14065_),
    .Y(_15905_));
 sg13g2_nand2b_1 _23247_ (.Y(_15906_),
    .B(_15905_),
    .A_N(_15904_));
 sg13g2_o21ai_1 _23248_ (.B1(net3829),
    .Y(_15907_),
    .A1(net4643),
    .A2(\u_inv.d_next[18] ));
 sg13g2_a21oi_1 _23249_ (.A1(net4644),
    .A2(_15906_),
    .Y(_15908_),
    .B1(_15907_));
 sg13g2_o21ai_1 _23250_ (.B1(_14098_),
    .Y(_15909_),
    .A1(_14033_),
    .A2(_14071_));
 sg13g2_a21oi_1 _23251_ (.A1(_14067_),
    .A2(_15909_),
    .Y(_15910_),
    .B1(_14065_));
 sg13g2_nand3_1 _23252_ (.B(_14067_),
    .C(_15909_),
    .A(_14065_),
    .Y(_15911_));
 sg13g2_nor2_1 _23253_ (.A(net3829),
    .B(_15910_),
    .Y(_15912_));
 sg13g2_a21oi_2 _23254_ (.B1(_15908_),
    .Y(_15913_),
    .A2(_15912_),
    .A1(_15911_));
 sg13g2_nor2_1 _23255_ (.A(net3469),
    .B(_15913_),
    .Y(_15914_));
 sg13g2_xnor2_1 _23256_ (.Y(_15915_),
    .A(net3469),
    .B(_15913_));
 sg13g2_o21ai_1 _23257_ (.B1(net3399),
    .Y(_15916_),
    .A1(_15878_),
    .A2(_15898_));
 sg13g2_nand2_1 _23258_ (.Y(_15917_),
    .A(_15887_),
    .B(_15899_));
 sg13g2_nand2_1 _23259_ (.Y(_15918_),
    .A(_15916_),
    .B(_15917_));
 sg13g2_a21oi_1 _23260_ (.A1(_15916_),
    .A2(_15917_),
    .Y(_15919_),
    .B1(_15915_));
 sg13g2_xnor2_1 _23261_ (.Y(_15920_),
    .A(_15915_),
    .B(_15918_));
 sg13g2_nor2_1 _23262_ (.A(net4291),
    .B(_15920_),
    .Y(_15921_));
 sg13g2_a21oi_1 _23263_ (.A1(net4290),
    .A2(_15913_),
    .Y(_15922_),
    .B1(_15921_));
 sg13g2_a22oi_1 _23264_ (.Y(_15923_),
    .B1(net3877),
    .B2(_15922_),
    .A2(net3921),
    .A1(net4805));
 sg13g2_inv_1 _23265_ (.Y(_00294_),
    .A(_15923_));
 sg13g2_a21oi_1 _23266_ (.A1(net4531),
    .A2(\u_inv.d_next[19] ),
    .Y(_15924_),
    .B1(net3746));
 sg13g2_a21oi_1 _23267_ (.A1(\u_inv.d_next[18] ),
    .A2(\u_inv.d_reg[18] ),
    .Y(_15925_),
    .B1(_15904_));
 sg13g2_xnor2_1 _23268_ (.Y(_15926_),
    .A(_14063_),
    .B(_15925_));
 sg13g2_nand2_1 _23269_ (.Y(_15927_),
    .A(net4644),
    .B(_15926_));
 sg13g2_nand2_1 _23270_ (.Y(_15928_),
    .A(_14100_),
    .B(_15911_));
 sg13g2_o21ai_1 _23271_ (.B1(net3746),
    .Y(_15929_),
    .A1(_14063_),
    .A2(_15928_));
 sg13g2_a21oi_1 _23272_ (.A1(_14063_),
    .A2(_15928_),
    .Y(_15930_),
    .B1(_15929_));
 sg13g2_a21oi_2 _23273_ (.B1(_15930_),
    .Y(_15931_),
    .A2(_15927_),
    .A1(_15924_));
 sg13g2_xnor2_1 _23274_ (.Y(_15932_),
    .A(net3399),
    .B(_15931_));
 sg13g2_nor2_1 _23275_ (.A(_15914_),
    .B(_15919_),
    .Y(_15933_));
 sg13g2_xnor2_1 _23276_ (.Y(_15934_),
    .A(_15932_),
    .B(_15933_));
 sg13g2_o21ai_1 _23277_ (.B1(net3877),
    .Y(_15935_),
    .A1(net4307),
    .A2(_15931_));
 sg13g2_a21oi_1 _23278_ (.A1(net4307),
    .A2(_15934_),
    .Y(_15936_),
    .B1(_15935_));
 sg13g2_a21o_1 _23279_ (.A2(net3922),
    .A1(net3191),
    .B1(_15936_),
    .X(_00295_));
 sg13g2_and3_1 _23280_ (.X(_15937_),
    .A(_15550_),
    .B(_15612_),
    .C(_15613_));
 sg13g2_nand2b_2 _23281_ (.Y(_15938_),
    .B(_15551_),
    .A_N(_15937_));
 sg13g2_xnor2_1 _23282_ (.Y(_15939_),
    .A(_14086_),
    .B(_15938_));
 sg13g2_o21ai_1 _23283_ (.B1(net3829),
    .Y(_15940_),
    .A1(net4644),
    .A2(\u_inv.d_next[20] ));
 sg13g2_a21o_1 _23284_ (.A2(_15939_),
    .A1(net4644),
    .B1(_15940_),
    .X(_15941_));
 sg13g2_o21ai_1 _23285_ (.B1(_14102_),
    .Y(_15942_),
    .A1(_14033_),
    .A2(_14073_));
 sg13g2_nand2b_1 _23286_ (.Y(_15943_),
    .B(_15942_),
    .A_N(_14086_));
 sg13g2_xor2_1 _23287_ (.B(_15942_),
    .A(_14086_),
    .X(_15944_));
 sg13g2_o21ai_1 _23288_ (.B1(_15941_),
    .Y(_15945_),
    .A1(net3829),
    .A2(_15944_));
 sg13g2_nand2_1 _23289_ (.Y(_15946_),
    .A(net3405),
    .B(_15945_));
 sg13g2_xnor2_1 _23290_ (.Y(_15947_),
    .A(net3405),
    .B(_15945_));
 sg13g2_a21o_1 _23291_ (.A2(_15931_),
    .A1(net3399),
    .B1(_15914_),
    .X(_15948_));
 sg13g2_nor2_1 _23292_ (.A(_15915_),
    .B(_15932_),
    .Y(_15949_));
 sg13g2_a21o_1 _23293_ (.A2(_15949_),
    .A1(_15918_),
    .B1(_15948_),
    .X(_15950_));
 sg13g2_nand2b_1 _23294_ (.Y(_15951_),
    .B(_15950_),
    .A_N(_15947_));
 sg13g2_xnor2_1 _23295_ (.Y(_15952_),
    .A(_15947_),
    .B(_15950_));
 sg13g2_nor2_1 _23296_ (.A(net4315),
    .B(_15945_),
    .Y(_15953_));
 sg13g2_o21ai_1 _23297_ (.B1(net3881),
    .Y(_15954_),
    .A1(net4294),
    .A2(_15952_));
 sg13g2_nand2_1 _23298_ (.Y(_15955_),
    .A(net2134),
    .B(net3922));
 sg13g2_o21ai_1 _23299_ (.B1(_15955_),
    .Y(_00296_),
    .A1(_15953_),
    .A2(_15954_));
 sg13g2_nand2_1 _23300_ (.Y(_15956_),
    .A(net2911),
    .B(net3922));
 sg13g2_a21oi_1 _23301_ (.A1(net4531),
    .A2(\u_inv.d_next[21] ),
    .Y(_15957_),
    .B1(net3751));
 sg13g2_a21oi_1 _23302_ (.A1(_14086_),
    .A2(_15938_),
    .Y(_15958_),
    .B1(_14085_));
 sg13g2_xnor2_1 _23303_ (.Y(_15959_),
    .A(_14084_),
    .B(_15958_));
 sg13g2_nand2_1 _23304_ (.Y(_15960_),
    .A(net4644),
    .B(_15959_));
 sg13g2_nand2_1 _23305_ (.Y(_15961_),
    .A(_14095_),
    .B(_15943_));
 sg13g2_or2_1 _23306_ (.X(_15962_),
    .B(_15961_),
    .A(_14084_));
 sg13g2_a21oi_1 _23307_ (.A1(_14084_),
    .A2(_15961_),
    .Y(_15963_),
    .B1(net3829));
 sg13g2_a22oi_1 _23308_ (.Y(_15964_),
    .B1(_15962_),
    .B2(_15963_),
    .A2(_15960_),
    .A1(_15957_));
 sg13g2_nor2_1 _23309_ (.A(net3405),
    .B(_15964_),
    .Y(_15965_));
 sg13g2_xnor2_1 _23310_ (.Y(_15966_),
    .A(net3405),
    .B(_15964_));
 sg13g2_nand2_1 _23311_ (.Y(_15967_),
    .A(_15946_),
    .B(_15951_));
 sg13g2_xnor2_1 _23312_ (.Y(_15968_),
    .A(_15966_),
    .B(_15967_));
 sg13g2_nor2_1 _23313_ (.A(net4294),
    .B(_15968_),
    .Y(_15969_));
 sg13g2_o21ai_1 _23314_ (.B1(net3881),
    .Y(_15970_),
    .A1(net4315),
    .A2(_15964_));
 sg13g2_o21ai_1 _23315_ (.B1(_15956_),
    .Y(_00297_),
    .A1(_15969_),
    .A2(_15970_));
 sg13g2_a21oi_1 _23316_ (.A1(_14087_),
    .A2(_15942_),
    .Y(_15971_),
    .B1(_14096_));
 sg13g2_xnor2_1 _23317_ (.Y(_15972_),
    .A(_14080_),
    .B(_15971_));
 sg13g2_a21oi_1 _23318_ (.A1(_15559_),
    .A2(_15938_),
    .Y(_15973_),
    .B1(_15564_));
 sg13g2_a21oi_1 _23319_ (.A1(_14081_),
    .A2(_15973_),
    .Y(_15974_),
    .B1(net4533));
 sg13g2_o21ai_1 _23320_ (.B1(_15974_),
    .Y(_15975_),
    .A1(_14081_),
    .A2(_15973_));
 sg13g2_a21oi_1 _23321_ (.A1(net4533),
    .A2(\u_inv.d_next[22] ),
    .Y(_15976_),
    .B1(net3746));
 sg13g2_a22oi_1 _23322_ (.Y(_15977_),
    .B1(_15975_),
    .B2(_15976_),
    .A2(_15972_),
    .A1(net3746));
 sg13g2_xnor2_1 _23323_ (.Y(_15978_),
    .A(net3405),
    .B(_15977_));
 sg13g2_o21ai_1 _23324_ (.B1(net3406),
    .Y(_15979_),
    .A1(_15945_),
    .A2(_15964_));
 sg13g2_a21oi_1 _23325_ (.A1(_15951_),
    .A2(_15979_),
    .Y(_15980_),
    .B1(_15965_));
 sg13g2_nor2b_1 _23326_ (.A(_15978_),
    .B_N(_15980_),
    .Y(_15981_));
 sg13g2_xor2_1 _23327_ (.B(_15980_),
    .A(_15978_),
    .X(_15982_));
 sg13g2_o21ai_1 _23328_ (.B1(net3881),
    .Y(_15983_),
    .A1(net4315),
    .A2(_15977_));
 sg13g2_a21oi_1 _23329_ (.A1(net4315),
    .A2(_15982_),
    .Y(_15984_),
    .B1(_15983_));
 sg13g2_a21o_1 _23330_ (.A2(net3922),
    .A1(net3085),
    .B1(_15984_),
    .X(_00298_));
 sg13g2_nand2_1 _23331_ (.Y(_15985_),
    .A(net2840),
    .B(net3925));
 sg13g2_a21oi_1 _23332_ (.A1(net4533),
    .A2(\u_inv.d_next[23] ),
    .Y(_15986_),
    .B1(net3749));
 sg13g2_o21ai_1 _23333_ (.B1(_14078_),
    .Y(_15987_),
    .A1(_14081_),
    .A2(_15973_));
 sg13g2_xnor2_1 _23334_ (.Y(_15988_),
    .A(_14076_),
    .B(_15987_));
 sg13g2_nand2_1 _23335_ (.Y(_15989_),
    .A(net4646),
    .B(_15988_));
 sg13g2_o21ai_1 _23336_ (.B1(_14092_),
    .Y(_15990_),
    .A1(_14080_),
    .A2(_15971_));
 sg13g2_o21ai_1 _23337_ (.B1(net3749),
    .Y(_15991_),
    .A1(_14077_),
    .A2(_15990_));
 sg13g2_a21oi_1 _23338_ (.A1(_14077_),
    .A2(_15990_),
    .Y(_15992_),
    .B1(_15991_));
 sg13g2_a21oi_2 _23339_ (.B1(_15992_),
    .Y(_15993_),
    .A2(_15989_),
    .A1(_15986_));
 sg13g2_xnor2_1 _23340_ (.Y(_15994_),
    .A(net3405),
    .B(_15993_));
 sg13g2_a21o_1 _23341_ (.A2(_15977_),
    .A1(net3405),
    .B1(_15981_),
    .X(_15995_));
 sg13g2_o21ai_1 _23342_ (.B1(net4315),
    .Y(_15996_),
    .A1(_15994_),
    .A2(_15995_));
 sg13g2_a21oi_1 _23343_ (.A1(_15994_),
    .A2(_15995_),
    .Y(_15997_),
    .B1(_15996_));
 sg13g2_o21ai_1 _23344_ (.B1(net3881),
    .Y(_15998_),
    .A1(net4315),
    .A2(_15993_));
 sg13g2_o21ai_1 _23345_ (.B1(_15985_),
    .Y(_00299_),
    .A1(_15997_),
    .A2(_15998_));
 sg13g2_a21oi_1 _23346_ (.A1(_14088_),
    .A2(_15942_),
    .Y(_15999_),
    .B1(_14103_));
 sg13g2_a21o_1 _23347_ (.A2(_15942_),
    .A1(_14088_),
    .B1(_14103_),
    .X(_16000_));
 sg13g2_xnor2_1 _23348_ (.Y(_16001_),
    .A(_14058_),
    .B(_16000_));
 sg13g2_o21ai_1 _23349_ (.B1(_15561_),
    .Y(_16002_),
    .A1(_15552_),
    .A2(_15937_));
 sg13g2_and2_1 _23350_ (.A(_15567_),
    .B(_16002_),
    .X(_16003_));
 sg13g2_a21oi_1 _23351_ (.A1(_14058_),
    .A2(_16003_),
    .Y(_16004_),
    .B1(net4533));
 sg13g2_o21ai_1 _23352_ (.B1(_16004_),
    .Y(_16005_),
    .A1(_14058_),
    .A2(_16003_));
 sg13g2_a21oi_1 _23353_ (.A1(net4533),
    .A2(\u_inv.d_next[24] ),
    .Y(_16006_),
    .B1(net3749));
 sg13g2_a22oi_1 _23354_ (.Y(_16007_),
    .B1(_16005_),
    .B2(_16006_),
    .A2(_16001_),
    .A1(net3749));
 sg13g2_nand2_1 _23355_ (.Y(_16008_),
    .A(net3401),
    .B(_16007_));
 sg13g2_xnor2_1 _23356_ (.Y(_16009_),
    .A(net3406),
    .B(_16007_));
 sg13g2_nor4_1 _23357_ (.A(_15947_),
    .B(_15966_),
    .C(_15978_),
    .D(_15994_),
    .Y(_16010_));
 sg13g2_nor3_1 _23358_ (.A(_15915_),
    .B(_15916_),
    .C(_15932_),
    .Y(_16011_));
 sg13g2_o21ai_1 _23359_ (.B1(_16010_),
    .Y(_16012_),
    .A1(_15948_),
    .A2(_16011_));
 sg13g2_o21ai_1 _23360_ (.B1(net3405),
    .Y(_16013_),
    .A1(_15977_),
    .A2(_15993_));
 sg13g2_nor3_1 _23361_ (.A(_15978_),
    .B(_15979_),
    .C(_15994_),
    .Y(_16014_));
 sg13g2_nor2b_1 _23362_ (.A(_16014_),
    .B_N(_16013_),
    .Y(_16015_));
 sg13g2_nand4_1 _23363_ (.B(_15899_),
    .C(_15949_),
    .A(_15879_),
    .Y(_16016_),
    .D(_16010_));
 sg13g2_nand2b_1 _23364_ (.Y(_16017_),
    .B(_15886_),
    .A_N(_16016_));
 sg13g2_nand3_1 _23365_ (.B(_16015_),
    .C(_16017_),
    .A(_16012_),
    .Y(_16018_));
 sg13g2_nand2b_1 _23366_ (.Y(_16019_),
    .B(_16018_),
    .A_N(_16009_));
 sg13g2_xor2_1 _23367_ (.B(_16018_),
    .A(_16009_),
    .X(_16020_));
 sg13g2_o21ai_1 _23368_ (.B1(net3880),
    .Y(_16021_),
    .A1(net4315),
    .A2(_16007_));
 sg13g2_a21oi_1 _23369_ (.A1(net4315),
    .A2(_16020_),
    .Y(_16022_),
    .B1(_16021_));
 sg13g2_a21o_1 _23370_ (.A2(net3924),
    .A1(net3258),
    .B1(_16022_),
    .X(_00300_));
 sg13g2_a21oi_1 _23371_ (.A1(net4533),
    .A2(\u_inv.d_next[25] ),
    .Y(_16023_),
    .B1(net3749));
 sg13g2_o21ai_1 _23372_ (.B1(_14057_),
    .Y(_16024_),
    .A1(_14058_),
    .A2(_16003_));
 sg13g2_xnor2_1 _23373_ (.Y(_16025_),
    .A(_14056_),
    .B(_16024_));
 sg13g2_nand2_1 _23374_ (.Y(_16026_),
    .A(net4646),
    .B(_16025_));
 sg13g2_a21oi_1 _23375_ (.A1(_14058_),
    .A2(_16000_),
    .Y(_16027_),
    .B1(_14113_));
 sg13g2_o21ai_1 _23376_ (.B1(net3749),
    .Y(_16028_),
    .A1(_14056_),
    .A2(_16027_));
 sg13g2_a21oi_1 _23377_ (.A1(_14056_),
    .A2(_16027_),
    .Y(_16029_),
    .B1(_16028_));
 sg13g2_a21oi_2 _23378_ (.B1(_16029_),
    .Y(_16030_),
    .A2(_16026_),
    .A1(_16023_));
 sg13g2_xnor2_1 _23379_ (.Y(_16031_),
    .A(net3401),
    .B(_16030_));
 sg13g2_and2_1 _23380_ (.A(_16008_),
    .B(_16019_),
    .X(_16032_));
 sg13g2_xnor2_1 _23381_ (.Y(_16033_),
    .A(_16031_),
    .B(_16032_));
 sg13g2_o21ai_1 _23382_ (.B1(net3879),
    .Y(_16034_),
    .A1(net4311),
    .A2(_16030_));
 sg13g2_a21oi_1 _23383_ (.A1(net4311),
    .A2(_16033_),
    .Y(_16035_),
    .B1(_16034_));
 sg13g2_a21o_1 _23384_ (.A2(net3924),
    .A1(net3115),
    .B1(_16035_),
    .X(_00301_));
 sg13g2_o21ai_1 _23385_ (.B1(net3406),
    .Y(_16036_),
    .A1(_16007_),
    .A2(_16030_));
 sg13g2_o21ai_1 _23386_ (.B1(_16036_),
    .Y(_16037_),
    .A1(_16019_),
    .A2(_16031_));
 sg13g2_o21ai_1 _23387_ (.B1(_14114_),
    .Y(_16038_),
    .A1(_14059_),
    .A2(_15999_));
 sg13g2_xnor2_1 _23388_ (.Y(_16039_),
    .A(_14052_),
    .B(_16038_));
 sg13g2_a21oi_1 _23389_ (.A1(_15567_),
    .A2(_16002_),
    .Y(_16040_),
    .B1(_15556_));
 sg13g2_nor3_1 _23390_ (.A(_14051_),
    .B(_15574_),
    .C(_16040_),
    .Y(_16041_));
 sg13g2_o21ai_1 _23391_ (.B1(_14051_),
    .Y(_16042_),
    .A1(_15574_),
    .A2(_16040_));
 sg13g2_nand3b_1 _23392_ (.B(_16042_),
    .C(net4646),
    .Y(_16043_),
    .A_N(_16041_));
 sg13g2_a21oi_1 _23393_ (.A1(net4534),
    .A2(\u_inv.d_next[26] ),
    .Y(_16044_),
    .B1(net3749));
 sg13g2_a22oi_1 _23394_ (.Y(_16045_),
    .B1(_16043_),
    .B2(_16044_),
    .A2(_16039_),
    .A1(net3749));
 sg13g2_xnor2_1 _23395_ (.Y(_16046_),
    .A(net3407),
    .B(_16045_));
 sg13g2_nor2b_1 _23396_ (.A(_16046_),
    .B_N(_16037_),
    .Y(_16047_));
 sg13g2_xnor2_1 _23397_ (.Y(_16048_),
    .A(_16037_),
    .B(_16046_));
 sg13g2_nor2_1 _23398_ (.A(net4316),
    .B(_16045_),
    .Y(_16049_));
 sg13g2_o21ai_1 _23399_ (.B1(net3879),
    .Y(_16050_),
    .A1(net4291),
    .A2(_16048_));
 sg13g2_nand2_1 _23400_ (.Y(_16051_),
    .A(net2465),
    .B(net3925));
 sg13g2_o21ai_1 _23401_ (.B1(_16051_),
    .Y(_00302_),
    .A1(_16049_),
    .A2(_16050_));
 sg13g2_a21oi_1 _23402_ (.A1(net3407),
    .A2(_16045_),
    .Y(_16052_),
    .B1(_16047_));
 sg13g2_a21oi_1 _23403_ (.A1(net4534),
    .A2(\u_inv.d_next[27] ),
    .Y(_16053_),
    .B1(net3750));
 sg13g2_a21o_1 _23404_ (.A2(_16042_),
    .A1(_14050_),
    .B1(_14048_),
    .X(_16054_));
 sg13g2_nand3_1 _23405_ (.B(_14050_),
    .C(_16042_),
    .A(_14048_),
    .Y(_16055_));
 sg13g2_nand3_1 _23406_ (.B(_16054_),
    .C(_16055_),
    .A(net4646),
    .Y(_16056_));
 sg13g2_a21oi_1 _23407_ (.A1(_14052_),
    .A2(_16038_),
    .Y(_16057_),
    .B1(_14115_));
 sg13g2_or2_1 _23408_ (.X(_16058_),
    .B(_16057_),
    .A(_14048_));
 sg13g2_a21oi_1 _23409_ (.A1(_14048_),
    .A2(_16057_),
    .Y(_16059_),
    .B1(net3830));
 sg13g2_a22oi_1 _23410_ (.Y(_16060_),
    .B1(_16058_),
    .B2(_16059_),
    .A2(_16056_),
    .A1(_16053_));
 sg13g2_xnor2_1 _23411_ (.Y(_16061_),
    .A(net3407),
    .B(_16060_));
 sg13g2_xnor2_1 _23412_ (.Y(_16062_),
    .A(_16052_),
    .B(_16061_));
 sg13g2_o21ai_1 _23413_ (.B1(net3880),
    .Y(_16063_),
    .A1(net4317),
    .A2(_16060_));
 sg13g2_a21oi_1 _23414_ (.A1(net4317),
    .A2(_16062_),
    .Y(_16064_),
    .B1(_16063_));
 sg13g2_a21o_1 _23415_ (.A2(net3925),
    .A1(net3143),
    .B1(_16064_),
    .X(_00303_));
 sg13g2_o21ai_1 _23416_ (.B1(_14117_),
    .Y(_16065_),
    .A1(_14060_),
    .A2(_15999_));
 sg13g2_xnor2_1 _23417_ (.Y(_16066_),
    .A(_14042_),
    .B(_16065_));
 sg13g2_a21oi_1 _23418_ (.A1(_15567_),
    .A2(_16002_),
    .Y(_16067_),
    .B1(_15557_));
 sg13g2_or3_1 _23419_ (.A(_14043_),
    .B(_15576_),
    .C(_16067_),
    .X(_16068_));
 sg13g2_o21ai_1 _23420_ (.B1(_14043_),
    .Y(_16069_),
    .A1(_15576_),
    .A2(_16067_));
 sg13g2_nand3_1 _23421_ (.B(_16068_),
    .C(_16069_),
    .A(net4645),
    .Y(_16070_));
 sg13g2_a21oi_1 _23422_ (.A1(net4534),
    .A2(\u_inv.d_next[28] ),
    .Y(_16071_),
    .B1(net3750));
 sg13g2_a22oi_1 _23423_ (.Y(_16072_),
    .B1(_16070_),
    .B2(_16071_),
    .A2(_16066_),
    .A1(net3750));
 sg13g2_nand2_1 _23424_ (.Y(_16073_),
    .A(net3407),
    .B(_16072_));
 sg13g2_xnor2_1 _23425_ (.Y(_16074_),
    .A(net3407),
    .B(_16072_));
 sg13g2_o21ai_1 _23426_ (.B1(net3407),
    .Y(_16075_),
    .A1(_16045_),
    .A2(_16060_));
 sg13g2_nor2_1 _23427_ (.A(_16046_),
    .B(_16061_),
    .Y(_16076_));
 sg13g2_nand2_1 _23428_ (.Y(_16077_),
    .A(_16037_),
    .B(_16076_));
 sg13g2_nand2_1 _23429_ (.Y(_16078_),
    .A(_16075_),
    .B(_16077_));
 sg13g2_nand2b_1 _23430_ (.Y(_16079_),
    .B(_16078_),
    .A_N(_16074_));
 sg13g2_xor2_1 _23431_ (.B(_16078_),
    .A(_16074_),
    .X(_16080_));
 sg13g2_o21ai_1 _23432_ (.B1(net3880),
    .Y(_16081_),
    .A1(net4316),
    .A2(_16072_));
 sg13g2_a21oi_1 _23433_ (.A1(net4316),
    .A2(_16080_),
    .Y(_16082_),
    .B1(_16081_));
 sg13g2_a21o_1 _23434_ (.A2(net3924),
    .A1(net2780),
    .B1(_16082_),
    .X(_00304_));
 sg13g2_a21oi_1 _23435_ (.A1(net4533),
    .A2(\u_inv.d_next[29] ),
    .Y(_16083_),
    .B1(net3750));
 sg13g2_nand3_1 _23436_ (.B(_14041_),
    .C(_16069_),
    .A(_14040_),
    .Y(_16084_));
 sg13g2_a21o_1 _23437_ (.A2(_16069_),
    .A1(_14041_),
    .B1(_14040_),
    .X(_16085_));
 sg13g2_nand3_1 _23438_ (.B(_16084_),
    .C(_16085_),
    .A(net4645),
    .Y(_16086_));
 sg13g2_a21oi_1 _23439_ (.A1(_14042_),
    .A2(_16065_),
    .Y(_16087_),
    .B1(_14106_));
 sg13g2_or2_1 _23440_ (.X(_16088_),
    .B(_16087_),
    .A(_14040_));
 sg13g2_a21oi_1 _23441_ (.A1(_14040_),
    .A2(_16087_),
    .Y(_16089_),
    .B1(net3829));
 sg13g2_a22oi_1 _23442_ (.Y(_16090_),
    .B1(_16088_),
    .B2(_16089_),
    .A2(_16086_),
    .A1(_16083_));
 sg13g2_nor2_1 _23443_ (.A(net3407),
    .B(_16090_),
    .Y(_16091_));
 sg13g2_xnor2_1 _23444_ (.Y(_16092_),
    .A(net3407),
    .B(_16090_));
 sg13g2_nand2_1 _23445_ (.Y(_16093_),
    .A(_16073_),
    .B(_16079_));
 sg13g2_xor2_1 _23446_ (.B(_16093_),
    .A(_16092_),
    .X(_16094_));
 sg13g2_o21ai_1 _23447_ (.B1(net3880),
    .Y(_16095_),
    .A1(net4316),
    .A2(_16090_));
 sg13g2_a21oi_1 _23448_ (.A1(net4316),
    .A2(_16094_),
    .Y(_16096_),
    .B1(_16095_));
 sg13g2_a21o_1 _23449_ (.A2(net3924),
    .A1(net2605),
    .B1(_16096_),
    .X(_00305_));
 sg13g2_a21oi_1 _23450_ (.A1(_14044_),
    .A2(_16065_),
    .Y(_16097_),
    .B1(_14108_));
 sg13g2_xnor2_1 _23451_ (.Y(_16098_),
    .A(_14037_),
    .B(_16097_));
 sg13g2_o21ai_1 _23452_ (.B1(_15553_),
    .Y(_16099_),
    .A1(_15576_),
    .A2(_16067_));
 sg13g2_nand3_1 _23453_ (.B(_15569_),
    .C(_16099_),
    .A(_14038_),
    .Y(_16100_));
 sg13g2_a21o_1 _23454_ (.A2(_16099_),
    .A1(_15569_),
    .B1(_14038_),
    .X(_16101_));
 sg13g2_nand3_1 _23455_ (.B(_16100_),
    .C(_16101_),
    .A(net4646),
    .Y(_16102_));
 sg13g2_a21oi_1 _23456_ (.A1(net4533),
    .A2(\u_inv.d_next[30] ),
    .Y(_16103_),
    .B1(net3750));
 sg13g2_a22oi_1 _23457_ (.Y(_16104_),
    .B1(_16102_),
    .B2(_16103_),
    .A2(_16098_),
    .A1(net3750));
 sg13g2_and2_1 _23458_ (.A(net3404),
    .B(_16104_),
    .X(_16105_));
 sg13g2_xnor2_1 _23459_ (.Y(_16106_),
    .A(net3471),
    .B(_16104_));
 sg13g2_o21ai_1 _23460_ (.B1(net3408),
    .Y(_16107_),
    .A1(_16072_),
    .A2(_16090_));
 sg13g2_a21oi_1 _23461_ (.A1(_16079_),
    .A2(_16107_),
    .Y(_16108_),
    .B1(_16091_));
 sg13g2_xnor2_1 _23462_ (.Y(_16109_),
    .A(_16106_),
    .B(_16108_));
 sg13g2_a21oi_1 _23463_ (.A1(net4316),
    .A2(_16109_),
    .Y(_16110_),
    .B1(net4233));
 sg13g2_o21ai_1 _23464_ (.B1(_16110_),
    .Y(_16111_),
    .A1(net4316),
    .A2(_16104_));
 sg13g2_o21ai_1 _23465_ (.B1(_16111_),
    .Y(_00306_),
    .A1(_10618_),
    .A2(net4013));
 sg13g2_a21oi_1 _23466_ (.A1(net4534),
    .A2(\u_inv.d_next[31] ),
    .Y(_16112_),
    .B1(net3750));
 sg13g2_nand3_1 _23467_ (.B(_14036_),
    .C(_16101_),
    .A(_14034_),
    .Y(_16113_));
 sg13g2_a21o_1 _23468_ (.A2(_16101_),
    .A1(_14036_),
    .B1(_14034_),
    .X(_16114_));
 sg13g2_nand3_1 _23469_ (.B(_16113_),
    .C(_16114_),
    .A(net4646),
    .Y(_16115_));
 sg13g2_o21ai_1 _23470_ (.B1(_14109_),
    .Y(_16116_),
    .A1(_14037_),
    .A2(_16097_));
 sg13g2_or2_1 _23471_ (.X(_16117_),
    .B(_16116_),
    .A(_14035_));
 sg13g2_a21oi_1 _23472_ (.A1(_14035_),
    .A2(_16116_),
    .Y(_16118_),
    .B1(net3829));
 sg13g2_a22oi_1 _23473_ (.Y(_16119_),
    .B1(_16117_),
    .B2(_16118_),
    .A2(_16115_),
    .A1(_16112_));
 sg13g2_xnor2_1 _23474_ (.Y(_16120_),
    .A(net3471),
    .B(_16119_));
 sg13g2_a21o_1 _23475_ (.A2(_16108_),
    .A1(_16106_),
    .B1(_16105_),
    .X(_16121_));
 sg13g2_xnor2_1 _23476_ (.Y(_16122_),
    .A(_16120_),
    .B(_16121_));
 sg13g2_o21ai_1 _23477_ (.B1(net3879),
    .Y(_16123_),
    .A1(net4314),
    .A2(_16119_));
 sg13g2_a21oi_1 _23478_ (.A1(net4314),
    .A2(_16122_),
    .Y(_16124_),
    .B1(_16123_));
 sg13g2_a21o_1 _23479_ (.A2(net3924),
    .A1(net3281),
    .B1(_16124_),
    .X(_00307_));
 sg13g2_nand2_1 _23480_ (.Y(_16125_),
    .A(_16106_),
    .B(_16120_));
 sg13g2_nor2_1 _23481_ (.A(_16074_),
    .B(_16092_),
    .Y(_16126_));
 sg13g2_nand3_1 _23482_ (.B(_16120_),
    .C(_16126_),
    .A(_16106_),
    .Y(_16127_));
 sg13g2_nor4_1 _23483_ (.A(_16009_),
    .B(_16031_),
    .C(_16046_),
    .D(_16061_),
    .Y(_16128_));
 sg13g2_nand4_1 _23484_ (.B(_16120_),
    .C(_16126_),
    .A(_16106_),
    .Y(_16129_),
    .D(_16128_));
 sg13g2_or2_1 _23485_ (.X(_16130_),
    .B(_16129_),
    .A(_16016_));
 sg13g2_a21oi_2 _23486_ (.B1(_16130_),
    .Y(_16131_),
    .A2(_15885_),
    .A1(_15883_));
 sg13g2_a21oi_1 _23487_ (.A1(_16012_),
    .A2(_16015_),
    .Y(_16132_),
    .B1(_16129_));
 sg13g2_o21ai_1 _23488_ (.B1(net3408),
    .Y(_16133_),
    .A1(_16104_),
    .A2(_16119_));
 sg13g2_o21ai_1 _23489_ (.B1(_16133_),
    .Y(_16134_),
    .A1(_16107_),
    .A2(_16125_));
 sg13g2_nand2b_1 _23490_ (.Y(_16135_),
    .B(_16076_),
    .A_N(_16036_));
 sg13g2_a21oi_1 _23491_ (.A1(_16075_),
    .A2(_16135_),
    .Y(_16136_),
    .B1(_16127_));
 sg13g2_or3_1 _23492_ (.A(_16132_),
    .B(_16134_),
    .C(_16136_),
    .X(_16137_));
 sg13g2_nor2_2 _23493_ (.A(_16131_),
    .B(_16137_),
    .Y(_16138_));
 sg13g2_xnor2_1 _23494_ (.Y(_16139_),
    .A(_14232_),
    .B(_15616_));
 sg13g2_o21ai_1 _23495_ (.B1(net3835),
    .Y(_16140_),
    .A1(net4658),
    .A2(\u_inv.d_next[32] ));
 sg13g2_a21oi_1 _23496_ (.A1(net4658),
    .A2(_16139_),
    .Y(_16141_),
    .B1(_16140_));
 sg13g2_nand2_1 _23497_ (.Y(_16142_),
    .A(_14121_),
    .B(_14232_));
 sg13g2_xnor2_1 _23498_ (.Y(_16143_),
    .A(_14121_),
    .B(_14231_));
 sg13g2_a21oi_2 _23499_ (.B1(_16141_),
    .Y(_16144_),
    .A2(_16143_),
    .A1(net3758));
 sg13g2_inv_1 _23500_ (.Y(_16145_),
    .A(_16144_));
 sg13g2_xnor2_1 _23501_ (.Y(_16146_),
    .A(net3472),
    .B(_16144_));
 sg13g2_o21ai_1 _23502_ (.B1(_16146_),
    .Y(_16147_),
    .A1(_16131_),
    .A2(_16137_));
 sg13g2_xor2_1 _23503_ (.B(_16146_),
    .A(_16138_),
    .X(_16148_));
 sg13g2_nand2_1 _23504_ (.Y(_16149_),
    .A(net4292),
    .B(_16144_));
 sg13g2_a21oi_1 _23505_ (.A1(net4319),
    .A2(_16148_),
    .Y(_16150_),
    .B1(net4234));
 sg13g2_a22oi_1 _23506_ (.Y(_16151_),
    .B1(_16149_),
    .B2(_16150_),
    .A2(net3933),
    .A1(net3303));
 sg13g2_inv_1 _23507_ (.Y(_00308_),
    .A(_16151_));
 sg13g2_o21ai_1 _23508_ (.B1(_16147_),
    .Y(_16152_),
    .A1(net3411),
    .A2(_16144_));
 sg13g2_a21o_1 _23509_ (.A2(_15617_),
    .A1(_14231_),
    .B1(_14230_),
    .X(_16153_));
 sg13g2_xnor2_1 _23510_ (.Y(_16154_),
    .A(_14228_),
    .B(_16153_));
 sg13g2_nand2_1 _23511_ (.Y(_16155_),
    .A(net4658),
    .B(_16154_));
 sg13g2_a21oi_1 _23512_ (.A1(net4542),
    .A2(\u_inv.d_next[33] ),
    .Y(_16156_),
    .B1(net3758));
 sg13g2_nand3_1 _23513_ (.B(_14240_),
    .C(_16142_),
    .A(_14228_),
    .Y(_16157_));
 sg13g2_a21oi_1 _23514_ (.A1(_14240_),
    .A2(_16142_),
    .Y(_16158_),
    .B1(_14228_));
 sg13g2_nor2_1 _23515_ (.A(net3835),
    .B(_16158_),
    .Y(_16159_));
 sg13g2_a22oi_1 _23516_ (.Y(_16160_),
    .B1(_16157_),
    .B2(_16159_),
    .A2(_16156_),
    .A1(_16155_));
 sg13g2_xnor2_1 _23517_ (.Y(_16161_),
    .A(net3472),
    .B(_16160_));
 sg13g2_xnor2_1 _23518_ (.Y(_16162_),
    .A(_16152_),
    .B(_16161_));
 sg13g2_o21ai_1 _23519_ (.B1(net3888),
    .Y(_16163_),
    .A1(net4323),
    .A2(_16160_));
 sg13g2_a21oi_1 _23520_ (.A1(net4323),
    .A2(_16162_),
    .Y(_16164_),
    .B1(_16163_));
 sg13g2_a21o_1 _23521_ (.A2(net3933),
    .A1(net3104),
    .B1(_16164_),
    .X(_00309_));
 sg13g2_a21oi_1 _23522_ (.A1(_14091_),
    .A2(_14119_),
    .Y(_16165_),
    .B1(_14234_));
 sg13g2_nor3_1 _23523_ (.A(_14224_),
    .B(_14241_),
    .C(_16165_),
    .Y(_16166_));
 sg13g2_o21ai_1 _23524_ (.B1(_14224_),
    .Y(_16167_),
    .A1(_14241_),
    .A2(_16165_));
 sg13g2_nor2b_1 _23525_ (.A(_16166_),
    .B_N(_16167_),
    .Y(_16168_));
 sg13g2_a21oi_1 _23526_ (.A1(_14229_),
    .A2(_16153_),
    .Y(_16169_),
    .B1(_15482_));
 sg13g2_xnor2_1 _23527_ (.Y(_16170_),
    .A(_14224_),
    .B(_16169_));
 sg13g2_a21oi_1 _23528_ (.A1(net4542),
    .A2(\u_inv.d_next[34] ),
    .Y(_16171_),
    .B1(net3758));
 sg13g2_o21ai_1 _23529_ (.B1(_16171_),
    .Y(_16172_),
    .A1(net4542),
    .A2(_16170_));
 sg13g2_o21ai_1 _23530_ (.B1(_16172_),
    .Y(_16173_),
    .A1(net3835),
    .A2(_16168_));
 sg13g2_a21oi_1 _23531_ (.A1(net3491),
    .A2(net3490),
    .Y(_16174_),
    .B1(_16173_));
 sg13g2_and3_1 _23532_ (.X(_16175_),
    .A(net3491),
    .B(net3490),
    .C(_16173_));
 sg13g2_or2_1 _23533_ (.X(_16176_),
    .B(_16175_),
    .A(_16174_));
 sg13g2_o21ai_1 _23534_ (.B1(_16160_),
    .Y(_16177_),
    .A1(net3411),
    .A2(_16145_));
 sg13g2_nand2b_2 _23535_ (.Y(_16178_),
    .B(_16161_),
    .A_N(_16147_));
 sg13g2_a21o_1 _23536_ (.A2(_16178_),
    .A1(_16177_),
    .B1(_16176_),
    .X(_16179_));
 sg13g2_nand3_1 _23537_ (.B(_16177_),
    .C(_16178_),
    .A(_16176_),
    .Y(_16180_));
 sg13g2_a21oi_1 _23538_ (.A1(_16179_),
    .A2(_16180_),
    .Y(_16181_),
    .B1(net4292));
 sg13g2_a21o_1 _23539_ (.A2(_16173_),
    .A1(net4292),
    .B1(net4234),
    .X(_16182_));
 sg13g2_nand2_1 _23540_ (.Y(_16183_),
    .A(net2864),
    .B(net3933));
 sg13g2_o21ai_1 _23541_ (.B1(_16183_),
    .Y(_00310_),
    .A1(_16181_),
    .A2(_16182_));
 sg13g2_nand2_1 _23542_ (.Y(_16184_),
    .A(net2889),
    .B(net3933));
 sg13g2_nand2b_1 _23543_ (.Y(_16185_),
    .B(net3835),
    .A_N(\u_inv.d_next[35] ));
 sg13g2_and2_1 _23544_ (.A(net3726),
    .B(_16185_),
    .X(_16186_));
 sg13g2_o21ai_1 _23545_ (.B1(_14222_),
    .Y(_16187_),
    .A1(_14224_),
    .A2(_16169_));
 sg13g2_xnor2_1 _23546_ (.Y(_16188_),
    .A(_14221_),
    .B(_16187_));
 sg13g2_a22oi_1 _23547_ (.Y(_16189_),
    .B1(_16188_),
    .B2(net4657),
    .A2(_16185_),
    .A1(net3726));
 sg13g2_a21o_1 _23548_ (.A2(_16188_),
    .A1(net4657),
    .B1(_16186_),
    .X(_16190_));
 sg13g2_a21o_1 _23549_ (.A2(_16167_),
    .A1(_14242_),
    .B1(_14221_),
    .X(_16191_));
 sg13g2_nand3_1 _23550_ (.B(_14242_),
    .C(_16167_),
    .A(_14221_),
    .Y(_16192_));
 sg13g2_and2_1 _23551_ (.A(net3755),
    .B(_16192_),
    .X(_16193_));
 sg13g2_nand3_1 _23552_ (.B(_16191_),
    .C(_16192_),
    .A(net3755),
    .Y(_16194_));
 sg13g2_and2_1 _23553_ (.A(_16190_),
    .B(_16194_),
    .X(_16195_));
 sg13g2_a221oi_1 _23554_ (.B2(_16193_),
    .C1(_16189_),
    .B1(_16191_),
    .A1(net3491),
    .Y(_16196_),
    .A2(net3490));
 sg13g2_a221oi_1 _23555_ (.B2(_16194_),
    .C1(_15646_),
    .B1(_16190_),
    .A1(_13598_),
    .Y(_16197_),
    .A2(_15033_));
 sg13g2_or2_1 _23556_ (.X(_16198_),
    .B(_16197_),
    .A(_16196_));
 sg13g2_nand2b_1 _23557_ (.Y(_16199_),
    .B(_16179_),
    .A_N(_16174_));
 sg13g2_o21ai_1 _23558_ (.B1(net4319),
    .Y(_16200_),
    .A1(_16198_),
    .A2(_16199_));
 sg13g2_a21oi_1 _23559_ (.A1(_16198_),
    .A2(_16199_),
    .Y(_16201_),
    .B1(_16200_));
 sg13g2_o21ai_1 _23560_ (.B1(net3882),
    .Y(_16202_),
    .A1(net4319),
    .A2(_16195_));
 sg13g2_o21ai_1 _23561_ (.B1(_16184_),
    .Y(_00311_),
    .A1(_16201_),
    .A2(_16202_));
 sg13g2_a21oi_1 _23562_ (.A1(_15617_),
    .A2(_15618_),
    .Y(_16203_),
    .B1(_15485_));
 sg13g2_a21o_1 _23563_ (.A2(_15618_),
    .A1(_15617_),
    .B1(_15485_),
    .X(_16204_));
 sg13g2_xnor2_1 _23564_ (.Y(_16205_),
    .A(_14216_),
    .B(_16203_));
 sg13g2_nor2_1 _23565_ (.A(net4656),
    .B(\u_inv.d_next[36] ),
    .Y(_16206_));
 sg13g2_a21oi_1 _23566_ (.A1(net4656),
    .A2(_16205_),
    .Y(_16207_),
    .B1(_16206_));
 sg13g2_o21ai_1 _23567_ (.B1(_14225_),
    .Y(_16208_),
    .A1(_14241_),
    .A2(_16165_));
 sg13g2_a21oi_1 _23568_ (.A1(_14243_),
    .A2(_16208_),
    .Y(_16209_),
    .B1(_14215_));
 sg13g2_a21o_1 _23569_ (.A2(_16208_),
    .A1(_14243_),
    .B1(_14215_),
    .X(_16210_));
 sg13g2_nand3_1 _23570_ (.B(_14243_),
    .C(_16208_),
    .A(_14215_),
    .Y(_16211_));
 sg13g2_and2_1 _23571_ (.A(net3756),
    .B(_16211_),
    .X(_16212_));
 sg13g2_a22oi_1 _23572_ (.Y(_16213_),
    .B1(_16210_),
    .B2(_16212_),
    .A2(_16207_),
    .A1(net3835));
 sg13g2_a21oi_1 _23573_ (.A1(net3491),
    .A2(net3490),
    .Y(_16214_),
    .B1(_16213_));
 sg13g2_and3_1 _23574_ (.X(_16215_),
    .A(_15034_),
    .B(_15647_),
    .C(_16213_));
 sg13g2_or2_1 _23575_ (.X(_16216_),
    .B(_16215_),
    .A(_16214_));
 sg13g2_nor2_1 _23576_ (.A(_16176_),
    .B(_16198_),
    .Y(_16217_));
 sg13g2_or4_1 _23577_ (.A(_16174_),
    .B(_16175_),
    .C(_16196_),
    .D(_16197_),
    .X(_16218_));
 sg13g2_nor2_1 _23578_ (.A(_16177_),
    .B(_16218_),
    .Y(_16219_));
 sg13g2_nor2_1 _23579_ (.A(_16174_),
    .B(_16196_),
    .Y(_16220_));
 sg13g2_nor2b_1 _23580_ (.A(_16219_),
    .B_N(_16220_),
    .Y(_16221_));
 sg13g2_o21ai_1 _23581_ (.B1(_16220_),
    .Y(_16222_),
    .A1(_16177_),
    .A2(_16218_));
 sg13g2_nand2b_1 _23582_ (.Y(_16223_),
    .B(_16217_),
    .A_N(_16178_));
 sg13g2_a21oi_1 _23583_ (.A1(_16221_),
    .A2(_16223_),
    .Y(_16224_),
    .B1(_16216_));
 sg13g2_nand3_1 _23584_ (.B(_16221_),
    .C(_16223_),
    .A(_16216_),
    .Y(_16225_));
 sg13g2_nand2b_1 _23585_ (.Y(_16226_),
    .B(_16225_),
    .A_N(_16224_));
 sg13g2_nand2_1 _23586_ (.Y(_16227_),
    .A(net4292),
    .B(_16213_));
 sg13g2_a21oi_1 _23587_ (.A1(net4319),
    .A2(_16226_),
    .Y(_16228_),
    .B1(net4234));
 sg13g2_a22oi_1 _23588_ (.Y(_16229_),
    .B1(_16227_),
    .B2(_16228_),
    .A2(net3933),
    .A1(net2844));
 sg13g2_inv_1 _23589_ (.Y(_00312_),
    .A(_16229_));
 sg13g2_a21oi_1 _23590_ (.A1(net4541),
    .A2(\u_inv.d_next[37] ),
    .Y(_16230_),
    .B1(net3755));
 sg13g2_o21ai_1 _23591_ (.B1(_14214_),
    .Y(_16231_),
    .A1(_14216_),
    .A2(_16203_));
 sg13g2_a21oi_1 _23592_ (.A1(_14212_),
    .A2(_16231_),
    .Y(_16232_),
    .B1(net4541));
 sg13g2_o21ai_1 _23593_ (.B1(_16232_),
    .Y(_16233_),
    .A1(_14212_),
    .A2(_16231_));
 sg13g2_nand2_1 _23594_ (.Y(_16234_),
    .A(_16230_),
    .B(_16233_));
 sg13g2_o21ai_1 _23595_ (.B1(_14212_),
    .Y(_16235_),
    .A1(_14249_),
    .A2(_16209_));
 sg13g2_or3_1 _23596_ (.A(_14212_),
    .B(_14249_),
    .C(_16209_),
    .X(_16236_));
 sg13g2_and3_1 _23597_ (.X(_16237_),
    .A(net3755),
    .B(_16235_),
    .C(_16236_));
 sg13g2_nand3_1 _23598_ (.B(_16235_),
    .C(_16236_),
    .A(net3755),
    .Y(_16238_));
 sg13g2_and2_1 _23599_ (.A(_16234_),
    .B(_16238_),
    .X(_16239_));
 sg13g2_a221oi_1 _23600_ (.B2(_16233_),
    .C1(_16237_),
    .B1(_16230_),
    .A1(_15034_),
    .Y(_16240_),
    .A2(_15647_));
 sg13g2_a221oi_1 _23601_ (.B2(_16238_),
    .C1(_15646_),
    .B1(_16234_),
    .A1(_13598_),
    .Y(_16241_),
    .A2(_15033_));
 sg13g2_or2_1 _23602_ (.X(_16242_),
    .B(_16241_),
    .A(_16240_));
 sg13g2_nor2_1 _23603_ (.A(_16214_),
    .B(_16224_),
    .Y(_16243_));
 sg13g2_xnor2_1 _23604_ (.Y(_16244_),
    .A(_16242_),
    .B(_16243_));
 sg13g2_o21ai_1 _23605_ (.B1(net3882),
    .Y(_16245_),
    .A1(net4319),
    .A2(_16239_));
 sg13g2_a21oi_1 _23606_ (.A1(net4319),
    .A2(_16244_),
    .Y(_16246_),
    .B1(_16245_));
 sg13g2_a21o_1 _23607_ (.A2(net3932),
    .A1(net3122),
    .B1(_16246_),
    .X(_00313_));
 sg13g2_a21oi_1 _23608_ (.A1(_14243_),
    .A2(_16208_),
    .Y(_16247_),
    .B1(_14217_));
 sg13g2_o21ai_1 _23609_ (.B1(_14208_),
    .Y(_16248_),
    .A1(_14250_),
    .A2(_16247_));
 sg13g2_or3_1 _23610_ (.A(_14208_),
    .B(_14250_),
    .C(_16247_),
    .X(_16249_));
 sg13g2_nand2_1 _23611_ (.Y(_16250_),
    .A(_16248_),
    .B(_16249_));
 sg13g2_a21oi_1 _23612_ (.A1(_15479_),
    .A2(_16204_),
    .Y(_16251_),
    .B1(_15486_));
 sg13g2_nor2_1 _23613_ (.A(_14208_),
    .B(_16251_),
    .Y(_16252_));
 sg13g2_a21oi_1 _23614_ (.A1(_14208_),
    .A2(_16251_),
    .Y(_16253_),
    .B1(net4540));
 sg13g2_nand2b_1 _23615_ (.Y(_16254_),
    .B(_16253_),
    .A_N(_16252_));
 sg13g2_a21oi_1 _23616_ (.A1(net4540),
    .A2(\u_inv.d_next[38] ),
    .Y(_16255_),
    .B1(net3755));
 sg13g2_a22oi_1 _23617_ (.Y(_16256_),
    .B1(_16254_),
    .B2(_16255_),
    .A2(_16250_),
    .A1(net3758));
 sg13g2_nand2_1 _23618_ (.Y(_16257_),
    .A(net3410),
    .B(_16256_));
 sg13g2_xnor2_1 _23619_ (.Y(_16258_),
    .A(net3410),
    .B(_16256_));
 sg13g2_or2_1 _23620_ (.X(_16259_),
    .B(_16240_),
    .A(_16214_));
 sg13g2_nor2_1 _23621_ (.A(_16224_),
    .B(_16259_),
    .Y(_16260_));
 sg13g2_or2_1 _23622_ (.X(_16261_),
    .B(_16260_),
    .A(_16241_));
 sg13g2_xnor2_1 _23623_ (.Y(_16262_),
    .A(_16258_),
    .B(_16261_));
 sg13g2_o21ai_1 _23624_ (.B1(net3882),
    .Y(_16263_),
    .A1(net4318),
    .A2(_16256_));
 sg13g2_a21oi_1 _23625_ (.A1(net4318),
    .A2(_16262_),
    .Y(_16264_),
    .B1(_16263_));
 sg13g2_a21o_1 _23626_ (.A2(net3932),
    .A1(net2922),
    .B1(_16264_),
    .X(_00314_));
 sg13g2_a21oi_1 _23627_ (.A1(net4543),
    .A2(\u_inv.d_next[39] ),
    .Y(_16265_),
    .B1(net3759));
 sg13g2_nor2_1 _23628_ (.A(_14206_),
    .B(_16252_),
    .Y(_16266_));
 sg13g2_xnor2_1 _23629_ (.Y(_16267_),
    .A(_14204_),
    .B(_16266_));
 sg13g2_o21ai_1 _23630_ (.B1(_16265_),
    .Y(_16268_),
    .A1(net4543),
    .A2(_16267_));
 sg13g2_a21o_1 _23631_ (.A2(_16248_),
    .A1(_14246_),
    .B1(_14204_),
    .X(_16269_));
 sg13g2_nand3_1 _23632_ (.B(_14246_),
    .C(_16248_),
    .A(_14204_),
    .Y(_16270_));
 sg13g2_nand3_1 _23633_ (.B(_16269_),
    .C(_16270_),
    .A(net3759),
    .Y(_16271_));
 sg13g2_nand2_1 _23634_ (.Y(_16272_),
    .A(_16268_),
    .B(_16271_));
 sg13g2_and3_1 _23635_ (.X(_16273_),
    .A(net3410),
    .B(_16268_),
    .C(_16271_));
 sg13g2_a21oi_1 _23636_ (.A1(_16268_),
    .A2(_16271_),
    .Y(_16274_),
    .B1(net3411));
 sg13g2_nor2_1 _23637_ (.A(_16273_),
    .B(_16274_),
    .Y(_16275_));
 sg13g2_o21ai_1 _23638_ (.B1(_16257_),
    .Y(_16276_),
    .A1(_16258_),
    .A2(_16261_));
 sg13g2_xor2_1 _23639_ (.B(_16276_),
    .A(_16275_),
    .X(_16277_));
 sg13g2_a21oi_1 _23640_ (.A1(net4292),
    .A2(_16272_),
    .Y(_16278_),
    .B1(net4234));
 sg13g2_o21ai_1 _23641_ (.B1(_16278_),
    .Y(_16279_),
    .A1(net4293),
    .A2(_16277_));
 sg13g2_o21ai_1 _23642_ (.B1(_16279_),
    .Y(_00315_),
    .A1(_10616_),
    .A2(net4014));
 sg13g2_o21ai_1 _23643_ (.B1(_15489_),
    .Y(_16280_),
    .A1(_15616_),
    .A2(_15619_));
 sg13g2_xnor2_1 _23644_ (.Y(_16281_),
    .A(_14198_),
    .B(_16280_));
 sg13g2_nor2_1 _23645_ (.A(net4659),
    .B(\u_inv.d_next[40] ),
    .Y(_16282_));
 sg13g2_a21oi_1 _23646_ (.A1(net4659),
    .A2(_16281_),
    .Y(_16283_),
    .B1(_16282_));
 sg13g2_o21ai_1 _23647_ (.B1(_14235_),
    .Y(_16284_),
    .A1(_14090_),
    .A2(_14120_));
 sg13g2_nand2_1 _23648_ (.Y(_16285_),
    .A(_14251_),
    .B(_16284_));
 sg13g2_inv_1 _23649_ (.Y(_16286_),
    .A(_16285_));
 sg13g2_nand2_1 _23650_ (.Y(_16287_),
    .A(_14199_),
    .B(_16285_));
 sg13g2_a21oi_1 _23651_ (.A1(_14198_),
    .A2(_16286_),
    .Y(_16288_),
    .B1(net3836));
 sg13g2_a22oi_1 _23652_ (.Y(_16289_),
    .B1(_16287_),
    .B2(_16288_),
    .A2(_16283_),
    .A1(net3836));
 sg13g2_nor2_1 _23653_ (.A(net3472),
    .B(_16289_),
    .Y(_16290_));
 sg13g2_xnor2_1 _23654_ (.Y(_16291_),
    .A(net3412),
    .B(_16289_));
 sg13g2_nor3_1 _23655_ (.A(_16258_),
    .B(_16273_),
    .C(_16274_),
    .Y(_16292_));
 sg13g2_or4_1 _23656_ (.A(_16214_),
    .B(_16215_),
    .C(_16240_),
    .D(_16241_),
    .X(_16293_));
 sg13g2_nor4_1 _23657_ (.A(_16258_),
    .B(_16273_),
    .C(_16274_),
    .D(_16293_),
    .Y(_16294_));
 sg13g2_o21ai_1 _23658_ (.B1(_16257_),
    .Y(_16295_),
    .A1(net3472),
    .A2(_16272_));
 sg13g2_a221oi_1 _23659_ (.B2(_16222_),
    .C1(_16295_),
    .B1(_16294_),
    .A1(_16259_),
    .Y(_16296_),
    .A2(_16292_));
 sg13g2_nand4_1 _23660_ (.B(_16161_),
    .C(_16217_),
    .A(_16146_),
    .Y(_16297_),
    .D(_16294_));
 sg13g2_o21ai_1 _23661_ (.B1(_16296_),
    .Y(_16298_),
    .A1(_16138_),
    .A2(_16297_));
 sg13g2_and2_1 _23662_ (.A(_16291_),
    .B(_16298_),
    .X(_16299_));
 sg13g2_nor2_1 _23663_ (.A(_16291_),
    .B(_16298_),
    .Y(_16300_));
 sg13g2_o21ai_1 _23664_ (.B1(net4320),
    .Y(_16301_),
    .A1(_16299_),
    .A2(_16300_));
 sg13g2_a21oi_1 _23665_ (.A1(net4292),
    .A2(_16289_),
    .Y(_16302_),
    .B1(net4234));
 sg13g2_a22oi_1 _23666_ (.Y(_16303_),
    .B1(_16301_),
    .B2(_16302_),
    .A2(net3934),
    .A1(net3168));
 sg13g2_inv_1 _23667_ (.Y(_00316_),
    .A(_16303_));
 sg13g2_a21oi_1 _23668_ (.A1(net4543),
    .A2(\u_inv.d_next[41] ),
    .Y(_16304_),
    .B1(net3759));
 sg13g2_a21oi_1 _23669_ (.A1(_14198_),
    .A2(_16280_),
    .Y(_16305_),
    .B1(_14197_));
 sg13g2_a21oi_1 _23670_ (.A1(_14196_),
    .A2(_16305_),
    .Y(_16306_),
    .B1(net4543));
 sg13g2_o21ai_1 _23671_ (.B1(_16306_),
    .Y(_16307_),
    .A1(_14196_),
    .A2(_16305_));
 sg13g2_nand3_1 _23672_ (.B(_14259_),
    .C(_16287_),
    .A(_14196_),
    .Y(_16308_));
 sg13g2_a21oi_1 _23673_ (.A1(_14259_),
    .A2(_16287_),
    .Y(_16309_),
    .B1(_14196_));
 sg13g2_nor2_1 _23674_ (.A(net3836),
    .B(_16309_),
    .Y(_16310_));
 sg13g2_a21oi_1 _23675_ (.A1(_14251_),
    .A2(_16284_),
    .Y(_16311_),
    .B1(_14200_));
 sg13g2_a22oi_1 _23676_ (.Y(_16312_),
    .B1(_16308_),
    .B2(_16310_),
    .A2(_16307_),
    .A1(_16304_));
 sg13g2_xnor2_1 _23677_ (.Y(_16313_),
    .A(net3472),
    .B(_16312_));
 sg13g2_nor2_1 _23678_ (.A(_16290_),
    .B(_16299_),
    .Y(_16314_));
 sg13g2_xor2_1 _23679_ (.B(_16314_),
    .A(_16313_),
    .X(_16315_));
 sg13g2_o21ai_1 _23680_ (.B1(net3882),
    .Y(_16316_),
    .A1(net4320),
    .A2(_16312_));
 sg13g2_a21oi_1 _23681_ (.A1(net4320),
    .A2(_16315_),
    .Y(_16317_),
    .B1(_16316_));
 sg13g2_a21o_1 _23682_ (.A2(net3934),
    .A1(net3117),
    .B1(_16317_),
    .X(_00317_));
 sg13g2_nand2b_1 _23683_ (.Y(_16318_),
    .B(_14261_),
    .A_N(_16311_));
 sg13g2_xnor2_1 _23684_ (.Y(_16319_),
    .A(_14191_),
    .B(_16318_));
 sg13g2_a221oi_1 _23685_ (.B2(_16280_),
    .C1(_14195_),
    .B1(_15493_),
    .A1(_14194_),
    .Y(_16320_),
    .A2(_14197_));
 sg13g2_a21oi_1 _23686_ (.A1(_14191_),
    .A2(_16320_),
    .Y(_16321_),
    .B1(net4543));
 sg13g2_o21ai_1 _23687_ (.B1(_16321_),
    .Y(_16322_),
    .A1(_14191_),
    .A2(_16320_));
 sg13g2_a21oi_1 _23688_ (.A1(net4543),
    .A2(\u_inv.d_next[42] ),
    .Y(_16323_),
    .B1(net3759));
 sg13g2_a22oi_1 _23689_ (.Y(_16324_),
    .B1(_16322_),
    .B2(_16323_),
    .A2(_16319_),
    .A1(net3759));
 sg13g2_nand2_1 _23690_ (.Y(_16325_),
    .A(net3412),
    .B(_16324_));
 sg13g2_xnor2_1 _23691_ (.Y(_16326_),
    .A(net3472),
    .B(_16324_));
 sg13g2_xnor2_1 _23692_ (.Y(_16327_),
    .A(net3412),
    .B(_16324_));
 sg13g2_a21o_1 _23693_ (.A2(_16312_),
    .A1(net3412),
    .B1(_16290_),
    .X(_16328_));
 sg13g2_a21oi_1 _23694_ (.A1(_16299_),
    .A2(_16313_),
    .Y(_16329_),
    .B1(_16328_));
 sg13g2_xnor2_1 _23695_ (.Y(_16330_),
    .A(_16327_),
    .B(_16329_));
 sg13g2_o21ai_1 _23696_ (.B1(net3882),
    .Y(_01828_),
    .A1(net4322),
    .A2(_16324_));
 sg13g2_a21oi_1 _23697_ (.A1(net4322),
    .A2(_16330_),
    .Y(_01829_),
    .B1(_01828_));
 sg13g2_a21o_1 _23698_ (.A2(net3934),
    .A1(net2970),
    .B1(_01829_),
    .X(_00318_));
 sg13g2_a21oi_1 _23699_ (.A1(net4543),
    .A2(\u_inv.d_next[43] ),
    .Y(_01830_),
    .B1(net3759));
 sg13g2_o21ai_1 _23700_ (.B1(_14190_),
    .Y(_01831_),
    .A1(_14191_),
    .A2(_16320_));
 sg13g2_o21ai_1 _23701_ (.B1(net4659),
    .Y(_01832_),
    .A1(_14189_),
    .A2(_01831_));
 sg13g2_a21o_1 _23702_ (.A2(_01831_),
    .A1(_14189_),
    .B1(_01832_),
    .X(_01833_));
 sg13g2_a21oi_1 _23703_ (.A1(_14191_),
    .A2(_16318_),
    .Y(_01834_),
    .B1(_14262_));
 sg13g2_or2_1 _23704_ (.X(_01835_),
    .B(_01834_),
    .A(_14188_));
 sg13g2_a21oi_1 _23705_ (.A1(_14188_),
    .A2(_01834_),
    .Y(_01836_),
    .B1(net3836));
 sg13g2_a22oi_1 _23706_ (.Y(_01837_),
    .B1(_01835_),
    .B2(_01836_),
    .A2(_01833_),
    .A1(_01830_));
 sg13g2_nand2_1 _23707_ (.Y(_01838_),
    .A(net3412),
    .B(_01837_));
 sg13g2_xnor2_1 _23708_ (.Y(_01839_),
    .A(net3473),
    .B(_01837_));
 sg13g2_o21ai_1 _23709_ (.B1(_16325_),
    .Y(_01840_),
    .A1(_16327_),
    .A2(_16329_));
 sg13g2_xnor2_1 _23710_ (.Y(_01841_),
    .A(_01839_),
    .B(_01840_));
 sg13g2_o21ai_1 _23711_ (.B1(net3884),
    .Y(_01842_),
    .A1(net4320),
    .A2(_01837_));
 sg13g2_a21oi_1 _23712_ (.A1(net4320),
    .A2(_01841_),
    .Y(_01843_),
    .B1(_01842_));
 sg13g2_a21o_1 _23713_ (.A2(net3934),
    .A1(net3094),
    .B1(_01843_),
    .X(_00319_));
 sg13g2_a21o_2 _23714_ (.A2(_16311_),
    .A1(_14193_),
    .B1(_14264_),
    .X(_01844_));
 sg13g2_xnor2_1 _23715_ (.Y(_01845_),
    .A(_14183_),
    .B(_01844_));
 sg13g2_a21oi_1 _23716_ (.A1(_15494_),
    .A2(_16280_),
    .Y(_01846_),
    .B1(_15499_));
 sg13g2_a21o_1 _23717_ (.A2(_16280_),
    .A1(_15494_),
    .B1(_15499_),
    .X(_01847_));
 sg13g2_a21oi_1 _23718_ (.A1(_14183_),
    .A2(_01846_),
    .Y(_01848_),
    .B1(net4545));
 sg13g2_o21ai_1 _23719_ (.B1(_01848_),
    .Y(_01849_),
    .A1(_14183_),
    .A2(_01846_));
 sg13g2_a21oi_1 _23720_ (.A1(net4545),
    .A2(\u_inv.d_next[44] ),
    .Y(_01850_),
    .B1(net3760));
 sg13g2_a22oi_1 _23721_ (.Y(_01851_),
    .B1(_01849_),
    .B2(_01850_),
    .A2(_01845_),
    .A1(net3761));
 sg13g2_xnor2_1 _23722_ (.Y(_01852_),
    .A(net3412),
    .B(_01851_));
 sg13g2_nand2_1 _23723_ (.Y(_01853_),
    .A(_16325_),
    .B(_01838_));
 sg13g2_o21ai_1 _23724_ (.B1(_01840_),
    .Y(_01854_),
    .A1(net3412),
    .A2(_01837_));
 sg13g2_and2_1 _23725_ (.A(_16326_),
    .B(_01839_),
    .X(_01855_));
 sg13g2_nand2_1 _23726_ (.Y(_01856_),
    .A(_01838_),
    .B(_01854_));
 sg13g2_nor2b_1 _23727_ (.A(_01852_),
    .B_N(_01856_),
    .Y(_01857_));
 sg13g2_xor2_1 _23728_ (.B(_01856_),
    .A(_01852_),
    .X(_01858_));
 sg13g2_o21ai_1 _23729_ (.B1(net3883),
    .Y(_01859_),
    .A1(net4320),
    .A2(_01851_));
 sg13g2_a21oi_1 _23730_ (.A1(net4321),
    .A2(_01858_),
    .Y(_01860_),
    .B1(_01859_));
 sg13g2_a21o_1 _23731_ (.A2(net3934),
    .A1(net3273),
    .B1(_01860_),
    .X(_00320_));
 sg13g2_a21oi_1 _23732_ (.A1(net4545),
    .A2(\u_inv.d_next[45] ),
    .Y(_01861_),
    .B1(net3761));
 sg13g2_o21ai_1 _23733_ (.B1(_14182_),
    .Y(_01862_),
    .A1(_14183_),
    .A2(_01846_));
 sg13g2_xnor2_1 _23734_ (.Y(_01863_),
    .A(_14181_),
    .B(_01862_));
 sg13g2_nand2_1 _23735_ (.Y(_01864_),
    .A(net4659),
    .B(_01863_));
 sg13g2_a21oi_1 _23736_ (.A1(_14183_),
    .A2(_01844_),
    .Y(_01865_),
    .B1(_14254_));
 sg13g2_or2_1 _23737_ (.X(_01866_),
    .B(_01865_),
    .A(_14181_));
 sg13g2_a21oi_1 _23738_ (.A1(_14181_),
    .A2(_01865_),
    .Y(_01867_),
    .B1(net3836));
 sg13g2_a22oi_1 _23739_ (.Y(_01868_),
    .B1(_01866_),
    .B2(_01867_),
    .A2(_01864_),
    .A1(_01861_));
 sg13g2_and2_1 _23740_ (.A(net3413),
    .B(_01868_),
    .X(_01869_));
 sg13g2_nand2b_1 _23741_ (.Y(_01870_),
    .B(net3473),
    .A_N(_01868_));
 sg13g2_xnor2_1 _23742_ (.Y(_01871_),
    .A(net3413),
    .B(_01868_));
 sg13g2_a21o_1 _23743_ (.A2(_01851_),
    .A1(net3413),
    .B1(_01857_),
    .X(_01872_));
 sg13g2_xor2_1 _23744_ (.B(_01872_),
    .A(_01871_),
    .X(_01873_));
 sg13g2_o21ai_1 _23745_ (.B1(net3884),
    .Y(_01874_),
    .A1(net4320),
    .A2(_01868_));
 sg13g2_a21oi_1 _23746_ (.A1(net4321),
    .A2(_01873_),
    .Y(_01875_),
    .B1(_01874_));
 sg13g2_a21o_1 _23747_ (.A2(net3935),
    .A1(net3146),
    .B1(_01875_),
    .X(_00321_));
 sg13g2_a21oi_1 _23748_ (.A1(_14184_),
    .A2(_01844_),
    .Y(_01876_),
    .B1(_14255_));
 sg13g2_xnor2_1 _23749_ (.Y(_01877_),
    .A(_14177_),
    .B(_01876_));
 sg13g2_a21oi_1 _23750_ (.A1(_15490_),
    .A2(_01847_),
    .Y(_01878_),
    .B1(_15501_));
 sg13g2_a21oi_1 _23751_ (.A1(_14178_),
    .A2(_01878_),
    .Y(_01879_),
    .B1(net4545));
 sg13g2_o21ai_1 _23752_ (.B1(_01879_),
    .Y(_01880_),
    .A1(_14178_),
    .A2(_01878_));
 sg13g2_a21oi_1 _23753_ (.A1(net4545),
    .A2(\u_inv.d_next[46] ),
    .Y(_01881_),
    .B1(net3760));
 sg13g2_a22oi_1 _23754_ (.Y(_01882_),
    .B1(_01880_),
    .B2(_01881_),
    .A2(_01877_),
    .A1(net3760));
 sg13g2_nand2_1 _23755_ (.Y(_01883_),
    .A(net3414),
    .B(_01882_));
 sg13g2_xnor2_1 _23756_ (.Y(_01884_),
    .A(net3414),
    .B(_01882_));
 sg13g2_inv_1 _23757_ (.Y(_01885_),
    .A(_01884_));
 sg13g2_a21o_1 _23758_ (.A2(_01851_),
    .A1(net3413),
    .B1(_01869_),
    .X(_01886_));
 sg13g2_o21ai_1 _23759_ (.B1(_01870_),
    .Y(_01887_),
    .A1(_01857_),
    .A2(_01886_));
 sg13g2_xnor2_1 _23760_ (.Y(_01888_),
    .A(_01884_),
    .B(_01887_));
 sg13g2_o21ai_1 _23761_ (.B1(net3883),
    .Y(_01889_),
    .A1(net4321),
    .A2(_01882_));
 sg13g2_a21oi_1 _23762_ (.A1(net4321),
    .A2(_01888_),
    .Y(_01890_),
    .B1(_01889_));
 sg13g2_a21o_1 _23763_ (.A2(net3935),
    .A1(net3023),
    .B1(_01890_),
    .X(_00322_));
 sg13g2_a21oi_1 _23764_ (.A1(net4545),
    .A2(\u_inv.d_next[47] ),
    .Y(_01891_),
    .B1(net3760));
 sg13g2_o21ai_1 _23765_ (.B1(_14176_),
    .Y(_01892_),
    .A1(_14178_),
    .A2(_01878_));
 sg13g2_o21ai_1 _23766_ (.B1(net4659),
    .Y(_01893_),
    .A1(_14175_),
    .A2(_01892_));
 sg13g2_a21o_1 _23767_ (.A2(_01892_),
    .A1(_14175_),
    .B1(_01893_),
    .X(_01894_));
 sg13g2_o21ai_1 _23768_ (.B1(_14256_),
    .Y(_01895_),
    .A1(_14177_),
    .A2(_01876_));
 sg13g2_or2_1 _23769_ (.X(_01896_),
    .B(_01895_),
    .A(_14175_));
 sg13g2_a21oi_1 _23770_ (.A1(_14175_),
    .A2(_01895_),
    .Y(_01897_),
    .B1(net3836));
 sg13g2_a22oi_1 _23771_ (.Y(_01898_),
    .B1(_01896_),
    .B2(_01897_),
    .A2(_01894_),
    .A1(_01891_));
 sg13g2_xnor2_1 _23772_ (.Y(_01899_),
    .A(net3473),
    .B(_01898_));
 sg13g2_o21ai_1 _23773_ (.B1(_01883_),
    .Y(_01900_),
    .A1(_01884_),
    .A2(_01887_));
 sg13g2_xnor2_1 _23774_ (.Y(_01901_),
    .A(_01899_),
    .B(_01900_));
 sg13g2_o21ai_1 _23775_ (.B1(net3883),
    .Y(_01902_),
    .A1(net4320),
    .A2(_01898_));
 sg13g2_a21oi_1 _23776_ (.A1(net4321),
    .A2(_01901_),
    .Y(_01903_),
    .B1(_01902_));
 sg13g2_a21o_1 _23777_ (.A2(net3935),
    .A1(net3182),
    .B1(_01903_),
    .X(_00323_));
 sg13g2_a21oi_1 _23778_ (.A1(_15617_),
    .A2(_15620_),
    .Y(_01904_),
    .B1(_15507_));
 sg13g2_a21o_2 _23779_ (.A2(_15620_),
    .A1(_15617_),
    .B1(_15507_),
    .X(_01905_));
 sg13g2_nand2_1 _23780_ (.Y(_01906_),
    .A(_14171_),
    .B(_01905_));
 sg13g2_xnor2_1 _23781_ (.Y(_01907_),
    .A(_14171_),
    .B(_01905_));
 sg13g2_nor2_1 _23782_ (.A(net4670),
    .B(\u_inv.d_next[48] ),
    .Y(_01908_));
 sg13g2_a21oi_1 _23783_ (.A1(net4672),
    .A2(_01907_),
    .Y(_01909_),
    .B1(_01908_));
 sg13g2_o21ai_1 _23784_ (.B1(_14236_),
    .Y(_01910_),
    .A1(_14090_),
    .A2(_14120_));
 sg13g2_and2_1 _23785_ (.A(_14267_),
    .B(_01910_),
    .X(_01911_));
 sg13g2_or2_1 _23786_ (.X(_01912_),
    .B(_01911_),
    .A(_14171_));
 sg13g2_a21oi_1 _23787_ (.A1(_14171_),
    .A2(_01911_),
    .Y(_01913_),
    .B1(net3841));
 sg13g2_a22oi_1 _23788_ (.Y(_01914_),
    .B1(_01912_),
    .B2(_01913_),
    .A2(_01909_),
    .A1(net3842));
 sg13g2_nor2_1 _23789_ (.A(net3474),
    .B(_01914_),
    .Y(_01915_));
 sg13g2_xnor2_1 _23790_ (.Y(_01916_),
    .A(net3418),
    .B(_01914_));
 sg13g2_nor2_1 _23791_ (.A(_01852_),
    .B(_01871_),
    .Y(_01917_));
 sg13g2_and4_1 _23792_ (.A(_16291_),
    .B(_16313_),
    .C(_16326_),
    .D(_01839_),
    .X(_01918_));
 sg13g2_nand4_1 _23793_ (.B(_01899_),
    .C(_01917_),
    .A(_01885_),
    .Y(_01919_),
    .D(_01918_));
 sg13g2_or2_1 _23794_ (.X(_01920_),
    .B(_01919_),
    .A(_16296_));
 sg13g2_nand3_1 _23795_ (.B(_01886_),
    .C(_01899_),
    .A(_01885_),
    .Y(_01921_));
 sg13g2_o21ai_1 _23796_ (.B1(net3412),
    .Y(_01922_),
    .A1(_01882_),
    .A2(_01898_));
 sg13g2_a21o_1 _23797_ (.A2(_01855_),
    .A1(_16328_),
    .B1(_01853_),
    .X(_01923_));
 sg13g2_nand4_1 _23798_ (.B(_01899_),
    .C(_01917_),
    .A(_01885_),
    .Y(_01924_),
    .D(_01923_));
 sg13g2_nand4_1 _23799_ (.B(_01921_),
    .C(_01922_),
    .A(_01920_),
    .Y(_01925_),
    .D(_01924_));
 sg13g2_or2_1 _23800_ (.X(_01926_),
    .B(_01919_),
    .A(_16297_));
 sg13g2_nor2_1 _23801_ (.A(_16138_),
    .B(_01926_),
    .Y(_01927_));
 sg13g2_or2_1 _23802_ (.X(_01928_),
    .B(_01927_),
    .A(_01925_));
 sg13g2_xnor2_1 _23803_ (.Y(_01929_),
    .A(_01916_),
    .B(_01928_));
 sg13g2_nand2_1 _23804_ (.Y(_01930_),
    .A(net4293),
    .B(_01914_));
 sg13g2_a21oi_1 _23805_ (.A1(net4327),
    .A2(_01929_),
    .Y(_01931_),
    .B1(net4235));
 sg13g2_a22oi_1 _23806_ (.Y(_01932_),
    .B1(_01930_),
    .B2(_01931_),
    .A2(net3946),
    .A1(net3225));
 sg13g2_inv_1 _23807_ (.Y(_00324_),
    .A(_01932_));
 sg13g2_nand2_1 _23808_ (.Y(_01933_),
    .A(net2215),
    .B(net3943));
 sg13g2_a21oi_1 _23809_ (.A1(_01916_),
    .A2(_01928_),
    .Y(_01934_),
    .B1(_01915_));
 sg13g2_nand3_1 _23810_ (.B(_14170_),
    .C(_01906_),
    .A(_14168_),
    .Y(_01935_));
 sg13g2_a21oi_1 _23811_ (.A1(_15511_),
    .A2(_01905_),
    .Y(_01936_),
    .B1(net4549));
 sg13g2_nand3_1 _23812_ (.B(_01935_),
    .C(_01936_),
    .A(_15533_),
    .Y(_01937_));
 sg13g2_a21oi_1 _23813_ (.A1(net4557),
    .A2(\u_inv.d_next[49] ),
    .Y(_01938_),
    .B1(net3767));
 sg13g2_nand2_1 _23814_ (.Y(_01939_),
    .A(_14285_),
    .B(_01912_));
 sg13g2_xnor2_1 _23815_ (.Y(_01940_),
    .A(_14168_),
    .B(_01939_));
 sg13g2_a22oi_1 _23816_ (.Y(_01941_),
    .B1(_01940_),
    .B2(net3767),
    .A2(_01938_),
    .A1(_01937_));
 sg13g2_nand2_1 _23817_ (.Y(_01942_),
    .A(net3418),
    .B(_01941_));
 sg13g2_nor2_1 _23818_ (.A(net3418),
    .B(_01941_),
    .Y(_01943_));
 sg13g2_xnor2_1 _23819_ (.Y(_01944_),
    .A(net3474),
    .B(_01941_));
 sg13g2_o21ai_1 _23820_ (.B1(net4327),
    .Y(_01945_),
    .A1(_01934_),
    .A2(_01944_));
 sg13g2_a21oi_1 _23821_ (.A1(_01934_),
    .A2(_01944_),
    .Y(_01946_),
    .B1(_01945_));
 sg13g2_o21ai_1 _23822_ (.B1(net3886),
    .Y(_01947_),
    .A1(net4327),
    .A2(_01941_));
 sg13g2_o21ai_1 _23823_ (.B1(_01933_),
    .Y(_00325_),
    .A1(_01946_),
    .A2(_01947_));
 sg13g2_o21ai_1 _23824_ (.B1(_14287_),
    .Y(_01948_),
    .A1(_14172_),
    .A2(_01911_));
 sg13g2_xnor2_1 _23825_ (.Y(_01949_),
    .A(_14165_),
    .B(_01948_));
 sg13g2_a21oi_1 _23826_ (.A1(_15511_),
    .A2(_01905_),
    .Y(_01950_),
    .B1(_15534_));
 sg13g2_a21o_1 _23827_ (.A2(_01905_),
    .A1(_15511_),
    .B1(_15534_),
    .X(_01951_));
 sg13g2_nand2b_1 _23828_ (.Y(_01952_),
    .B(_01951_),
    .A_N(_14165_));
 sg13g2_a21oi_1 _23829_ (.A1(_14165_),
    .A2(_01950_),
    .Y(_01953_),
    .B1(net4549));
 sg13g2_nand2_1 _23830_ (.Y(_01954_),
    .A(_01952_),
    .B(_01953_));
 sg13g2_a21oi_1 _23831_ (.A1(net4549),
    .A2(\u_inv.d_next[50] ),
    .Y(_01955_),
    .B1(net3767));
 sg13g2_a22oi_1 _23832_ (.Y(_01956_),
    .B1(_01954_),
    .B2(_01955_),
    .A2(_01949_),
    .A1(net3767));
 sg13g2_xnor2_1 _23833_ (.Y(_01957_),
    .A(net3418),
    .B(_01956_));
 sg13g2_nor2b_1 _23834_ (.A(_01915_),
    .B_N(_01942_),
    .Y(_01958_));
 sg13g2_o21ai_1 _23835_ (.B1(_01942_),
    .Y(_01959_),
    .A1(_01934_),
    .A2(_01943_));
 sg13g2_nor2b_1 _23836_ (.A(_01957_),
    .B_N(_01959_),
    .Y(_01960_));
 sg13g2_xor2_1 _23837_ (.B(_01959_),
    .A(_01957_),
    .X(_01961_));
 sg13g2_a21oi_1 _23838_ (.A1(net4327),
    .A2(_01961_),
    .Y(_01962_),
    .B1(net4235));
 sg13g2_o21ai_1 _23839_ (.B1(_01962_),
    .Y(_01963_),
    .A1(net4327),
    .A2(_01956_));
 sg13g2_o21ai_1 _23840_ (.B1(_01963_),
    .Y(_00326_),
    .A1(_10614_),
    .A2(net4025));
 sg13g2_nand2_1 _23841_ (.Y(_01964_),
    .A(net2064),
    .B(net3946));
 sg13g2_nand3_1 _23842_ (.B(_14164_),
    .C(_01952_),
    .A(_14163_),
    .Y(_01965_));
 sg13g2_a21o_1 _23843_ (.A2(_01952_),
    .A1(_14164_),
    .B1(_14163_),
    .X(_01966_));
 sg13g2_nand3_1 _23844_ (.B(_01965_),
    .C(_01966_),
    .A(net4670),
    .Y(_01967_));
 sg13g2_a21oi_1 _23845_ (.A1(net4549),
    .A2(\u_inv.d_next[51] ),
    .Y(_01968_),
    .B1(net3767));
 sg13g2_a21oi_1 _23846_ (.A1(_14165_),
    .A2(_01948_),
    .Y(_01969_),
    .B1(_14289_));
 sg13g2_or2_1 _23847_ (.X(_01970_),
    .B(_01969_),
    .A(_14163_));
 sg13g2_a21oi_1 _23848_ (.A1(_14163_),
    .A2(_01969_),
    .Y(_01971_),
    .B1(net3842));
 sg13g2_a22oi_1 _23849_ (.Y(_01972_),
    .B1(_01970_),
    .B2(_01971_),
    .A2(_01968_),
    .A1(_01967_));
 sg13g2_xnor2_1 _23850_ (.Y(_01973_),
    .A(net3422),
    .B(_01972_));
 sg13g2_a21o_1 _23851_ (.A2(_01956_),
    .A1(net3418),
    .B1(_01960_),
    .X(_01974_));
 sg13g2_o21ai_1 _23852_ (.B1(net4327),
    .Y(_01975_),
    .A1(_01973_),
    .A2(_01974_));
 sg13g2_a21oi_1 _23853_ (.A1(_01973_),
    .A2(_01974_),
    .Y(_01976_),
    .B1(_01975_));
 sg13g2_o21ai_1 _23854_ (.B1(net3888),
    .Y(_01977_),
    .A1(net4331),
    .A2(_01972_));
 sg13g2_o21ai_1 _23855_ (.B1(_01964_),
    .Y(_00327_),
    .A1(_01976_),
    .A2(_01977_));
 sg13g2_a21oi_2 _23856_ (.B1(_14291_),
    .Y(_01978_),
    .A2(_01948_),
    .A1(_14166_));
 sg13g2_xnor2_1 _23857_ (.Y(_01979_),
    .A(_14159_),
    .B(_01978_));
 sg13g2_a21oi_1 _23858_ (.A1(_15510_),
    .A2(_01951_),
    .Y(_01980_),
    .B1(_15532_));
 sg13g2_a21o_2 _23859_ (.A2(_01951_),
    .A1(_15510_),
    .B1(_15532_),
    .X(_01981_));
 sg13g2_a21oi_1 _23860_ (.A1(_14159_),
    .A2(_01981_),
    .Y(_01982_),
    .B1(net4552));
 sg13g2_o21ai_1 _23861_ (.B1(_01982_),
    .Y(_01983_),
    .A1(_14159_),
    .A2(_01981_));
 sg13g2_a21oi_1 _23862_ (.A1(net4552),
    .A2(\u_inv.d_next[52] ),
    .Y(_01984_),
    .B1(net3771));
 sg13g2_a22oi_1 _23863_ (.Y(_01985_),
    .B1(_01983_),
    .B2(_01984_),
    .A2(_01979_),
    .A1(net3771));
 sg13g2_nand2_1 _23864_ (.Y(_01986_),
    .A(net3419),
    .B(_01985_));
 sg13g2_xnor2_1 _23865_ (.Y(_01987_),
    .A(net3420),
    .B(_01985_));
 sg13g2_nor2_1 _23866_ (.A(_01957_),
    .B(_01973_),
    .Y(_01988_));
 sg13g2_or2_1 _23867_ (.X(_01989_),
    .B(_01973_),
    .A(_01957_));
 sg13g2_o21ai_1 _23868_ (.B1(net3418),
    .Y(_01990_),
    .A1(_01956_),
    .A2(_01972_));
 sg13g2_o21ai_1 _23869_ (.B1(_01990_),
    .Y(_01991_),
    .A1(_01958_),
    .A2(_01989_));
 sg13g2_nand3_1 _23870_ (.B(_01944_),
    .C(_01988_),
    .A(_01916_),
    .Y(_01992_));
 sg13g2_inv_1 _23871_ (.Y(_01993_),
    .A(_01992_));
 sg13g2_a21oi_1 _23872_ (.A1(_01928_),
    .A2(_01993_),
    .Y(_01994_),
    .B1(_01991_));
 sg13g2_xnor2_1 _23873_ (.Y(_01995_),
    .A(_01987_),
    .B(_01994_));
 sg13g2_a21oi_1 _23874_ (.A1(net4329),
    .A2(_01995_),
    .Y(_01996_),
    .B1(net4235));
 sg13g2_o21ai_1 _23875_ (.B1(_01996_),
    .Y(_01997_),
    .A1(net4332),
    .A2(_01985_));
 sg13g2_o21ai_1 _23876_ (.B1(_01997_),
    .Y(_00328_),
    .A1(_10613_),
    .A2(net4025));
 sg13g2_nand2_1 _23877_ (.Y(_01998_),
    .A(net2447),
    .B(net3945));
 sg13g2_a21oi_1 _23878_ (.A1(net4552),
    .A2(\u_inv.d_next[53] ),
    .Y(_01999_),
    .B1(net3771));
 sg13g2_o21ai_1 _23879_ (.B1(_14158_),
    .Y(_02000_),
    .A1(_14160_),
    .A2(_01980_));
 sg13g2_o21ai_1 _23880_ (.B1(net4672),
    .Y(_02001_),
    .A1(_14156_),
    .A2(_02000_));
 sg13g2_a21o_1 _23881_ (.A2(_02000_),
    .A1(_14156_),
    .B1(_02001_),
    .X(_02002_));
 sg13g2_o21ai_1 _23882_ (.B1(_14295_),
    .Y(_02003_),
    .A1(_14159_),
    .A2(_01978_));
 sg13g2_nand2b_1 _23883_ (.Y(_02004_),
    .B(_14157_),
    .A_N(_02003_));
 sg13g2_a21oi_1 _23884_ (.A1(_14156_),
    .A2(_02003_),
    .Y(_02005_),
    .B1(net3842));
 sg13g2_a22oi_1 _23885_ (.Y(_02006_),
    .B1(_02004_),
    .B2(_02005_),
    .A2(_02002_),
    .A1(_01999_));
 sg13g2_nand2_1 _23886_ (.Y(_02007_),
    .A(net3419),
    .B(_02006_));
 sg13g2_xnor2_1 _23887_ (.Y(_02008_),
    .A(net3419),
    .B(_02006_));
 sg13g2_o21ai_1 _23888_ (.B1(_01986_),
    .Y(_02009_),
    .A1(_01987_),
    .A2(_01994_));
 sg13g2_o21ai_1 _23889_ (.B1(net4329),
    .Y(_02010_),
    .A1(_02008_),
    .A2(_02009_));
 sg13g2_a21oi_1 _23890_ (.A1(_02008_),
    .A2(_02009_),
    .Y(_02011_),
    .B1(_02010_));
 sg13g2_o21ai_1 _23891_ (.B1(net3888),
    .Y(_02012_),
    .A1(net4331),
    .A2(_02006_));
 sg13g2_o21ai_1 _23892_ (.B1(_01998_),
    .Y(_00329_),
    .A1(_02011_),
    .A2(_02012_));
 sg13g2_o21ai_1 _23893_ (.B1(_14297_),
    .Y(_02013_),
    .A1(_14161_),
    .A2(_01978_));
 sg13g2_xnor2_1 _23894_ (.Y(_02014_),
    .A(_14152_),
    .B(_02013_));
 sg13g2_a21oi_1 _23895_ (.A1(_15508_),
    .A2(_01981_),
    .Y(_02015_),
    .B1(_15536_));
 sg13g2_a21oi_1 _23896_ (.A1(_14152_),
    .A2(_02015_),
    .Y(_02016_),
    .B1(net4552));
 sg13g2_o21ai_1 _23897_ (.B1(_02016_),
    .Y(_02017_),
    .A1(_14152_),
    .A2(_02015_));
 sg13g2_a21oi_1 _23898_ (.A1(net4552),
    .A2(\u_inv.d_next[54] ),
    .Y(_02018_),
    .B1(net3771));
 sg13g2_a22oi_1 _23899_ (.Y(_02019_),
    .B1(_02017_),
    .B2(_02018_),
    .A2(_02014_),
    .A1(net3771));
 sg13g2_and2_1 _23900_ (.A(net3419),
    .B(_02019_),
    .X(_02020_));
 sg13g2_xnor2_1 _23901_ (.Y(_02021_),
    .A(net3420),
    .B(_02019_));
 sg13g2_inv_2 _23902_ (.Y(_02022_),
    .A(_02021_));
 sg13g2_nand2_1 _23903_ (.Y(_02023_),
    .A(_01986_),
    .B(_02007_));
 sg13g2_nor2_1 _23904_ (.A(_01987_),
    .B(_02008_),
    .Y(_02024_));
 sg13g2_or2_1 _23905_ (.X(_02025_),
    .B(_02008_),
    .A(_01987_));
 sg13g2_nor2_1 _23906_ (.A(_01994_),
    .B(_02025_),
    .Y(_02026_));
 sg13g2_or2_1 _23907_ (.X(_02027_),
    .B(_02026_),
    .A(_02023_));
 sg13g2_xnor2_1 _23908_ (.Y(_02028_),
    .A(_02022_),
    .B(_02027_));
 sg13g2_o21ai_1 _23909_ (.B1(net3886),
    .Y(_02029_),
    .A1(net4329),
    .A2(_02019_));
 sg13g2_a21oi_1 _23910_ (.A1(net4329),
    .A2(_02028_),
    .Y(_02030_),
    .B1(_02029_));
 sg13g2_a21o_1 _23911_ (.A2(net3945),
    .A1(net3079),
    .B1(_02030_),
    .X(_00330_));
 sg13g2_a21oi_1 _23912_ (.A1(net4552),
    .A2(\u_inv.d_next[55] ),
    .Y(_02031_),
    .B1(net3771));
 sg13g2_o21ai_1 _23913_ (.B1(_14150_),
    .Y(_02032_),
    .A1(_14152_),
    .A2(_02015_));
 sg13g2_o21ai_1 _23914_ (.B1(net4672),
    .Y(_02033_),
    .A1(_14149_),
    .A2(_02032_));
 sg13g2_a21o_1 _23915_ (.A2(_02032_),
    .A1(_14149_),
    .B1(_02033_),
    .X(_02034_));
 sg13g2_a21oi_1 _23916_ (.A1(_14152_),
    .A2(_02013_),
    .Y(_02035_),
    .B1(_14293_));
 sg13g2_or2_1 _23917_ (.X(_02036_),
    .B(_02035_),
    .A(_14148_));
 sg13g2_a21oi_1 _23918_ (.A1(_14148_),
    .A2(_02035_),
    .Y(_02037_),
    .B1(net3842));
 sg13g2_a22oi_1 _23919_ (.Y(_02038_),
    .B1(_02036_),
    .B2(_02037_),
    .A2(_02034_),
    .A1(_02031_));
 sg13g2_xnor2_1 _23920_ (.Y(_02039_),
    .A(net3475),
    .B(_02038_));
 sg13g2_xnor2_1 _23921_ (.Y(_02040_),
    .A(net3420),
    .B(_02038_));
 sg13g2_a21oi_1 _23922_ (.A1(_02022_),
    .A2(_02027_),
    .Y(_02041_),
    .B1(_02020_));
 sg13g2_xnor2_1 _23923_ (.Y(_02042_),
    .A(_02040_),
    .B(_02041_));
 sg13g2_o21ai_1 _23924_ (.B1(net3885),
    .Y(_02043_),
    .A1(net4329),
    .A2(_02038_));
 sg13g2_a21oi_1 _23925_ (.A1(net4329),
    .A2(_02042_),
    .Y(_02044_),
    .B1(_02043_));
 sg13g2_a21o_1 _23926_ (.A2(net3945),
    .A1(net3026),
    .B1(_02044_),
    .X(_00331_));
 sg13g2_a21o_2 _23927_ (.A2(_01910_),
    .A1(_14267_),
    .B1(_14173_),
    .X(_02045_));
 sg13g2_a21oi_1 _23928_ (.A1(_14299_),
    .A2(_02045_),
    .Y(_02046_),
    .B1(_14142_));
 sg13g2_nand3_1 _23929_ (.B(_14299_),
    .C(_02045_),
    .A(_14142_),
    .Y(_02047_));
 sg13g2_nand2b_1 _23930_ (.Y(_02048_),
    .B(_02047_),
    .A_N(_02046_));
 sg13g2_o21ai_1 _23931_ (.B1(_15540_),
    .Y(_02049_),
    .A1(_15512_),
    .A2(_01904_));
 sg13g2_nand2_1 _23932_ (.Y(_02050_),
    .A(_14142_),
    .B(_02049_));
 sg13g2_o21ai_1 _23933_ (.B1(net4671),
    .Y(_02051_),
    .A1(_14142_),
    .A2(_02049_));
 sg13g2_nand2b_1 _23934_ (.Y(_02052_),
    .B(_02050_),
    .A_N(_02051_));
 sg13g2_a21oi_1 _23935_ (.A1(net4553),
    .A2(\u_inv.d_next[56] ),
    .Y(_02053_),
    .B1(net3772));
 sg13g2_a22oi_1 _23936_ (.Y(_02054_),
    .B1(_02052_),
    .B2(_02053_),
    .A2(_02048_),
    .A1(net3772));
 sg13g2_nand2_1 _23937_ (.Y(_02055_),
    .A(net3421),
    .B(_02054_));
 sg13g2_xnor2_1 _23938_ (.Y(_02056_),
    .A(net3421),
    .B(_02054_));
 sg13g2_nand4_1 _23939_ (.B(_02022_),
    .C(_02024_),
    .A(_01991_),
    .Y(_02057_),
    .D(_02039_));
 sg13g2_nand3_1 _23940_ (.B(_02023_),
    .C(_02039_),
    .A(_02022_),
    .Y(_02058_));
 sg13g2_a21oi_1 _23941_ (.A1(net3420),
    .A2(_02038_),
    .Y(_02059_),
    .B1(_02020_));
 sg13g2_nand3_1 _23942_ (.B(_02058_),
    .C(_02059_),
    .A(_02057_),
    .Y(_02060_));
 sg13g2_or4_1 _23943_ (.A(_01992_),
    .B(_02021_),
    .C(_02025_),
    .D(_02040_),
    .X(_02061_));
 sg13g2_inv_1 _23944_ (.Y(_02062_),
    .A(_02061_));
 sg13g2_a21oi_1 _23945_ (.A1(_01928_),
    .A2(_02062_),
    .Y(_02063_),
    .B1(_02060_));
 sg13g2_or2_1 _23946_ (.X(_02064_),
    .B(_02063_),
    .A(_02056_));
 sg13g2_xnor2_1 _23947_ (.Y(_02065_),
    .A(_02056_),
    .B(_02063_));
 sg13g2_o21ai_1 _23948_ (.B1(net3888),
    .Y(_02066_),
    .A1(net4331),
    .A2(_02054_));
 sg13g2_a21oi_1 _23949_ (.A1(net4330),
    .A2(_02065_),
    .Y(_02067_),
    .B1(_02066_));
 sg13g2_a21o_1 _23950_ (.A2(net3945),
    .A1(net2458),
    .B1(_02067_),
    .X(_00332_));
 sg13g2_nand2_1 _23951_ (.Y(_02068_),
    .A(net2112),
    .B(net3945));
 sg13g2_nand2_1 _23952_ (.Y(_02069_),
    .A(_02055_),
    .B(_02064_));
 sg13g2_a21oi_1 _23953_ (.A1(_15517_),
    .A2(_02049_),
    .Y(_02070_),
    .B1(_15519_));
 sg13g2_nor2_1 _23954_ (.A(_14140_),
    .B(_14141_),
    .Y(_02071_));
 sg13g2_a21oi_1 _23955_ (.A1(_02050_),
    .A2(_02071_),
    .Y(_02072_),
    .B1(net4553));
 sg13g2_nand2_1 _23956_ (.Y(_02073_),
    .A(_02070_),
    .B(_02072_));
 sg13g2_a21oi_1 _23957_ (.A1(net4552),
    .A2(\u_inv.d_next[57] ),
    .Y(_02074_),
    .B1(net3772));
 sg13g2_nor2_1 _23958_ (.A(_14269_),
    .B(_02046_),
    .Y(_02075_));
 sg13g2_xnor2_1 _23959_ (.Y(_02076_),
    .A(_14140_),
    .B(_02075_));
 sg13g2_a22oi_1 _23960_ (.Y(_02077_),
    .B1(_02076_),
    .B2(net3772),
    .A2(_02074_),
    .A1(_02073_));
 sg13g2_xnor2_1 _23961_ (.Y(_02078_),
    .A(net3421),
    .B(_02077_));
 sg13g2_o21ai_1 _23962_ (.B1(net4331),
    .Y(_02079_),
    .A1(_02069_),
    .A2(_02078_));
 sg13g2_a21oi_1 _23963_ (.A1(_02069_),
    .A2(_02078_),
    .Y(_02080_),
    .B1(_02079_));
 sg13g2_o21ai_1 _23964_ (.B1(net3887),
    .Y(_02081_),
    .A1(net4331),
    .A2(_02077_));
 sg13g2_o21ai_1 _23965_ (.B1(_02068_),
    .Y(_00333_),
    .A1(_02080_),
    .A2(_02081_));
 sg13g2_a21oi_1 _23966_ (.A1(_14299_),
    .A2(_02045_),
    .Y(_02082_),
    .B1(_14144_));
 sg13g2_o21ai_1 _23967_ (.B1(_14138_),
    .Y(_02083_),
    .A1(_14271_),
    .A2(_02082_));
 sg13g2_or3_1 _23968_ (.A(_14138_),
    .B(_14271_),
    .C(_02082_),
    .X(_02084_));
 sg13g2_nand2_1 _23969_ (.Y(_02085_),
    .A(_02083_),
    .B(_02084_));
 sg13g2_a221oi_1 _23970_ (.B2(_02049_),
    .C1(_15519_),
    .B1(_15517_),
    .A1(\u_inv.d_next[57] ),
    .Y(_02086_),
    .A2(\u_inv.d_reg[57] ));
 sg13g2_nand2b_1 _23971_ (.Y(_02087_),
    .B(_14137_),
    .A_N(_02086_));
 sg13g2_a21oi_1 _23972_ (.A1(_14138_),
    .A2(_02086_),
    .Y(_02088_),
    .B1(net4552));
 sg13g2_a221oi_1 _23973_ (.B2(_02088_),
    .C1(net3771),
    .B1(_02087_),
    .A1(net4553),
    .Y(_02089_),
    .A2(net4804));
 sg13g2_a21oi_2 _23974_ (.B1(_02089_),
    .Y(_02090_),
    .A2(_02085_),
    .A1(net3772));
 sg13g2_nand2_1 _23975_ (.Y(_02091_),
    .A(net3421),
    .B(_02090_));
 sg13g2_xnor2_1 _23976_ (.Y(_02092_),
    .A(net3475),
    .B(_02090_));
 sg13g2_o21ai_1 _23977_ (.B1(net3421),
    .Y(_02093_),
    .A1(_02054_),
    .A2(_02077_));
 sg13g2_inv_1 _23978_ (.Y(_02094_),
    .A(_02093_));
 sg13g2_nor2_1 _23979_ (.A(_02056_),
    .B(_02078_),
    .Y(_02095_));
 sg13g2_o21ai_1 _23980_ (.B1(_02093_),
    .Y(_02096_),
    .A1(_02064_),
    .A2(_02078_));
 sg13g2_nand2_1 _23981_ (.Y(_02097_),
    .A(_02092_),
    .B(_02096_));
 sg13g2_xnor2_1 _23982_ (.Y(_02098_),
    .A(_02092_),
    .B(_02096_));
 sg13g2_a21oi_1 _23983_ (.A1(net4331),
    .A2(_02098_),
    .Y(_02099_),
    .B1(net4235));
 sg13g2_o21ai_1 _23984_ (.B1(_02099_),
    .Y(_02100_),
    .A1(net4331),
    .A2(_02090_));
 sg13g2_o21ai_1 _23985_ (.B1(_02100_),
    .Y(_00334_),
    .A1(_10612_),
    .A2(net4025));
 sg13g2_nand2_1 _23986_ (.Y(_02101_),
    .A(_02091_),
    .B(_02097_));
 sg13g2_nand2b_1 _23987_ (.Y(_02102_),
    .B(net3842),
    .A_N(\u_inv.d_next[59] ));
 sg13g2_o21ai_1 _23988_ (.B1(_14136_),
    .Y(_02103_),
    .A1(_14138_),
    .A2(_02086_));
 sg13g2_xnor2_1 _23989_ (.Y(_02104_),
    .A(_14134_),
    .B(_02103_));
 sg13g2_a22oi_1 _23990_ (.Y(_02105_),
    .B1(_02104_),
    .B2(net4671),
    .A2(_02102_),
    .A1(net3728));
 sg13g2_a21oi_1 _23991_ (.A1(_14273_),
    .A2(_02083_),
    .Y(_02106_),
    .B1(_14134_));
 sg13g2_and3_1 _23992_ (.X(_02107_),
    .A(_14134_),
    .B(_14273_),
    .C(_02083_));
 sg13g2_nor3_1 _23993_ (.A(net3842),
    .B(_02106_),
    .C(_02107_),
    .Y(_02108_));
 sg13g2_or3_1 _23994_ (.A(net3479),
    .B(_02105_),
    .C(_02108_),
    .X(_02109_));
 sg13g2_o21ai_1 _23995_ (.B1(net3479),
    .Y(_02110_),
    .A1(_02105_),
    .A2(_02108_));
 sg13g2_nand2_1 _23996_ (.Y(_02111_),
    .A(_02109_),
    .B(_02110_));
 sg13g2_xor2_1 _23997_ (.B(_02111_),
    .A(_02101_),
    .X(_02112_));
 sg13g2_o21ai_1 _23998_ (.B1(net4295),
    .Y(_02113_),
    .A1(_02105_),
    .A2(_02108_));
 sg13g2_nand2_1 _23999_ (.Y(_02114_),
    .A(net3887),
    .B(_02113_));
 sg13g2_a21oi_1 _24000_ (.A1(net4331),
    .A2(_02112_),
    .Y(_02115_),
    .B1(_02114_));
 sg13g2_a21o_1 _24001_ (.A2(net3945),
    .A1(net4804),
    .B1(_02115_),
    .X(_00335_));
 sg13g2_a221oi_1 _24002_ (.B2(_14139_),
    .C1(_14274_),
    .B1(_02082_),
    .A1(_14132_),
    .Y(_02116_),
    .A2(_14272_));
 sg13g2_xnor2_1 _24003_ (.Y(_02117_),
    .A(_14129_),
    .B(_02116_));
 sg13g2_and3_2 _24004_ (.X(_02118_),
    .A(_15516_),
    .B(_15517_),
    .C(_02049_));
 sg13g2_o21ai_1 _24005_ (.B1(_14129_),
    .Y(_02119_),
    .A1(_15523_),
    .A2(_02118_));
 sg13g2_or3_1 _24006_ (.A(_14129_),
    .B(_15523_),
    .C(_02118_),
    .X(_02120_));
 sg13g2_nand3_1 _24007_ (.B(_02119_),
    .C(_02120_),
    .A(net4671),
    .Y(_02121_));
 sg13g2_a21oi_1 _24008_ (.A1(net4562),
    .A2(\u_inv.d_next[60] ),
    .Y(_02122_),
    .B1(net3780));
 sg13g2_a22oi_1 _24009_ (.Y(_02123_),
    .B1(_02121_),
    .B2(_02122_),
    .A2(_02117_),
    .A1(net3780));
 sg13g2_nand2_1 _24010_ (.Y(_02124_),
    .A(net3434),
    .B(_02123_));
 sg13g2_xnor2_1 _24011_ (.Y(_02125_),
    .A(net3434),
    .B(_02123_));
 sg13g2_nand2_1 _24012_ (.Y(_02126_),
    .A(_02091_),
    .B(_02109_));
 sg13g2_and3_2 _24013_ (.X(_02127_),
    .A(_02092_),
    .B(_02109_),
    .C(_02110_));
 sg13g2_a21oi_2 _24014_ (.B1(_02126_),
    .Y(_02128_),
    .A2(_02127_),
    .A1(_02096_));
 sg13g2_xnor2_1 _24015_ (.Y(_02129_),
    .A(_02125_),
    .B(_02128_));
 sg13g2_o21ai_1 _24016_ (.B1(net3887),
    .Y(_02130_),
    .A1(net4344),
    .A2(_02123_));
 sg13g2_a21oi_1 _24017_ (.A1(net4344),
    .A2(_02129_),
    .Y(_02131_),
    .B1(_02130_));
 sg13g2_a21o_1 _24018_ (.A2(net3954),
    .A1(net3219),
    .B1(_02131_),
    .X(_00336_));
 sg13g2_nand2_1 _24019_ (.Y(_02132_),
    .A(net2094),
    .B(net3954));
 sg13g2_o21ai_1 _24020_ (.B1(_02124_),
    .Y(_02133_),
    .A1(_02125_),
    .A2(_02128_));
 sg13g2_nand3_1 _24021_ (.B(_14128_),
    .C(_02119_),
    .A(_14127_),
    .Y(_02134_));
 sg13g2_o21ai_1 _24022_ (.B1(_15514_),
    .Y(_02135_),
    .A1(_15523_),
    .A2(_02118_));
 sg13g2_nor2_1 _24023_ (.A(net4553),
    .B(_15525_),
    .Y(_02136_));
 sg13g2_nand3_1 _24024_ (.B(_02135_),
    .C(_02136_),
    .A(_02134_),
    .Y(_02137_));
 sg13g2_a21oi_1 _24025_ (.A1(net4562),
    .A2(\u_inv.d_next[61] ),
    .Y(_02138_),
    .B1(net3780));
 sg13g2_o21ai_1 _24026_ (.B1(_14277_),
    .Y(_02139_),
    .A1(_14129_),
    .A2(_02116_));
 sg13g2_xnor2_1 _24027_ (.Y(_02140_),
    .A(_14127_),
    .B(_02139_));
 sg13g2_a22oi_1 _24028_ (.Y(_02141_),
    .B1(_02140_),
    .B2(net3780),
    .A2(_02138_),
    .A1(_02137_));
 sg13g2_nand2_1 _24029_ (.Y(_02142_),
    .A(net3434),
    .B(_02141_));
 sg13g2_xnor2_1 _24030_ (.Y(_02143_),
    .A(net3434),
    .B(_02141_));
 sg13g2_o21ai_1 _24031_ (.B1(net4344),
    .Y(_02144_),
    .A1(_02133_),
    .A2(_02143_));
 sg13g2_a21oi_1 _24032_ (.A1(_02133_),
    .A2(_02143_),
    .Y(_02145_),
    .B1(_02144_));
 sg13g2_o21ai_1 _24033_ (.B1(net3887),
    .Y(_02146_),
    .A1(net4344),
    .A2(_02141_));
 sg13g2_o21ai_1 _24034_ (.B1(_02132_),
    .Y(_00337_),
    .A1(_02145_),
    .A2(_02146_));
 sg13g2_o21ai_1 _24035_ (.B1(_14279_),
    .Y(_02147_),
    .A1(_14130_),
    .A2(_02116_));
 sg13g2_xnor2_1 _24036_ (.Y(_02148_),
    .A(_14125_),
    .B(_02147_));
 sg13g2_a21o_1 _24037_ (.A2(_02135_),
    .A1(_15526_),
    .B1(_14125_),
    .X(_02149_));
 sg13g2_nand3_1 _24038_ (.B(_15526_),
    .C(_02135_),
    .A(_14125_),
    .Y(_02150_));
 sg13g2_nand3_1 _24039_ (.B(_02149_),
    .C(_02150_),
    .A(net4671),
    .Y(_02151_));
 sg13g2_a21oi_1 _24040_ (.A1(net4553),
    .A2(\u_inv.d_next[62] ),
    .Y(_02152_),
    .B1(net3772));
 sg13g2_a22oi_1 _24041_ (.Y(_02153_),
    .B1(_02151_),
    .B2(_02152_),
    .A2(_02148_),
    .A1(net3771));
 sg13g2_nand2_1 _24042_ (.Y(_02154_),
    .A(net3426),
    .B(_02153_));
 sg13g2_inv_1 _24043_ (.Y(_02155_),
    .A(_02154_));
 sg13g2_xnor2_1 _24044_ (.Y(_02156_),
    .A(net3477),
    .B(_02153_));
 sg13g2_nand2_1 _24045_ (.Y(_02157_),
    .A(_02124_),
    .B(_02142_));
 sg13g2_nor2_1 _24046_ (.A(_02125_),
    .B(_02143_),
    .Y(_02158_));
 sg13g2_nor2b_1 _24047_ (.A(_02128_),
    .B_N(_02158_),
    .Y(_02159_));
 sg13g2_or2_1 _24048_ (.X(_02160_),
    .B(_02159_),
    .A(_02157_));
 sg13g2_xnor2_1 _24049_ (.Y(_02161_),
    .A(_02156_),
    .B(_02160_));
 sg13g2_a21oi_1 _24050_ (.A1(net4329),
    .A2(_02161_),
    .Y(_02162_),
    .B1(net4235));
 sg13g2_o21ai_1 _24051_ (.B1(_02162_),
    .Y(_02163_),
    .A1(net4329),
    .A2(_02153_));
 sg13g2_o21ai_1 _24052_ (.B1(_02163_),
    .Y(_00338_),
    .A1(_10611_),
    .A2(net4025));
 sg13g2_a21oi_1 _24053_ (.A1(net4562),
    .A2(\u_inv.d_next[63] ),
    .Y(_02164_),
    .B1(net3780));
 sg13g2_nand3_1 _24054_ (.B(_14124_),
    .C(_02149_),
    .A(_14123_),
    .Y(_02165_));
 sg13g2_a21o_1 _24055_ (.A2(_02149_),
    .A1(_14124_),
    .B1(_14123_),
    .X(_02166_));
 sg13g2_nand3_1 _24056_ (.B(_02165_),
    .C(_02166_),
    .A(net4680),
    .Y(_02167_));
 sg13g2_a21oi_1 _24057_ (.A1(_14125_),
    .A2(_02147_),
    .Y(_02168_),
    .B1(_14281_));
 sg13g2_or2_1 _24058_ (.X(_02169_),
    .B(_02168_),
    .A(_14123_));
 sg13g2_a21oi_1 _24059_ (.A1(_14123_),
    .A2(_02168_),
    .Y(_02170_),
    .B1(net3849));
 sg13g2_a22oi_1 _24060_ (.Y(_02171_),
    .B1(_02169_),
    .B2(_02170_),
    .A2(_02167_),
    .A1(_02164_));
 sg13g2_nand2_1 _24061_ (.Y(_02172_),
    .A(net3426),
    .B(_02171_));
 sg13g2_xnor2_1 _24062_ (.Y(_02173_),
    .A(net3478),
    .B(_02171_));
 sg13g2_a21oi_1 _24063_ (.A1(_02156_),
    .A2(_02160_),
    .Y(_02174_),
    .B1(_02155_));
 sg13g2_xor2_1 _24064_ (.B(_02174_),
    .A(_02173_),
    .X(_02175_));
 sg13g2_o21ai_1 _24065_ (.B1(net3886),
    .Y(_02176_),
    .A1(net4330),
    .A2(_02171_));
 sg13g2_a21oi_1 _24066_ (.A1(net4330),
    .A2(_02175_),
    .Y(_02177_),
    .B1(_02176_));
 sg13g2_a21o_1 _24067_ (.A2(net3945),
    .A1(net2665),
    .B1(_02177_),
    .X(_00339_));
 sg13g2_xnor2_1 _24068_ (.Y(_02178_),
    .A(_14530_),
    .B(_15622_));
 sg13g2_o21ai_1 _24069_ (.B1(net3849),
    .Y(_02179_),
    .A1(net4680),
    .A2(\u_inv.d_next[64] ));
 sg13g2_a21oi_1 _24070_ (.A1(net4680),
    .A2(_02178_),
    .Y(_02180_),
    .B1(_02179_));
 sg13g2_a21oi_1 _24071_ (.A1(_14239_),
    .A2(_14301_),
    .Y(_02181_),
    .B1(_14529_));
 sg13g2_nor3_1 _24072_ (.A(_14238_),
    .B(_14302_),
    .C(_14530_),
    .Y(_02182_));
 sg13g2_nor3_1 _24073_ (.A(net3849),
    .B(_02181_),
    .C(_02182_),
    .Y(_02183_));
 sg13g2_nor2_2 _24074_ (.A(_02180_),
    .B(_02183_),
    .Y(_02184_));
 sg13g2_nor2_1 _24075_ (.A(net3478),
    .B(_02184_),
    .Y(_02185_));
 sg13g2_xnor2_1 _24076_ (.Y(_02186_),
    .A(net3431),
    .B(_02184_));
 sg13g2_and2_1 _24077_ (.A(_02095_),
    .B(_02127_),
    .X(_02187_));
 sg13g2_nand4_1 _24078_ (.B(_02158_),
    .C(_02173_),
    .A(_02156_),
    .Y(_02188_),
    .D(_02187_));
 sg13g2_inv_1 _24079_ (.Y(_02189_),
    .A(_02188_));
 sg13g2_nor2_1 _24080_ (.A(_02061_),
    .B(_02188_),
    .Y(_02190_));
 sg13g2_nor3_1 _24081_ (.A(_01926_),
    .B(_02061_),
    .C(_02188_),
    .Y(_02191_));
 sg13g2_o21ai_1 _24082_ (.B1(_02191_),
    .Y(_02192_),
    .A1(_16131_),
    .A2(_16137_));
 sg13g2_a21o_1 _24083_ (.A2(_02127_),
    .A1(_02094_),
    .B1(_02126_),
    .X(_02193_));
 sg13g2_nand4_1 _24084_ (.B(_02158_),
    .C(_02173_),
    .A(_02156_),
    .Y(_02194_),
    .D(_02193_));
 sg13g2_nand3_1 _24085_ (.B(_02157_),
    .C(_02173_),
    .A(_02156_),
    .Y(_02195_));
 sg13g2_nand4_1 _24086_ (.B(_02172_),
    .C(_02194_),
    .A(_02154_),
    .Y(_02196_),
    .D(_02195_));
 sg13g2_a221oi_1 _24087_ (.B2(_01925_),
    .C1(_02196_),
    .B1(_02190_),
    .A1(_02060_),
    .Y(_02197_),
    .A2(_02189_));
 sg13g2_nand2_2 _24088_ (.Y(_02198_),
    .A(_02192_),
    .B(_02197_));
 sg13g2_xor2_1 _24089_ (.B(_02198_),
    .A(_02186_),
    .X(_02199_));
 sg13g2_o21ai_1 _24090_ (.B1(net3890),
    .Y(_02200_),
    .A1(net4295),
    .A2(_02199_));
 sg13g2_a21oi_1 _24091_ (.A1(net4295),
    .A2(_02184_),
    .Y(_02201_),
    .B1(_02200_));
 sg13g2_a21o_1 _24092_ (.A2(net3954),
    .A1(net3114),
    .B1(_02201_),
    .X(_00340_));
 sg13g2_a21oi_1 _24093_ (.A1(_02186_),
    .A2(_02198_),
    .Y(_02202_),
    .B1(_02185_));
 sg13g2_nand3_1 _24094_ (.B(_14529_),
    .C(_15623_),
    .A(_14526_),
    .Y(_02203_));
 sg13g2_nand2_1 _24095_ (.Y(_02204_),
    .A(_14525_),
    .B(_14528_));
 sg13g2_a21oi_1 _24096_ (.A1(_14529_),
    .A2(_15623_),
    .Y(_02205_),
    .B1(_02204_));
 sg13g2_nor3_1 _24097_ (.A(net4562),
    .B(_15364_),
    .C(_02205_),
    .Y(_02206_));
 sg13g2_a22oi_1 _24098_ (.Y(_02207_),
    .B1(_02203_),
    .B2(_02206_),
    .A2(\u_inv.d_next[65] ),
    .A1(net4562));
 sg13g2_nor2_1 _24099_ (.A(_14538_),
    .B(_02181_),
    .Y(_02208_));
 sg13g2_o21ai_1 _24100_ (.B1(net3781),
    .Y(_02209_),
    .A1(_14525_),
    .A2(_02208_));
 sg13g2_a21oi_1 _24101_ (.A1(_14525_),
    .A2(_02208_),
    .Y(_02210_),
    .B1(_02209_));
 sg13g2_a21oi_2 _24102_ (.B1(_02210_),
    .Y(_02211_),
    .A2(_02207_),
    .A1(net3849));
 sg13g2_nand2_1 _24103_ (.Y(_02212_),
    .A(net3431),
    .B(_02211_));
 sg13g2_nor2_1 _24104_ (.A(net3431),
    .B(_02211_),
    .Y(_02213_));
 sg13g2_xnor2_1 _24105_ (.Y(_02214_),
    .A(net3478),
    .B(_02211_));
 sg13g2_xor2_1 _24106_ (.B(_02214_),
    .A(_02202_),
    .X(_02215_));
 sg13g2_o21ai_1 _24107_ (.B1(net3891),
    .Y(_02216_),
    .A1(net4336),
    .A2(_02211_));
 sg13g2_a21oi_1 _24108_ (.A1(net4336),
    .A2(_02215_),
    .Y(_02217_),
    .B1(_02216_));
 sg13g2_a21o_1 _24109_ (.A2(net3954),
    .A1(net3241),
    .B1(_02217_),
    .X(_00341_));
 sg13g2_o21ai_1 _24110_ (.B1(_14539_),
    .Y(_02218_),
    .A1(_14303_),
    .A2(_14531_));
 sg13g2_xor2_1 _24111_ (.B(_02218_),
    .A(_14520_),
    .X(_02219_));
 sg13g2_nor2_1 _24112_ (.A(net3849),
    .B(_02219_),
    .Y(_02220_));
 sg13g2_a21o_1 _24113_ (.A2(_02203_),
    .A1(_15365_),
    .B1(_14520_),
    .X(_02221_));
 sg13g2_nand3_1 _24114_ (.B(_15365_),
    .C(_02203_),
    .A(_14520_),
    .Y(_02222_));
 sg13g2_nand3_1 _24115_ (.B(_02221_),
    .C(_02222_),
    .A(net4680),
    .Y(_02223_));
 sg13g2_a21oi_1 _24116_ (.A1(net4562),
    .A2(\u_inv.d_next[66] ),
    .Y(_02224_),
    .B1(net3781));
 sg13g2_a21o_2 _24117_ (.A2(_02224_),
    .A1(_02223_),
    .B1(_02220_),
    .X(_02225_));
 sg13g2_nor2_1 _24118_ (.A(net3477),
    .B(_02225_),
    .Y(_02226_));
 sg13g2_nand2_1 _24119_ (.Y(_02227_),
    .A(net3477),
    .B(_02225_));
 sg13g2_xnor2_1 _24120_ (.Y(_02228_),
    .A(net3478),
    .B(_02225_));
 sg13g2_nand2b_1 _24121_ (.Y(_02229_),
    .B(_02212_),
    .A_N(_02185_));
 sg13g2_o21ai_1 _24122_ (.B1(_02212_),
    .Y(_02230_),
    .A1(_02202_),
    .A2(_02213_));
 sg13g2_xnor2_1 _24123_ (.Y(_02231_),
    .A(_02228_),
    .B(_02230_));
 sg13g2_o21ai_1 _24124_ (.B1(net3891),
    .Y(_02232_),
    .A1(net4295),
    .A2(_02231_));
 sg13g2_a21oi_1 _24125_ (.A1(net4295),
    .A2(_02225_),
    .Y(_02233_),
    .B1(_02232_));
 sg13g2_a21o_1 _24126_ (.A2(net3954),
    .A1(net2607),
    .B1(_02233_),
    .X(_00342_));
 sg13g2_a21oi_1 _24127_ (.A1(_02227_),
    .A2(_02230_),
    .Y(_02234_),
    .B1(_02226_));
 sg13g2_a21oi_1 _24128_ (.A1(net4567),
    .A2(\u_inv.d_next[67] ),
    .Y(_02235_),
    .B1(net3781));
 sg13g2_a21o_1 _24129_ (.A2(_02221_),
    .A1(_14518_),
    .B1(_14517_),
    .X(_02236_));
 sg13g2_nand3_1 _24130_ (.B(_14518_),
    .C(_02221_),
    .A(_14517_),
    .Y(_02237_));
 sg13g2_nand3_1 _24131_ (.B(_02236_),
    .C(_02237_),
    .A(net4688),
    .Y(_02238_));
 sg13g2_and2_1 _24132_ (.A(_02235_),
    .B(_02238_),
    .X(_02239_));
 sg13g2_a21oi_1 _24133_ (.A1(_14520_),
    .A2(_02218_),
    .Y(_02240_),
    .B1(_14541_));
 sg13g2_or2_1 _24134_ (.X(_02241_),
    .B(_02240_),
    .A(_14517_));
 sg13g2_a21oi_1 _24135_ (.A1(_14517_),
    .A2(_02240_),
    .Y(_02242_),
    .B1(net3850));
 sg13g2_a22oi_1 _24136_ (.Y(_02243_),
    .B1(_02241_),
    .B2(_02242_),
    .A2(_02238_),
    .A1(_02235_));
 sg13g2_a21o_1 _24137_ (.A2(_02242_),
    .A1(_02241_),
    .B1(_02239_),
    .X(_02244_));
 sg13g2_xnor2_1 _24138_ (.Y(_02245_),
    .A(net3434),
    .B(_02243_));
 sg13g2_xnor2_1 _24139_ (.Y(_02246_),
    .A(_02234_),
    .B(_02245_));
 sg13g2_nand2_1 _24140_ (.Y(_02247_),
    .A(net4336),
    .B(_02246_));
 sg13g2_a21oi_1 _24141_ (.A1(net4295),
    .A2(_02244_),
    .Y(_02248_),
    .B1(net4237));
 sg13g2_a22oi_1 _24142_ (.Y(_02249_),
    .B1(_02247_),
    .B2(_02248_),
    .A2(net3954),
    .A1(net2948));
 sg13g2_inv_1 _24143_ (.Y(_00343_),
    .A(_02249_));
 sg13g2_a21oi_2 _24144_ (.B1(_14543_),
    .Y(_02250_),
    .A2(_02218_),
    .A1(_14521_));
 sg13g2_xnor2_1 _24145_ (.Y(_02251_),
    .A(_14514_),
    .B(_02250_));
 sg13g2_a21oi_1 _24146_ (.A1(_15623_),
    .A2(_15624_),
    .Y(_02252_),
    .B1(_15368_));
 sg13g2_nor2b_1 _24147_ (.A(_02252_),
    .B_N(_14514_),
    .Y(_02253_));
 sg13g2_nand2b_1 _24148_ (.Y(_02254_),
    .B(_02252_),
    .A_N(_14514_));
 sg13g2_nand3b_1 _24149_ (.B(_02254_),
    .C(net4680),
    .Y(_02255_),
    .A_N(_02253_));
 sg13g2_a21oi_1 _24150_ (.A1(net4562),
    .A2(\u_inv.d_next[68] ),
    .Y(_02256_),
    .B1(net3780));
 sg13g2_a22oi_1 _24151_ (.Y(_02257_),
    .B1(_02255_),
    .B2(_02256_),
    .A2(_02251_),
    .A1(net3780));
 sg13g2_nand2_1 _24152_ (.Y(_02258_),
    .A(net3433),
    .B(_02257_));
 sg13g2_xnor2_1 _24153_ (.Y(_02259_),
    .A(net3433),
    .B(_02257_));
 sg13g2_a21oi_1 _24154_ (.A1(_02225_),
    .A2(_02244_),
    .Y(_02260_),
    .B1(net3477));
 sg13g2_nor2_1 _24155_ (.A(_02228_),
    .B(_02245_),
    .Y(_02261_));
 sg13g2_a21o_2 _24156_ (.A2(_02261_),
    .A1(_02230_),
    .B1(_02260_),
    .X(_02262_));
 sg13g2_nand2b_1 _24157_ (.Y(_02263_),
    .B(_02262_),
    .A_N(_02259_));
 sg13g2_xor2_1 _24158_ (.B(_02262_),
    .A(_02259_),
    .X(_02264_));
 sg13g2_a21oi_1 _24159_ (.A1(net4343),
    .A2(_02264_),
    .Y(_02265_),
    .B1(net4237));
 sg13g2_o21ai_1 _24160_ (.B1(_02265_),
    .Y(_02266_),
    .A1(net4344),
    .A2(_02257_));
 sg13g2_o21ai_1 _24161_ (.B1(_02266_),
    .Y(_00344_),
    .A1(_10610_),
    .A2(net4029));
 sg13g2_a21oi_1 _24162_ (.A1(net4562),
    .A2(net4803),
    .Y(_02267_),
    .B1(net3781));
 sg13g2_a21o_1 _24163_ (.A2(\u_inv.d_reg[68] ),
    .A1(\u_inv.d_next[68] ),
    .B1(_02253_),
    .X(_02268_));
 sg13g2_o21ai_1 _24164_ (.B1(net4680),
    .Y(_02269_),
    .A1(_14512_),
    .A2(_02268_));
 sg13g2_a21o_1 _24165_ (.A2(_02268_),
    .A1(_14512_),
    .B1(_02269_),
    .X(_02270_));
 sg13g2_o21ai_1 _24166_ (.B1(_14547_),
    .Y(_02271_),
    .A1(_14514_),
    .A2(_02250_));
 sg13g2_nand2b_1 _24167_ (.Y(_02272_),
    .B(_14513_),
    .A_N(_02271_));
 sg13g2_a21oi_1 _24168_ (.A1(_14512_),
    .A2(_02271_),
    .Y(_02273_),
    .B1(net3849));
 sg13g2_a22oi_1 _24169_ (.Y(_02274_),
    .B1(_02272_),
    .B2(_02273_),
    .A2(_02270_),
    .A1(_02267_));
 sg13g2_nand2_1 _24170_ (.Y(_02275_),
    .A(net3433),
    .B(_02274_));
 sg13g2_xnor2_1 _24171_ (.Y(_02276_),
    .A(net3479),
    .B(_02274_));
 sg13g2_nand2_1 _24172_ (.Y(_02277_),
    .A(_02258_),
    .B(_02263_));
 sg13g2_xnor2_1 _24173_ (.Y(_02278_),
    .A(_02276_),
    .B(_02277_));
 sg13g2_o21ai_1 _24174_ (.B1(net3894),
    .Y(_02279_),
    .A1(net4343),
    .A2(_02274_));
 sg13g2_a21oi_1 _24175_ (.A1(net4344),
    .A2(_02278_),
    .Y(_02280_),
    .B1(_02279_));
 sg13g2_a21o_1 _24176_ (.A2(net3953),
    .A1(net3150),
    .B1(_02280_),
    .X(_00345_));
 sg13g2_o21ai_1 _24177_ (.B1(_14549_),
    .Y(_02281_),
    .A1(_14515_),
    .A2(_02250_));
 sg13g2_xnor2_1 _24178_ (.Y(_02282_),
    .A(_14509_),
    .B(_02281_));
 sg13g2_nor2_1 _24179_ (.A(_15360_),
    .B(_02252_),
    .Y(_02283_));
 sg13g2_nor2_1 _24180_ (.A(_15370_),
    .B(_02283_),
    .Y(_02284_));
 sg13g2_a21oi_1 _24181_ (.A1(_14509_),
    .A2(_02284_),
    .Y(_02285_),
    .B1(net4566));
 sg13g2_o21ai_1 _24182_ (.B1(_02285_),
    .Y(_02286_),
    .A1(_14509_),
    .A2(_02284_));
 sg13g2_a21oi_1 _24183_ (.A1(net4566),
    .A2(\u_inv.d_next[70] ),
    .Y(_02287_),
    .B1(net3785));
 sg13g2_a22oi_1 _24184_ (.Y(_02288_),
    .B1(_02286_),
    .B2(_02287_),
    .A2(_02282_),
    .A1(net3785));
 sg13g2_and2_1 _24185_ (.A(net3433),
    .B(_02288_),
    .X(_02289_));
 sg13g2_xnor2_1 _24186_ (.Y(_02290_),
    .A(net3479),
    .B(_02288_));
 sg13g2_nand2_1 _24187_ (.Y(_02291_),
    .A(_02258_),
    .B(_02275_));
 sg13g2_nor2b_1 _24188_ (.A(_02259_),
    .B_N(_02276_),
    .Y(_02292_));
 sg13g2_a21oi_1 _24189_ (.A1(_02262_),
    .A2(_02292_),
    .Y(_02293_),
    .B1(_02291_));
 sg13g2_inv_1 _24190_ (.Y(_02294_),
    .A(_02293_));
 sg13g2_xnor2_1 _24191_ (.Y(_02295_),
    .A(_02290_),
    .B(_02293_));
 sg13g2_nor2_1 _24192_ (.A(net4343),
    .B(_02288_),
    .Y(_02296_));
 sg13g2_o21ai_1 _24193_ (.B1(net3890),
    .Y(_02297_),
    .A1(net4295),
    .A2(_02295_));
 sg13g2_nand2_1 _24194_ (.Y(_02298_),
    .A(net4803),
    .B(net3954));
 sg13g2_o21ai_1 _24195_ (.B1(_02298_),
    .Y(_00346_),
    .A1(_02296_),
    .A2(_02297_));
 sg13g2_nand2_1 _24196_ (.Y(_02299_),
    .A(net2374),
    .B(net3956));
 sg13g2_a21oi_1 _24197_ (.A1(net4566),
    .A2(\u_inv.d_next[71] ),
    .Y(_02300_),
    .B1(net3785));
 sg13g2_o21ai_1 _24198_ (.B1(_14507_),
    .Y(_02301_),
    .A1(_14509_),
    .A2(_02284_));
 sg13g2_xnor2_1 _24199_ (.Y(_02302_),
    .A(_14506_),
    .B(_02301_));
 sg13g2_nand2_1 _24200_ (.Y(_02303_),
    .A(net4682),
    .B(_02302_));
 sg13g2_a21oi_1 _24201_ (.A1(_14509_),
    .A2(_02281_),
    .Y(_02304_),
    .B1(_14546_));
 sg13g2_or2_1 _24202_ (.X(_02305_),
    .B(_02304_),
    .A(_14506_));
 sg13g2_a21oi_1 _24203_ (.A1(_14506_),
    .A2(_02304_),
    .Y(_02306_),
    .B1(net3858));
 sg13g2_a22oi_1 _24204_ (.Y(_02307_),
    .B1(_02305_),
    .B2(_02306_),
    .A2(_02303_),
    .A1(_02300_));
 sg13g2_xnor2_1 _24205_ (.Y(_02308_),
    .A(net3479),
    .B(_02307_));
 sg13g2_a21oi_1 _24206_ (.A1(_02290_),
    .A2(_02294_),
    .Y(_02309_),
    .B1(_02289_));
 sg13g2_o21ai_1 _24207_ (.B1(net4341),
    .Y(_02310_),
    .A1(_02308_),
    .A2(_02309_));
 sg13g2_a21oi_1 _24208_ (.A1(_02308_),
    .A2(_02309_),
    .Y(_02311_),
    .B1(_02310_));
 sg13g2_o21ai_1 _24209_ (.B1(net3894),
    .Y(_02312_),
    .A1(net4343),
    .A2(_02307_));
 sg13g2_o21ai_1 _24210_ (.B1(_02299_),
    .Y(_00347_),
    .A1(_02311_),
    .A2(_02312_));
 sg13g2_a21o_1 _24211_ (.A2(_14301_),
    .A1(_14239_),
    .B1(_14532_),
    .X(_02313_));
 sg13g2_nand2_1 _24212_ (.Y(_02314_),
    .A(_14552_),
    .B(_02313_));
 sg13g2_xnor2_1 _24213_ (.Y(_02315_),
    .A(_14500_),
    .B(_02314_));
 sg13g2_a21o_2 _24214_ (.A2(_15625_),
    .A1(_15623_),
    .B1(_15375_),
    .X(_02316_));
 sg13g2_nor2b_1 _24215_ (.A(_14500_),
    .B_N(_02316_),
    .Y(_02317_));
 sg13g2_nand2b_1 _24216_ (.Y(_02318_),
    .B(_14500_),
    .A_N(_02316_));
 sg13g2_nand3b_1 _24217_ (.B(_02318_),
    .C(net4682),
    .Y(_02319_),
    .A_N(_02317_));
 sg13g2_a21oi_1 _24218_ (.A1(net4566),
    .A2(\u_inv.d_next[72] ),
    .Y(_02320_),
    .B1(net3785));
 sg13g2_a22oi_1 _24219_ (.Y(_02321_),
    .B1(_02319_),
    .B2(_02320_),
    .A2(_02315_),
    .A1(net3785));
 sg13g2_xnor2_1 _24220_ (.Y(_02322_),
    .A(net3434),
    .B(_02321_));
 sg13g2_a21o_1 _24221_ (.A2(_02261_),
    .A1(_02229_),
    .B1(_02260_),
    .X(_02323_));
 sg13g2_nand4_1 _24222_ (.B(_02292_),
    .C(_02308_),
    .A(_02290_),
    .Y(_02324_),
    .D(_02323_));
 sg13g2_a21oi_1 _24223_ (.A1(net3433),
    .A2(_02307_),
    .Y(_02325_),
    .B1(_02289_));
 sg13g2_nand3_1 _24224_ (.B(_02291_),
    .C(_02308_),
    .A(_02290_),
    .Y(_02326_));
 sg13g2_nand3_1 _24225_ (.B(_02325_),
    .C(_02326_),
    .A(_02324_),
    .Y(_02327_));
 sg13g2_and3_1 _24226_ (.X(_02328_),
    .A(_02186_),
    .B(_02214_),
    .C(_02261_));
 sg13g2_and4_1 _24227_ (.A(_02290_),
    .B(_02292_),
    .C(_02308_),
    .D(_02328_),
    .X(_02329_));
 sg13g2_a21oi_1 _24228_ (.A1(_02198_),
    .A2(_02329_),
    .Y(_02330_),
    .B1(_02327_));
 sg13g2_nor2_1 _24229_ (.A(_02322_),
    .B(_02330_),
    .Y(_02331_));
 sg13g2_xnor2_1 _24230_ (.Y(_02332_),
    .A(_02322_),
    .B(_02330_));
 sg13g2_o21ai_1 _24231_ (.B1(net3894),
    .Y(_02333_),
    .A1(net4343),
    .A2(_02321_));
 sg13g2_a21oi_1 _24232_ (.A1(net4343),
    .A2(_02332_),
    .Y(_02334_),
    .B1(_02333_));
 sg13g2_a21o_1 _24233_ (.A2(net3956),
    .A1(net2787),
    .B1(_02334_),
    .X(_00348_));
 sg13g2_a21oi_1 _24234_ (.A1(net4566),
    .A2(\u_inv.d_next[73] ),
    .Y(_02335_),
    .B1(net3785));
 sg13g2_a21oi_1 _24235_ (.A1(\u_inv.d_next[72] ),
    .A2(\u_inv.d_reg[72] ),
    .Y(_02336_),
    .B1(_02317_));
 sg13g2_xnor2_1 _24236_ (.Y(_02337_),
    .A(_14499_),
    .B(_02336_));
 sg13g2_nand2_1 _24237_ (.Y(_02338_),
    .A(net4682),
    .B(_02337_));
 sg13g2_a21o_1 _24238_ (.A2(_02314_),
    .A1(_14500_),
    .B1(_14561_),
    .X(_02339_));
 sg13g2_o21ai_1 _24239_ (.B1(net3785),
    .Y(_02340_),
    .A1(_14499_),
    .A2(_02339_));
 sg13g2_a21oi_1 _24240_ (.A1(_14499_),
    .A2(_02339_),
    .Y(_02341_),
    .B1(_02340_));
 sg13g2_a21oi_2 _24241_ (.B1(_02341_),
    .Y(_02342_),
    .A2(_02338_),
    .A1(_02335_));
 sg13g2_xnor2_1 _24242_ (.Y(_02343_),
    .A(net3433),
    .B(_02342_));
 sg13g2_a21oi_1 _24243_ (.A1(net3433),
    .A2(_02321_),
    .Y(_02344_),
    .B1(_02331_));
 sg13g2_xnor2_1 _24244_ (.Y(_02345_),
    .A(_02343_),
    .B(_02344_));
 sg13g2_o21ai_1 _24245_ (.B1(net3894),
    .Y(_02346_),
    .A1(net4343),
    .A2(_02342_));
 sg13g2_a21oi_1 _24246_ (.A1(net4344),
    .A2(_02345_),
    .Y(_02347_),
    .B1(_02346_));
 sg13g2_a21o_1 _24247_ (.A2(net3956),
    .A1(net3058),
    .B1(_02347_),
    .X(_00349_));
 sg13g2_a21oi_2 _24248_ (.B1(_14501_),
    .Y(_02348_),
    .A2(_02313_),
    .A1(_14552_));
 sg13g2_nor2_1 _24249_ (.A(_14563_),
    .B(_02348_),
    .Y(_02349_));
 sg13g2_o21ai_1 _24250_ (.B1(_14495_),
    .Y(_02350_),
    .A1(_14563_),
    .A2(_02348_));
 sg13g2_xnor2_1 _24251_ (.Y(_02351_),
    .A(_14494_),
    .B(_02349_));
 sg13g2_a21oi_1 _24252_ (.A1(_15356_),
    .A2(_02316_),
    .Y(_02352_),
    .B1(_15382_));
 sg13g2_a21oi_1 _24253_ (.A1(_14495_),
    .A2(_02352_),
    .Y(_02353_),
    .B1(net4566));
 sg13g2_o21ai_1 _24254_ (.B1(_02353_),
    .Y(_02354_),
    .A1(_14495_),
    .A2(_02352_));
 sg13g2_a21oi_1 _24255_ (.A1(net4566),
    .A2(\u_inv.d_next[74] ),
    .Y(_02355_),
    .B1(net3785));
 sg13g2_a22oi_1 _24256_ (.Y(_02356_),
    .B1(_02354_),
    .B2(_02355_),
    .A2(_02351_),
    .A1(net3786));
 sg13g2_nand2_1 _24257_ (.Y(_02357_),
    .A(net3442),
    .B(_02356_));
 sg13g2_nor2_1 _24258_ (.A(net3442),
    .B(_02356_),
    .Y(_02358_));
 sg13g2_xnor2_1 _24259_ (.Y(_02359_),
    .A(net3482),
    .B(_02356_));
 sg13g2_o21ai_1 _24260_ (.B1(net3433),
    .Y(_02360_),
    .A1(_02321_),
    .A2(_02342_));
 sg13g2_nor3_1 _24261_ (.A(_02322_),
    .B(_02330_),
    .C(_02343_),
    .Y(_02361_));
 sg13g2_nor2b_1 _24262_ (.A(_02361_),
    .B_N(_02360_),
    .Y(_02362_));
 sg13g2_xnor2_1 _24263_ (.Y(_02363_),
    .A(_02359_),
    .B(_02362_));
 sg13g2_nor2_1 _24264_ (.A(net4343),
    .B(_02356_),
    .Y(_02364_));
 sg13g2_o21ai_1 _24265_ (.B1(net3894),
    .Y(_02365_),
    .A1(net4296),
    .A2(_02363_));
 sg13g2_nand2_1 _24266_ (.Y(_02366_),
    .A(net2315),
    .B(net3956));
 sg13g2_o21ai_1 _24267_ (.B1(_02366_),
    .Y(_00350_),
    .A1(_02364_),
    .A2(_02365_));
 sg13g2_o21ai_1 _24268_ (.B1(_02357_),
    .Y(_02367_),
    .A1(_02358_),
    .A2(_02362_));
 sg13g2_nand2_1 _24269_ (.Y(_02368_),
    .A(_10609_),
    .B(net3850));
 sg13g2_o21ai_1 _24270_ (.B1(_14492_),
    .Y(_02369_),
    .A1(_14495_),
    .A2(_02352_));
 sg13g2_xnor2_1 _24271_ (.Y(_02370_),
    .A(_14490_),
    .B(_02369_));
 sg13g2_a22oi_1 _24272_ (.Y(_02371_),
    .B1(_02370_),
    .B2(net4682),
    .A2(_02368_),
    .A1(net3730));
 sg13g2_a21oi_1 _24273_ (.A1(_14564_),
    .A2(_02350_),
    .Y(_02372_),
    .B1(_14490_));
 sg13g2_and3_1 _24274_ (.X(_02373_),
    .A(_14490_),
    .B(_14564_),
    .C(_02350_));
 sg13g2_nor3_1 _24275_ (.A(net3850),
    .B(_02372_),
    .C(_02373_),
    .Y(_02374_));
 sg13g2_or3_1 _24276_ (.A(net3482),
    .B(_02371_),
    .C(_02374_),
    .X(_02375_));
 sg13g2_inv_1 _24277_ (.Y(_02376_),
    .A(_02375_));
 sg13g2_o21ai_1 _24278_ (.B1(net3482),
    .Y(_02377_),
    .A1(_02371_),
    .A2(_02374_));
 sg13g2_nand2_1 _24279_ (.Y(_02378_),
    .A(_02375_),
    .B(_02377_));
 sg13g2_xor2_1 _24280_ (.B(_02378_),
    .A(_02367_),
    .X(_02379_));
 sg13g2_o21ai_1 _24281_ (.B1(net4296),
    .Y(_02380_),
    .A1(_02371_),
    .A2(_02374_));
 sg13g2_nand2_1 _24282_ (.Y(_02381_),
    .A(net3894),
    .B(_02380_));
 sg13g2_a21oi_1 _24283_ (.A1(net4354),
    .A2(_02379_),
    .Y(_02382_),
    .B1(_02381_));
 sg13g2_a21o_1 _24284_ (.A2(net3956),
    .A1(net3211),
    .B1(_02382_),
    .X(_00351_));
 sg13g2_a21oi_2 _24285_ (.B1(_14567_),
    .Y(_02383_),
    .A2(_02348_),
    .A1(_14496_));
 sg13g2_xnor2_1 _24286_ (.Y(_02384_),
    .A(_14486_),
    .B(_02383_));
 sg13g2_a21oi_1 _24287_ (.A1(_15358_),
    .A2(_02316_),
    .Y(_02385_),
    .B1(_15385_));
 sg13g2_a21o_1 _24288_ (.A2(_02316_),
    .A1(_15358_),
    .B1(_15385_),
    .X(_02386_));
 sg13g2_a21oi_1 _24289_ (.A1(_14487_),
    .A2(_02385_),
    .Y(_02387_),
    .B1(net4572));
 sg13g2_o21ai_1 _24290_ (.B1(_02387_),
    .Y(_02388_),
    .A1(_14487_),
    .A2(_02385_));
 sg13g2_a21oi_1 _24291_ (.A1(net4572),
    .A2(\u_inv.d_next[76] ),
    .Y(_02389_),
    .B1(net3790));
 sg13g2_a22oi_1 _24292_ (.Y(_02390_),
    .B1(_02388_),
    .B2(_02389_),
    .A2(_02384_),
    .A1(net3790));
 sg13g2_nand2_1 _24293_ (.Y(_02391_),
    .A(net3442),
    .B(_02390_));
 sg13g2_xnor2_1 _24294_ (.Y(_02392_),
    .A(net3442),
    .B(_02390_));
 sg13g2_and2_1 _24295_ (.A(_02357_),
    .B(_02375_),
    .X(_02393_));
 sg13g2_nand3_1 _24296_ (.B(_02375_),
    .C(_02377_),
    .A(_02359_),
    .Y(_02394_));
 sg13g2_a21oi_1 _24297_ (.A1(_02367_),
    .A2(_02377_),
    .Y(_02395_),
    .B1(_02376_));
 sg13g2_xnor2_1 _24298_ (.Y(_02396_),
    .A(_02392_),
    .B(_02395_));
 sg13g2_a21oi_1 _24299_ (.A1(net4354),
    .A2(_02396_),
    .Y(_02397_),
    .B1(net4237));
 sg13g2_o21ai_1 _24300_ (.B1(_02397_),
    .Y(_02398_),
    .A1(net4354),
    .A2(_02390_));
 sg13g2_o21ai_1 _24301_ (.B1(_02398_),
    .Y(_00352_),
    .A1(_10609_),
    .A2(net4029));
 sg13g2_nand2_1 _24302_ (.Y(_02399_),
    .A(net2716),
    .B(net3956));
 sg13g2_a21oi_1 _24303_ (.A1(net4572),
    .A2(\u_inv.d_next[77] ),
    .Y(_02400_),
    .B1(net3790));
 sg13g2_o21ai_1 _24304_ (.B1(_14485_),
    .Y(_02401_),
    .A1(_14487_),
    .A2(_02385_));
 sg13g2_a21oi_1 _24305_ (.A1(_14483_),
    .A2(_02401_),
    .Y(_02402_),
    .B1(net4572));
 sg13g2_o21ai_1 _24306_ (.B1(_02402_),
    .Y(_02403_),
    .A1(_14483_),
    .A2(_02401_));
 sg13g2_o21ai_1 _24307_ (.B1(_14555_),
    .Y(_02404_),
    .A1(_14486_),
    .A2(_02383_));
 sg13g2_nand2b_1 _24308_ (.Y(_02405_),
    .B(_14484_),
    .A_N(_02404_));
 sg13g2_a21oi_1 _24309_ (.A1(_14483_),
    .A2(_02404_),
    .Y(_02406_),
    .B1(net3854));
 sg13g2_a22oi_1 _24310_ (.Y(_02407_),
    .B1(_02405_),
    .B2(_02406_),
    .A2(_02403_),
    .A1(_02400_));
 sg13g2_and2_1 _24311_ (.A(net3442),
    .B(_02407_),
    .X(_02408_));
 sg13g2_nand2b_1 _24312_ (.Y(_02409_),
    .B(net3482),
    .A_N(_02407_));
 sg13g2_xnor2_1 _24313_ (.Y(_02410_),
    .A(net3442),
    .B(_02407_));
 sg13g2_o21ai_1 _24314_ (.B1(_02391_),
    .Y(_02411_),
    .A1(_02392_),
    .A2(_02395_));
 sg13g2_o21ai_1 _24315_ (.B1(net4354),
    .Y(_02412_),
    .A1(_02410_),
    .A2(_02411_));
 sg13g2_a21oi_1 _24316_ (.A1(_02410_),
    .A2(_02411_),
    .Y(_02413_),
    .B1(_02412_));
 sg13g2_o21ai_1 _24317_ (.B1(net3894),
    .Y(_02414_),
    .A1(net4354),
    .A2(_02407_));
 sg13g2_o21ai_1 _24318_ (.B1(_02399_),
    .Y(_00353_),
    .A1(_02413_),
    .A2(_02414_));
 sg13g2_o21ai_1 _24319_ (.B1(_14557_),
    .Y(_02415_),
    .A1(_14488_),
    .A2(_02383_));
 sg13g2_xnor2_1 _24320_ (.Y(_02416_),
    .A(_14480_),
    .B(_02415_));
 sg13g2_a21oi_1 _24321_ (.A1(_15353_),
    .A2(_02386_),
    .Y(_02417_),
    .B1(_15377_));
 sg13g2_a21oi_1 _24322_ (.A1(_14480_),
    .A2(_02417_),
    .Y(_02418_),
    .B1(net4572));
 sg13g2_o21ai_1 _24323_ (.B1(_02418_),
    .Y(_02419_),
    .A1(_14480_),
    .A2(_02417_));
 sg13g2_a21oi_1 _24324_ (.A1(net4572),
    .A2(\u_inv.d_next[78] ),
    .Y(_02420_),
    .B1(net3790));
 sg13g2_a22oi_1 _24325_ (.Y(_02421_),
    .B1(_02419_),
    .B2(_02420_),
    .A2(_02416_),
    .A1(net3790));
 sg13g2_xnor2_1 _24326_ (.Y(_02422_),
    .A(net3482),
    .B(_02421_));
 sg13g2_a21o_1 _24327_ (.A2(_02390_),
    .A1(net3442),
    .B1(_02408_),
    .X(_02423_));
 sg13g2_a21o_1 _24328_ (.A2(_02411_),
    .A1(_02409_),
    .B1(_02408_),
    .X(_02424_));
 sg13g2_and2_1 _24329_ (.A(_02422_),
    .B(_02424_),
    .X(_02425_));
 sg13g2_xnor2_1 _24330_ (.Y(_02426_),
    .A(_02422_),
    .B(_02424_));
 sg13g2_o21ai_1 _24331_ (.B1(net3894),
    .Y(_02427_),
    .A1(net4354),
    .A2(_02421_));
 sg13g2_a21oi_1 _24332_ (.A1(net4354),
    .A2(_02426_),
    .Y(_02428_),
    .B1(_02427_));
 sg13g2_a21o_1 _24333_ (.A2(net3966),
    .A1(net3267),
    .B1(_02428_),
    .X(_00354_));
 sg13g2_a21oi_1 _24334_ (.A1(net4572),
    .A2(\u_inv.d_next[79] ),
    .Y(_02429_),
    .B1(net3790));
 sg13g2_o21ai_1 _24335_ (.B1(_14479_),
    .Y(_02430_),
    .A1(_14480_),
    .A2(_02417_));
 sg13g2_xnor2_1 _24336_ (.Y(_02431_),
    .A(_14477_),
    .B(_02430_));
 sg13g2_nand2_1 _24337_ (.Y(_02432_),
    .A(net4692),
    .B(_02431_));
 sg13g2_a21oi_1 _24338_ (.A1(_14480_),
    .A2(_02415_),
    .Y(_02433_),
    .B1(_14558_));
 sg13g2_or2_1 _24339_ (.X(_02434_),
    .B(_02433_),
    .A(_14477_));
 sg13g2_a21oi_1 _24340_ (.A1(_14477_),
    .A2(_02433_),
    .Y(_02435_),
    .B1(net3853));
 sg13g2_a22oi_1 _24341_ (.Y(_02436_),
    .B1(_02434_),
    .B2(_02435_),
    .A2(_02432_),
    .A1(_02429_));
 sg13g2_xnor2_1 _24342_ (.Y(_02437_),
    .A(net3482),
    .B(_02436_));
 sg13g2_a21o_1 _24343_ (.A2(_02421_),
    .A1(net3442),
    .B1(_02425_),
    .X(_02438_));
 sg13g2_xnor2_1 _24344_ (.Y(_02439_),
    .A(_02437_),
    .B(_02438_));
 sg13g2_o21ai_1 _24345_ (.B1(net3895),
    .Y(_02440_),
    .A1(net4354),
    .A2(_02436_));
 sg13g2_a21oi_1 _24346_ (.A1(net4346),
    .A2(_02439_),
    .Y(_02441_),
    .B1(_02440_));
 sg13g2_a21o_1 _24347_ (.A2(net3966),
    .A1(net2829),
    .B1(_02441_),
    .X(_00355_));
 sg13g2_a21o_2 _24348_ (.A2(_14301_),
    .A1(_14239_),
    .B1(_14533_),
    .X(_02442_));
 sg13g2_nand2_1 _24349_ (.Y(_02443_),
    .A(_14569_),
    .B(_02442_));
 sg13g2_xnor2_1 _24350_ (.Y(_02444_),
    .A(_14469_),
    .B(_02443_));
 sg13g2_o21ai_1 _24351_ (.B1(_15387_),
    .Y(_02445_),
    .A1(_15622_),
    .A2(_15626_));
 sg13g2_nand2_1 _24352_ (.Y(_02446_),
    .A(_14468_),
    .B(_02445_));
 sg13g2_o21ai_1 _24353_ (.B1(net4681),
    .Y(_02447_),
    .A1(_14468_),
    .A2(_02445_));
 sg13g2_nand2b_1 _24354_ (.Y(_02448_),
    .B(_02446_),
    .A_N(_02447_));
 sg13g2_a21oi_1 _24355_ (.A1(net4566),
    .A2(\u_inv.d_next[80] ),
    .Y(_02449_),
    .B1(net3786));
 sg13g2_a22oi_1 _24356_ (.Y(_02450_),
    .B1(_02448_),
    .B2(_02449_),
    .A2(_02444_),
    .A1(net3786));
 sg13g2_nand2_1 _24357_ (.Y(_02451_),
    .A(net3429),
    .B(_02450_));
 sg13g2_xnor2_1 _24358_ (.Y(_02452_),
    .A(net3429),
    .B(_02450_));
 sg13g2_nor2_1 _24359_ (.A(_02392_),
    .B(_02410_),
    .Y(_02453_));
 sg13g2_nor3_1 _24360_ (.A(_02322_),
    .B(_02343_),
    .C(_02394_),
    .Y(_02454_));
 sg13g2_and4_1 _24361_ (.A(_02422_),
    .B(_02437_),
    .C(_02453_),
    .D(_02454_),
    .X(_02455_));
 sg13g2_o21ai_1 _24362_ (.B1(_02393_),
    .Y(_02456_),
    .A1(_02360_),
    .A2(_02394_));
 sg13g2_nand4_1 _24363_ (.B(_02437_),
    .C(_02453_),
    .A(_02422_),
    .Y(_02457_),
    .D(_02456_));
 sg13g2_o21ai_1 _24364_ (.B1(net3446),
    .Y(_02458_),
    .A1(_02421_),
    .A2(_02436_));
 sg13g2_nand3_1 _24365_ (.B(_02423_),
    .C(_02437_),
    .A(_02422_),
    .Y(_02459_));
 sg13g2_nand3_1 _24366_ (.B(_02458_),
    .C(_02459_),
    .A(_02457_),
    .Y(_02460_));
 sg13g2_a21o_1 _24367_ (.A2(_02455_),
    .A1(_02327_),
    .B1(_02460_),
    .X(_02461_));
 sg13g2_and2_1 _24368_ (.A(_02329_),
    .B(_02455_),
    .X(_02462_));
 sg13g2_a21oi_1 _24369_ (.A1(_02198_),
    .A2(_02462_),
    .Y(_02463_),
    .B1(_02461_));
 sg13g2_or2_1 _24370_ (.X(_02464_),
    .B(_02463_),
    .A(_02452_));
 sg13g2_xnor2_1 _24371_ (.Y(_02465_),
    .A(_02452_),
    .B(_02463_));
 sg13g2_o21ai_1 _24372_ (.B1(net3893),
    .Y(_02466_),
    .A1(net4341),
    .A2(_02450_));
 sg13g2_a21oi_1 _24373_ (.A1(net4341),
    .A2(_02465_),
    .Y(_02467_),
    .B1(_02466_));
 sg13g2_a21o_1 _24374_ (.A2(net3956),
    .A1(net2848),
    .B1(_02467_),
    .X(_00356_));
 sg13g2_nand2_1 _24375_ (.Y(_02468_),
    .A(net1997),
    .B(net3957));
 sg13g2_nand2_1 _24376_ (.Y(_02469_),
    .A(_02451_),
    .B(_02464_));
 sg13g2_nand3_1 _24377_ (.B(_14467_),
    .C(_02446_),
    .A(_14466_),
    .Y(_02470_));
 sg13g2_nand2_1 _24378_ (.Y(_02471_),
    .A(_15398_),
    .B(_02445_));
 sg13g2_nand4_1 _24379_ (.B(_15410_),
    .C(_02470_),
    .A(net4681),
    .Y(_02472_),
    .D(_02471_));
 sg13g2_a21oi_1 _24380_ (.A1(net4567),
    .A2(\u_inv.d_next[81] ),
    .Y(_02473_),
    .B1(net3786));
 sg13g2_a21oi_1 _24381_ (.A1(_14469_),
    .A2(_02443_),
    .Y(_02474_),
    .B1(_14579_));
 sg13g2_xor2_1 _24382_ (.B(_02474_),
    .A(_14466_),
    .X(_02475_));
 sg13g2_a22oi_1 _24383_ (.Y(_02476_),
    .B1(_02475_),
    .B2(net3786),
    .A2(_02473_),
    .A1(_02472_));
 sg13g2_xnor2_1 _24384_ (.Y(_02477_),
    .A(net3429),
    .B(_02476_));
 sg13g2_o21ai_1 _24385_ (.B1(net4341),
    .Y(_02478_),
    .A1(_02469_),
    .A2(_02477_));
 sg13g2_a21oi_1 _24386_ (.A1(_02469_),
    .A2(_02477_),
    .Y(_02479_),
    .B1(_02478_));
 sg13g2_o21ai_1 _24387_ (.B1(net3893),
    .Y(_02480_),
    .A1(net4342),
    .A2(_02476_));
 sg13g2_o21ai_1 _24388_ (.B1(_02468_),
    .Y(_00357_),
    .A1(_02479_),
    .A2(_02480_));
 sg13g2_o21ai_1 _24389_ (.B1(net3429),
    .Y(_02481_),
    .A1(_02450_),
    .A2(_02476_));
 sg13g2_o21ai_1 _24390_ (.B1(_02481_),
    .Y(_02482_),
    .A1(_02464_),
    .A2(_02477_));
 sg13g2_a21oi_2 _24391_ (.B1(_14471_),
    .Y(_02483_),
    .A2(_02442_),
    .A1(_14569_));
 sg13g2_nor2_1 _24392_ (.A(_14580_),
    .B(_02483_),
    .Y(_02484_));
 sg13g2_o21ai_1 _24393_ (.B1(_14462_),
    .Y(_02485_),
    .A1(_14580_),
    .A2(_02483_));
 sg13g2_xnor2_1 _24394_ (.Y(_02486_),
    .A(_14461_),
    .B(_02484_));
 sg13g2_a21oi_1 _24395_ (.A1(_15398_),
    .A2(_02445_),
    .Y(_02487_),
    .B1(_15412_));
 sg13g2_a21oi_1 _24396_ (.A1(_14462_),
    .A2(_02487_),
    .Y(_02488_),
    .B1(net4564));
 sg13g2_o21ai_1 _24397_ (.B1(_02488_),
    .Y(_02489_),
    .A1(_14462_),
    .A2(_02487_));
 sg13g2_a21oi_1 _24398_ (.A1(net4564),
    .A2(\u_inv.d_next[82] ),
    .Y(_02490_),
    .B1(net3783));
 sg13g2_a22oi_1 _24399_ (.Y(_02491_),
    .B1(_02489_),
    .B2(_02490_),
    .A2(_02486_),
    .A1(net3783));
 sg13g2_nand2_1 _24400_ (.Y(_02492_),
    .A(net3429),
    .B(_02491_));
 sg13g2_inv_1 _24401_ (.Y(_02493_),
    .A(_02492_));
 sg13g2_xnor2_1 _24402_ (.Y(_02494_),
    .A(net3429),
    .B(_02491_));
 sg13g2_nor2b_1 _24403_ (.A(_02494_),
    .B_N(_02482_),
    .Y(_02495_));
 sg13g2_xnor2_1 _24404_ (.Y(_02496_),
    .A(_02482_),
    .B(_02494_));
 sg13g2_nor2_1 _24405_ (.A(net4342),
    .B(_02491_),
    .Y(_02497_));
 sg13g2_o21ai_1 _24406_ (.B1(net3893),
    .Y(_02498_),
    .A1(net4296),
    .A2(_02496_));
 sg13g2_nand2_1 _24407_ (.Y(_02499_),
    .A(net2241),
    .B(net3956));
 sg13g2_o21ai_1 _24408_ (.B1(_02499_),
    .Y(_00358_),
    .A1(_02497_),
    .A2(_02498_));
 sg13g2_nor2_1 _24409_ (.A(_02493_),
    .B(_02495_),
    .Y(_02500_));
 sg13g2_a21oi_1 _24410_ (.A1(net4564),
    .A2(\u_inv.d_next[83] ),
    .Y(_02501_),
    .B1(net3784));
 sg13g2_o21ai_1 _24411_ (.B1(_14460_),
    .Y(_02502_),
    .A1(_14462_),
    .A2(_02487_));
 sg13g2_xnor2_1 _24412_ (.Y(_02503_),
    .A(_14459_),
    .B(_02502_));
 sg13g2_nand2_1 _24413_ (.Y(_02504_),
    .A(net4681),
    .B(_02503_));
 sg13g2_a21oi_1 _24414_ (.A1(_14581_),
    .A2(_02485_),
    .Y(_02505_),
    .B1(_14459_));
 sg13g2_nand3_1 _24415_ (.B(_14581_),
    .C(_02485_),
    .A(_14459_),
    .Y(_02506_));
 sg13g2_nor2_1 _24416_ (.A(net3850),
    .B(_02505_),
    .Y(_02507_));
 sg13g2_a22oi_1 _24417_ (.Y(_02508_),
    .B1(_02506_),
    .B2(_02507_),
    .A2(_02504_),
    .A1(_02501_));
 sg13g2_xnor2_1 _24418_ (.Y(_02509_),
    .A(net3429),
    .B(_02508_));
 sg13g2_xnor2_1 _24419_ (.Y(_02510_),
    .A(_02500_),
    .B(_02509_));
 sg13g2_o21ai_1 _24420_ (.B1(net3893),
    .Y(_02511_),
    .A1(net4346),
    .A2(_02508_));
 sg13g2_a21oi_1 _24421_ (.A1(net4346),
    .A2(_02510_),
    .Y(_02512_),
    .B1(_02511_));
 sg13g2_a21o_1 _24422_ (.A2(net3957),
    .A1(net2862),
    .B1(_02512_),
    .X(_00359_));
 sg13g2_a21oi_2 _24423_ (.B1(_14583_),
    .Y(_02513_),
    .A2(_02483_),
    .A1(_14463_));
 sg13g2_xnor2_1 _24424_ (.Y(_02514_),
    .A(_14454_),
    .B(_02513_));
 sg13g2_nand3_1 _24425_ (.B(_15398_),
    .C(_02445_),
    .A(_15390_),
    .Y(_02515_));
 sg13g2_nand2_1 _24426_ (.Y(_02516_),
    .A(_15414_),
    .B(_02515_));
 sg13g2_o21ai_1 _24427_ (.B1(net4681),
    .Y(_02517_),
    .A1(_14454_),
    .A2(_02516_));
 sg13g2_a21o_1 _24428_ (.A2(_02516_),
    .A1(_14454_),
    .B1(_02517_),
    .X(_02518_));
 sg13g2_a21oi_1 _24429_ (.A1(net4565),
    .A2(\u_inv.d_next[84] ),
    .Y(_02519_),
    .B1(net3784));
 sg13g2_a22oi_1 _24430_ (.Y(_02520_),
    .B1(_02518_),
    .B2(_02519_),
    .A2(_02514_),
    .A1(net3784));
 sg13g2_nand2_1 _24431_ (.Y(_02521_),
    .A(net3430),
    .B(_02520_));
 sg13g2_xnor2_1 _24432_ (.Y(_02522_),
    .A(net3430),
    .B(_02520_));
 sg13g2_o21ai_1 _24433_ (.B1(net3429),
    .Y(_02523_),
    .A1(_02491_),
    .A2(_02508_));
 sg13g2_or2_1 _24434_ (.X(_02524_),
    .B(_02509_),
    .A(_02494_));
 sg13g2_inv_1 _24435_ (.Y(_02525_),
    .A(_02524_));
 sg13g2_a221oi_1 _24436_ (.B2(_02482_),
    .C1(_02493_),
    .B1(_02525_),
    .A1(net3431),
    .Y(_02526_),
    .A2(_02508_));
 sg13g2_xnor2_1 _24437_ (.Y(_02527_),
    .A(_02522_),
    .B(_02526_));
 sg13g2_o21ai_1 _24438_ (.B1(net3890),
    .Y(_02528_),
    .A1(net4341),
    .A2(_02520_));
 sg13g2_a21oi_1 _24439_ (.A1(net4341),
    .A2(_02527_),
    .Y(_02529_),
    .B1(_02528_));
 sg13g2_a21o_1 _24440_ (.A2(net3957),
    .A1(net2662),
    .B1(_02529_),
    .X(_00360_));
 sg13g2_nand2_1 _24441_ (.Y(_02530_),
    .A(net2615),
    .B(net3955));
 sg13g2_a21oi_1 _24442_ (.A1(net4565),
    .A2(\u_inv.d_next[85] ),
    .Y(_02531_),
    .B1(net3784));
 sg13g2_a21oi_1 _24443_ (.A1(_14454_),
    .A2(_02516_),
    .Y(_02532_),
    .B1(_14453_));
 sg13g2_xnor2_1 _24444_ (.Y(_02533_),
    .A(_14452_),
    .B(_02532_));
 sg13g2_nand2_1 _24445_ (.Y(_02534_),
    .A(net4681),
    .B(_02533_));
 sg13g2_o21ai_1 _24446_ (.B1(_14585_),
    .Y(_02535_),
    .A1(_14454_),
    .A2(_02513_));
 sg13g2_o21ai_1 _24447_ (.B1(net3784),
    .Y(_02536_),
    .A1(_14452_),
    .A2(_02535_));
 sg13g2_a21oi_1 _24448_ (.A1(_14452_),
    .A2(_02535_),
    .Y(_02537_),
    .B1(_02536_));
 sg13g2_a21oi_2 _24449_ (.B1(_02537_),
    .Y(_02538_),
    .A2(_02534_),
    .A1(_02531_));
 sg13g2_nand2_1 _24450_ (.Y(_02539_),
    .A(net3430),
    .B(_02538_));
 sg13g2_xnor2_1 _24451_ (.Y(_02540_),
    .A(net3431),
    .B(_02538_));
 sg13g2_o21ai_1 _24452_ (.B1(_02521_),
    .Y(_02541_),
    .A1(_02522_),
    .A2(_02526_));
 sg13g2_o21ai_1 _24453_ (.B1(net4341),
    .Y(_02542_),
    .A1(_02540_),
    .A2(_02541_));
 sg13g2_a21oi_1 _24454_ (.A1(_02540_),
    .A2(_02541_),
    .Y(_02543_),
    .B1(_02542_));
 sg13g2_o21ai_1 _24455_ (.B1(net3890),
    .Y(_02544_),
    .A1(net4341),
    .A2(_02538_));
 sg13g2_o21ai_1 _24456_ (.B1(_02530_),
    .Y(_00361_),
    .A1(_02543_),
    .A2(_02544_));
 sg13g2_o21ai_1 _24457_ (.B1(_14587_),
    .Y(_02545_),
    .A1(_14455_),
    .A2(_02513_));
 sg13g2_xnor2_1 _24458_ (.Y(_02546_),
    .A(_14449_),
    .B(_02545_));
 sg13g2_a21o_1 _24459_ (.A2(_02515_),
    .A1(_15414_),
    .B1(_15388_),
    .X(_02547_));
 sg13g2_a21o_1 _24460_ (.A2(_02547_),
    .A1(_15416_),
    .B1(_14449_),
    .X(_02548_));
 sg13g2_nand3_1 _24461_ (.B(_15416_),
    .C(_02547_),
    .A(_14449_),
    .Y(_02549_));
 sg13g2_nand3_1 _24462_ (.B(_02548_),
    .C(_02549_),
    .A(net4681),
    .Y(_02550_));
 sg13g2_a21oi_1 _24463_ (.A1(net4565),
    .A2(\u_inv.d_next[86] ),
    .Y(_02551_),
    .B1(net3783));
 sg13g2_a22oi_1 _24464_ (.Y(_02552_),
    .B1(_02550_),
    .B2(_02551_),
    .A2(_02546_),
    .A1(net3783));
 sg13g2_nand2_1 _24465_ (.Y(_02553_),
    .A(net3430),
    .B(_02552_));
 sg13g2_xnor2_1 _24466_ (.Y(_02554_),
    .A(net3430),
    .B(_02552_));
 sg13g2_nand2_1 _24467_ (.Y(_02555_),
    .A(_02521_),
    .B(_02539_));
 sg13g2_o21ai_1 _24468_ (.B1(_02541_),
    .Y(_02556_),
    .A1(net3430),
    .A2(_02538_));
 sg13g2_a21o_1 _24469_ (.A2(_02556_),
    .A1(_02539_),
    .B1(_02554_),
    .X(_02557_));
 sg13g2_nand3_1 _24470_ (.B(_02554_),
    .C(_02556_),
    .A(_02539_),
    .Y(_02558_));
 sg13g2_and2_1 _24471_ (.A(_02557_),
    .B(_02558_),
    .X(_02559_));
 sg13g2_nor2_1 _24472_ (.A(net4339),
    .B(_02552_),
    .Y(_02560_));
 sg13g2_o21ai_1 _24473_ (.B1(net3892),
    .Y(_02561_),
    .A1(net4296),
    .A2(_02559_));
 sg13g2_nand2_1 _24474_ (.Y(_02562_),
    .A(net2695),
    .B(net3955));
 sg13g2_o21ai_1 _24475_ (.B1(_02562_),
    .Y(_00362_),
    .A1(_02560_),
    .A2(_02561_));
 sg13g2_a21oi_1 _24476_ (.A1(net4564),
    .A2(\u_inv.d_next[87] ),
    .Y(_02563_),
    .B1(net3783));
 sg13g2_a21o_1 _24477_ (.A2(_02548_),
    .A1(_14447_),
    .B1(_14446_),
    .X(_02564_));
 sg13g2_nand3_1 _24478_ (.B(_14447_),
    .C(_02548_),
    .A(_14446_),
    .Y(_02565_));
 sg13g2_nand3_1 _24479_ (.B(_02564_),
    .C(_02565_),
    .A(net4682),
    .Y(_02566_));
 sg13g2_a21oi_1 _24480_ (.A1(_14449_),
    .A2(_02545_),
    .Y(_02567_),
    .B1(_14584_));
 sg13g2_or2_1 _24481_ (.X(_02568_),
    .B(_02567_),
    .A(_14446_));
 sg13g2_a21oi_1 _24482_ (.A1(_14446_),
    .A2(_02567_),
    .Y(_02569_),
    .B1(net3850));
 sg13g2_a22oi_1 _24483_ (.Y(_02570_),
    .B1(_02568_),
    .B2(_02569_),
    .A2(_02566_),
    .A1(_02563_));
 sg13g2_nand2_1 _24484_ (.Y(_02571_),
    .A(net3430),
    .B(_02570_));
 sg13g2_xnor2_1 _24485_ (.Y(_02572_),
    .A(net3430),
    .B(_02570_));
 sg13g2_nand2_1 _24486_ (.Y(_02573_),
    .A(_02553_),
    .B(_02557_));
 sg13g2_xor2_1 _24487_ (.B(_02573_),
    .A(_02572_),
    .X(_02574_));
 sg13g2_o21ai_1 _24488_ (.B1(net3892),
    .Y(_02575_),
    .A1(net4339),
    .A2(_02570_));
 sg13g2_a21oi_1 _24489_ (.A1(net4339),
    .A2(_02574_),
    .Y(_02576_),
    .B1(_02575_));
 sg13g2_a21o_1 _24490_ (.A2(net3955),
    .A1(net3174),
    .B1(_02576_),
    .X(_00363_));
 sg13g2_a21oi_1 _24491_ (.A1(_14569_),
    .A2(_02442_),
    .Y(_02577_),
    .B1(_14473_));
 sg13g2_nor2_1 _24492_ (.A(_14589_),
    .B(_02577_),
    .Y(_02578_));
 sg13g2_nor2_1 _24493_ (.A(_14440_),
    .B(_02578_),
    .Y(_02579_));
 sg13g2_xnor2_1 _24494_ (.Y(_02580_),
    .A(_14440_),
    .B(_02578_));
 sg13g2_a21o_2 _24495_ (.A2(_02445_),
    .A1(_15422_),
    .B1(_15420_),
    .X(_02581_));
 sg13g2_o21ai_1 _24496_ (.B1(net4681),
    .Y(_02582_),
    .A1(_14440_),
    .A2(_02581_));
 sg13g2_a21o_1 _24497_ (.A2(_02581_),
    .A1(_14440_),
    .B1(_02582_),
    .X(_02583_));
 sg13g2_a21oi_1 _24498_ (.A1(net4563),
    .A2(\u_inv.d_next[88] ),
    .Y(_02584_),
    .B1(net3782));
 sg13g2_a22oi_1 _24499_ (.Y(_02585_),
    .B1(_02583_),
    .B2(_02584_),
    .A2(_02580_),
    .A1(net3782));
 sg13g2_nand2_1 _24500_ (.Y(_02586_),
    .A(net3428),
    .B(_02585_));
 sg13g2_xnor2_1 _24501_ (.Y(_02587_),
    .A(net3428),
    .B(_02585_));
 sg13g2_nor2_1 _24502_ (.A(_02554_),
    .B(_02572_),
    .Y(_02588_));
 sg13g2_nor4_1 _24503_ (.A(_02522_),
    .B(_02540_),
    .C(_02554_),
    .D(_02572_),
    .Y(_02589_));
 sg13g2_o21ai_1 _24504_ (.B1(_02523_),
    .Y(_02590_),
    .A1(_02481_),
    .A2(_02524_));
 sg13g2_nand2_1 _24505_ (.Y(_02591_),
    .A(_02553_),
    .B(_02571_));
 sg13g2_a221oi_1 _24506_ (.B2(_02590_),
    .C1(_02591_),
    .B1(_02589_),
    .A1(_02555_),
    .Y(_02592_),
    .A2(_02588_));
 sg13g2_inv_1 _24507_ (.Y(_02593_),
    .A(_02592_));
 sg13g2_nor3_1 _24508_ (.A(_02452_),
    .B(_02477_),
    .C(_02524_),
    .Y(_02594_));
 sg13g2_and2_1 _24509_ (.A(_02589_),
    .B(_02594_),
    .X(_02595_));
 sg13g2_nand2b_1 _24510_ (.Y(_02596_),
    .B(_02595_),
    .A_N(_02463_));
 sg13g2_nand2_1 _24511_ (.Y(_02597_),
    .A(_02592_),
    .B(_02596_));
 sg13g2_nand2b_1 _24512_ (.Y(_02598_),
    .B(_02597_),
    .A_N(_02587_));
 sg13g2_nand3_1 _24513_ (.B(_02592_),
    .C(_02596_),
    .A(_02587_),
    .Y(_02599_));
 sg13g2_a21oi_1 _24514_ (.A1(_02598_),
    .A2(_02599_),
    .Y(_02600_),
    .B1(net4296));
 sg13g2_o21ai_1 _24515_ (.B1(net3892),
    .Y(_02601_),
    .A1(net4339),
    .A2(_02585_));
 sg13g2_nand2_1 _24516_ (.Y(_02602_),
    .A(net2815),
    .B(net3955));
 sg13g2_o21ai_1 _24517_ (.B1(_02602_),
    .Y(_00364_),
    .A1(_02600_),
    .A2(_02601_));
 sg13g2_nand2_1 _24518_ (.Y(_02603_),
    .A(net3098),
    .B(net3955));
 sg13g2_nand2_1 _24519_ (.Y(_02604_),
    .A(_02586_),
    .B(_02598_));
 sg13g2_a21o_1 _24520_ (.A2(_02581_),
    .A1(_14440_),
    .B1(_14438_),
    .X(_02605_));
 sg13g2_a221oi_1 _24521_ (.B2(_02581_),
    .C1(net4563),
    .B1(_15395_),
    .A1(_14438_),
    .Y(_02606_),
    .A2(_14439_));
 sg13g2_o21ai_1 _24522_ (.B1(_02606_),
    .Y(_02607_),
    .A1(_14439_),
    .A2(_02605_));
 sg13g2_a21oi_1 _24523_ (.A1(net4563),
    .A2(\u_inv.d_next[89] ),
    .Y(_02608_),
    .B1(net3782));
 sg13g2_or2_1 _24524_ (.X(_02609_),
    .B(_02579_),
    .A(_14570_));
 sg13g2_xnor2_1 _24525_ (.Y(_02610_),
    .A(_14437_),
    .B(_02609_));
 sg13g2_a22oi_1 _24526_ (.Y(_02611_),
    .B1(_02610_),
    .B2(net3782),
    .A2(_02608_),
    .A1(_02607_));
 sg13g2_nor2_1 _24527_ (.A(net3427),
    .B(_02611_),
    .Y(_02612_));
 sg13g2_xnor2_1 _24528_ (.Y(_02613_),
    .A(net3428),
    .B(_02611_));
 sg13g2_o21ai_1 _24529_ (.B1(net4338),
    .Y(_02614_),
    .A1(_02604_),
    .A2(_02613_));
 sg13g2_a21oi_1 _24530_ (.A1(_02604_),
    .A2(_02613_),
    .Y(_02615_),
    .B1(_02614_));
 sg13g2_o21ai_1 _24531_ (.B1(net3892),
    .Y(_02616_),
    .A1(net4338),
    .A2(_02611_));
 sg13g2_o21ai_1 _24532_ (.B1(_02603_),
    .Y(_00365_),
    .A1(_02615_),
    .A2(_02616_));
 sg13g2_o21ai_1 _24533_ (.B1(_14442_),
    .Y(_02617_),
    .A1(_14589_),
    .A2(_02577_));
 sg13g2_a21oi_1 _24534_ (.A1(_14571_),
    .A2(_02617_),
    .Y(_02618_),
    .B1(_14433_));
 sg13g2_nand3_1 _24535_ (.B(_14571_),
    .C(_02617_),
    .A(_14433_),
    .Y(_02619_));
 sg13g2_nand2b_1 _24536_ (.Y(_02620_),
    .B(_02619_),
    .A_N(_02618_));
 sg13g2_a221oi_1 _24537_ (.B2(_02581_),
    .C1(_15401_),
    .B1(_15395_),
    .A1(_14438_),
    .Y(_02621_),
    .A2(_14439_));
 sg13g2_a21oi_1 _24538_ (.A1(_14432_),
    .A2(_02621_),
    .Y(_02622_),
    .B1(net4563));
 sg13g2_o21ai_1 _24539_ (.B1(_02622_),
    .Y(_02623_),
    .A1(_14432_),
    .A2(_02621_));
 sg13g2_a21oi_1 _24540_ (.A1(net4563),
    .A2(\u_inv.d_next[90] ),
    .Y(_02624_),
    .B1(net3782));
 sg13g2_a22oi_1 _24541_ (.Y(_02625_),
    .B1(_02623_),
    .B2(_02624_),
    .A2(_02620_),
    .A1(net3782));
 sg13g2_nand2_1 _24542_ (.Y(_02626_),
    .A(net3428),
    .B(_02625_));
 sg13g2_xnor2_1 _24543_ (.Y(_02627_),
    .A(net3428),
    .B(_02625_));
 sg13g2_o21ai_1 _24544_ (.B1(net3428),
    .Y(_02628_),
    .A1(_02585_),
    .A2(_02611_));
 sg13g2_a21o_1 _24545_ (.A2(_02628_),
    .A1(_02598_),
    .B1(_02612_),
    .X(_02629_));
 sg13g2_xnor2_1 _24546_ (.Y(_02630_),
    .A(_02627_),
    .B(_02629_));
 sg13g2_o21ai_1 _24547_ (.B1(net3892),
    .Y(_02631_),
    .A1(net4338),
    .A2(_02625_));
 sg13g2_a21oi_1 _24548_ (.A1(net4338),
    .A2(_02630_),
    .Y(_02632_),
    .B1(_02631_));
 sg13g2_a21o_1 _24549_ (.A2(net3955),
    .A1(net2351),
    .B1(_02632_),
    .X(_00366_));
 sg13g2_nand2_1 _24550_ (.Y(_02633_),
    .A(net2708),
    .B(net3955));
 sg13g2_nand2b_1 _24551_ (.Y(_02634_),
    .B(net3850),
    .A_N(\u_inv.d_next[91] ));
 sg13g2_o21ai_1 _24552_ (.B1(_14431_),
    .Y(_02635_),
    .A1(_14432_),
    .A2(_02621_));
 sg13g2_xnor2_1 _24553_ (.Y(_02636_),
    .A(_14429_),
    .B(_02635_));
 sg13g2_a22oi_1 _24554_ (.Y(_02637_),
    .B1(_02636_),
    .B2(net4681),
    .A2(_02634_),
    .A1(net3730));
 sg13g2_o21ai_1 _24555_ (.B1(_14430_),
    .Y(_02638_),
    .A1(_14572_),
    .A2(_02618_));
 sg13g2_or3_1 _24556_ (.A(_14430_),
    .B(_14572_),
    .C(_02618_),
    .X(_02639_));
 sg13g2_and3_2 _24557_ (.X(_02640_),
    .A(net3782),
    .B(_02638_),
    .C(_02639_));
 sg13g2_nor2_1 _24558_ (.A(_02637_),
    .B(_02640_),
    .Y(_02641_));
 sg13g2_or3_1 _24559_ (.A(net3478),
    .B(_02637_),
    .C(_02640_),
    .X(_02642_));
 sg13g2_o21ai_1 _24560_ (.B1(net3478),
    .Y(_02643_),
    .A1(_02637_),
    .A2(_02640_));
 sg13g2_nand2_1 _24561_ (.Y(_02644_),
    .A(_02642_),
    .B(_02643_));
 sg13g2_o21ai_1 _24562_ (.B1(_02626_),
    .Y(_02645_),
    .A1(_02627_),
    .A2(_02629_));
 sg13g2_o21ai_1 _24563_ (.B1(net4338),
    .Y(_02646_),
    .A1(_02644_),
    .A2(_02645_));
 sg13g2_a21oi_1 _24564_ (.A1(_02644_),
    .A2(_02645_),
    .Y(_02647_),
    .B1(_02646_));
 sg13g2_o21ai_1 _24565_ (.B1(net3892),
    .Y(_02648_),
    .A1(net4338),
    .A2(_02641_));
 sg13g2_o21ai_1 _24566_ (.B1(_02633_),
    .Y(_00367_),
    .A1(_02647_),
    .A2(_02648_));
 sg13g2_o21ai_1 _24567_ (.B1(_14574_),
    .Y(_02649_),
    .A1(_14434_),
    .A2(_02617_));
 sg13g2_xnor2_1 _24568_ (.Y(_02650_),
    .A(_14424_),
    .B(_02649_));
 sg13g2_a21oi_2 _24569_ (.B1(_15404_),
    .Y(_02651_),
    .A2(_02581_),
    .A1(_15396_));
 sg13g2_a21oi_1 _24570_ (.A1(_14424_),
    .A2(_02651_),
    .Y(_02652_),
    .B1(net4563));
 sg13g2_o21ai_1 _24571_ (.B1(_02652_),
    .Y(_02653_),
    .A1(_14424_),
    .A2(_02651_));
 sg13g2_a21oi_1 _24572_ (.A1(net4563),
    .A2(\u_inv.d_next[92] ),
    .Y(_02654_),
    .B1(net3782));
 sg13g2_a22oi_1 _24573_ (.Y(_02655_),
    .B1(_02653_),
    .B2(_02654_),
    .A2(_02650_),
    .A1(net3783));
 sg13g2_nand2_1 _24574_ (.Y(_02656_),
    .A(net3435),
    .B(_02655_));
 sg13g2_xnor2_1 _24575_ (.Y(_02657_),
    .A(net3435),
    .B(_02655_));
 sg13g2_nand3b_1 _24576_ (.B(_02642_),
    .C(_02643_),
    .Y(_02658_),
    .A_N(_02627_));
 sg13g2_and2_1 _24577_ (.A(_02626_),
    .B(_02642_),
    .X(_02659_));
 sg13g2_o21ai_1 _24578_ (.B1(_02659_),
    .Y(_02660_),
    .A1(_02628_),
    .A2(_02658_));
 sg13g2_nor3_2 _24579_ (.A(_02587_),
    .B(_02613_),
    .C(_02658_),
    .Y(_02661_));
 sg13g2_a21oi_2 _24580_ (.B1(_02660_),
    .Y(_02662_),
    .A2(_02661_),
    .A1(_02597_));
 sg13g2_xnor2_1 _24581_ (.Y(_02663_),
    .A(_02657_),
    .B(_02662_));
 sg13g2_o21ai_1 _24582_ (.B1(net3892),
    .Y(_02664_),
    .A1(net4338),
    .A2(_02655_));
 sg13g2_a21oi_1 _24583_ (.A1(net4338),
    .A2(_02663_),
    .Y(_02665_),
    .B1(_02664_));
 sg13g2_a21o_1 _24584_ (.A2(net3955),
    .A1(net2732),
    .B1(_02665_),
    .X(_00368_));
 sg13g2_nand2_1 _24585_ (.Y(_02666_),
    .A(net2198),
    .B(net3957));
 sg13g2_nor2_1 _24586_ (.A(_14422_),
    .B(_14423_),
    .Y(_02667_));
 sg13g2_o21ai_1 _24587_ (.B1(_02667_),
    .Y(_02668_),
    .A1(_14424_),
    .A2(_02651_));
 sg13g2_or3_1 _24588_ (.A(_14421_),
    .B(_14424_),
    .C(_02651_),
    .X(_02669_));
 sg13g2_a21oi_1 _24589_ (.A1(_14422_),
    .A2(_14423_),
    .Y(_02670_),
    .B1(net4571));
 sg13g2_nand3_1 _24590_ (.B(_02669_),
    .C(_02670_),
    .A(_02668_),
    .Y(_02671_));
 sg13g2_a21oi_1 _24591_ (.A1(net4571),
    .A2(\u_inv.d_next[93] ),
    .Y(_02672_),
    .B1(net3789));
 sg13g2_a21oi_1 _24592_ (.A1(_14424_),
    .A2(_02649_),
    .Y(_02673_),
    .B1(_14575_));
 sg13g2_xnor2_1 _24593_ (.Y(_02674_),
    .A(_14422_),
    .B(_02673_));
 sg13g2_a22oi_1 _24594_ (.Y(_02675_),
    .B1(_02674_),
    .B2(net3789),
    .A2(_02672_),
    .A1(_02671_));
 sg13g2_nand2_1 _24595_ (.Y(_02676_),
    .A(net3435),
    .B(_02675_));
 sg13g2_xnor2_1 _24596_ (.Y(_02677_),
    .A(net3435),
    .B(_02675_));
 sg13g2_o21ai_1 _24597_ (.B1(_02656_),
    .Y(_02678_),
    .A1(_02657_),
    .A2(_02662_));
 sg13g2_o21ai_1 _24598_ (.B1(net4345),
    .Y(_02679_),
    .A1(_02677_),
    .A2(_02678_));
 sg13g2_a21oi_1 _24599_ (.A1(_02677_),
    .A2(_02678_),
    .Y(_02680_),
    .B1(_02679_));
 sg13g2_o21ai_1 _24600_ (.B1(net3893),
    .Y(_02681_),
    .A1(net4345),
    .A2(_02675_));
 sg13g2_o21ai_1 _24601_ (.B1(_02666_),
    .Y(_00369_),
    .A1(_02680_),
    .A2(_02681_));
 sg13g2_a21oi_1 _24602_ (.A1(_14425_),
    .A2(_02649_),
    .Y(_02682_),
    .B1(_14576_));
 sg13g2_xnor2_1 _24603_ (.Y(_02683_),
    .A(_14416_),
    .B(_02682_));
 sg13g2_a21o_1 _24604_ (.A2(_02669_),
    .A1(_15406_),
    .B1(_14417_),
    .X(_02684_));
 sg13g2_nand3_1 _24605_ (.B(_15406_),
    .C(_02669_),
    .A(_14417_),
    .Y(_02685_));
 sg13g2_nand3_1 _24606_ (.B(_02684_),
    .C(_02685_),
    .A(net4692),
    .Y(_02686_));
 sg13g2_a21oi_1 _24607_ (.A1(net4571),
    .A2(\u_inv.d_next[94] ),
    .Y(_02687_),
    .B1(net3789));
 sg13g2_a22oi_1 _24608_ (.Y(_02688_),
    .B1(_02686_),
    .B2(_02687_),
    .A2(_02683_),
    .A1(net3789));
 sg13g2_nand2_1 _24609_ (.Y(_02689_),
    .A(net3435),
    .B(_02688_));
 sg13g2_xnor2_1 _24610_ (.Y(_02690_),
    .A(net3481),
    .B(_02688_));
 sg13g2_nand2_1 _24611_ (.Y(_02691_),
    .A(_02656_),
    .B(_02676_));
 sg13g2_o21ai_1 _24612_ (.B1(_02678_),
    .Y(_02692_),
    .A1(net3435),
    .A2(_02675_));
 sg13g2_nor2_1 _24613_ (.A(_02657_),
    .B(_02677_),
    .Y(_02693_));
 sg13g2_nand2_1 _24614_ (.Y(_02694_),
    .A(_02676_),
    .B(_02692_));
 sg13g2_nand2_1 _24615_ (.Y(_02695_),
    .A(_02690_),
    .B(_02694_));
 sg13g2_xnor2_1 _24616_ (.Y(_02696_),
    .A(_02690_),
    .B(_02694_));
 sg13g2_o21ai_1 _24617_ (.B1(net3893),
    .Y(_02697_),
    .A1(net4345),
    .A2(_02688_));
 sg13g2_a21oi_1 _24618_ (.A1(net4345),
    .A2(_02696_),
    .Y(_02698_),
    .B1(_02697_));
 sg13g2_a21o_1 _24619_ (.A2(net3965),
    .A1(net2631),
    .B1(_02698_),
    .X(_00370_));
 sg13g2_nand2_1 _24620_ (.Y(_02699_),
    .A(net2210),
    .B(net3957));
 sg13g2_a21oi_1 _24621_ (.A1(net4563),
    .A2(\u_inv.d_next[95] ),
    .Y(_02700_),
    .B1(net3783));
 sg13g2_nand3_1 _24622_ (.B(_14415_),
    .C(_02684_),
    .A(_14414_),
    .Y(_02701_));
 sg13g2_a21o_1 _24623_ (.A2(_02684_),
    .A1(_14415_),
    .B1(_14414_),
    .X(_02702_));
 sg13g2_nand3_1 _24624_ (.B(_02701_),
    .C(_02702_),
    .A(net4692),
    .Y(_02703_));
 sg13g2_o21ai_1 _24625_ (.B1(_14577_),
    .Y(_02704_),
    .A1(_14416_),
    .A2(_02682_));
 sg13g2_nand2b_1 _24626_ (.Y(_02705_),
    .B(_14414_),
    .A_N(_02704_));
 sg13g2_a21oi_1 _24627_ (.A1(_14413_),
    .A2(_02704_),
    .Y(_02706_),
    .B1(net3850));
 sg13g2_a22oi_1 _24628_ (.Y(_02707_),
    .B1(_02705_),
    .B2(_02706_),
    .A2(_02703_),
    .A1(_02700_));
 sg13g2_xnor2_1 _24629_ (.Y(_02708_),
    .A(net3481),
    .B(_02707_));
 sg13g2_a21oi_1 _24630_ (.A1(_02689_),
    .A2(_02695_),
    .Y(_02709_),
    .B1(_02708_));
 sg13g2_and3_1 _24631_ (.X(_02710_),
    .A(_02689_),
    .B(_02695_),
    .C(_02708_));
 sg13g2_nor3_1 _24632_ (.A(net4296),
    .B(_02709_),
    .C(_02710_),
    .Y(_02711_));
 sg13g2_o21ai_1 _24633_ (.B1(net3892),
    .Y(_02712_),
    .A1(net4345),
    .A2(_02707_));
 sg13g2_o21ai_1 _24634_ (.B1(_02699_),
    .Y(_00371_),
    .A1(_02711_),
    .A2(_02712_));
 sg13g2_o21ai_1 _24635_ (.B1(_14534_),
    .Y(_02713_),
    .A1(_14238_),
    .A2(_14302_));
 sg13g2_nand2_1 _24636_ (.Y(_02714_),
    .A(_14594_),
    .B(_02713_));
 sg13g2_xnor2_1 _24637_ (.Y(_02715_),
    .A(_14405_),
    .B(_02714_));
 sg13g2_a21oi_2 _24638_ (.B1(_15423_),
    .Y(_02716_),
    .A2(_15627_),
    .A1(_15623_));
 sg13g2_a21o_2 _24639_ (.A2(_15627_),
    .A1(_15623_),
    .B1(_15423_),
    .X(_02717_));
 sg13g2_nand2b_1 _24640_ (.Y(_02718_),
    .B(_02717_),
    .A_N(_14405_));
 sg13g2_a21oi_1 _24641_ (.A1(_14405_),
    .A2(_02716_),
    .Y(_02719_),
    .B1(net4570));
 sg13g2_nand2_1 _24642_ (.Y(_02720_),
    .A(_02718_),
    .B(_02719_));
 sg13g2_a21oi_1 _24643_ (.A1(net4570),
    .A2(\u_inv.d_next[96] ),
    .Y(_02721_),
    .B1(net3788));
 sg13g2_a22oi_1 _24644_ (.Y(_02722_),
    .B1(_02720_),
    .B2(_02721_),
    .A2(_02715_),
    .A1(net3788));
 sg13g2_and2_1 _24645_ (.A(net3438),
    .B(_02722_),
    .X(_02723_));
 sg13g2_xnor2_1 _24646_ (.Y(_02724_),
    .A(net3480),
    .B(_02722_));
 sg13g2_and4_1 _24647_ (.A(_02661_),
    .B(_02690_),
    .C(_02693_),
    .D(_02708_),
    .X(_02725_));
 sg13g2_and2_1 _24648_ (.A(_02595_),
    .B(_02725_),
    .X(_02726_));
 sg13g2_nand3_1 _24649_ (.B(_02595_),
    .C(_02725_),
    .A(_02462_),
    .Y(_02727_));
 sg13g2_a21o_2 _24650_ (.A2(_02197_),
    .A1(_02192_),
    .B1(_02727_),
    .X(_02728_));
 sg13g2_nand4_1 _24651_ (.B(_02690_),
    .C(_02693_),
    .A(_02660_),
    .Y(_02729_),
    .D(_02708_));
 sg13g2_nand3_1 _24652_ (.B(_02691_),
    .C(_02708_),
    .A(_02690_),
    .Y(_02730_));
 sg13g2_o21ai_1 _24653_ (.B1(net3435),
    .Y(_02731_),
    .A1(_02688_),
    .A2(_02707_));
 sg13g2_nand3_1 _24654_ (.B(_02730_),
    .C(_02731_),
    .A(_02729_),
    .Y(_02732_));
 sg13g2_a221oi_1 _24655_ (.B2(_02461_),
    .C1(_02732_),
    .B1(_02726_),
    .A1(_02593_),
    .Y(_02733_),
    .A2(_02725_));
 sg13g2_nand2_2 _24656_ (.Y(_02734_),
    .A(_02728_),
    .B(_02733_));
 sg13g2_xnor2_1 _24657_ (.Y(_02735_),
    .A(_02724_),
    .B(_02734_));
 sg13g2_o21ai_1 _24658_ (.B1(net3896),
    .Y(_02736_),
    .A1(net4349),
    .A2(_02722_));
 sg13g2_a21oi_1 _24659_ (.A1(net4349),
    .A2(_02735_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_a21o_1 _24660_ (.A2(net3965),
    .A1(net4955),
    .B1(_02737_),
    .X(_00372_));
 sg13g2_nand2_1 _24661_ (.Y(_02738_),
    .A(net2139),
    .B(net3965));
 sg13g2_a21oi_2 _24662_ (.B1(_02723_),
    .Y(_02739_),
    .A2(_02734_),
    .A1(_02724_));
 sg13g2_nor2_1 _24663_ (.A(_14403_),
    .B(_14404_),
    .Y(_02740_));
 sg13g2_a21oi_1 _24664_ (.A1(_14403_),
    .A2(_14404_),
    .Y(_02741_),
    .B1(net4570));
 sg13g2_o21ai_1 _24665_ (.B1(_02741_),
    .Y(_02742_),
    .A1(_15344_),
    .A2(_02716_));
 sg13g2_a21o_1 _24666_ (.A2(_02740_),
    .A1(_02718_),
    .B1(_02742_),
    .X(_02743_));
 sg13g2_a21oi_1 _24667_ (.A1(net4570),
    .A2(\u_inv.d_next[97] ),
    .Y(_02744_),
    .B1(net3788));
 sg13g2_a21oi_1 _24668_ (.A1(_14405_),
    .A2(_02714_),
    .Y(_02745_),
    .B1(_14627_));
 sg13g2_xnor2_1 _24669_ (.Y(_02746_),
    .A(_14403_),
    .B(_02745_));
 sg13g2_a22oi_1 _24670_ (.Y(_02747_),
    .B1(_02746_),
    .B2(net3788),
    .A2(_02744_),
    .A1(_02743_));
 sg13g2_nand2_1 _24671_ (.Y(_02748_),
    .A(net3438),
    .B(_02747_));
 sg13g2_nand2b_1 _24672_ (.Y(_02749_),
    .B(net3480),
    .A_N(_02747_));
 sg13g2_inv_1 _24673_ (.Y(_02750_),
    .A(_02749_));
 sg13g2_and2_1 _24674_ (.A(_02748_),
    .B(_02749_),
    .X(_02751_));
 sg13g2_o21ai_1 _24675_ (.B1(net4349),
    .Y(_02752_),
    .A1(_02739_),
    .A2(_02751_));
 sg13g2_a21oi_1 _24676_ (.A1(_02739_),
    .A2(_02751_),
    .Y(_02753_),
    .B1(_02752_));
 sg13g2_o21ai_1 _24677_ (.B1(net3896),
    .Y(_02754_),
    .A1(net4349),
    .A2(_02747_));
 sg13g2_o21ai_1 _24678_ (.B1(_02738_),
    .Y(_00373_),
    .A1(_02753_),
    .A2(_02754_));
 sg13g2_nor2_1 _24679_ (.A(_02739_),
    .B(_02750_),
    .Y(_02755_));
 sg13g2_nand2b_1 _24680_ (.Y(_02756_),
    .B(_02748_),
    .A_N(_02723_));
 sg13g2_a21oi_1 _24681_ (.A1(net3438),
    .A2(_02747_),
    .Y(_02757_),
    .B1(_02755_));
 sg13g2_o21ai_1 _24682_ (.B1(_02748_),
    .Y(_02758_),
    .A1(_02739_),
    .A2(_02750_));
 sg13g2_a21o_1 _24683_ (.A2(_02713_),
    .A1(_14594_),
    .B1(_14406_),
    .X(_02759_));
 sg13g2_and2_1 _24684_ (.A(_14628_),
    .B(_02759_),
    .X(_02760_));
 sg13g2_a21oi_1 _24685_ (.A1(_14628_),
    .A2(_02759_),
    .Y(_02761_),
    .B1(_14399_));
 sg13g2_xnor2_1 _24686_ (.Y(_02762_),
    .A(_14399_),
    .B(_02760_));
 sg13g2_a221oi_1 _24687_ (.B2(_02717_),
    .C1(_15451_),
    .B1(_15343_),
    .A1(_14403_),
    .Y(_02763_),
    .A2(_14404_));
 sg13g2_o21ai_1 _24688_ (.B1(_15452_),
    .Y(_02764_),
    .A1(_15344_),
    .A2(_02716_));
 sg13g2_xnor2_1 _24689_ (.Y(_02765_),
    .A(_14399_),
    .B(_02763_));
 sg13g2_nand2_1 _24690_ (.Y(_02766_),
    .A(net4692),
    .B(_02765_));
 sg13g2_a21oi_1 _24691_ (.A1(net4570),
    .A2(\u_inv.d_next[98] ),
    .Y(_02767_),
    .B1(net3788));
 sg13g2_a22oi_1 _24692_ (.Y(_02768_),
    .B1(_02766_),
    .B2(_02767_),
    .A2(_02762_),
    .A1(net3788));
 sg13g2_nand2_1 _24693_ (.Y(_02769_),
    .A(net3438),
    .B(_02768_));
 sg13g2_xnor2_1 _24694_ (.Y(_02770_),
    .A(net3438),
    .B(_02768_));
 sg13g2_xor2_1 _24695_ (.B(_02770_),
    .A(_02758_),
    .X(_02771_));
 sg13g2_o21ai_1 _24696_ (.B1(net3896),
    .Y(_02772_),
    .A1(net4349),
    .A2(_02768_));
 sg13g2_a21oi_1 _24697_ (.A1(net4349),
    .A2(_02771_),
    .Y(_02773_),
    .B1(_02772_));
 sg13g2_a21o_1 _24698_ (.A2(net3965),
    .A1(net2782),
    .B1(_02773_),
    .X(_00374_));
 sg13g2_o21ai_1 _24699_ (.B1(_02769_),
    .Y(_02774_),
    .A1(_02757_),
    .A2(_02770_));
 sg13g2_nand2_1 _24700_ (.Y(_02775_),
    .A(_14396_),
    .B(_14398_));
 sg13g2_a21oi_1 _24701_ (.A1(_14399_),
    .A2(_02764_),
    .Y(_02776_),
    .B1(_02775_));
 sg13g2_nor2_1 _24702_ (.A(_15348_),
    .B(_02763_),
    .Y(_02777_));
 sg13g2_nor4_1 _24703_ (.A(net4570),
    .B(_15458_),
    .C(_02776_),
    .D(_02777_),
    .Y(_02778_));
 sg13g2_a21oi_1 _24704_ (.A1(net4570),
    .A2(\u_inv.d_next[99] ),
    .Y(_02779_),
    .B1(net3788));
 sg13g2_nor2b_1 _24705_ (.A(_02778_),
    .B_N(_02779_),
    .Y(_02780_));
 sg13g2_o21ai_1 _24706_ (.B1(_14397_),
    .Y(_02781_),
    .A1(_14629_),
    .A2(_02761_));
 sg13g2_nor3_1 _24707_ (.A(_14397_),
    .B(_14629_),
    .C(_02761_),
    .Y(_02782_));
 sg13g2_nor2_1 _24708_ (.A(net3853),
    .B(_02782_),
    .Y(_02783_));
 sg13g2_a21oi_2 _24709_ (.B1(_02780_),
    .Y(_02784_),
    .A2(_02783_),
    .A1(_02781_));
 sg13g2_nand2_1 _24710_ (.Y(_02785_),
    .A(net3438),
    .B(_02784_));
 sg13g2_xnor2_1 _24711_ (.Y(_02786_),
    .A(net3438),
    .B(_02784_));
 sg13g2_xor2_1 _24712_ (.B(_02786_),
    .A(_02774_),
    .X(_02787_));
 sg13g2_o21ai_1 _24713_ (.B1(net3896),
    .Y(_02788_),
    .A1(net4345),
    .A2(_02784_));
 sg13g2_a21oi_1 _24714_ (.A1(net4349),
    .A2(_02787_),
    .Y(_02789_),
    .B1(_02788_));
 sg13g2_a21o_1 _24715_ (.A2(net3965),
    .A1(net2724),
    .B1(_02789_),
    .X(_00375_));
 sg13g2_o21ai_1 _24716_ (.B1(_14630_),
    .Y(_02790_),
    .A1(_14400_),
    .A2(_02760_));
 sg13g2_xnor2_1 _24717_ (.Y(_02791_),
    .A(_14391_),
    .B(_02790_));
 sg13g2_a21oi_1 _24718_ (.A1(_15347_),
    .A2(_02764_),
    .Y(_02792_),
    .B1(_15459_));
 sg13g2_a21o_1 _24719_ (.A2(_02764_),
    .A1(_15347_),
    .B1(_15459_),
    .X(_02793_));
 sg13g2_a21oi_1 _24720_ (.A1(_14391_),
    .A2(_02792_),
    .Y(_02794_),
    .B1(net4571));
 sg13g2_o21ai_1 _24721_ (.B1(_02794_),
    .Y(_02795_),
    .A1(_14391_),
    .A2(_02792_));
 sg13g2_a21oi_1 _24722_ (.A1(net4571),
    .A2(\u_inv.d_next[100] ),
    .Y(_02796_),
    .B1(net3789));
 sg13g2_a22oi_1 _24723_ (.Y(_02797_),
    .B1(_02795_),
    .B2(_02796_),
    .A2(_02791_),
    .A1(net3789));
 sg13g2_and2_1 _24724_ (.A(net3435),
    .B(_02797_),
    .X(_02798_));
 sg13g2_xnor2_1 _24725_ (.Y(_02799_),
    .A(net3441),
    .B(_02797_));
 sg13g2_nand2_1 _24726_ (.Y(_02800_),
    .A(_02769_),
    .B(_02785_));
 sg13g2_nor2_1 _24727_ (.A(_02770_),
    .B(_02786_),
    .Y(_02801_));
 sg13g2_a21oi_2 _24728_ (.B1(_02800_),
    .Y(_02802_),
    .A2(_02801_),
    .A1(_02758_));
 sg13g2_nor2_1 _24729_ (.A(_02799_),
    .B(_02802_),
    .Y(_02803_));
 sg13g2_xor2_1 _24730_ (.B(_02802_),
    .A(_02799_),
    .X(_02804_));
 sg13g2_nor2_1 _24731_ (.A(net4345),
    .B(_02797_),
    .Y(_02805_));
 sg13g2_o21ai_1 _24732_ (.B1(net3896),
    .Y(_02806_),
    .A1(net4296),
    .A2(_02804_));
 sg13g2_nand2_1 _24733_ (.Y(_02807_),
    .A(net2612),
    .B(net3965));
 sg13g2_o21ai_1 _24734_ (.B1(_02807_),
    .Y(_00376_),
    .A1(_02805_),
    .A2(_02806_));
 sg13g2_nor2_1 _24735_ (.A(_02798_),
    .B(_02803_),
    .Y(_02808_));
 sg13g2_nand2_1 _24736_ (.Y(_02809_),
    .A(_10608_),
    .B(net3853));
 sg13g2_o21ai_1 _24737_ (.B1(_14390_),
    .Y(_02810_),
    .A1(_14391_),
    .A2(_02792_));
 sg13g2_xnor2_1 _24738_ (.Y(_02811_),
    .A(_14389_),
    .B(_02810_));
 sg13g2_a22oi_1 _24739_ (.Y(_02812_),
    .B1(_02811_),
    .B2(net4692),
    .A2(_02809_),
    .A1(net3731));
 sg13g2_a21oi_1 _24740_ (.A1(_14391_),
    .A2(_02790_),
    .Y(_02813_),
    .B1(_14635_));
 sg13g2_or2_1 _24741_ (.X(_02814_),
    .B(_02813_),
    .A(_14389_));
 sg13g2_a21oi_1 _24742_ (.A1(_14389_),
    .A2(_02813_),
    .Y(_02815_),
    .B1(net3853));
 sg13g2_a21oi_2 _24743_ (.B1(_02812_),
    .Y(_02816_),
    .A2(_02815_),
    .A1(_02814_));
 sg13g2_xnor2_1 _24744_ (.Y(_02817_),
    .A(net3481),
    .B(_02816_));
 sg13g2_xor2_1 _24745_ (.B(_02817_),
    .A(_02808_),
    .X(_02818_));
 sg13g2_o21ai_1 _24746_ (.B1(net3896),
    .Y(_02819_),
    .A1(net4346),
    .A2(_02816_));
 sg13g2_a21oi_1 _24747_ (.A1(net4346),
    .A2(_02818_),
    .Y(_02820_),
    .B1(_02819_));
 sg13g2_a21o_1 _24748_ (.A2(net3965),
    .A1(net3066),
    .B1(_02820_),
    .X(_00377_));
 sg13g2_a21oi_1 _24749_ (.A1(_14392_),
    .A2(_02790_),
    .Y(_02821_),
    .B1(_14637_));
 sg13g2_xnor2_1 _24750_ (.Y(_02822_),
    .A(_14385_),
    .B(_02821_));
 sg13g2_a21oi_1 _24751_ (.A1(_15345_),
    .A2(_02793_),
    .Y(_02823_),
    .B1(_15454_));
 sg13g2_a21oi_1 _24752_ (.A1(_14386_),
    .A2(_02823_),
    .Y(_02824_),
    .B1(net4571));
 sg13g2_o21ai_1 _24753_ (.B1(_02824_),
    .Y(_02825_),
    .A1(_14386_),
    .A2(_02823_));
 sg13g2_a21oi_1 _24754_ (.A1(net4570),
    .A2(\u_inv.d_next[102] ),
    .Y(_02826_),
    .B1(net3789));
 sg13g2_a22oi_1 _24755_ (.Y(_02827_),
    .B1(_02825_),
    .B2(_02826_),
    .A2(_02822_),
    .A1(net3788));
 sg13g2_and2_1 _24756_ (.A(net3439),
    .B(_02827_),
    .X(_02828_));
 sg13g2_xnor2_1 _24757_ (.Y(_02829_),
    .A(net3439),
    .B(_02827_));
 sg13g2_a21oi_2 _24758_ (.B1(_02798_),
    .Y(_02830_),
    .A2(_02816_),
    .A1(net3441));
 sg13g2_nand2b_2 _24759_ (.Y(_02831_),
    .B(_02817_),
    .A_N(_02799_));
 sg13g2_o21ai_1 _24760_ (.B1(_02830_),
    .Y(_02832_),
    .A1(_02802_),
    .A2(_02831_));
 sg13g2_nor2b_1 _24761_ (.A(_02829_),
    .B_N(_02832_),
    .Y(_02833_));
 sg13g2_xor2_1 _24762_ (.B(_02832_),
    .A(_02829_),
    .X(_02834_));
 sg13g2_a21oi_1 _24763_ (.A1(net4350),
    .A2(_02834_),
    .Y(_02835_),
    .B1(net4236));
 sg13g2_o21ai_1 _24764_ (.B1(_02835_),
    .Y(_02836_),
    .A1(net4350),
    .A2(_02827_));
 sg13g2_o21ai_1 _24765_ (.B1(_02836_),
    .Y(_00378_),
    .A1(_10608_),
    .A2(net4034));
 sg13g2_nand2_1 _24766_ (.Y(_02837_),
    .A(_10607_),
    .B(net3853));
 sg13g2_o21ai_1 _24767_ (.B1(_14384_),
    .Y(_02838_),
    .A1(_14386_),
    .A2(_02823_));
 sg13g2_xnor2_1 _24768_ (.Y(_02839_),
    .A(_14382_),
    .B(_02838_));
 sg13g2_a22oi_1 _24769_ (.Y(_02840_),
    .B1(_02839_),
    .B2(net4692),
    .A2(_02837_),
    .A1(net3731));
 sg13g2_o21ai_1 _24770_ (.B1(_14633_),
    .Y(_02841_),
    .A1(_14385_),
    .A2(_02821_));
 sg13g2_or2_1 _24771_ (.X(_02842_),
    .B(_02841_),
    .A(_14383_));
 sg13g2_a21oi_1 _24772_ (.A1(_14383_),
    .A2(_02841_),
    .Y(_02843_),
    .B1(net3853));
 sg13g2_a21oi_2 _24773_ (.B1(_02840_),
    .Y(_02844_),
    .A2(_02843_),
    .A1(_02842_));
 sg13g2_and2_1 _24774_ (.A(net3439),
    .B(_02844_),
    .X(_02845_));
 sg13g2_xnor2_1 _24775_ (.Y(_02846_),
    .A(net3439),
    .B(_02844_));
 sg13g2_nor2_1 _24776_ (.A(_02828_),
    .B(_02833_),
    .Y(_02847_));
 sg13g2_xnor2_1 _24777_ (.Y(_02848_),
    .A(_02846_),
    .B(_02847_));
 sg13g2_o21ai_1 _24778_ (.B1(net3899),
    .Y(_02849_),
    .A1(net4350),
    .A2(_02844_));
 sg13g2_a21oi_1 _24779_ (.A1(net4350),
    .A2(_02848_),
    .Y(_02850_),
    .B1(_02849_));
 sg13g2_a21o_1 _24780_ (.A2(net3965),
    .A1(net3068),
    .B1(_02850_),
    .X(_00379_));
 sg13g2_a21oi_1 _24781_ (.A1(_14594_),
    .A2(_02713_),
    .Y(_02851_),
    .B1(_14408_));
 sg13g2_nor2_1 _24782_ (.A(_14639_),
    .B(_02851_),
    .Y(_02852_));
 sg13g2_xnor2_1 _24783_ (.Y(_02853_),
    .A(_14378_),
    .B(_02852_));
 sg13g2_a21oi_2 _24784_ (.B1(_15462_),
    .Y(_02854_),
    .A2(_02717_),
    .A1(_15350_));
 sg13g2_a21oi_1 _24785_ (.A1(_14379_),
    .A2(_02854_),
    .Y(_02855_),
    .B1(net4573));
 sg13g2_o21ai_1 _24786_ (.B1(_02855_),
    .Y(_02856_),
    .A1(_14379_),
    .A2(_02854_));
 sg13g2_a21oi_1 _24787_ (.A1(net4573),
    .A2(\u_inv.d_next[104] ),
    .Y(_02857_),
    .B1(net3790));
 sg13g2_a22oi_1 _24788_ (.Y(_02858_),
    .B1(_02856_),
    .B2(_02857_),
    .A2(_02853_),
    .A1(net3791));
 sg13g2_and2_1 _24789_ (.A(net3439),
    .B(_02858_),
    .X(_02859_));
 sg13g2_xnor2_1 _24790_ (.Y(_02860_),
    .A(net3439),
    .B(_02858_));
 sg13g2_a21oi_1 _24791_ (.A1(_02756_),
    .A2(_02801_),
    .Y(_02861_),
    .B1(_02800_));
 sg13g2_nor4_1 _24792_ (.A(_02829_),
    .B(_02831_),
    .C(_02846_),
    .D(_02861_),
    .Y(_02862_));
 sg13g2_nor3_1 _24793_ (.A(_02829_),
    .B(_02830_),
    .C(_02846_),
    .Y(_02863_));
 sg13g2_or4_1 _24794_ (.A(_02828_),
    .B(_02845_),
    .C(_02862_),
    .D(_02863_),
    .X(_02864_));
 sg13g2_nand3_1 _24795_ (.B(_02751_),
    .C(_02801_),
    .A(_02724_),
    .Y(_02865_));
 sg13g2_nor4_1 _24796_ (.A(_02829_),
    .B(_02831_),
    .C(_02846_),
    .D(_02865_),
    .Y(_02866_));
 sg13g2_a21oi_1 _24797_ (.A1(_02734_),
    .A2(_02866_),
    .Y(_02867_),
    .B1(_02864_));
 sg13g2_or2_1 _24798_ (.X(_02868_),
    .B(_02867_),
    .A(_02860_));
 sg13g2_xnor2_1 _24799_ (.Y(_02869_),
    .A(_02860_),
    .B(_02867_));
 sg13g2_o21ai_1 _24800_ (.B1(net3899),
    .Y(_02870_),
    .A1(net4350),
    .A2(_02858_));
 sg13g2_a21oi_1 _24801_ (.A1(net4350),
    .A2(_02869_),
    .Y(_02871_),
    .B1(_02870_));
 sg13g2_a21o_1 _24802_ (.A2(net3966),
    .A1(net2834),
    .B1(_02871_),
    .X(_00380_));
 sg13g2_nand2_1 _24803_ (.Y(_02872_),
    .A(net2796),
    .B(net3966));
 sg13g2_nand2b_1 _24804_ (.Y(_02873_),
    .B(_02868_),
    .A_N(_02859_));
 sg13g2_nor2_1 _24805_ (.A(_14376_),
    .B(_14377_),
    .Y(_02874_));
 sg13g2_o21ai_1 _24806_ (.B1(_02874_),
    .Y(_02875_),
    .A1(_14379_),
    .A2(_02854_));
 sg13g2_a21oi_1 _24807_ (.A1(_14376_),
    .A2(_14377_),
    .Y(_02876_),
    .B1(net4572));
 sg13g2_o21ai_1 _24808_ (.B1(_02876_),
    .Y(_02877_),
    .A1(_15338_),
    .A2(_02854_));
 sg13g2_nand2b_1 _24809_ (.Y(_02878_),
    .B(_02875_),
    .A_N(_02877_));
 sg13g2_a21oi_1 _24810_ (.A1(net4573),
    .A2(\u_inv.d_next[105] ),
    .Y(_02879_),
    .B1(net3791));
 sg13g2_o21ai_1 _24811_ (.B1(_14641_),
    .Y(_02880_),
    .A1(_14378_),
    .A2(_02852_));
 sg13g2_xor2_1 _24812_ (.B(_02880_),
    .A(_14376_),
    .X(_02881_));
 sg13g2_a22oi_1 _24813_ (.Y(_02882_),
    .B1(_02881_),
    .B2(net3790),
    .A2(_02879_),
    .A1(_02878_));
 sg13g2_xnor2_1 _24814_ (.Y(_02883_),
    .A(net3439),
    .B(_02882_));
 sg13g2_o21ai_1 _24815_ (.B1(net4350),
    .Y(_02884_),
    .A1(_02873_),
    .A2(_02883_));
 sg13g2_a21oi_1 _24816_ (.A1(_02873_),
    .A2(_02883_),
    .Y(_02885_),
    .B1(_02884_));
 sg13g2_o21ai_1 _24817_ (.B1(net3896),
    .Y(_02886_),
    .A1(net4345),
    .A2(_02882_));
 sg13g2_o21ai_1 _24818_ (.B1(_02872_),
    .Y(_00381_),
    .A1(_02885_),
    .A2(_02886_));
 sg13g2_o21ai_1 _24819_ (.B1(_14380_),
    .Y(_02887_),
    .A1(_14639_),
    .A2(_02851_));
 sg13g2_a21oi_1 _24820_ (.A1(_14643_),
    .A2(_02887_),
    .Y(_02888_),
    .B1(_14374_));
 sg13g2_nand3_1 _24821_ (.B(_14643_),
    .C(_02887_),
    .A(_14374_),
    .Y(_02889_));
 sg13g2_nand2b_1 _24822_ (.Y(_02890_),
    .B(_02889_),
    .A_N(_02888_));
 sg13g2_o21ai_1 _24823_ (.B1(_15468_),
    .Y(_02891_),
    .A1(_15338_),
    .A2(_02854_));
 sg13g2_o21ai_1 _24824_ (.B1(net4692),
    .Y(_02892_),
    .A1(_14374_),
    .A2(_02891_));
 sg13g2_a21o_1 _24825_ (.A2(_02891_),
    .A1(_14374_),
    .B1(_02892_),
    .X(_02893_));
 sg13g2_a21oi_1 _24826_ (.A1(net4573),
    .A2(\u_inv.d_next[106] ),
    .Y(_02894_),
    .B1(net3791));
 sg13g2_a22oi_1 _24827_ (.Y(_02895_),
    .B1(_02893_),
    .B2(_02894_),
    .A2(_02890_),
    .A1(net3791));
 sg13g2_nand2_1 _24828_ (.Y(_02896_),
    .A(net3440),
    .B(_02895_));
 sg13g2_xnor2_1 _24829_ (.Y(_02897_),
    .A(net3480),
    .B(_02895_));
 sg13g2_inv_1 _24830_ (.Y(_02898_),
    .A(_02897_));
 sg13g2_a21o_1 _24831_ (.A2(_02882_),
    .A1(net3439),
    .B1(_02859_),
    .X(_02899_));
 sg13g2_nor2_1 _24832_ (.A(_02868_),
    .B(_02883_),
    .Y(_02900_));
 sg13g2_nor2_1 _24833_ (.A(_02899_),
    .B(_02900_),
    .Y(_02901_));
 sg13g2_xnor2_1 _24834_ (.Y(_02902_),
    .A(_02898_),
    .B(_02901_));
 sg13g2_a21oi_1 _24835_ (.A1(net4350),
    .A2(_02902_),
    .Y(_02903_),
    .B1(net4236));
 sg13g2_o21ai_1 _24836_ (.B1(_02903_),
    .Y(_02904_),
    .A1(net4357),
    .A2(_02895_));
 sg13g2_o21ai_1 _24837_ (.B1(_02904_),
    .Y(_00382_),
    .A1(_10606_),
    .A2(net4034));
 sg13g2_nand2_1 _24838_ (.Y(_02905_),
    .A(net2445),
    .B(net3966));
 sg13g2_nand2b_1 _24839_ (.Y(_02906_),
    .B(net3853),
    .A_N(\u_inv.d_next[107] ));
 sg13g2_a21oi_1 _24840_ (.A1(_14374_),
    .A2(_02891_),
    .Y(_02907_),
    .B1(_14372_));
 sg13g2_xnor2_1 _24841_ (.Y(_02908_),
    .A(_14371_),
    .B(_02907_));
 sg13g2_a22oi_1 _24842_ (.Y(_02909_),
    .B1(_02908_),
    .B2(net4692),
    .A2(_02906_),
    .A1(net3731));
 sg13g2_o21ai_1 _24843_ (.B1(_14371_),
    .Y(_02910_),
    .A1(_14644_),
    .A2(_02888_));
 sg13g2_or3_1 _24844_ (.A(_14371_),
    .B(_14644_),
    .C(_02888_),
    .X(_02911_));
 sg13g2_and3_1 _24845_ (.X(_02912_),
    .A(net3791),
    .B(_02910_),
    .C(_02911_));
 sg13g2_nor2_1 _24846_ (.A(_02909_),
    .B(_02912_),
    .Y(_02913_));
 sg13g2_or3_1 _24847_ (.A(net3482),
    .B(_02909_),
    .C(_02912_),
    .X(_02914_));
 sg13g2_o21ai_1 _24848_ (.B1(net3482),
    .Y(_02915_),
    .A1(_02909_),
    .A2(_02912_));
 sg13g2_nand2_1 _24849_ (.Y(_02916_),
    .A(_02914_),
    .B(_02915_));
 sg13g2_o21ai_1 _24850_ (.B1(_02896_),
    .Y(_02917_),
    .A1(_02898_),
    .A2(_02901_));
 sg13g2_o21ai_1 _24851_ (.B1(net4352),
    .Y(_02918_),
    .A1(_02916_),
    .A2(_02917_));
 sg13g2_a21oi_1 _24852_ (.A1(_02916_),
    .A2(_02917_),
    .Y(_02919_),
    .B1(_02918_));
 sg13g2_o21ai_1 _24853_ (.B1(net3902),
    .Y(_02920_),
    .A1(net4357),
    .A2(_02913_));
 sg13g2_o21ai_1 _24854_ (.B1(_02905_),
    .Y(_00383_),
    .A1(_02919_),
    .A2(_02920_));
 sg13g2_o21ai_1 _24855_ (.B1(_14646_),
    .Y(_02921_),
    .A1(_14375_),
    .A2(_02887_));
 sg13g2_xnor2_1 _24856_ (.Y(_02922_),
    .A(_14366_),
    .B(_02921_));
 sg13g2_o21ai_1 _24857_ (.B1(_15471_),
    .Y(_02923_),
    .A1(_15339_),
    .A2(_02854_));
 sg13g2_nand2b_1 _24858_ (.Y(_02924_),
    .B(_02923_),
    .A_N(_14366_));
 sg13g2_nand2b_1 _24859_ (.Y(_02925_),
    .B(_14366_),
    .A_N(_02923_));
 sg13g2_nand3_1 _24860_ (.B(_02924_),
    .C(_02925_),
    .A(net4690),
    .Y(_02926_));
 sg13g2_a21oi_1 _24861_ (.A1(net4576),
    .A2(\u_inv.d_next[108] ),
    .Y(_02927_),
    .B1(net3796));
 sg13g2_a22oi_1 _24862_ (.Y(_02928_),
    .B1(_02926_),
    .B2(_02927_),
    .A2(_02922_),
    .A1(net3796));
 sg13g2_nand2_1 _24863_ (.Y(_02929_),
    .A(net3445),
    .B(_02928_));
 sg13g2_xnor2_1 _24864_ (.Y(_02930_),
    .A(net3445),
    .B(_02928_));
 sg13g2_nand4_1 _24865_ (.B(_02899_),
    .C(_02914_),
    .A(_02897_),
    .Y(_02931_),
    .D(_02915_));
 sg13g2_nand3_1 _24866_ (.B(_02914_),
    .C(_02931_),
    .A(_02896_),
    .Y(_02932_));
 sg13g2_nor4_1 _24867_ (.A(_02860_),
    .B(_02883_),
    .C(_02898_),
    .D(_02916_),
    .Y(_02933_));
 sg13g2_nor2b_1 _24868_ (.A(_02867_),
    .B_N(_02933_),
    .Y(_02934_));
 sg13g2_or2_1 _24869_ (.X(_02935_),
    .B(_02934_),
    .A(_02932_));
 sg13g2_nand2b_1 _24870_ (.Y(_02936_),
    .B(_02935_),
    .A_N(_02930_));
 sg13g2_xnor2_1 _24871_ (.Y(_02937_),
    .A(_02930_),
    .B(_02935_));
 sg13g2_nor2_1 _24872_ (.A(net4356),
    .B(_02928_),
    .Y(_02938_));
 sg13g2_o21ai_1 _24873_ (.B1(net3900),
    .Y(_02939_),
    .A1(net4297),
    .A2(_02937_));
 sg13g2_nand2_1 _24874_ (.Y(_02940_),
    .A(net2292),
    .B(net3968));
 sg13g2_o21ai_1 _24875_ (.B1(_02940_),
    .Y(_00384_),
    .A1(_02938_),
    .A2(_02939_));
 sg13g2_nand2_1 _24876_ (.Y(_02941_),
    .A(net2237),
    .B(net3969));
 sg13g2_nand2_1 _24877_ (.Y(_02942_),
    .A(_15340_),
    .B(_02923_));
 sg13g2_nand3_1 _24878_ (.B(_14365_),
    .C(_02924_),
    .A(_14364_),
    .Y(_02943_));
 sg13g2_nor2_1 _24879_ (.A(net4576),
    .B(_15473_),
    .Y(_02944_));
 sg13g2_nand3_1 _24880_ (.B(_02943_),
    .C(_02944_),
    .A(_02942_),
    .Y(_02945_));
 sg13g2_a21oi_1 _24881_ (.A1(net4576),
    .A2(\u_inv.d_next[109] ),
    .Y(_02946_),
    .B1(net3796));
 sg13g2_a21oi_1 _24882_ (.A1(_14366_),
    .A2(_02921_),
    .Y(_02947_),
    .B1(_14648_));
 sg13g2_xor2_1 _24883_ (.B(_02947_),
    .A(_14364_),
    .X(_02948_));
 sg13g2_a22oi_1 _24884_ (.Y(_02949_),
    .B1(_02948_),
    .B2(net3796),
    .A2(_02946_),
    .A1(_02945_));
 sg13g2_nand2_1 _24885_ (.Y(_02950_),
    .A(net3445),
    .B(_02949_));
 sg13g2_xnor2_1 _24886_ (.Y(_02951_),
    .A(net3445),
    .B(_02949_));
 sg13g2_nand2_1 _24887_ (.Y(_02952_),
    .A(_02929_),
    .B(_02936_));
 sg13g2_o21ai_1 _24888_ (.B1(net4356),
    .Y(_02953_),
    .A1(_02951_),
    .A2(_02952_));
 sg13g2_a21oi_1 _24889_ (.A1(_02951_),
    .A2(_02952_),
    .Y(_02954_),
    .B1(_02953_));
 sg13g2_o21ai_1 _24890_ (.B1(net3900),
    .Y(_02955_),
    .A1(net4356),
    .A2(_02949_));
 sg13g2_o21ai_1 _24891_ (.B1(_02941_),
    .Y(_00385_),
    .A1(_02954_),
    .A2(_02955_));
 sg13g2_a21oi_1 _24892_ (.A1(_14367_),
    .A2(_02921_),
    .Y(_02956_),
    .B1(_14650_));
 sg13g2_xnor2_1 _24893_ (.Y(_02957_),
    .A(_14361_),
    .B(_02956_));
 sg13g2_a21oi_1 _24894_ (.A1(_15474_),
    .A2(_02942_),
    .Y(_02958_),
    .B1(_14362_));
 sg13g2_nand3_1 _24895_ (.B(_15474_),
    .C(_02942_),
    .A(_14362_),
    .Y(_02959_));
 sg13g2_nand3b_1 _24896_ (.B(_02959_),
    .C(net4690),
    .Y(_02960_),
    .A_N(_02958_));
 sg13g2_a21oi_1 _24897_ (.A1(net4576),
    .A2(\u_inv.d_next[110] ),
    .Y(_02961_),
    .B1(net3796));
 sg13g2_a22oi_1 _24898_ (.Y(_02962_),
    .B1(_02960_),
    .B2(_02961_),
    .A2(_02957_),
    .A1(net3796));
 sg13g2_nand2_1 _24899_ (.Y(_02963_),
    .A(net3440),
    .B(_02962_));
 sg13g2_xnor2_1 _24900_ (.Y(_02964_),
    .A(net3480),
    .B(_02962_));
 sg13g2_inv_1 _24901_ (.Y(_02965_),
    .A(_02964_));
 sg13g2_nand2_1 _24902_ (.Y(_02966_),
    .A(_02929_),
    .B(_02950_));
 sg13g2_nor2_1 _24903_ (.A(_02930_),
    .B(_02951_),
    .Y(_02967_));
 sg13g2_a21oi_1 _24904_ (.A1(_02935_),
    .A2(_02967_),
    .Y(_02968_),
    .B1(_02966_));
 sg13g2_xnor2_1 _24905_ (.Y(_02969_),
    .A(_02965_),
    .B(_02968_));
 sg13g2_a21oi_1 _24906_ (.A1(net4351),
    .A2(_02969_),
    .Y(_02970_),
    .B1(net4236));
 sg13g2_o21ai_1 _24907_ (.B1(_02970_),
    .Y(_02971_),
    .A1(net4351),
    .A2(_02962_));
 sg13g2_o21ai_1 _24908_ (.B1(_02971_),
    .Y(_00386_),
    .A1(_10605_),
    .A2(net4034));
 sg13g2_a21oi_1 _24909_ (.A1(net4573),
    .A2(\u_inv.d_next[111] ),
    .Y(_02972_),
    .B1(net3796));
 sg13g2_or3_1 _24910_ (.A(_14359_),
    .B(_14360_),
    .C(_02958_),
    .X(_02973_));
 sg13g2_o21ai_1 _24911_ (.B1(_14359_),
    .Y(_02974_),
    .A1(_14360_),
    .A2(_02958_));
 sg13g2_nand3_1 _24912_ (.B(_02973_),
    .C(_02974_),
    .A(net4690),
    .Y(_02975_));
 sg13g2_o21ai_1 _24913_ (.B1(_14651_),
    .Y(_02976_),
    .A1(_14361_),
    .A2(_02956_));
 sg13g2_or2_1 _24914_ (.X(_02977_),
    .B(_02976_),
    .A(_14359_));
 sg13g2_a21oi_1 _24915_ (.A1(_14359_),
    .A2(_02976_),
    .Y(_02978_),
    .B1(net3853));
 sg13g2_a22oi_1 _24916_ (.Y(_02979_),
    .B1(_02977_),
    .B2(_02978_),
    .A2(_02975_),
    .A1(_02972_));
 sg13g2_xnor2_1 _24917_ (.Y(_02980_),
    .A(net3481),
    .B(_02979_));
 sg13g2_o21ai_1 _24918_ (.B1(_02963_),
    .Y(_02981_),
    .A1(_02965_),
    .A2(_02968_));
 sg13g2_xnor2_1 _24919_ (.Y(_02982_),
    .A(_02980_),
    .B(_02981_));
 sg13g2_o21ai_1 _24920_ (.B1(net3898),
    .Y(_02983_),
    .A1(net4351),
    .A2(_02979_));
 sg13g2_a21oi_1 _24921_ (.A1(net4352),
    .A2(_02982_),
    .Y(_02984_),
    .B1(_02983_));
 sg13g2_a21o_1 _24922_ (.A2(net3969),
    .A1(net3217),
    .B1(_02984_),
    .X(_00387_));
 sg13g2_a21oi_2 _24923_ (.B1(_14410_),
    .Y(_02985_),
    .A2(_02713_),
    .A1(_14594_));
 sg13g2_nor2_1 _24924_ (.A(_14654_),
    .B(_02985_),
    .Y(_02986_));
 sg13g2_o21ai_1 _24925_ (.B1(_14354_),
    .Y(_02987_),
    .A1(_14654_),
    .A2(_02985_));
 sg13g2_xnor2_1 _24926_ (.Y(_02988_),
    .A(_14353_),
    .B(_02986_));
 sg13g2_o21ai_1 _24927_ (.B1(_15476_),
    .Y(_02989_),
    .A1(_15351_),
    .A2(_02716_));
 sg13g2_a21oi_1 _24928_ (.A1(_14353_),
    .A2(_02989_),
    .Y(_02990_),
    .B1(net4574));
 sg13g2_o21ai_1 _24929_ (.B1(_02990_),
    .Y(_02991_),
    .A1(_14353_),
    .A2(_02989_));
 sg13g2_a21oi_1 _24930_ (.A1(net4574),
    .A2(\u_inv.d_next[112] ),
    .Y(_02992_),
    .B1(net3794));
 sg13g2_a22oi_1 _24931_ (.Y(_02993_),
    .B1(_02991_),
    .B2(_02992_),
    .A2(_02988_),
    .A1(net3794));
 sg13g2_nand2_1 _24932_ (.Y(_02994_),
    .A(net3437),
    .B(_02993_));
 sg13g2_xnor2_1 _24933_ (.Y(_02995_),
    .A(net3480),
    .B(_02993_));
 sg13g2_inv_1 _24934_ (.Y(_02996_),
    .A(_02995_));
 sg13g2_and4_1 _24935_ (.A(_02933_),
    .B(_02964_),
    .C(_02967_),
    .D(_02980_),
    .X(_02997_));
 sg13g2_nand4_1 _24936_ (.B(_02964_),
    .C(_02967_),
    .A(_02932_),
    .Y(_02998_),
    .D(_02980_));
 sg13g2_nand3_1 _24937_ (.B(_02966_),
    .C(_02980_),
    .A(_02964_),
    .Y(_02999_));
 sg13g2_o21ai_1 _24938_ (.B1(net3440),
    .Y(_03000_),
    .A1(_02962_),
    .A2(_02979_));
 sg13g2_nand3_1 _24939_ (.B(_02999_),
    .C(_03000_),
    .A(_02998_),
    .Y(_03001_));
 sg13g2_a21o_1 _24940_ (.A2(_02997_),
    .A1(_02864_),
    .B1(_03001_),
    .X(_03002_));
 sg13g2_and2_1 _24941_ (.A(_02866_),
    .B(_02997_),
    .X(_03003_));
 sg13g2_a21o_2 _24942_ (.A2(_03003_),
    .A1(_02734_),
    .B1(_03002_),
    .X(_03004_));
 sg13g2_nand2_1 _24943_ (.Y(_03005_),
    .A(_02995_),
    .B(_03004_));
 sg13g2_xnor2_1 _24944_ (.Y(_03006_),
    .A(_02995_),
    .B(_03004_));
 sg13g2_a21oi_1 _24945_ (.A1(net4348),
    .A2(_03006_),
    .Y(_03007_),
    .B1(net4236));
 sg13g2_o21ai_1 _24946_ (.B1(_03007_),
    .Y(_03008_),
    .A1(net4351),
    .A2(_02993_));
 sg13g2_o21ai_1 _24947_ (.B1(_03008_),
    .Y(_00388_),
    .A1(_10604_),
    .A2(net4034));
 sg13g2_nand2_1 _24948_ (.Y(_03009_),
    .A(_02994_),
    .B(_03005_));
 sg13g2_a21oi_1 _24949_ (.A1(_14353_),
    .A2(_02989_),
    .Y(_03010_),
    .B1(_14351_));
 sg13g2_nand3_1 _24950_ (.B(_14353_),
    .C(_02989_),
    .A(_14351_),
    .Y(_03011_));
 sg13g2_a21oi_1 _24951_ (.A1(_14352_),
    .A2(_03010_),
    .Y(_03012_),
    .B1(_15426_));
 sg13g2_nand3_1 _24952_ (.B(_03011_),
    .C(_03012_),
    .A(net4689),
    .Y(_03013_));
 sg13g2_a21oi_1 _24953_ (.A1(net4574),
    .A2(\u_inv.d_next[113] ),
    .Y(_03014_),
    .B1(net3794));
 sg13g2_nand2b_1 _24954_ (.Y(_03015_),
    .B(_02987_),
    .A_N(_14596_));
 sg13g2_xnor2_1 _24955_ (.Y(_03016_),
    .A(_14350_),
    .B(_03015_));
 sg13g2_a22oi_1 _24956_ (.Y(_03017_),
    .B1(_03016_),
    .B2(net3794),
    .A2(_03014_),
    .A1(_03013_));
 sg13g2_nand2_1 _24957_ (.Y(_03018_),
    .A(net3437),
    .B(_03017_));
 sg13g2_xnor2_1 _24958_ (.Y(_03019_),
    .A(net3437),
    .B(_03017_));
 sg13g2_xor2_1 _24959_ (.B(_03019_),
    .A(_03009_),
    .X(_03020_));
 sg13g2_o21ai_1 _24960_ (.B1(net3896),
    .Y(_03021_),
    .A1(net4348),
    .A2(_03017_));
 sg13g2_a21oi_1 _24961_ (.A1(net4348),
    .A2(_03020_),
    .Y(_03022_),
    .B1(_03021_));
 sg13g2_a21o_1 _24962_ (.A2(net3967),
    .A1(net2876),
    .B1(_03022_),
    .X(_00389_));
 sg13g2_o21ai_1 _24963_ (.B1(_14355_),
    .Y(_03023_),
    .A1(_14654_),
    .A2(_02985_));
 sg13g2_a21oi_1 _24964_ (.A1(_14597_),
    .A2(_03023_),
    .Y(_03024_),
    .B1(_14346_));
 sg13g2_and3_1 _24965_ (.X(_03025_),
    .A(_14346_),
    .B(_14597_),
    .C(_03023_));
 sg13g2_o21ai_1 _24966_ (.B1(net3792),
    .Y(_03026_),
    .A1(_03024_),
    .A2(_03025_));
 sg13g2_a21o_1 _24967_ (.A2(_03011_),
    .A1(_15427_),
    .B1(_14345_),
    .X(_03027_));
 sg13g2_nand3_1 _24968_ (.B(_15427_),
    .C(_03011_),
    .A(_14345_),
    .Y(_03028_));
 sg13g2_nand3_1 _24969_ (.B(_03027_),
    .C(_03028_),
    .A(net4689),
    .Y(_03029_));
 sg13g2_o21ai_1 _24970_ (.B1(_03029_),
    .Y(_03030_),
    .A1(net4689),
    .A2(_10603_));
 sg13g2_o21ai_1 _24971_ (.B1(_03026_),
    .Y(_03031_),
    .A1(net3794),
    .A2(_03030_));
 sg13g2_nor2_1 _24972_ (.A(net3480),
    .B(_03031_),
    .Y(_03032_));
 sg13g2_xnor2_1 _24973_ (.Y(_03033_),
    .A(net3480),
    .B(_03031_));
 sg13g2_nand2_1 _24974_ (.Y(_03034_),
    .A(_02994_),
    .B(_03018_));
 sg13g2_nand2b_1 _24975_ (.Y(_03035_),
    .B(_03005_),
    .A_N(_03034_));
 sg13g2_o21ai_1 _24976_ (.B1(_03035_),
    .Y(_03036_),
    .A1(net3437),
    .A2(_03017_));
 sg13g2_nor2_1 _24977_ (.A(_03033_),
    .B(_03036_),
    .Y(_03037_));
 sg13g2_xnor2_1 _24978_ (.Y(_03038_),
    .A(_03033_),
    .B(_03036_));
 sg13g2_nand2_1 _24979_ (.Y(_03039_),
    .A(net4297),
    .B(_03031_));
 sg13g2_a21oi_1 _24980_ (.A1(net4348),
    .A2(_03038_),
    .Y(_03040_),
    .B1(net4236));
 sg13g2_a22oi_1 _24981_ (.Y(_03041_),
    .B1(_03039_),
    .B2(_03040_),
    .A2(net3967),
    .A1(net2917));
 sg13g2_inv_1 _24982_ (.Y(_00390_),
    .A(_03041_));
 sg13g2_nand2_1 _24983_ (.Y(_03042_),
    .A(net2540),
    .B(net3967));
 sg13g2_a21oi_1 _24984_ (.A1(net4574),
    .A2(\u_inv.d_next[115] ),
    .Y(_03043_),
    .B1(net3794));
 sg13g2_a21o_1 _24985_ (.A2(_03027_),
    .A1(_14344_),
    .B1(_14342_),
    .X(_03044_));
 sg13g2_nand3_1 _24986_ (.B(_14344_),
    .C(_03027_),
    .A(_14342_),
    .Y(_03045_));
 sg13g2_nand3_1 _24987_ (.B(_03044_),
    .C(_03045_),
    .A(net4689),
    .Y(_03046_));
 sg13g2_o21ai_1 _24988_ (.B1(_14343_),
    .Y(_03047_),
    .A1(_14598_),
    .A2(_03024_));
 sg13g2_nor3_1 _24989_ (.A(_14343_),
    .B(_14598_),
    .C(_03024_),
    .Y(_03048_));
 sg13g2_nor2_1 _24990_ (.A(net3854),
    .B(_03048_),
    .Y(_03049_));
 sg13g2_a22oi_1 _24991_ (.Y(_03050_),
    .B1(_03047_),
    .B2(_03049_),
    .A2(_03046_),
    .A1(_03043_));
 sg13g2_xnor2_1 _24992_ (.Y(_03051_),
    .A(net3480),
    .B(_03050_));
 sg13g2_nor2_1 _24993_ (.A(_03032_),
    .B(_03037_),
    .Y(_03052_));
 sg13g2_o21ai_1 _24994_ (.B1(net4348),
    .Y(_03053_),
    .A1(_03051_),
    .A2(_03052_));
 sg13g2_a21oi_1 _24995_ (.A1(_03051_),
    .A2(_03052_),
    .Y(_03054_),
    .B1(_03053_));
 sg13g2_o21ai_1 _24996_ (.B1(net3897),
    .Y(_03055_),
    .A1(net4347),
    .A2(_03050_));
 sg13g2_o21ai_1 _24997_ (.B1(_03042_),
    .Y(_00391_),
    .A1(_03054_),
    .A2(_03055_));
 sg13g2_o21ai_1 _24998_ (.B1(_14600_),
    .Y(_03056_),
    .A1(_14347_),
    .A2(_03023_));
 sg13g2_nand2_1 _24999_ (.Y(_03057_),
    .A(_14332_),
    .B(_03056_));
 sg13g2_xnor2_1 _25000_ (.Y(_03058_),
    .A(_14332_),
    .B(_03056_));
 sg13g2_a21oi_1 _25001_ (.A1(_15334_),
    .A2(_02989_),
    .Y(_03059_),
    .B1(_15430_));
 sg13g2_or2_1 _25002_ (.X(_03060_),
    .B(_03059_),
    .A(_14332_));
 sg13g2_a21oi_1 _25003_ (.A1(_14332_),
    .A2(_03059_),
    .Y(_03061_),
    .B1(net4574));
 sg13g2_nand2_1 _25004_ (.Y(_03062_),
    .A(_03060_),
    .B(_03061_));
 sg13g2_a21oi_1 _25005_ (.A1(net4574),
    .A2(\u_inv.d_next[116] ),
    .Y(_03063_),
    .B1(net3792));
 sg13g2_a22oi_1 _25006_ (.Y(_03064_),
    .B1(_03062_),
    .B2(_03063_),
    .A2(_03058_),
    .A1(net3792));
 sg13g2_nand2_1 _25007_ (.Y(_03065_),
    .A(net3436),
    .B(_03064_));
 sg13g2_xnor2_1 _25008_ (.Y(_03066_),
    .A(net3436),
    .B(_03064_));
 sg13g2_nand2b_1 _25009_ (.Y(_03067_),
    .B(_03051_),
    .A_N(_03033_));
 sg13g2_nand3b_1 _25010_ (.B(_03034_),
    .C(_03051_),
    .Y(_03068_),
    .A_N(_03033_));
 sg13g2_a21oi_1 _25011_ (.A1(net3436),
    .A2(_03050_),
    .Y(_03069_),
    .B1(_03032_));
 sg13g2_nand2_1 _25012_ (.Y(_03070_),
    .A(_03068_),
    .B(_03069_));
 sg13g2_nor3_1 _25013_ (.A(_02996_),
    .B(_03019_),
    .C(_03067_),
    .Y(_03071_));
 sg13g2_a21oi_1 _25014_ (.A1(_03004_),
    .A2(_03071_),
    .Y(_03072_),
    .B1(_03070_));
 sg13g2_or2_1 _25015_ (.X(_03073_),
    .B(_03072_),
    .A(_03066_));
 sg13g2_xnor2_1 _25016_ (.Y(_03074_),
    .A(_03066_),
    .B(_03072_));
 sg13g2_o21ai_1 _25017_ (.B1(net3897),
    .Y(_03075_),
    .A1(net4347),
    .A2(_03064_));
 sg13g2_a21oi_1 _25018_ (.A1(net4347),
    .A2(_03074_),
    .Y(_03076_),
    .B1(_03075_));
 sg13g2_a21o_1 _25019_ (.A2(net3967),
    .A1(net3201),
    .B1(_03076_),
    .X(_00392_));
 sg13g2_nand2_1 _25020_ (.Y(_03077_),
    .A(net2344),
    .B(net3967));
 sg13g2_nand3_1 _25021_ (.B(_14331_),
    .C(_03060_),
    .A(_14330_),
    .Y(_03078_));
 sg13g2_or3_1 _25022_ (.A(_14330_),
    .B(_14332_),
    .C(_03059_),
    .X(_03079_));
 sg13g2_nand4_1 _25023_ (.B(_15432_),
    .C(_03078_),
    .A(net4689),
    .Y(_03080_),
    .D(_03079_));
 sg13g2_a21oi_1 _25024_ (.A1(net4575),
    .A2(\u_inv.d_next[117] ),
    .Y(_03081_),
    .B1(net3792));
 sg13g2_and2_1 _25025_ (.A(_14602_),
    .B(_03057_),
    .X(_03082_));
 sg13g2_xor2_1 _25026_ (.B(_03082_),
    .A(_14330_),
    .X(_03083_));
 sg13g2_a22oi_1 _25027_ (.Y(_03084_),
    .B1(_03083_),
    .B2(net3792),
    .A2(_03081_),
    .A1(_03080_));
 sg13g2_nor2_1 _25028_ (.A(net3436),
    .B(_03084_),
    .Y(_03085_));
 sg13g2_xnor2_1 _25029_ (.Y(_03086_),
    .A(net3436),
    .B(_03084_));
 sg13g2_nand2_1 _25030_ (.Y(_03087_),
    .A(_03065_),
    .B(_03073_));
 sg13g2_o21ai_1 _25031_ (.B1(net4347),
    .Y(_03088_),
    .A1(_03086_),
    .A2(_03087_));
 sg13g2_a21oi_1 _25032_ (.A1(_03086_),
    .A2(_03087_),
    .Y(_03089_),
    .B1(_03088_));
 sg13g2_o21ai_1 _25033_ (.B1(net3897),
    .Y(_03090_),
    .A1(net4347),
    .A2(_03084_));
 sg13g2_o21ai_1 _25034_ (.B1(_03077_),
    .Y(_00393_),
    .A1(_03089_),
    .A2(_03090_));
 sg13g2_a21oi_1 _25035_ (.A1(_14333_),
    .A2(_03056_),
    .Y(_03091_),
    .B1(_14603_));
 sg13g2_xnor2_1 _25036_ (.Y(_03092_),
    .A(_14336_),
    .B(_03091_));
 sg13g2_a21oi_1 _25037_ (.A1(_15433_),
    .A2(_03079_),
    .Y(_03093_),
    .B1(_14337_));
 sg13g2_nand3_1 _25038_ (.B(_15433_),
    .C(_03079_),
    .A(_14337_),
    .Y(_03094_));
 sg13g2_nand3b_1 _25039_ (.B(_03094_),
    .C(net4689),
    .Y(_03095_),
    .A_N(_03093_));
 sg13g2_a21oi_1 _25040_ (.A1(net4575),
    .A2(\u_inv.d_next[118] ),
    .Y(_03096_),
    .B1(net3792));
 sg13g2_a22oi_1 _25041_ (.Y(_03097_),
    .B1(_03095_),
    .B2(_03096_),
    .A2(_03092_),
    .A1(net3792));
 sg13g2_nand2_1 _25042_ (.Y(_03098_),
    .A(net3449),
    .B(_03097_));
 sg13g2_xnor2_1 _25043_ (.Y(_03099_),
    .A(net3436),
    .B(_03097_));
 sg13g2_o21ai_1 _25044_ (.B1(net3436),
    .Y(_03100_),
    .A1(_03064_),
    .A2(_03084_));
 sg13g2_a21oi_1 _25045_ (.A1(_03073_),
    .A2(_03100_),
    .Y(_03101_),
    .B1(_03085_));
 sg13g2_nand2b_1 _25046_ (.Y(_03102_),
    .B(_03101_),
    .A_N(_03099_));
 sg13g2_xor2_1 _25047_ (.B(_03101_),
    .A(_03099_),
    .X(_03103_));
 sg13g2_o21ai_1 _25048_ (.B1(net3897),
    .Y(_03104_),
    .A1(net4347),
    .A2(_03097_));
 sg13g2_a21oi_1 _25049_ (.A1(net4347),
    .A2(_03103_),
    .Y(_03105_),
    .B1(_03104_));
 sg13g2_a21o_1 _25050_ (.A2(net3967),
    .A1(net3081),
    .B1(_03105_),
    .X(_00394_));
 sg13g2_nand2_1 _25051_ (.Y(_03106_),
    .A(net2598),
    .B(net3967));
 sg13g2_a21oi_1 _25052_ (.A1(net4574),
    .A2(\u_inv.d_next[119] ),
    .Y(_03107_),
    .B1(net3792));
 sg13g2_or3_1 _25053_ (.A(_14334_),
    .B(_14335_),
    .C(_03093_),
    .X(_03108_));
 sg13g2_o21ai_1 _25054_ (.B1(_14334_),
    .Y(_03109_),
    .A1(_14335_),
    .A2(_03093_));
 sg13g2_nand3_1 _25055_ (.B(_03108_),
    .C(_03109_),
    .A(net4689),
    .Y(_03110_));
 sg13g2_o21ai_1 _25056_ (.B1(_14605_),
    .Y(_03111_),
    .A1(_14336_),
    .A2(_03091_));
 sg13g2_or2_1 _25057_ (.X(_03112_),
    .B(_03111_),
    .A(_14334_));
 sg13g2_a21oi_1 _25058_ (.A1(_14334_),
    .A2(_03111_),
    .Y(_03113_),
    .B1(net3854));
 sg13g2_a22oi_1 _25059_ (.Y(_03114_),
    .B1(_03112_),
    .B2(_03113_),
    .A2(_03110_),
    .A1(_03107_));
 sg13g2_xnor2_1 _25060_ (.Y(_03115_),
    .A(net3436),
    .B(_03114_));
 sg13g2_nand2_1 _25061_ (.Y(_03116_),
    .A(_03098_),
    .B(_03102_));
 sg13g2_o21ai_1 _25062_ (.B1(net4347),
    .Y(_03117_),
    .A1(_03115_),
    .A2(_03116_));
 sg13g2_a21oi_1 _25063_ (.A1(_03115_),
    .A2(_03116_),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_o21ai_1 _25064_ (.B1(net3897),
    .Y(_03119_),
    .A1(net4359),
    .A2(_03114_));
 sg13g2_o21ai_1 _25065_ (.B1(_03106_),
    .Y(_00395_),
    .A1(_03118_),
    .A2(_03119_));
 sg13g2_o21ai_1 _25066_ (.B1(_14357_),
    .Y(_03120_),
    .A1(_14654_),
    .A2(_02985_));
 sg13g2_nand2_1 _25067_ (.Y(_03121_),
    .A(_14608_),
    .B(_03120_));
 sg13g2_xnor2_1 _25068_ (.Y(_03122_),
    .A(_14325_),
    .B(_03121_));
 sg13g2_a21oi_2 _25069_ (.B1(_15437_),
    .Y(_03123_),
    .A2(_02989_),
    .A1(_15335_));
 sg13g2_a21oi_1 _25070_ (.A1(_14325_),
    .A2(_03123_),
    .Y(_03124_),
    .B1(net4575));
 sg13g2_o21ai_1 _25071_ (.B1(_03124_),
    .Y(_03125_),
    .A1(_14325_),
    .A2(_03123_));
 sg13g2_a21oi_1 _25072_ (.A1(net4574),
    .A2(\u_inv.d_next[120] ),
    .Y(_03126_),
    .B1(net3793));
 sg13g2_a22oi_1 _25073_ (.Y(_03127_),
    .B1(_03125_),
    .B2(_03126_),
    .A2(_03122_),
    .A1(net3793));
 sg13g2_nand2_1 _25074_ (.Y(_03128_),
    .A(net3440),
    .B(_03127_));
 sg13g2_xnor2_1 _25075_ (.Y(_03129_),
    .A(net3440),
    .B(_03127_));
 sg13g2_nor4_1 _25076_ (.A(_03066_),
    .B(_03086_),
    .C(_03099_),
    .D(_03115_),
    .Y(_03130_));
 sg13g2_nand2_1 _25077_ (.Y(_03131_),
    .A(_03070_),
    .B(_03130_));
 sg13g2_or3_1 _25078_ (.A(_03099_),
    .B(_03100_),
    .C(_03115_),
    .X(_03132_));
 sg13g2_o21ai_1 _25079_ (.B1(net3449),
    .Y(_03133_),
    .A1(_03097_),
    .A2(_03114_));
 sg13g2_nand3_1 _25080_ (.B(_03132_),
    .C(_03133_),
    .A(_03131_),
    .Y(_03134_));
 sg13g2_and2_1 _25081_ (.A(_03071_),
    .B(_03130_),
    .X(_03135_));
 sg13g2_a21oi_1 _25082_ (.A1(_03004_),
    .A2(_03135_),
    .Y(_03136_),
    .B1(_03134_));
 sg13g2_xnor2_1 _25083_ (.Y(_03137_),
    .A(_03129_),
    .B(_03136_));
 sg13g2_o21ai_1 _25084_ (.B1(net3897),
    .Y(_03138_),
    .A1(net4351),
    .A2(_03127_));
 sg13g2_a21oi_1 _25085_ (.A1(net4351),
    .A2(_03137_),
    .Y(_03139_),
    .B1(_03138_));
 sg13g2_a21o_1 _25086_ (.A2(net3968),
    .A1(net2926),
    .B1(_03139_),
    .X(_00396_));
 sg13g2_and2_1 _25087_ (.A(_14323_),
    .B(_14324_),
    .X(_03140_));
 sg13g2_o21ai_1 _25088_ (.B1(_03140_),
    .Y(_03141_),
    .A1(_14325_),
    .A2(_03123_));
 sg13g2_nor2_1 _25089_ (.A(_15331_),
    .B(_03123_),
    .Y(_03142_));
 sg13g2_nor3_1 _25090_ (.A(net4575),
    .B(_15439_),
    .C(_03142_),
    .Y(_03143_));
 sg13g2_a221oi_1 _25091_ (.B2(_03143_),
    .C1(net3793),
    .B1(_03141_),
    .A1(net4575),
    .Y(_03144_),
    .A2(\u_inv.d_next[121] ));
 sg13g2_a21oi_1 _25092_ (.A1(_14325_),
    .A2(_03121_),
    .Y(_03145_),
    .B1(_14610_));
 sg13g2_xor2_1 _25093_ (.B(_03145_),
    .A(_14323_),
    .X(_03146_));
 sg13g2_a21oi_2 _25094_ (.B1(_03144_),
    .Y(_03147_),
    .A2(_03146_),
    .A1(net3793));
 sg13g2_nand2_1 _25095_ (.Y(_03148_),
    .A(net3448),
    .B(_03147_));
 sg13g2_xnor2_1 _25096_ (.Y(_03149_),
    .A(net3440),
    .B(_03147_));
 sg13g2_o21ai_1 _25097_ (.B1(_03128_),
    .Y(_03150_),
    .A1(_03129_),
    .A2(_03136_));
 sg13g2_xor2_1 _25098_ (.B(_03150_),
    .A(_03149_),
    .X(_03151_));
 sg13g2_o21ai_1 _25099_ (.B1(net3897),
    .Y(_03152_),
    .A1(net4351),
    .A2(_03147_));
 sg13g2_a21oi_1 _25100_ (.A1(net4351),
    .A2(_03151_),
    .Y(_03153_),
    .B1(_03152_));
 sg13g2_a21o_1 _25101_ (.A2(net3967),
    .A1(net3060),
    .B1(_03153_),
    .X(_00397_));
 sg13g2_a21oi_2 _25102_ (.B1(_14326_),
    .Y(_03154_),
    .A2(_03120_),
    .A1(_14608_));
 sg13g2_nor2_1 _25103_ (.A(_14612_),
    .B(_03154_),
    .Y(_03155_));
 sg13g2_o21ai_1 _25104_ (.B1(_14318_),
    .Y(_03156_),
    .A1(_14612_),
    .A2(_03154_));
 sg13g2_xnor2_1 _25105_ (.Y(_03157_),
    .A(_14317_),
    .B(_03155_));
 sg13g2_o21ai_1 _25106_ (.B1(_15440_),
    .Y(_03158_),
    .A1(_15331_),
    .A2(_03123_));
 sg13g2_o21ai_1 _25107_ (.B1(net4689),
    .Y(_03159_),
    .A1(_14317_),
    .A2(_03158_));
 sg13g2_a21o_1 _25108_ (.A2(_03158_),
    .A1(_14317_),
    .B1(_03159_),
    .X(_03160_));
 sg13g2_a21oi_1 _25109_ (.A1(net4575),
    .A2(\u_inv.d_next[122] ),
    .Y(_03161_),
    .B1(net3793));
 sg13g2_a22oi_1 _25110_ (.Y(_03162_),
    .B1(_03160_),
    .B2(_03161_),
    .A2(_03157_),
    .A1(net3793));
 sg13g2_and2_1 _25111_ (.A(net3448),
    .B(_03162_),
    .X(_03163_));
 sg13g2_xnor2_1 _25112_ (.Y(_03164_),
    .A(net3484),
    .B(_03162_));
 sg13g2_o21ai_1 _25113_ (.B1(_03150_),
    .Y(_03165_),
    .A1(net3448),
    .A2(_03147_));
 sg13g2_o21ai_1 _25114_ (.B1(net3448),
    .Y(_03166_),
    .A1(_03127_),
    .A2(_03147_));
 sg13g2_nand2_1 _25115_ (.Y(_03167_),
    .A(_03148_),
    .B(_03165_));
 sg13g2_xnor2_1 _25116_ (.Y(_03168_),
    .A(_03164_),
    .B(_03167_));
 sg13g2_o21ai_1 _25117_ (.B1(net3898),
    .Y(_03169_),
    .A1(net4360),
    .A2(_03162_));
 sg13g2_a21oi_1 _25118_ (.A1(net4364),
    .A2(_03168_),
    .Y(_03170_),
    .B1(_03169_));
 sg13g2_a21o_1 _25119_ (.A2(net3968),
    .A1(net2756),
    .B1(_03170_),
    .X(_00398_));
 sg13g2_nand2b_1 _25120_ (.Y(_03171_),
    .B(net3854),
    .A_N(\u_inv.d_next[123] ));
 sg13g2_a21oi_1 _25121_ (.A1(_14317_),
    .A2(_03158_),
    .Y(_03172_),
    .B1(_14316_));
 sg13g2_xnor2_1 _25122_ (.Y(_03173_),
    .A(_14320_),
    .B(_03172_));
 sg13g2_a22oi_1 _25123_ (.Y(_03174_),
    .B1(_03173_),
    .B2(net4691),
    .A2(_03171_),
    .A1(net3731));
 sg13g2_a21oi_1 _25124_ (.A1(_14614_),
    .A2(_03156_),
    .Y(_03175_),
    .B1(_14321_));
 sg13g2_and3_1 _25125_ (.X(_03176_),
    .A(_14321_),
    .B(_14614_),
    .C(_03156_));
 sg13g2_nor3_2 _25126_ (.A(net3854),
    .B(_03175_),
    .C(_03176_),
    .Y(_03177_));
 sg13g2_nor3_1 _25127_ (.A(net3484),
    .B(_03174_),
    .C(_03177_),
    .Y(_03178_));
 sg13g2_o21ai_1 _25128_ (.B1(net3484),
    .Y(_03179_),
    .A1(_03174_),
    .A2(_03177_));
 sg13g2_nand2b_1 _25129_ (.Y(_03180_),
    .B(_03179_),
    .A_N(_03178_));
 sg13g2_a21oi_1 _25130_ (.A1(_03164_),
    .A2(_03167_),
    .Y(_03181_),
    .B1(_03163_));
 sg13g2_xnor2_1 _25131_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_o21ai_1 _25132_ (.B1(net4297),
    .Y(_03183_),
    .A1(_03174_),
    .A2(_03177_));
 sg13g2_nand2_1 _25133_ (.Y(_03184_),
    .A(net3897),
    .B(_03183_));
 sg13g2_a21oi_1 _25134_ (.A1(net4360),
    .A2(_03182_),
    .Y(_03185_),
    .B1(_03184_));
 sg13g2_a21o_1 _25135_ (.A2(net3968),
    .A1(net3230),
    .B1(_03185_),
    .X(_00399_));
 sg13g2_a21oi_2 _25136_ (.B1(_14616_),
    .Y(_03186_),
    .A2(_03154_),
    .A1(_14322_));
 sg13g2_xnor2_1 _25137_ (.Y(_03187_),
    .A(_14312_),
    .B(_03186_));
 sg13g2_nor3_1 _25138_ (.A(_15329_),
    .B(_15331_),
    .C(_03123_),
    .Y(_03188_));
 sg13g2_o21ai_1 _25139_ (.B1(_14312_),
    .Y(_03189_),
    .A1(_15443_),
    .A2(_03188_));
 sg13g2_or3_1 _25140_ (.A(_14312_),
    .B(_15443_),
    .C(_03188_),
    .X(_03190_));
 sg13g2_nand3_1 _25141_ (.B(_03189_),
    .C(_03190_),
    .A(net4690),
    .Y(_03191_));
 sg13g2_a21oi_1 _25142_ (.A1(net4577),
    .A2(\u_inv.d_next[124] ),
    .Y(_03192_),
    .B1(net3811));
 sg13g2_a22oi_1 _25143_ (.Y(_03193_),
    .B1(_03191_),
    .B2(_03192_),
    .A2(_03187_),
    .A1(net3795));
 sg13g2_nand2_1 _25144_ (.Y(_03194_),
    .A(net3448),
    .B(_03193_));
 sg13g2_xnor2_1 _25145_ (.Y(_03195_),
    .A(net3448),
    .B(_03193_));
 sg13g2_nor2_1 _25146_ (.A(_03163_),
    .B(_03178_),
    .Y(_03196_));
 sg13g2_nand3b_1 _25147_ (.B(_03179_),
    .C(_03164_),
    .Y(_03197_),
    .A_N(_03178_));
 sg13g2_a21oi_1 _25148_ (.A1(_03148_),
    .A2(_03165_),
    .Y(_03198_),
    .B1(_03197_));
 sg13g2_nor2b_2 _25149_ (.A(_03198_),
    .B_N(_03196_),
    .Y(_03199_));
 sg13g2_xnor2_1 _25150_ (.Y(_03200_),
    .A(_03195_),
    .B(_03199_));
 sg13g2_o21ai_1 _25151_ (.B1(net3898),
    .Y(_03201_),
    .A1(net4360),
    .A2(_03193_));
 sg13g2_a21oi_1 _25152_ (.A1(net4360),
    .A2(_03200_),
    .Y(_03202_),
    .B1(_03201_));
 sg13g2_a21o_1 _25153_ (.A2(net3968),
    .A1(net3235),
    .B1(_03202_),
    .X(_00400_));
 sg13g2_a21oi_1 _25154_ (.A1(net4577),
    .A2(\u_inv.d_next[125] ),
    .Y(_03203_),
    .B1(net3811));
 sg13g2_nand3_1 _25155_ (.B(_14311_),
    .C(_03189_),
    .A(_14309_),
    .Y(_03204_));
 sg13g2_a21o_1 _25156_ (.A2(_03189_),
    .A1(_14311_),
    .B1(_14309_),
    .X(_03205_));
 sg13g2_nand3_1 _25157_ (.B(_03204_),
    .C(_03205_),
    .A(net4702),
    .Y(_03206_));
 sg13g2_o21ai_1 _25158_ (.B1(_14619_),
    .Y(_03207_),
    .A1(_14312_),
    .A2(_03186_));
 sg13g2_nand2b_1 _25159_ (.Y(_03208_),
    .B(_14309_),
    .A_N(_03207_));
 sg13g2_a21oi_1 _25160_ (.A1(_14310_),
    .A2(_03207_),
    .Y(_03209_),
    .B1(net3854));
 sg13g2_a22oi_1 _25161_ (.Y(_03210_),
    .B1(_03208_),
    .B2(_03209_),
    .A2(_03206_),
    .A1(_03203_));
 sg13g2_xnor2_1 _25162_ (.Y(_03211_),
    .A(net3449),
    .B(_03210_));
 sg13g2_o21ai_1 _25163_ (.B1(_03194_),
    .Y(_03212_),
    .A1(_03195_),
    .A2(_03199_));
 sg13g2_xor2_1 _25164_ (.B(_03212_),
    .A(_03211_),
    .X(_03213_));
 sg13g2_o21ai_1 _25165_ (.B1(net3898),
    .Y(_03214_),
    .A1(net4360),
    .A2(_03210_));
 sg13g2_a21oi_1 _25166_ (.A1(net4360),
    .A2(_03213_),
    .Y(_03215_),
    .B1(_03214_));
 sg13g2_a21o_1 _25167_ (.A2(net3977),
    .A1(net2955),
    .B1(_03215_),
    .X(_00401_));
 sg13g2_o21ai_1 _25168_ (.B1(_14620_),
    .Y(_03216_),
    .A1(_14314_),
    .A2(_03186_));
 sg13g2_xnor2_1 _25169_ (.Y(_03217_),
    .A(_14306_),
    .B(_03216_));
 sg13g2_o21ai_1 _25170_ (.B1(_15326_),
    .Y(_03218_),
    .A1(_15443_),
    .A2(_03188_));
 sg13g2_a21o_1 _25171_ (.A2(_03218_),
    .A1(_15447_),
    .B1(_14306_),
    .X(_03219_));
 sg13g2_nand3_1 _25172_ (.B(_15447_),
    .C(_03218_),
    .A(_14306_),
    .Y(_03220_));
 sg13g2_nand3_1 _25173_ (.B(_03219_),
    .C(_03220_),
    .A(net4690),
    .Y(_03221_));
 sg13g2_a21oi_1 _25174_ (.A1(net4577),
    .A2(\u_inv.d_next[126] ),
    .Y(_03222_),
    .B1(net3795));
 sg13g2_a22oi_1 _25175_ (.Y(_03223_),
    .B1(_03221_),
    .B2(_03222_),
    .A2(_03217_),
    .A1(net3795));
 sg13g2_nand2_1 _25176_ (.Y(_03224_),
    .A(net3459),
    .B(_03223_));
 sg13g2_xnor2_1 _25177_ (.Y(_03225_),
    .A(net3484),
    .B(_03223_));
 sg13g2_o21ai_1 _25178_ (.B1(net3448),
    .Y(_03226_),
    .A1(_03193_),
    .A2(_03210_));
 sg13g2_nor2_1 _25179_ (.A(_03195_),
    .B(_03211_),
    .Y(_03227_));
 sg13g2_or2_1 _25180_ (.X(_03228_),
    .B(_03211_),
    .A(_03195_));
 sg13g2_o21ai_1 _25181_ (.B1(_03226_),
    .Y(_03229_),
    .A1(_03199_),
    .A2(_03228_));
 sg13g2_nand2_1 _25182_ (.Y(_03230_),
    .A(_03225_),
    .B(_03229_));
 sg13g2_xnor2_1 _25183_ (.Y(_03231_),
    .A(_03225_),
    .B(_03229_));
 sg13g2_o21ai_1 _25184_ (.B1(net3900),
    .Y(_03232_),
    .A1(net4367),
    .A2(_03223_));
 sg13g2_a21oi_1 _25185_ (.A1(net4367),
    .A2(_03231_),
    .Y(_03233_),
    .B1(_03232_));
 sg13g2_a21o_1 _25186_ (.A2(net3968),
    .A1(net3126),
    .B1(_03233_),
    .X(_00402_));
 sg13g2_nand2_1 _25187_ (.Y(_03234_),
    .A(net2030),
    .B(net3968));
 sg13g2_a21oi_1 _25188_ (.A1(net4577),
    .A2(\u_inv.d_next[127] ),
    .Y(_03235_),
    .B1(net3795));
 sg13g2_a21o_1 _25189_ (.A2(_03219_),
    .A1(_14305_),
    .B1(_14304_),
    .X(_03236_));
 sg13g2_nand3_1 _25190_ (.B(_14305_),
    .C(_03219_),
    .A(_14304_),
    .Y(_03237_));
 sg13g2_nand3_1 _25191_ (.B(_03236_),
    .C(_03237_),
    .A(net4690),
    .Y(_03238_));
 sg13g2_a21oi_1 _25192_ (.A1(_14306_),
    .A2(_03216_),
    .Y(_03239_),
    .B1(_14621_));
 sg13g2_or2_1 _25193_ (.X(_03240_),
    .B(_03239_),
    .A(_14304_));
 sg13g2_a21oi_1 _25194_ (.A1(_14304_),
    .A2(_03239_),
    .Y(_03241_),
    .B1(net3854));
 sg13g2_a22oi_1 _25195_ (.Y(_03242_),
    .B1(_03240_),
    .B2(_03241_),
    .A2(_03238_),
    .A1(_03235_));
 sg13g2_xnor2_1 _25196_ (.Y(_03243_),
    .A(net3485),
    .B(_03242_));
 sg13g2_a21oi_1 _25197_ (.A1(_03224_),
    .A2(_03230_),
    .Y(_03244_),
    .B1(_03243_));
 sg13g2_and3_1 _25198_ (.X(_03245_),
    .A(_03224_),
    .B(_03230_),
    .C(_03243_));
 sg13g2_nor3_1 _25199_ (.A(net4297),
    .B(_03244_),
    .C(_03245_),
    .Y(_03246_));
 sg13g2_o21ai_1 _25200_ (.B1(net3900),
    .Y(_03247_),
    .A1(net4367),
    .A2(_03242_));
 sg13g2_o21ai_1 _25201_ (.B1(_03234_),
    .Y(_00403_),
    .A1(_03246_),
    .A2(_03247_));
 sg13g2_xnor2_1 _25202_ (.Y(_03248_),
    .A(_14658_),
    .B(_14892_));
 sg13g2_a21oi_1 _25203_ (.A1(_14892_),
    .A2(_15629_),
    .Y(_03249_),
    .B1(net4585));
 sg13g2_o21ai_1 _25204_ (.B1(_03249_),
    .Y(_03250_),
    .A1(_14892_),
    .A2(_15629_));
 sg13g2_a21oi_1 _25205_ (.A1(net4585),
    .A2(\u_inv.d_next[128] ),
    .Y(_03251_),
    .B1(net3805));
 sg13g2_a22oi_1 _25206_ (.Y(_03252_),
    .B1(_03250_),
    .B2(_03251_),
    .A2(_03248_),
    .A1(net3805));
 sg13g2_and2_1 _25207_ (.A(net3449),
    .B(_03252_),
    .X(_03253_));
 sg13g2_xnor2_1 _25208_ (.Y(_03254_),
    .A(net3484),
    .B(_03252_));
 sg13g2_nor3_1 _25209_ (.A(_03129_),
    .B(_03149_),
    .C(_03197_),
    .Y(_03255_));
 sg13g2_and4_1 _25210_ (.A(_03225_),
    .B(_03227_),
    .C(_03243_),
    .D(_03255_),
    .X(_03256_));
 sg13g2_and2_1 _25211_ (.A(_03135_),
    .B(_03256_),
    .X(_03257_));
 sg13g2_nand3_1 _25212_ (.B(_03135_),
    .C(_03256_),
    .A(_03003_),
    .Y(_03258_));
 sg13g2_a21o_2 _25213_ (.A2(_02733_),
    .A1(_02728_),
    .B1(_03258_),
    .X(_03259_));
 sg13g2_nand3b_1 _25214_ (.B(_03243_),
    .C(_03225_),
    .Y(_03260_),
    .A_N(_03226_));
 sg13g2_o21ai_1 _25215_ (.B1(net3448),
    .Y(_03261_),
    .A1(_03223_),
    .A2(_03242_));
 sg13g2_o21ai_1 _25216_ (.B1(_03196_),
    .Y(_03262_),
    .A1(_03166_),
    .A2(_03197_));
 sg13g2_nand4_1 _25217_ (.B(_03227_),
    .C(_03243_),
    .A(_03225_),
    .Y(_03263_),
    .D(_03262_));
 sg13g2_nand3_1 _25218_ (.B(_03261_),
    .C(_03263_),
    .A(_03260_),
    .Y(_03264_));
 sg13g2_a221oi_1 _25219_ (.B2(_03002_),
    .C1(_03264_),
    .B1(_03257_),
    .A1(_03134_),
    .Y(_03265_),
    .A2(_03256_));
 sg13g2_nand2_2 _25220_ (.Y(_03266_),
    .A(_03259_),
    .B(_03265_));
 sg13g2_xnor2_1 _25221_ (.Y(_03267_),
    .A(_03254_),
    .B(_03266_));
 sg13g2_a21oi_1 _25222_ (.A1(net4359),
    .A2(_03267_),
    .Y(_03268_),
    .B1(net4238));
 sg13g2_o21ai_1 _25223_ (.B1(_03268_),
    .Y(_03269_),
    .A1(net4359),
    .A2(_03252_));
 sg13g2_o21ai_1 _25224_ (.B1(_03269_),
    .Y(_00404_),
    .A1(_10601_),
    .A2(net4034));
 sg13g2_a21o_1 _25225_ (.A2(_03266_),
    .A1(_03254_),
    .B1(_03253_),
    .X(_03270_));
 sg13g2_o21ai_1 _25226_ (.B1(_14889_),
    .Y(_03271_),
    .A1(_14892_),
    .A2(_15629_));
 sg13g2_a221oi_1 _25227_ (.B2(_15631_),
    .C1(net4585),
    .B1(net3586),
    .A1(_14890_),
    .Y(_03272_),
    .A2(_14891_));
 sg13g2_o21ai_1 _25228_ (.B1(_03272_),
    .Y(_03273_),
    .A1(_14891_),
    .A2(_03271_));
 sg13g2_a21oi_1 _25229_ (.A1(net4585),
    .A2(\u_inv.d_next[129] ),
    .Y(_03274_),
    .B1(net3805));
 sg13g2_a21oi_1 _25230_ (.A1(_14658_),
    .A2(_14892_),
    .Y(_03275_),
    .B1(_14903_));
 sg13g2_or2_1 _25231_ (.X(_03276_),
    .B(_03275_),
    .A(_14889_));
 sg13g2_a21oi_1 _25232_ (.A1(_14889_),
    .A2(_03275_),
    .Y(_03277_),
    .B1(net3859));
 sg13g2_a22oi_1 _25233_ (.Y(_03278_),
    .B1(_03276_),
    .B2(_03277_),
    .A2(_03274_),
    .A1(_03273_));
 sg13g2_nand2b_1 _25234_ (.Y(_03279_),
    .B(net3484),
    .A_N(_03278_));
 sg13g2_nand2_1 _25235_ (.Y(_03280_),
    .A(net3449),
    .B(_03278_));
 sg13g2_inv_1 _25236_ (.Y(_03281_),
    .A(_03280_));
 sg13g2_and2_1 _25237_ (.A(_03279_),
    .B(_03280_),
    .X(_03282_));
 sg13g2_xnor2_1 _25238_ (.Y(_03283_),
    .A(_03270_),
    .B(_03282_));
 sg13g2_o21ai_1 _25239_ (.B1(net3903),
    .Y(_03284_),
    .A1(net4359),
    .A2(_03278_));
 sg13g2_a21oi_1 _25240_ (.A1(net4360),
    .A2(_03283_),
    .Y(_03285_),
    .B1(_03284_));
 sg13g2_a21o_1 _25241_ (.A2(net3976),
    .A1(net2580),
    .B1(_03285_),
    .X(_00405_));
 sg13g2_o21ai_1 _25242_ (.B1(_14893_),
    .Y(_03286_),
    .A1(_14536_),
    .A2(_14657_));
 sg13g2_and2_1 _25243_ (.A(_14904_),
    .B(_03286_),
    .X(_03287_));
 sg13g2_xnor2_1 _25244_ (.Y(_03288_),
    .A(_14884_),
    .B(_03287_));
 sg13g2_a221oi_1 _25245_ (.B2(_15631_),
    .C1(_15270_),
    .B1(net3586),
    .A1(_14890_),
    .Y(_03289_),
    .A2(_14891_));
 sg13g2_a21oi_1 _25246_ (.A1(_14885_),
    .A2(_03289_),
    .Y(_03290_),
    .B1(net4585));
 sg13g2_o21ai_1 _25247_ (.B1(_03290_),
    .Y(_03291_),
    .A1(_14885_),
    .A2(_03289_));
 sg13g2_a21oi_1 _25248_ (.A1(net4585),
    .A2(net4802),
    .Y(_03292_),
    .B1(net3805));
 sg13g2_a22oi_1 _25249_ (.Y(_03293_),
    .B1(_03291_),
    .B2(_03292_),
    .A2(_03288_),
    .A1(net3805));
 sg13g2_nand2_1 _25250_ (.Y(_03294_),
    .A(net3449),
    .B(_03293_));
 sg13g2_xnor2_1 _25251_ (.Y(_03295_),
    .A(net3449),
    .B(_03293_));
 sg13g2_inv_1 _25252_ (.Y(_03296_),
    .A(_03295_));
 sg13g2_nand2b_1 _25253_ (.Y(_03297_),
    .B(_03280_),
    .A_N(_03253_));
 sg13g2_a21oi_1 _25254_ (.A1(_03270_),
    .A2(_03279_),
    .Y(_03298_),
    .B1(_03281_));
 sg13g2_xnor2_1 _25255_ (.Y(_03299_),
    .A(_03295_),
    .B(_03298_));
 sg13g2_o21ai_1 _25256_ (.B1(net3903),
    .Y(_03300_),
    .A1(net4359),
    .A2(_03293_));
 sg13g2_a21oi_1 _25257_ (.A1(net4359),
    .A2(_03299_),
    .Y(_03301_),
    .B1(_03300_));
 sg13g2_a21o_1 _25258_ (.A2(net3976),
    .A1(net2934),
    .B1(_03301_),
    .X(_00406_));
 sg13g2_a21oi_1 _25259_ (.A1(net4585),
    .A2(\u_inv.d_next[131] ),
    .Y(_03302_),
    .B1(net3805));
 sg13g2_o21ai_1 _25260_ (.B1(_14883_),
    .Y(_03303_),
    .A1(_14885_),
    .A2(_03289_));
 sg13g2_o21ai_1 _25261_ (.B1(net4702),
    .Y(_03304_),
    .A1(_14882_),
    .A2(_03303_));
 sg13g2_a21o_1 _25262_ (.A2(_03303_),
    .A1(_14882_),
    .B1(_03304_),
    .X(_03305_));
 sg13g2_o21ai_1 _25263_ (.B1(_14905_),
    .Y(_03306_),
    .A1(_14884_),
    .A2(_03287_));
 sg13g2_or2_1 _25264_ (.X(_03307_),
    .B(_03306_),
    .A(_14882_));
 sg13g2_a21oi_1 _25265_ (.A1(_14882_),
    .A2(_03306_),
    .Y(_03308_),
    .B1(net3859));
 sg13g2_a22oi_1 _25266_ (.Y(_03309_),
    .B1(_03307_),
    .B2(_03308_),
    .A2(_03305_),
    .A1(_03302_));
 sg13g2_nand2_1 _25267_ (.Y(_03310_),
    .A(net3449),
    .B(_03309_));
 sg13g2_xnor2_1 _25268_ (.Y(_03311_),
    .A(net3484),
    .B(_03309_));
 sg13g2_o21ai_1 _25269_ (.B1(_03294_),
    .Y(_03312_),
    .A1(_03295_),
    .A2(_03298_));
 sg13g2_xnor2_1 _25270_ (.Y(_03313_),
    .A(_03311_),
    .B(_03312_));
 sg13g2_o21ai_1 _25271_ (.B1(net3903),
    .Y(_03314_),
    .A1(net4359),
    .A2(_03309_));
 sg13g2_a21oi_1 _25272_ (.A1(net4359),
    .A2(_03313_),
    .Y(_03315_),
    .B1(_03314_));
 sg13g2_a21o_1 _25273_ (.A2(net3976),
    .A1(net4802),
    .B1(_03315_),
    .X(_00407_));
 sg13g2_a21oi_1 _25274_ (.A1(_14904_),
    .A2(_03286_),
    .Y(_03316_),
    .B1(_14886_));
 sg13g2_a21o_1 _25275_ (.A2(_03286_),
    .A1(_14904_),
    .B1(_14886_),
    .X(_03317_));
 sg13g2_o21ai_1 _25276_ (.B1(_14875_),
    .Y(_03318_),
    .A1(_14907_),
    .A2(_03316_));
 sg13g2_nand3b_1 _25277_ (.B(_14906_),
    .C(_03317_),
    .Y(_03319_),
    .A_N(_14875_));
 sg13g2_nand2_1 _25278_ (.Y(_03320_),
    .A(_03318_),
    .B(_03319_));
 sg13g2_a21oi_1 _25279_ (.A1(net3586),
    .A2(_15632_),
    .Y(_03321_),
    .B1(_15273_));
 sg13g2_a21o_1 _25280_ (.A2(_15632_),
    .A1(net3586),
    .B1(_15273_),
    .X(_03322_));
 sg13g2_a21oi_1 _25281_ (.A1(_14875_),
    .A2(_03321_),
    .Y(_03323_),
    .B1(net4584));
 sg13g2_o21ai_1 _25282_ (.B1(_03323_),
    .Y(_03324_),
    .A1(_14875_),
    .A2(_03321_));
 sg13g2_a21oi_1 _25283_ (.A1(net4584),
    .A2(\u_inv.d_next[132] ),
    .Y(_03325_),
    .B1(net3804));
 sg13g2_a22oi_1 _25284_ (.Y(_03326_),
    .B1(_03324_),
    .B2(_03325_),
    .A2(_03320_),
    .A1(net3804));
 sg13g2_and2_1 _25285_ (.A(net3450),
    .B(_03326_),
    .X(_03327_));
 sg13g2_xnor2_1 _25286_ (.Y(_03328_),
    .A(net3450),
    .B(_03326_));
 sg13g2_nand3_1 _25287_ (.B(_03297_),
    .C(_03311_),
    .A(_03296_),
    .Y(_03329_));
 sg13g2_and3_1 _25288_ (.X(_03330_),
    .A(_03294_),
    .B(_03310_),
    .C(_03329_));
 sg13g2_nand3_1 _25289_ (.B(_03310_),
    .C(_03329_),
    .A(_03294_),
    .Y(_03331_));
 sg13g2_nand4_1 _25290_ (.B(_03282_),
    .C(_03296_),
    .A(_03254_),
    .Y(_03332_),
    .D(_03311_));
 sg13g2_nand2b_1 _25291_ (.Y(_03333_),
    .B(_03266_),
    .A_N(_03332_));
 sg13g2_nand2_1 _25292_ (.Y(_03334_),
    .A(_03330_),
    .B(_03333_));
 sg13g2_a21oi_1 _25293_ (.A1(_03330_),
    .A2(_03333_),
    .Y(_03335_),
    .B1(_03328_));
 sg13g2_xor2_1 _25294_ (.B(_03334_),
    .A(_03328_),
    .X(_03336_));
 sg13g2_o21ai_1 _25295_ (.B1(net3903),
    .Y(_03337_),
    .A1(net4362),
    .A2(_03326_));
 sg13g2_a21oi_1 _25296_ (.A1(net4361),
    .A2(_03336_),
    .Y(_03338_),
    .B1(_03337_));
 sg13g2_a21o_1 _25297_ (.A2(net3976),
    .A1(net3274),
    .B1(_03338_),
    .X(_00408_));
 sg13g2_a21oi_1 _25298_ (.A1(net4584),
    .A2(\u_inv.d_next[133] ),
    .Y(_03339_),
    .B1(net3804));
 sg13g2_o21ai_1 _25299_ (.B1(_14874_),
    .Y(_03340_),
    .A1(_14875_),
    .A2(_03321_));
 sg13g2_xnor2_1 _25300_ (.Y(_03341_),
    .A(_14872_),
    .B(_03340_));
 sg13g2_o21ai_1 _25301_ (.B1(_03339_),
    .Y(_03342_),
    .A1(net4586),
    .A2(_03341_));
 sg13g2_nand3_1 _25302_ (.B(_14912_),
    .C(_03318_),
    .A(_14873_),
    .Y(_03343_));
 sg13g2_a21o_1 _25303_ (.A2(_03318_),
    .A1(_14912_),
    .B1(_14873_),
    .X(_03344_));
 sg13g2_nand3_1 _25304_ (.B(_03343_),
    .C(_03344_),
    .A(net3804),
    .Y(_03345_));
 sg13g2_and3_1 _25305_ (.X(_03346_),
    .A(net3450),
    .B(_03342_),
    .C(_03345_));
 sg13g2_a21oi_1 _25306_ (.A1(_03342_),
    .A2(_03345_),
    .Y(_03347_),
    .B1(net3450));
 sg13g2_nor2_1 _25307_ (.A(_03346_),
    .B(_03347_),
    .Y(_03348_));
 sg13g2_nor2_1 _25308_ (.A(_03327_),
    .B(_03335_),
    .Y(_03349_));
 sg13g2_a21oi_1 _25309_ (.A1(_03348_),
    .A2(_03349_),
    .Y(_03350_),
    .B1(net4298));
 sg13g2_o21ai_1 _25310_ (.B1(_03350_),
    .Y(_03351_),
    .A1(_03348_),
    .A2(_03349_));
 sg13g2_a21oi_1 _25311_ (.A1(_03342_),
    .A2(_03345_),
    .Y(_03352_),
    .B1(net4361));
 sg13g2_nor2_1 _25312_ (.A(net4238),
    .B(_03352_),
    .Y(_03353_));
 sg13g2_a22oi_1 _25313_ (.Y(_03354_),
    .B1(_03351_),
    .B2(_03353_),
    .A2(net3976),
    .A1(net2825));
 sg13g2_inv_1 _25314_ (.Y(_00409_),
    .A(_03354_));
 sg13g2_a21oi_1 _25315_ (.A1(_14906_),
    .A2(_03317_),
    .Y(_03355_),
    .B1(_14877_));
 sg13g2_o21ai_1 _25316_ (.B1(_14868_),
    .Y(_03356_),
    .A1(_14913_),
    .A2(_03355_));
 sg13g2_or3_1 _25317_ (.A(_14868_),
    .B(_14913_),
    .C(_03355_),
    .X(_03357_));
 sg13g2_nand2_1 _25318_ (.Y(_03358_),
    .A(_03356_),
    .B(_03357_));
 sg13g2_a21oi_1 _25319_ (.A1(_15267_),
    .A2(_03322_),
    .Y(_03359_),
    .B1(_15274_));
 sg13g2_nor2_1 _25320_ (.A(_14868_),
    .B(_03359_),
    .Y(_03360_));
 sg13g2_a21oi_1 _25321_ (.A1(_14868_),
    .A2(_03359_),
    .Y(_03361_),
    .B1(net4586));
 sg13g2_nand2b_1 _25322_ (.Y(_03362_),
    .B(_03361_),
    .A_N(_03360_));
 sg13g2_a21oi_1 _25323_ (.A1(net4584),
    .A2(\u_inv.d_next[134] ),
    .Y(_03363_),
    .B1(net3806));
 sg13g2_a22oi_1 _25324_ (.Y(_03364_),
    .B1(_03362_),
    .B2(_03363_),
    .A2(_03358_),
    .A1(net3806));
 sg13g2_nand2_1 _25325_ (.Y(_03365_),
    .A(net3450),
    .B(_03364_));
 sg13g2_xnor2_1 _25326_ (.Y(_03366_),
    .A(net3450),
    .B(_03364_));
 sg13g2_or2_1 _25327_ (.X(_03367_),
    .B(_03346_),
    .A(_03327_));
 sg13g2_nor2_1 _25328_ (.A(_03347_),
    .B(_03349_),
    .Y(_03368_));
 sg13g2_or3_1 _25329_ (.A(_03328_),
    .B(_03346_),
    .C(_03347_),
    .X(_03369_));
 sg13g2_nor2_1 _25330_ (.A(_03346_),
    .B(_03368_),
    .Y(_03370_));
 sg13g2_xnor2_1 _25331_ (.Y(_03371_),
    .A(_03366_),
    .B(_03370_));
 sg13g2_o21ai_1 _25332_ (.B1(net3903),
    .Y(_03372_),
    .A1(net4361),
    .A2(_03364_));
 sg13g2_a21oi_1 _25333_ (.A1(net4361),
    .A2(_03371_),
    .Y(_03373_),
    .B1(_03372_));
 sg13g2_a21o_1 _25334_ (.A2(net3976),
    .A1(net2909),
    .B1(_03373_),
    .X(_00410_));
 sg13g2_a21oi_1 _25335_ (.A1(net4584),
    .A2(\u_inv.d_next[135] ),
    .Y(_03374_),
    .B1(net3804));
 sg13g2_nor2_1 _25336_ (.A(_14866_),
    .B(_03360_),
    .Y(_03375_));
 sg13g2_xnor2_1 _25337_ (.Y(_03376_),
    .A(_14864_),
    .B(_03375_));
 sg13g2_o21ai_1 _25338_ (.B1(_03374_),
    .Y(_03377_),
    .A1(net4584),
    .A2(_03376_));
 sg13g2_a21o_1 _25339_ (.A2(_03356_),
    .A1(_14909_),
    .B1(_14864_),
    .X(_03378_));
 sg13g2_nand3_1 _25340_ (.B(_14909_),
    .C(_03356_),
    .A(_14864_),
    .Y(_03379_));
 sg13g2_nand3_1 _25341_ (.B(_03378_),
    .C(_03379_),
    .A(net3805),
    .Y(_03380_));
 sg13g2_nand2_1 _25342_ (.Y(_03381_),
    .A(_03377_),
    .B(_03380_));
 sg13g2_and3_1 _25343_ (.X(_03382_),
    .A(net3451),
    .B(_03377_),
    .C(_03380_));
 sg13g2_a21oi_1 _25344_ (.A1(_03377_),
    .A2(_03380_),
    .Y(_03383_),
    .B1(net3451));
 sg13g2_nor2_1 _25345_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sg13g2_o21ai_1 _25346_ (.B1(_03365_),
    .Y(_03385_),
    .A1(_03366_),
    .A2(_03370_));
 sg13g2_xor2_1 _25347_ (.B(_03385_),
    .A(_03384_),
    .X(_03386_));
 sg13g2_a21oi_1 _25348_ (.A1(net4298),
    .A2(_03381_),
    .Y(_03387_),
    .B1(net4238));
 sg13g2_o21ai_1 _25349_ (.B1(_03387_),
    .Y(_03388_),
    .A1(net4298),
    .A2(_03386_));
 sg13g2_o21ai_1 _25350_ (.B1(_03388_),
    .Y(_00411_),
    .A1(_10600_),
    .A2(net4038));
 sg13g2_o21ai_1 _25351_ (.B1(_14895_),
    .Y(_03389_),
    .A1(_14536_),
    .A2(_14657_));
 sg13g2_a21oi_1 _25352_ (.A1(_14914_),
    .A2(_03389_),
    .Y(_03390_),
    .B1(_14858_));
 sg13g2_nand3_1 _25353_ (.B(_14914_),
    .C(_03389_),
    .A(_14858_),
    .Y(_03391_));
 sg13g2_nand2b_1 _25354_ (.Y(_03392_),
    .B(_03391_),
    .A_N(_03390_));
 sg13g2_o21ai_1 _25355_ (.B1(_15277_),
    .Y(_03393_),
    .A1(_15629_),
    .A2(_15633_));
 sg13g2_o21ai_1 _25356_ (.B1(net4702),
    .Y(_03394_),
    .A1(_14858_),
    .A2(_03393_));
 sg13g2_a21o_1 _25357_ (.A2(_03393_),
    .A1(_14858_),
    .B1(_03394_),
    .X(_03395_));
 sg13g2_a21oi_1 _25358_ (.A1(net4584),
    .A2(\u_inv.d_next[136] ),
    .Y(_03396_),
    .B1(net3804));
 sg13g2_a22oi_1 _25359_ (.Y(_03397_),
    .B1(_03395_),
    .B2(_03396_),
    .A2(_03392_),
    .A1(net3804));
 sg13g2_nand2_1 _25360_ (.Y(_03398_),
    .A(net3451),
    .B(_03397_));
 sg13g2_xnor2_1 _25361_ (.Y(_03399_),
    .A(net3450),
    .B(_03397_));
 sg13g2_nor3_1 _25362_ (.A(_03366_),
    .B(_03382_),
    .C(_03383_),
    .Y(_03400_));
 sg13g2_nor4_1 _25363_ (.A(_03366_),
    .B(_03369_),
    .C(_03382_),
    .D(_03383_),
    .Y(_03401_));
 sg13g2_and2_1 _25364_ (.A(_03331_),
    .B(_03401_),
    .X(_03402_));
 sg13g2_o21ai_1 _25365_ (.B1(_03365_),
    .Y(_03403_),
    .A1(net3484),
    .A2(_03381_));
 sg13g2_a21o_1 _25366_ (.A2(_03400_),
    .A1(_03367_),
    .B1(_03403_),
    .X(_03404_));
 sg13g2_nor2b_1 _25367_ (.A(_03332_),
    .B_N(_03401_),
    .Y(_03405_));
 sg13g2_a221oi_1 _25368_ (.B2(_03266_),
    .C1(_03404_),
    .B1(_03405_),
    .A1(_03331_),
    .Y(_03406_),
    .A2(_03401_));
 sg13g2_xnor2_1 _25369_ (.Y(_03407_),
    .A(_03399_),
    .B(_03406_));
 sg13g2_o21ai_1 _25370_ (.B1(net3903),
    .Y(_03408_),
    .A1(net4361),
    .A2(_03397_));
 sg13g2_a21oi_1 _25371_ (.A1(net4361),
    .A2(_03407_),
    .Y(_03409_),
    .B1(_03408_));
 sg13g2_a21o_1 _25372_ (.A2(net3976),
    .A1(net3090),
    .B1(_03409_),
    .X(_00412_));
 sg13g2_nand2_1 _25373_ (.Y(_03410_),
    .A(net2565),
    .B(net3977));
 sg13g2_o21ai_1 _25374_ (.B1(_03398_),
    .Y(_03411_),
    .A1(_03399_),
    .A2(_03406_));
 sg13g2_a21oi_1 _25375_ (.A1(net4584),
    .A2(\u_inv.d_next[137] ),
    .Y(_03412_),
    .B1(net3804));
 sg13g2_a21oi_1 _25376_ (.A1(_14858_),
    .A2(_03393_),
    .Y(_03413_),
    .B1(_14857_));
 sg13g2_o21ai_1 _25377_ (.B1(net4702),
    .Y(_03414_),
    .A1(_14856_),
    .A2(_03413_));
 sg13g2_a21o_1 _25378_ (.A2(_03413_),
    .A1(_14856_),
    .B1(_03414_),
    .X(_03415_));
 sg13g2_o21ai_1 _25379_ (.B1(_14855_),
    .Y(_03416_),
    .A1(_14923_),
    .A2(_03390_));
 sg13g2_nor3_1 _25380_ (.A(_14855_),
    .B(_14923_),
    .C(_03390_),
    .Y(_03417_));
 sg13g2_nor2_1 _25381_ (.A(net3859),
    .B(_03417_),
    .Y(_03418_));
 sg13g2_a22oi_1 _25382_ (.Y(_03419_),
    .B1(_03416_),
    .B2(_03418_),
    .A2(_03415_),
    .A1(_03412_));
 sg13g2_nand2_1 _25383_ (.Y(_03420_),
    .A(net3451),
    .B(_03419_));
 sg13g2_xnor2_1 _25384_ (.Y(_03421_),
    .A(net3450),
    .B(_03419_));
 sg13g2_o21ai_1 _25385_ (.B1(net4361),
    .Y(_03422_),
    .A1(_03411_),
    .A2(_03421_));
 sg13g2_a21oi_1 _25386_ (.A1(_03411_),
    .A2(_03421_),
    .Y(_03423_),
    .B1(_03422_));
 sg13g2_o21ai_1 _25387_ (.B1(net3904),
    .Y(_03424_),
    .A1(net4361),
    .A2(_03419_));
 sg13g2_o21ai_1 _25388_ (.B1(_03410_),
    .Y(_00413_),
    .A1(_03423_),
    .A2(_03424_));
 sg13g2_a21oi_1 _25389_ (.A1(_14914_),
    .A2(_03389_),
    .Y(_03425_),
    .B1(_14860_));
 sg13g2_a21o_1 _25390_ (.A2(_03389_),
    .A1(_14914_),
    .B1(_14860_),
    .X(_03426_));
 sg13g2_a21oi_1 _25391_ (.A1(_14924_),
    .A2(_03426_),
    .Y(_03427_),
    .B1(_14850_));
 sg13g2_nand3_1 _25392_ (.B(_14924_),
    .C(_03426_),
    .A(_14850_),
    .Y(_03428_));
 sg13g2_nand2b_1 _25393_ (.Y(_03429_),
    .B(_03428_),
    .A_N(_03427_));
 sg13g2_a221oi_1 _25394_ (.B2(_03393_),
    .C1(_14854_),
    .B1(_15264_),
    .A1(_14853_),
    .Y(_03430_),
    .A2(_14857_));
 sg13g2_a21oi_1 _25395_ (.A1(_14849_),
    .A2(_03430_),
    .Y(_03431_),
    .B1(net4587));
 sg13g2_o21ai_1 _25396_ (.B1(_03431_),
    .Y(_03432_),
    .A1(_14849_),
    .A2(_03430_));
 sg13g2_a21oi_1 _25397_ (.A1(net4587),
    .A2(\u_inv.d_next[138] ),
    .Y(_03433_),
    .B1(net3809));
 sg13g2_a22oi_1 _25398_ (.Y(_03434_),
    .B1(_03432_),
    .B2(_03433_),
    .A2(_03429_),
    .A1(net3809));
 sg13g2_nand2_1 _25399_ (.Y(_03435_),
    .A(net3451),
    .B(_03434_));
 sg13g2_xnor2_1 _25400_ (.Y(_03436_),
    .A(net3451),
    .B(_03434_));
 sg13g2_nand2_1 _25401_ (.Y(_03437_),
    .A(_03398_),
    .B(_03420_));
 sg13g2_nor2_1 _25402_ (.A(_03399_),
    .B(_03421_),
    .Y(_03438_));
 sg13g2_nor2b_1 _25403_ (.A(_03406_),
    .B_N(_03438_),
    .Y(_03439_));
 sg13g2_or2_1 _25404_ (.X(_03440_),
    .B(_03439_),
    .A(_03437_));
 sg13g2_nand2b_1 _25405_ (.Y(_03441_),
    .B(_03440_),
    .A_N(_03436_));
 sg13g2_xor2_1 _25406_ (.B(_03440_),
    .A(_03436_),
    .X(_03442_));
 sg13g2_o21ai_1 _25407_ (.B1(net3903),
    .Y(_03443_),
    .A1(net4362),
    .A2(_03434_));
 sg13g2_a21oi_1 _25408_ (.A1(net4362),
    .A2(_03442_),
    .Y(_03444_),
    .B1(_03443_));
 sg13g2_a21o_1 _25409_ (.A2(net3976),
    .A1(net3292),
    .B1(_03444_),
    .X(_00414_));
 sg13g2_nand2_1 _25410_ (.Y(_03445_),
    .A(_03435_),
    .B(_03441_));
 sg13g2_nand2b_1 _25411_ (.Y(_03446_),
    .B(net3859),
    .A_N(\u_inv.d_next[139] ));
 sg13g2_o21ai_1 _25412_ (.B1(_14848_),
    .Y(_03447_),
    .A1(_14849_),
    .A2(_03430_));
 sg13g2_xnor2_1 _25413_ (.Y(_03448_),
    .A(_14846_),
    .B(_03447_));
 sg13g2_a22oi_1 _25414_ (.Y(_03449_),
    .B1(_03448_),
    .B2(net4700),
    .A2(_03446_),
    .A1(net3735));
 sg13g2_o21ai_1 _25415_ (.B1(_14847_),
    .Y(_03450_),
    .A1(_14925_),
    .A2(_03427_));
 sg13g2_nor3_1 _25416_ (.A(_14847_),
    .B(_14925_),
    .C(_03427_),
    .Y(_03451_));
 sg13g2_nor2_1 _25417_ (.A(net3859),
    .B(_03451_),
    .Y(_03452_));
 sg13g2_a21oi_1 _25418_ (.A1(_03450_),
    .A2(_03452_),
    .Y(_03453_),
    .B1(_03449_));
 sg13g2_a21o_1 _25419_ (.A2(_03452_),
    .A1(_03450_),
    .B1(_03449_),
    .X(_03454_));
 sg13g2_xnor2_1 _25420_ (.Y(_03455_),
    .A(net3486),
    .B(_03453_));
 sg13g2_xnor2_1 _25421_ (.Y(_03456_),
    .A(_03445_),
    .B(_03455_));
 sg13g2_o21ai_1 _25422_ (.B1(net3903),
    .Y(_03457_),
    .A1(net4362),
    .A2(_03453_));
 sg13g2_a21oi_1 _25423_ (.A1(net4362),
    .A2(_03456_),
    .Y(_03458_),
    .B1(_03457_));
 sg13g2_a21o_1 _25424_ (.A2(net3978),
    .A1(net3291),
    .B1(_03458_),
    .X(_00415_));
 sg13g2_a21o_2 _25425_ (.A2(_03425_),
    .A1(_14851_),
    .B1(_14927_),
    .X(_03459_));
 sg13g2_xnor2_1 _25426_ (.Y(_03460_),
    .A(net4429),
    .B(_03459_));
 sg13g2_a21oi_1 _25427_ (.A1(_15265_),
    .A2(_03393_),
    .Y(_03461_),
    .B1(_15280_));
 sg13g2_a21o_1 _25428_ (.A2(_03393_),
    .A1(_15265_),
    .B1(_15280_),
    .X(_03462_));
 sg13g2_a21oi_1 _25429_ (.A1(net4429),
    .A2(_03461_),
    .Y(_03463_),
    .B1(net4587));
 sg13g2_o21ai_1 _25430_ (.B1(_03463_),
    .Y(_03464_),
    .A1(net4429),
    .A2(_03461_));
 sg13g2_a21oi_1 _25431_ (.A1(net4587),
    .A2(\u_inv.d_next[140] ),
    .Y(_03465_),
    .B1(net3807));
 sg13g2_a22oi_1 _25432_ (.Y(_03466_),
    .B1(_03464_),
    .B2(_03465_),
    .A2(_03460_),
    .A1(net3807));
 sg13g2_xnor2_1 _25433_ (.Y(_03467_),
    .A(net3460),
    .B(_03466_));
 sg13g2_o21ai_1 _25434_ (.B1(_03435_),
    .Y(_03468_),
    .A1(net3486),
    .A2(_03454_));
 sg13g2_nor2b_1 _25435_ (.A(_03436_),
    .B_N(_03455_),
    .Y(_03469_));
 sg13g2_a21o_1 _25436_ (.A2(_03469_),
    .A1(_03440_),
    .B1(_03468_),
    .X(_03470_));
 sg13g2_nor2b_1 _25437_ (.A(_03467_),
    .B_N(_03470_),
    .Y(_03471_));
 sg13g2_xor2_1 _25438_ (.B(_03470_),
    .A(_03467_),
    .X(_03472_));
 sg13g2_o21ai_1 _25439_ (.B1(net3905),
    .Y(_03473_),
    .A1(net4371),
    .A2(_03466_));
 sg13g2_a21oi_1 _25440_ (.A1(net4371),
    .A2(_03472_),
    .Y(_03474_),
    .B1(_03473_));
 sg13g2_a21o_1 _25441_ (.A2(net3978),
    .A1(net3207),
    .B1(_03474_),
    .X(_00416_));
 sg13g2_a21oi_1 _25442_ (.A1(net4588),
    .A2(\u_inv.d_next[141] ),
    .Y(_03475_),
    .B1(net3807));
 sg13g2_o21ai_1 _25443_ (.B1(_14839_),
    .Y(_03476_),
    .A1(net4429),
    .A2(_03461_));
 sg13g2_xnor2_1 _25444_ (.Y(_03477_),
    .A(net4430),
    .B(_03476_));
 sg13g2_nand2_1 _25445_ (.Y(_03478_),
    .A(net4700),
    .B(_03477_));
 sg13g2_a21oi_1 _25446_ (.A1(net4429),
    .A2(_03459_),
    .Y(_03479_),
    .B1(_14916_));
 sg13g2_or2_1 _25447_ (.X(_03480_),
    .B(_03479_),
    .A(net4430));
 sg13g2_a21oi_1 _25448_ (.A1(net4430),
    .A2(_03479_),
    .Y(_03481_),
    .B1(net3859));
 sg13g2_a22oi_1 _25449_ (.Y(_03482_),
    .B1(_03480_),
    .B2(_03481_),
    .A2(_03478_),
    .A1(_03475_));
 sg13g2_and2_1 _25450_ (.A(net3460),
    .B(_03482_),
    .X(_03483_));
 sg13g2_nand2b_1 _25451_ (.Y(_03484_),
    .B(net3487),
    .A_N(_03482_));
 sg13g2_xnor2_1 _25452_ (.Y(_03485_),
    .A(net3460),
    .B(_03482_));
 sg13g2_a21o_1 _25453_ (.A2(_03466_),
    .A1(net3460),
    .B1(_03471_),
    .X(_03486_));
 sg13g2_xor2_1 _25454_ (.B(_03486_),
    .A(_03485_),
    .X(_03487_));
 sg13g2_o21ai_1 _25455_ (.B1(net3905),
    .Y(_03488_),
    .A1(net4371),
    .A2(_03482_));
 sg13g2_a21oi_1 _25456_ (.A1(net4371),
    .A2(_03487_),
    .Y(_03489_),
    .B1(_03488_));
 sg13g2_a21o_1 _25457_ (.A2(net3978),
    .A1(net2852),
    .B1(_03489_),
    .X(_00417_));
 sg13g2_a221oi_1 _25458_ (.B2(_14841_),
    .C1(_14915_),
    .B1(_03459_),
    .A1(net4430),
    .Y(_03490_),
    .A2(_14916_));
 sg13g2_xnor2_1 _25459_ (.Y(_03491_),
    .A(_14835_),
    .B(_03490_));
 sg13g2_a21oi_1 _25460_ (.A1(_15261_),
    .A2(_03462_),
    .Y(_03492_),
    .B1(_15282_));
 sg13g2_a21oi_1 _25461_ (.A1(_14834_),
    .A2(_03492_),
    .Y(_03493_),
    .B1(net4588));
 sg13g2_o21ai_1 _25462_ (.B1(_03493_),
    .Y(_03494_),
    .A1(_14834_),
    .A2(_03492_));
 sg13g2_a21oi_1 _25463_ (.A1(net4588),
    .A2(\u_inv.d_next[142] ),
    .Y(_03495_),
    .B1(net3807));
 sg13g2_a22oi_1 _25464_ (.Y(_03496_),
    .B1(_03494_),
    .B2(_03495_),
    .A2(_03491_),
    .A1(net3807));
 sg13g2_nand2_1 _25465_ (.Y(_03497_),
    .A(net3460),
    .B(_03496_));
 sg13g2_xnor2_1 _25466_ (.Y(_03498_),
    .A(net3460),
    .B(_03496_));
 sg13g2_a21o_1 _25467_ (.A2(_03466_),
    .A1(net3460),
    .B1(_03483_),
    .X(_03499_));
 sg13g2_o21ai_1 _25468_ (.B1(_03484_),
    .Y(_03500_),
    .A1(_03471_),
    .A2(_03499_));
 sg13g2_xnor2_1 _25469_ (.Y(_03501_),
    .A(_03498_),
    .B(_03500_));
 sg13g2_o21ai_1 _25470_ (.B1(net3905),
    .Y(_03502_),
    .A1(net4371),
    .A2(_03496_));
 sg13g2_a21oi_1 _25471_ (.A1(net4371),
    .A2(_03501_),
    .Y(_03503_),
    .B1(_03502_));
 sg13g2_a21o_1 _25472_ (.A2(net3978),
    .A1(net2899),
    .B1(_03503_),
    .X(_00418_));
 sg13g2_a21oi_1 _25473_ (.A1(net4587),
    .A2(\u_inv.d_next[143] ),
    .Y(_03504_),
    .B1(net3807));
 sg13g2_o21ai_1 _25474_ (.B1(_14833_),
    .Y(_03505_),
    .A1(_14834_),
    .A2(_03492_));
 sg13g2_o21ai_1 _25475_ (.B1(net4700),
    .Y(_03506_),
    .A1(_14832_),
    .A2(_03505_));
 sg13g2_a21o_1 _25476_ (.A2(_03505_),
    .A1(_14832_),
    .B1(_03506_),
    .X(_03507_));
 sg13g2_o21ai_1 _25477_ (.B1(_14919_),
    .Y(_03508_),
    .A1(_14835_),
    .A2(_03490_));
 sg13g2_or2_1 _25478_ (.X(_03509_),
    .B(_03508_),
    .A(_14832_));
 sg13g2_a21oi_1 _25479_ (.A1(_14832_),
    .A2(_03508_),
    .Y(_03510_),
    .B1(net3859));
 sg13g2_a22oi_1 _25480_ (.Y(_03511_),
    .B1(_03509_),
    .B2(_03510_),
    .A2(_03507_),
    .A1(_03504_));
 sg13g2_nand2_1 _25481_ (.Y(_03512_),
    .A(net3461),
    .B(_03511_));
 sg13g2_xnor2_1 _25482_ (.Y(_03513_),
    .A(net3487),
    .B(_03511_));
 sg13g2_xnor2_1 _25483_ (.Y(_03514_),
    .A(net3460),
    .B(_03511_));
 sg13g2_o21ai_1 _25484_ (.B1(_03497_),
    .Y(_03515_),
    .A1(_03498_),
    .A2(_03500_));
 sg13g2_xnor2_1 _25485_ (.Y(_03516_),
    .A(_03513_),
    .B(_03515_));
 sg13g2_o21ai_1 _25486_ (.B1(net3905),
    .Y(_03517_),
    .A1(net4371),
    .A2(_03511_));
 sg13g2_a21oi_1 _25487_ (.A1(net4371),
    .A2(_03516_),
    .Y(_03518_),
    .B1(_03517_));
 sg13g2_a21o_1 _25488_ (.A2(net3978),
    .A1(net2641),
    .B1(_03518_),
    .X(_00419_));
 sg13g2_a21oi_2 _25489_ (.B1(_14897_),
    .Y(_03519_),
    .A2(_14656_),
    .A1(_14537_));
 sg13g2_nor2_1 _25490_ (.A(_14929_),
    .B(_03519_),
    .Y(_03520_));
 sg13g2_nor2_1 _25491_ (.A(_14824_),
    .B(_03520_),
    .Y(_03521_));
 sg13g2_xnor2_1 _25492_ (.Y(_03522_),
    .A(_14824_),
    .B(_03520_));
 sg13g2_a21oi_2 _25493_ (.B1(_15286_),
    .Y(_03523_),
    .A2(_15634_),
    .A1(net3586));
 sg13g2_a21oi_1 _25494_ (.A1(_14823_),
    .A2(_03523_),
    .Y(_03524_),
    .B1(net4594));
 sg13g2_o21ai_1 _25495_ (.B1(_03524_),
    .Y(_03525_),
    .A1(_14823_),
    .A2(_03523_));
 sg13g2_a21oi_1 _25496_ (.A1(net4594),
    .A2(\u_inv.d_next[144] ),
    .Y(_03526_),
    .B1(net3816));
 sg13g2_a22oi_1 _25497_ (.Y(_03527_),
    .B1(_03525_),
    .B2(_03526_),
    .A2(_03522_),
    .A1(net3816));
 sg13g2_nand2_1 _25498_ (.Y(_03528_),
    .A(net3462),
    .B(_03527_));
 sg13g2_xnor2_1 _25499_ (.Y(_03529_),
    .A(net3462),
    .B(_03527_));
 sg13g2_or2_1 _25500_ (.X(_03530_),
    .B(_03485_),
    .A(_03467_));
 sg13g2_nand3b_1 _25501_ (.B(_03438_),
    .C(_03455_),
    .Y(_03531_),
    .A_N(_03436_));
 sg13g2_nor4_2 _25502_ (.A(_03498_),
    .B(_03514_),
    .C(_03530_),
    .Y(_03532_),
    .D(_03531_));
 sg13g2_o21ai_1 _25503_ (.B1(_03532_),
    .Y(_03533_),
    .A1(_03402_),
    .A2(_03404_));
 sg13g2_nand3b_1 _25504_ (.B(_03499_),
    .C(_03513_),
    .Y(_03534_),
    .A_N(_03498_));
 sg13g2_and3_1 _25505_ (.X(_03535_),
    .A(_03497_),
    .B(_03512_),
    .C(_03534_));
 sg13g2_a21oi_1 _25506_ (.A1(_03437_),
    .A2(_03469_),
    .Y(_03536_),
    .B1(_03468_));
 sg13g2_or4_1 _25507_ (.A(_03498_),
    .B(_03514_),
    .C(_03530_),
    .D(_03536_),
    .X(_03537_));
 sg13g2_and3_2 _25508_ (.X(_03538_),
    .A(_03533_),
    .B(_03535_),
    .C(_03537_));
 sg13g2_nand3_1 _25509_ (.B(_03535_),
    .C(_03537_),
    .A(_03533_),
    .Y(_03539_));
 sg13g2_nand2_2 _25510_ (.Y(_03540_),
    .A(_03405_),
    .B(_03532_));
 sg13g2_a21o_2 _25511_ (.A2(_03265_),
    .A1(_03259_),
    .B1(_03540_),
    .X(_03541_));
 sg13g2_a21oi_2 _25512_ (.B1(_03529_),
    .Y(_03542_),
    .A2(_03541_),
    .A1(_03538_));
 sg13g2_nand3_1 _25513_ (.B(_03538_),
    .C(_03541_),
    .A(_03529_),
    .Y(_03543_));
 sg13g2_nor2b_1 _25514_ (.A(_03542_),
    .B_N(_03543_),
    .Y(_03544_));
 sg13g2_nor2_1 _25515_ (.A(net4373),
    .B(_03527_),
    .Y(_03545_));
 sg13g2_o21ai_1 _25516_ (.B1(net3909),
    .Y(_03546_),
    .A1(net4298),
    .A2(_03544_));
 sg13g2_nand2_1 _25517_ (.Y(_03547_),
    .A(net2567),
    .B(net3985));
 sg13g2_o21ai_1 _25518_ (.B1(_03547_),
    .Y(_00420_),
    .A1(_03545_),
    .A2(_03546_));
 sg13g2_nand2_1 _25519_ (.Y(_03548_),
    .A(net2150),
    .B(net3985));
 sg13g2_a21o_1 _25520_ (.A2(_03527_),
    .A1(net3462),
    .B1(_03542_),
    .X(_03549_));
 sg13g2_nand2b_1 _25521_ (.Y(_03550_),
    .B(_15256_),
    .A_N(_03523_));
 sg13g2_and2_1 _25522_ (.A(_14821_),
    .B(_14822_),
    .X(_03551_));
 sg13g2_o21ai_1 _25523_ (.B1(_03551_),
    .Y(_03552_),
    .A1(_14823_),
    .A2(_03523_));
 sg13g2_nor2b_1 _25524_ (.A(_15244_),
    .B_N(_03552_),
    .Y(_03553_));
 sg13g2_nand3_1 _25525_ (.B(_03550_),
    .C(_03553_),
    .A(net4713),
    .Y(_03554_));
 sg13g2_a21oi_1 _25526_ (.A1(net4595),
    .A2(\u_inv.d_next[145] ),
    .Y(_03555_),
    .B1(net3816));
 sg13g2_or2_1 _25527_ (.X(_03556_),
    .B(_03521_),
    .A(_14931_));
 sg13g2_xnor2_1 _25528_ (.Y(_03557_),
    .A(_14821_),
    .B(_03556_));
 sg13g2_a22oi_1 _25529_ (.Y(_03558_),
    .B1(_03557_),
    .B2(net3816),
    .A2(_03555_),
    .A1(_03554_));
 sg13g2_nand2_1 _25530_ (.Y(_03559_),
    .A(net3462),
    .B(_03558_));
 sg13g2_xnor2_1 _25531_ (.Y(_03560_),
    .A(net3462),
    .B(_03558_));
 sg13g2_inv_1 _25532_ (.Y(_03561_),
    .A(_03560_));
 sg13g2_o21ai_1 _25533_ (.B1(net4373),
    .Y(_03562_),
    .A1(_03549_),
    .A2(_03560_));
 sg13g2_a21oi_1 _25534_ (.A1(_03549_),
    .A2(_03560_),
    .Y(_03563_),
    .B1(_03562_));
 sg13g2_o21ai_1 _25535_ (.B1(net3909),
    .Y(_03564_),
    .A1(net4373),
    .A2(_03558_));
 sg13g2_o21ai_1 _25536_ (.B1(_03548_),
    .Y(_00421_),
    .A1(_03563_),
    .A2(_03564_));
 sg13g2_o21ai_1 _25537_ (.B1(_14825_),
    .Y(_03565_),
    .A1(_14929_),
    .A2(_03519_));
 sg13g2_a21oi_1 _25538_ (.A1(_14932_),
    .A2(_03565_),
    .Y(_03566_),
    .B1(_14817_));
 sg13g2_nand3_1 _25539_ (.B(_14932_),
    .C(_03565_),
    .A(_14817_),
    .Y(_03567_));
 sg13g2_nand2b_1 _25540_ (.Y(_03568_),
    .B(_03567_),
    .A_N(_03566_));
 sg13g2_a21oi_1 _25541_ (.A1(_15245_),
    .A2(_03550_),
    .Y(_03569_),
    .B1(_14816_));
 sg13g2_nand3_1 _25542_ (.B(_15245_),
    .C(_03550_),
    .A(_14816_),
    .Y(_03570_));
 sg13g2_nand3b_1 _25543_ (.B(_03570_),
    .C(net4713),
    .Y(_03571_),
    .A_N(_03569_));
 sg13g2_a21oi_1 _25544_ (.A1(net4595),
    .A2(\u_inv.d_next[146] ),
    .Y(_03572_),
    .B1(net3816));
 sg13g2_a22oi_1 _25545_ (.Y(_03573_),
    .B1(_03571_),
    .B2(_03572_),
    .A2(_03568_),
    .A1(net3816));
 sg13g2_nand2_1 _25546_ (.Y(_03574_),
    .A(net3464),
    .B(_03573_));
 sg13g2_xnor2_1 _25547_ (.Y(_03575_),
    .A(net3464),
    .B(_03573_));
 sg13g2_nand2_1 _25548_ (.Y(_03576_),
    .A(_03528_),
    .B(_03559_));
 sg13g2_a21oi_2 _25549_ (.B1(_03576_),
    .Y(_03577_),
    .A2(_03561_),
    .A1(_03542_));
 sg13g2_xnor2_1 _25550_ (.Y(_03578_),
    .A(_03575_),
    .B(_03577_));
 sg13g2_o21ai_1 _25551_ (.B1(net3909),
    .Y(_03579_),
    .A1(net4375),
    .A2(_03573_));
 sg13g2_a21oi_1 _25552_ (.A1(net4373),
    .A2(_03578_),
    .Y(_03580_),
    .B1(_03579_));
 sg13g2_a21o_1 _25553_ (.A2(net3996),
    .A1(net2959),
    .B1(_03580_),
    .X(_00422_));
 sg13g2_a21oi_1 _25554_ (.A1(net4595),
    .A2(\u_inv.d_next[147] ),
    .Y(_03581_),
    .B1(net3816));
 sg13g2_o21ai_1 _25555_ (.B1(_14813_),
    .Y(_03582_),
    .A1(_14814_),
    .A2(_03569_));
 sg13g2_nand3b_1 _25556_ (.B(_14812_),
    .C(_14815_),
    .Y(_03583_),
    .A_N(_03569_));
 sg13g2_nand3_1 _25557_ (.B(_03582_),
    .C(_03583_),
    .A(net4713),
    .Y(_03584_));
 sg13g2_o21ai_1 _25558_ (.B1(_14813_),
    .Y(_03585_),
    .A1(_14933_),
    .A2(_03566_));
 sg13g2_nor3_1 _25559_ (.A(_14813_),
    .B(_14933_),
    .C(_03566_),
    .Y(_03586_));
 sg13g2_nor2_1 _25560_ (.A(net3868),
    .B(_03586_),
    .Y(_03587_));
 sg13g2_a22oi_1 _25561_ (.Y(_03588_),
    .B1(_03585_),
    .B2(_03587_),
    .A2(_03584_),
    .A1(_03581_));
 sg13g2_xnor2_1 _25562_ (.Y(_03589_),
    .A(net3464),
    .B(_03588_));
 sg13g2_o21ai_1 _25563_ (.B1(_03574_),
    .Y(_03590_),
    .A1(_03575_),
    .A2(_03577_));
 sg13g2_xor2_1 _25564_ (.B(_03590_),
    .A(_03589_),
    .X(_03591_));
 sg13g2_o21ai_1 _25565_ (.B1(net3909),
    .Y(_03592_),
    .A1(net4375),
    .A2(_03588_));
 sg13g2_a21oi_1 _25566_ (.A1(net4375),
    .A2(_03591_),
    .Y(_03593_),
    .B1(_03592_));
 sg13g2_a21o_1 _25567_ (.A2(net3985),
    .A1(net2881),
    .B1(_03593_),
    .X(_00423_));
 sg13g2_o21ai_1 _25568_ (.B1(_14936_),
    .Y(_03594_),
    .A1(_14818_),
    .A2(_03565_));
 sg13g2_xnor2_1 _25569_ (.Y(_03595_),
    .A(_14807_),
    .B(_03594_));
 sg13g2_o21ai_1 _25570_ (.B1(_15249_),
    .Y(_03596_),
    .A1(_15257_),
    .A2(_03523_));
 sg13g2_xnor2_1 _25571_ (.Y(_03597_),
    .A(_14807_),
    .B(_03596_));
 sg13g2_nand2_1 _25572_ (.Y(_03598_),
    .A(net4709),
    .B(_03597_));
 sg13g2_a21oi_1 _25573_ (.A1(net4596),
    .A2(\u_inv.d_next[148] ),
    .Y(_03599_),
    .B1(net3818));
 sg13g2_a22oi_1 _25574_ (.Y(_03600_),
    .B1(_03598_),
    .B2(_03599_),
    .A2(_03595_),
    .A1(net3818));
 sg13g2_nand2_1 _25575_ (.Y(_03601_),
    .A(net3464),
    .B(_03600_));
 sg13g2_xnor2_1 _25576_ (.Y(_03602_),
    .A(net3487),
    .B(_03600_));
 sg13g2_inv_1 _25577_ (.Y(_03603_),
    .A(_03602_));
 sg13g2_o21ai_1 _25578_ (.B1(net3464),
    .Y(_03604_),
    .A1(_03573_),
    .A2(_03588_));
 sg13g2_or2_1 _25579_ (.X(_03605_),
    .B(_03589_),
    .A(_03575_));
 sg13g2_o21ai_1 _25580_ (.B1(_03604_),
    .Y(_03606_),
    .A1(_03577_),
    .A2(_03605_));
 sg13g2_nand2_1 _25581_ (.Y(_03607_),
    .A(_03602_),
    .B(_03606_));
 sg13g2_xnor2_1 _25582_ (.Y(_03608_),
    .A(_03602_),
    .B(_03606_));
 sg13g2_o21ai_1 _25583_ (.B1(net3907),
    .Y(_03609_),
    .A1(net4375),
    .A2(_03600_));
 sg13g2_a21oi_1 _25584_ (.A1(net4375),
    .A2(_03608_),
    .Y(_03610_),
    .B1(_03609_));
 sg13g2_a21o_1 _25585_ (.A2(net3986),
    .A1(net3197),
    .B1(_03610_),
    .X(_00424_));
 sg13g2_a21oi_1 _25586_ (.A1(net4600),
    .A2(\u_inv.d_next[149] ),
    .Y(_03611_),
    .B1(net3818));
 sg13g2_a21oi_1 _25587_ (.A1(_14806_),
    .A2(_03596_),
    .Y(_03612_),
    .B1(_14805_));
 sg13g2_o21ai_1 _25588_ (.B1(net4709),
    .Y(_03613_),
    .A1(_14804_),
    .A2(_03612_));
 sg13g2_a21o_1 _25589_ (.A2(_03612_),
    .A1(_14804_),
    .B1(_03613_),
    .X(_03614_));
 sg13g2_a21oi_1 _25590_ (.A1(_14807_),
    .A2(_03594_),
    .Y(_03615_),
    .B1(_14942_));
 sg13g2_or2_1 _25591_ (.X(_03616_),
    .B(_03615_),
    .A(_14804_));
 sg13g2_a21oi_1 _25592_ (.A1(_14804_),
    .A2(_03615_),
    .Y(_03617_),
    .B1(net3865));
 sg13g2_a22oi_1 _25593_ (.Y(_03618_),
    .B1(_03616_),
    .B2(_03617_),
    .A2(_03614_),
    .A1(_03611_));
 sg13g2_nand2_1 _25594_ (.Y(_03619_),
    .A(net3464),
    .B(_03618_));
 sg13g2_nor2_1 _25595_ (.A(net3465),
    .B(_03618_),
    .Y(_03620_));
 sg13g2_xnor2_1 _25596_ (.Y(_03621_),
    .A(net3464),
    .B(_03618_));
 sg13g2_nand2_1 _25597_ (.Y(_03622_),
    .A(_03601_),
    .B(_03607_));
 sg13g2_xor2_1 _25598_ (.B(_03622_),
    .A(_03621_),
    .X(_03623_));
 sg13g2_o21ai_1 _25599_ (.B1(net3907),
    .Y(_03624_),
    .A1(net4375),
    .A2(_03618_));
 sg13g2_a21oi_1 _25600_ (.A1(net4376),
    .A2(_03623_),
    .Y(_03625_),
    .B1(_03624_));
 sg13g2_a21o_1 _25601_ (.A2(net3986),
    .A1(net2837),
    .B1(_03625_),
    .X(_00425_));
 sg13g2_a21oi_1 _25602_ (.A1(_14808_),
    .A2(_03594_),
    .Y(_03626_),
    .B1(_14943_));
 sg13g2_xnor2_1 _25603_ (.Y(_03627_),
    .A(_14801_),
    .B(_03626_));
 sg13g2_a21oi_1 _25604_ (.A1(net4595),
    .A2(\u_inv.d_next[150] ),
    .Y(_03628_),
    .B1(net3818));
 sg13g2_a21oi_1 _25605_ (.A1(_15242_),
    .A2(_03596_),
    .Y(_03629_),
    .B1(_15252_));
 sg13g2_xnor2_1 _25606_ (.Y(_03630_),
    .A(_14801_),
    .B(_03629_));
 sg13g2_nand2_1 _25607_ (.Y(_03631_),
    .A(net4713),
    .B(_03630_));
 sg13g2_a22oi_1 _25608_ (.Y(_03632_),
    .B1(_03628_),
    .B2(_03631_),
    .A2(_03627_),
    .A1(net3818));
 sg13g2_nand2_1 _25609_ (.Y(_03633_),
    .A(net3465),
    .B(_03632_));
 sg13g2_xnor2_1 _25610_ (.Y(_03634_),
    .A(net3465),
    .B(_03632_));
 sg13g2_nand2_1 _25611_ (.Y(_03635_),
    .A(_03601_),
    .B(_03619_));
 sg13g2_a21oi_1 _25612_ (.A1(_03602_),
    .A2(_03606_),
    .Y(_03636_),
    .B1(_03635_));
 sg13g2_nor2_1 _25613_ (.A(_03620_),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_nand2b_1 _25614_ (.Y(_03638_),
    .B(_03637_),
    .A_N(_03634_));
 sg13g2_xor2_1 _25615_ (.B(_03637_),
    .A(_03634_),
    .X(_03639_));
 sg13g2_o21ai_1 _25616_ (.B1(net3907),
    .Y(_03640_),
    .A1(net4375),
    .A2(_03632_));
 sg13g2_a21oi_1 _25617_ (.A1(net4375),
    .A2(_03639_),
    .Y(_03641_),
    .B1(_03640_));
 sg13g2_a21o_1 _25618_ (.A2(net3986),
    .A1(net2972),
    .B1(_03641_),
    .X(_00426_));
 sg13g2_a21oi_1 _25619_ (.A1(net4595),
    .A2(\u_inv.d_next[151] ),
    .Y(_03642_),
    .B1(net3816));
 sg13g2_o21ai_1 _25620_ (.B1(_14798_),
    .Y(_03643_),
    .A1(_14799_),
    .A2(_03629_));
 sg13g2_o21ai_1 _25621_ (.B1(net4713),
    .Y(_03644_),
    .A1(_14797_),
    .A2(_03643_));
 sg13g2_a21o_1 _25622_ (.A2(_03643_),
    .A1(_14797_),
    .B1(_03644_),
    .X(_03645_));
 sg13g2_o21ai_1 _25623_ (.B1(_14938_),
    .Y(_03646_),
    .A1(_14801_),
    .A2(_03626_));
 sg13g2_or2_1 _25624_ (.X(_03647_),
    .B(_03646_),
    .A(_14797_));
 sg13g2_a21oi_1 _25625_ (.A1(_14797_),
    .A2(_03646_),
    .Y(_03648_),
    .B1(net3868));
 sg13g2_a22oi_1 _25626_ (.Y(_03649_),
    .B1(_03647_),
    .B2(_03648_),
    .A2(_03645_),
    .A1(_03642_));
 sg13g2_xnor2_1 _25627_ (.Y(_03650_),
    .A(net3488),
    .B(_03649_));
 sg13g2_nand2_1 _25628_ (.Y(_03651_),
    .A(_03633_),
    .B(_03638_));
 sg13g2_xnor2_1 _25629_ (.Y(_03652_),
    .A(_03650_),
    .B(_03651_));
 sg13g2_o21ai_1 _25630_ (.B1(net3909),
    .Y(_03653_),
    .A1(net4376),
    .A2(_03649_));
 sg13g2_a21oi_1 _25631_ (.A1(net4376),
    .A2(_03652_),
    .Y(_03654_),
    .B1(_03653_));
 sg13g2_a21o_1 _25632_ (.A2(net3985),
    .A1(net3152),
    .B1(_03654_),
    .X(_00427_));
 sg13g2_o21ai_1 _25633_ (.B1(_14827_),
    .Y(_03655_),
    .A1(_14929_),
    .A2(_03519_));
 sg13g2_a21oi_1 _25634_ (.A1(_14945_),
    .A2(_03655_),
    .Y(_03656_),
    .B1(_14792_));
 sg13g2_nand3_1 _25635_ (.B(_14945_),
    .C(_03655_),
    .A(_14792_),
    .Y(_03657_));
 sg13g2_nand2b_1 _25636_ (.Y(_03658_),
    .B(_03657_),
    .A_N(_03656_));
 sg13g2_o21ai_1 _25637_ (.B1(_15255_),
    .Y(_03659_),
    .A1(_15259_),
    .A2(_03523_));
 sg13g2_a21oi_1 _25638_ (.A1(_14792_),
    .A2(_03659_),
    .Y(_03660_),
    .B1(net4594));
 sg13g2_o21ai_1 _25639_ (.B1(_03660_),
    .Y(_03661_),
    .A1(_14792_),
    .A2(_03659_));
 sg13g2_a21oi_1 _25640_ (.A1(net4595),
    .A2(\u_inv.d_next[152] ),
    .Y(_03662_),
    .B1(net3819));
 sg13g2_a22oi_1 _25641_ (.Y(_03663_),
    .B1(_03661_),
    .B2(_03662_),
    .A2(_03658_),
    .A1(net3817));
 sg13g2_nand2_1 _25642_ (.Y(_03664_),
    .A(net3462),
    .B(_03663_));
 sg13g2_xnor2_1 _25643_ (.Y(_03665_),
    .A(net3487),
    .B(_03663_));
 sg13g2_inv_2 _25644_ (.Y(_03666_),
    .A(_03665_));
 sg13g2_nor2_1 _25645_ (.A(_03603_),
    .B(_03621_),
    .Y(_03667_));
 sg13g2_nand3b_1 _25646_ (.B(_03650_),
    .C(_03667_),
    .Y(_03668_),
    .A_N(_03634_));
 sg13g2_nand2b_1 _25647_ (.Y(_03669_),
    .B(_03576_),
    .A_N(_03605_));
 sg13g2_a21o_1 _25648_ (.A2(_03669_),
    .A1(_03604_),
    .B1(_03668_),
    .X(_03670_));
 sg13g2_o21ai_1 _25649_ (.B1(net3464),
    .Y(_03671_),
    .A1(_03632_),
    .A2(_03649_));
 sg13g2_nand3b_1 _25650_ (.B(_03635_),
    .C(_03650_),
    .Y(_03672_),
    .A_N(_03634_));
 sg13g2_nand3_1 _25651_ (.B(_03671_),
    .C(_03672_),
    .A(_03670_),
    .Y(_03673_));
 sg13g2_or4_1 _25652_ (.A(_03529_),
    .B(_03560_),
    .C(_03605_),
    .D(_03668_),
    .X(_03674_));
 sg13g2_a21oi_1 _25653_ (.A1(_03538_),
    .A2(_03541_),
    .Y(_03675_),
    .B1(_03674_));
 sg13g2_nor2_2 _25654_ (.A(_03673_),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_xnor2_1 _25655_ (.Y(_03677_),
    .A(_03666_),
    .B(_03676_));
 sg13g2_a21oi_1 _25656_ (.A1(net4374),
    .A2(_03677_),
    .Y(_03678_),
    .B1(net4239));
 sg13g2_o21ai_1 _25657_ (.B1(_03678_),
    .Y(_03679_),
    .A1(net4373),
    .A2(_03663_));
 sg13g2_o21ai_1 _25658_ (.B1(_03679_),
    .Y(_00428_),
    .A1(_10599_),
    .A2(net4043));
 sg13g2_nand2_1 _25659_ (.Y(_03680_),
    .A(net2501),
    .B(net3985));
 sg13g2_o21ai_1 _25660_ (.B1(_03664_),
    .Y(_03681_),
    .A1(_03666_),
    .A2(_03676_));
 sg13g2_a21oi_1 _25661_ (.A1(_14792_),
    .A2(_03659_),
    .Y(_03682_),
    .B1(_14791_));
 sg13g2_nand2b_1 _25662_ (.Y(_03683_),
    .B(_03682_),
    .A_N(_14790_));
 sg13g2_a221oi_1 _25663_ (.B2(_03659_),
    .C1(net4594),
    .B1(_15239_),
    .A1(_14790_),
    .Y(_03684_),
    .A2(_14791_));
 sg13g2_a221oi_1 _25664_ (.B2(_03684_),
    .C1(net3817),
    .B1(_03683_),
    .A1(net4595),
    .Y(_03685_),
    .A2(\u_inv.d_next[153] ));
 sg13g2_nor2_1 _25665_ (.A(_14948_),
    .B(_03656_),
    .Y(_03686_));
 sg13g2_xnor2_1 _25666_ (.Y(_03687_),
    .A(_14790_),
    .B(_03686_));
 sg13g2_a21oi_2 _25667_ (.B1(_03685_),
    .Y(_03688_),
    .A2(_03687_),
    .A1(net3817));
 sg13g2_xnor2_1 _25668_ (.Y(_03689_),
    .A(net3462),
    .B(_03688_));
 sg13g2_o21ai_1 _25669_ (.B1(net4374),
    .Y(_03690_),
    .A1(_03681_),
    .A2(_03689_));
 sg13g2_a21oi_1 _25670_ (.A1(_03681_),
    .A2(_03689_),
    .Y(_03691_),
    .B1(_03690_));
 sg13g2_o21ai_1 _25671_ (.B1(net3909),
    .Y(_03692_),
    .A1(net4373),
    .A2(_03688_));
 sg13g2_o21ai_1 _25672_ (.B1(_03680_),
    .Y(_00429_),
    .A1(_03691_),
    .A2(_03692_));
 sg13g2_a21oi_2 _25673_ (.B1(_14794_),
    .Y(_03693_),
    .A2(_03655_),
    .A1(_14945_));
 sg13g2_o21ai_1 _25674_ (.B1(_14786_),
    .Y(_03694_),
    .A1(_14949_),
    .A2(_03693_));
 sg13g2_or3_1 _25675_ (.A(_14786_),
    .B(_14949_),
    .C(_03693_),
    .X(_03695_));
 sg13g2_nand2_1 _25676_ (.Y(_03696_),
    .A(_03694_),
    .B(_03695_));
 sg13g2_a21oi_1 _25677_ (.A1(_15239_),
    .A2(_03659_),
    .Y(_03697_),
    .B1(_15289_));
 sg13g2_a21oi_1 _25678_ (.A1(_14786_),
    .A2(_03697_),
    .Y(_03698_),
    .B1(net4594));
 sg13g2_o21ai_1 _25679_ (.B1(_03698_),
    .Y(_03699_),
    .A1(_14786_),
    .A2(_03697_));
 sg13g2_a21oi_1 _25680_ (.A1(net4594),
    .A2(\u_inv.d_next[154] ),
    .Y(_03700_),
    .B1(net3817));
 sg13g2_a22oi_1 _25681_ (.Y(_03701_),
    .B1(_03699_),
    .B2(_03700_),
    .A2(_03696_),
    .A1(net3817));
 sg13g2_and2_1 _25682_ (.A(net3462),
    .B(_03701_),
    .X(_03702_));
 sg13g2_xnor2_1 _25683_ (.Y(_03703_),
    .A(net3463),
    .B(_03701_));
 sg13g2_o21ai_1 _25684_ (.B1(net3463),
    .Y(_03704_),
    .A1(_03663_),
    .A2(_03688_));
 sg13g2_or3_1 _25685_ (.A(_03666_),
    .B(_03676_),
    .C(_03689_),
    .X(_03705_));
 sg13g2_a21oi_1 _25686_ (.A1(_03704_),
    .A2(_03705_),
    .Y(_03706_),
    .B1(_03703_));
 sg13g2_nand3_1 _25687_ (.B(_03704_),
    .C(_03705_),
    .A(_03703_),
    .Y(_03707_));
 sg13g2_nand2b_1 _25688_ (.Y(_03708_),
    .B(_03707_),
    .A_N(_03706_));
 sg13g2_o21ai_1 _25689_ (.B1(net3909),
    .Y(_03709_),
    .A1(net4373),
    .A2(_03701_));
 sg13g2_a21oi_1 _25690_ (.A1(net4373),
    .A2(_03708_),
    .Y(_03710_),
    .B1(_03709_));
 sg13g2_a21o_1 _25691_ (.A2(net3985),
    .A1(net2870),
    .B1(_03710_),
    .X(_00430_));
 sg13g2_a21oi_1 _25692_ (.A1(net4594),
    .A2(\u_inv.d_next[155] ),
    .Y(_03711_),
    .B1(net3817));
 sg13g2_o21ai_1 _25693_ (.B1(_14785_),
    .Y(_03712_),
    .A1(_14786_),
    .A2(_03697_));
 sg13g2_xor2_1 _25694_ (.B(_03712_),
    .A(_14784_),
    .X(_03713_));
 sg13g2_o21ai_1 _25695_ (.B1(_03711_),
    .Y(_03714_),
    .A1(net4594),
    .A2(_03713_));
 sg13g2_a21o_1 _25696_ (.A2(_03694_),
    .A1(_14950_),
    .B1(_14784_),
    .X(_03715_));
 sg13g2_nand3_1 _25697_ (.B(_14950_),
    .C(_03694_),
    .A(_14784_),
    .Y(_03716_));
 sg13g2_nand3_1 _25698_ (.B(_03715_),
    .C(_03716_),
    .A(net3817),
    .Y(_03717_));
 sg13g2_and2_1 _25699_ (.A(_03714_),
    .B(_03717_),
    .X(_03718_));
 sg13g2_and3_1 _25700_ (.X(_03719_),
    .A(net3463),
    .B(_03714_),
    .C(_03717_));
 sg13g2_a21oi_1 _25701_ (.A1(_03714_),
    .A2(_03717_),
    .Y(_03720_),
    .B1(net3463));
 sg13g2_or2_1 _25702_ (.X(_03721_),
    .B(_03720_),
    .A(_03719_));
 sg13g2_nor2_1 _25703_ (.A(_03702_),
    .B(_03706_),
    .Y(_03722_));
 sg13g2_xnor2_1 _25704_ (.Y(_03723_),
    .A(_03721_),
    .B(_03722_));
 sg13g2_o21ai_1 _25705_ (.B1(net3909),
    .Y(_03724_),
    .A1(net4374),
    .A2(_03718_));
 sg13g2_a21oi_1 _25706_ (.A1(net4374),
    .A2(_03723_),
    .Y(_03725_),
    .B1(_03724_));
 sg13g2_a21o_1 _25707_ (.A2(net3985),
    .A1(net2747),
    .B1(_03725_),
    .X(_00431_));
 sg13g2_a21oi_2 _25708_ (.B1(_14952_),
    .Y(_03726_),
    .A2(_03693_),
    .A1(_14787_));
 sg13g2_xnor2_1 _25709_ (.Y(_03727_),
    .A(_14779_),
    .B(_03726_));
 sg13g2_nand3_1 _25710_ (.B(_15240_),
    .C(_03659_),
    .A(_15239_),
    .Y(_03728_));
 sg13g2_a21oi_1 _25711_ (.A1(_15291_),
    .A2(_03728_),
    .Y(_03729_),
    .B1(_14780_));
 sg13g2_nand3_1 _25712_ (.B(_15291_),
    .C(_03728_),
    .A(_14780_),
    .Y(_03730_));
 sg13g2_nand3b_1 _25713_ (.B(_03730_),
    .C(net4700),
    .Y(_03731_),
    .A_N(_03729_));
 sg13g2_a21oi_1 _25714_ (.A1(net4588),
    .A2(\u_inv.d_next[156] ),
    .Y(_03732_),
    .B1(net3808));
 sg13g2_a22oi_1 _25715_ (.Y(_03733_),
    .B1(_03731_),
    .B2(_03732_),
    .A2(_03727_),
    .A1(net3808));
 sg13g2_nand2_1 _25716_ (.Y(_03734_),
    .A(net3461),
    .B(_03733_));
 sg13g2_xnor2_1 _25717_ (.Y(_03735_),
    .A(net3461),
    .B(_03733_));
 sg13g2_nor4_1 _25718_ (.A(_03703_),
    .B(_03704_),
    .C(_03719_),
    .D(_03720_),
    .Y(_03736_));
 sg13g2_or3_1 _25719_ (.A(_03702_),
    .B(_03719_),
    .C(_03736_),
    .X(_03737_));
 sg13g2_nor4_1 _25720_ (.A(_03666_),
    .B(_03689_),
    .C(_03703_),
    .D(_03721_),
    .Y(_03738_));
 sg13g2_o21ai_1 _25721_ (.B1(_03738_),
    .Y(_03739_),
    .A1(_03673_),
    .A2(_03675_));
 sg13g2_nand2b_1 _25722_ (.Y(_03740_),
    .B(_03739_),
    .A_N(_03737_));
 sg13g2_nand2b_1 _25723_ (.Y(_03741_),
    .B(_03740_),
    .A_N(_03735_));
 sg13g2_xor2_1 _25724_ (.B(_03740_),
    .A(_03735_),
    .X(_03742_));
 sg13g2_o21ai_1 _25725_ (.B1(net3905),
    .Y(_03743_),
    .A1(net4372),
    .A2(_03733_));
 sg13g2_a21oi_1 _25726_ (.A1(net4377),
    .A2(_03742_),
    .Y(_03744_),
    .B1(_03743_));
 sg13g2_a21o_1 _25727_ (.A2(net3985),
    .A1(net2966),
    .B1(_03744_),
    .X(_00432_));
 sg13g2_a21oi_1 _25728_ (.A1(net4588),
    .A2(\u_inv.d_next[157] ),
    .Y(_03745_),
    .B1(net3807));
 sg13g2_nand3b_1 _25729_ (.B(_14775_),
    .C(_14778_),
    .Y(_03746_),
    .A_N(_03729_));
 sg13g2_o21ai_1 _25730_ (.B1(_14776_),
    .Y(_03747_),
    .A1(_14777_),
    .A2(_03729_));
 sg13g2_nand3_1 _25731_ (.B(_03746_),
    .C(_03747_),
    .A(net4700),
    .Y(_03748_));
 sg13g2_o21ai_1 _25732_ (.B1(_14953_),
    .Y(_03749_),
    .A1(_14779_),
    .A2(_03726_));
 sg13g2_or2_1 _25733_ (.X(_03750_),
    .B(_03749_),
    .A(_14776_));
 sg13g2_a21oi_1 _25734_ (.A1(_14776_),
    .A2(_03749_),
    .Y(_03751_),
    .B1(net3864));
 sg13g2_a22oi_1 _25735_ (.Y(_03752_),
    .B1(_03750_),
    .B2(_03751_),
    .A2(_03748_),
    .A1(_03745_));
 sg13g2_nor2_1 _25736_ (.A(net3461),
    .B(_03752_),
    .Y(_03753_));
 sg13g2_xnor2_1 _25737_ (.Y(_03754_),
    .A(net3487),
    .B(_03752_));
 sg13g2_nand2_1 _25738_ (.Y(_03755_),
    .A(_03734_),
    .B(_03741_));
 sg13g2_xnor2_1 _25739_ (.Y(_03756_),
    .A(_03754_),
    .B(_03755_));
 sg13g2_o21ai_1 _25740_ (.B1(net3905),
    .Y(_03757_),
    .A1(net4372),
    .A2(_03752_));
 sg13g2_a21oi_1 _25741_ (.A1(net4372),
    .A2(_03756_),
    .Y(_03758_),
    .B1(_03757_));
 sg13g2_a21o_1 _25742_ (.A2(net3978),
    .A1(net3190),
    .B1(_03758_),
    .X(_00433_));
 sg13g2_o21ai_1 _25743_ (.B1(_14955_),
    .Y(_03759_),
    .A1(_14781_),
    .A2(_03726_));
 sg13g2_xnor2_1 _25744_ (.Y(_03760_),
    .A(_14773_),
    .B(_03759_));
 sg13g2_a21oi_1 _25745_ (.A1(_15291_),
    .A2(_03728_),
    .Y(_03761_),
    .B1(_15237_));
 sg13g2_or3_1 _25746_ (.A(_14772_),
    .B(_15294_),
    .C(_03761_),
    .X(_03762_));
 sg13g2_o21ai_1 _25747_ (.B1(_14772_),
    .Y(_03763_),
    .A1(_15294_),
    .A2(_03761_));
 sg13g2_nand3_1 _25748_ (.B(_03762_),
    .C(_03763_),
    .A(net4700),
    .Y(_03764_));
 sg13g2_a21oi_1 _25749_ (.A1(net4588),
    .A2(\u_inv.d_next[158] ),
    .Y(_03765_),
    .B1(net3807));
 sg13g2_a22oi_1 _25750_ (.Y(_03766_),
    .B1(_03764_),
    .B2(_03765_),
    .A2(_03760_),
    .A1(net3808));
 sg13g2_and2_1 _25751_ (.A(net3461),
    .B(_03766_),
    .X(_03767_));
 sg13g2_xnor2_1 _25752_ (.Y(_03768_),
    .A(net3487),
    .B(_03766_));
 sg13g2_o21ai_1 _25753_ (.B1(net3461),
    .Y(_03769_),
    .A1(_03733_),
    .A2(_03752_));
 sg13g2_a21oi_1 _25754_ (.A1(_03741_),
    .A2(_03769_),
    .Y(_03770_),
    .B1(_03753_));
 sg13g2_xnor2_1 _25755_ (.Y(_03771_),
    .A(_03768_),
    .B(_03770_));
 sg13g2_a21oi_1 _25756_ (.A1(net4372),
    .A2(_03771_),
    .Y(_03772_),
    .B1(net4238));
 sg13g2_o21ai_1 _25757_ (.B1(_03772_),
    .Y(_03773_),
    .A1(net4372),
    .A2(_03766_));
 sg13g2_o21ai_1 _25758_ (.B1(_03773_),
    .Y(_00434_),
    .A1(_10598_),
    .A2(net4038));
 sg13g2_nand2_1 _25759_ (.Y(_03774_),
    .A(net2460),
    .B(net3978));
 sg13g2_a21oi_1 _25760_ (.A1(net4588),
    .A2(\u_inv.d_next[159] ),
    .Y(_03775_),
    .B1(net3808));
 sg13g2_nand3_1 _25761_ (.B(_14771_),
    .C(_03763_),
    .A(_14770_),
    .Y(_03776_));
 sg13g2_a21o_1 _25762_ (.A2(_03763_),
    .A1(_14771_),
    .B1(_14770_),
    .X(_03777_));
 sg13g2_nand3_1 _25763_ (.B(_03776_),
    .C(_03777_),
    .A(net4700),
    .Y(_03778_));
 sg13g2_a21oi_1 _25764_ (.A1(_14773_),
    .A2(_03759_),
    .Y(_03779_),
    .B1(_14956_));
 sg13g2_or2_1 _25765_ (.X(_03780_),
    .B(_03779_),
    .A(_14770_));
 sg13g2_a21oi_1 _25766_ (.A1(_14770_),
    .A2(_03779_),
    .Y(_03781_),
    .B1(net3859));
 sg13g2_a22oi_1 _25767_ (.Y(_03782_),
    .B1(_03780_),
    .B2(_03781_),
    .A2(_03778_),
    .A1(_03775_));
 sg13g2_xnor2_1 _25768_ (.Y(_03783_),
    .A(net3487),
    .B(_03782_));
 sg13g2_a21oi_1 _25769_ (.A1(_03768_),
    .A2(_03770_),
    .Y(_03784_),
    .B1(_03767_));
 sg13g2_o21ai_1 _25770_ (.B1(net4372),
    .Y(_03785_),
    .A1(_03783_),
    .A2(_03784_));
 sg13g2_a21oi_1 _25771_ (.A1(_03783_),
    .A2(_03784_),
    .Y(_03786_),
    .B1(_03785_));
 sg13g2_o21ai_1 _25772_ (.B1(net3905),
    .Y(_03787_),
    .A1(net4372),
    .A2(_03782_));
 sg13g2_o21ai_1 _25773_ (.B1(_03774_),
    .Y(_00435_),
    .A1(_03786_),
    .A2(_03787_));
 sg13g2_a21oi_2 _25774_ (.B1(_14899_),
    .Y(_03788_),
    .A2(_14656_),
    .A1(_14537_));
 sg13g2_nor2_1 _25775_ (.A(_14962_),
    .B(_03788_),
    .Y(_03789_));
 sg13g2_nor2_1 _25776_ (.A(_14762_),
    .B(_03789_),
    .Y(_03790_));
 sg13g2_xnor2_1 _25777_ (.Y(_03791_),
    .A(_14762_),
    .B(_03789_));
 sg13g2_a21oi_2 _25778_ (.B1(_15298_),
    .Y(_03792_),
    .A2(_15635_),
    .A1(net3586));
 sg13g2_a21o_2 _25779_ (.A2(_15635_),
    .A1(_15630_),
    .B1(_15298_),
    .X(_03793_));
 sg13g2_a21oi_1 _25780_ (.A1(_14763_),
    .A2(_03792_),
    .Y(_03794_),
    .B1(net4587));
 sg13g2_o21ai_1 _25781_ (.B1(_03794_),
    .Y(_03795_),
    .A1(_14763_),
    .A2(_03792_));
 sg13g2_a21oi_1 _25782_ (.A1(net4587),
    .A2(\u_inv.d_next[160] ),
    .Y(_03796_),
    .B1(net3809));
 sg13g2_a22oi_1 _25783_ (.Y(_03797_),
    .B1(_03795_),
    .B2(_03796_),
    .A2(_03791_),
    .A1(net3809));
 sg13g2_nand2_1 _25784_ (.Y(_03798_),
    .A(net3452),
    .B(_03797_));
 sg13g2_xnor2_1 _25785_ (.Y(_03799_),
    .A(net3452),
    .B(_03797_));
 sg13g2_nor2b_1 _25786_ (.A(_03735_),
    .B_N(_03754_),
    .Y(_03800_));
 sg13g2_nand4_1 _25787_ (.B(_03768_),
    .C(_03783_),
    .A(_03738_),
    .Y(_03801_),
    .D(_03800_));
 sg13g2_inv_1 _25788_ (.Y(_03802_),
    .A(_03801_));
 sg13g2_nor2_1 _25789_ (.A(_03674_),
    .B(_03801_),
    .Y(_03803_));
 sg13g2_nand4_1 _25790_ (.B(_03768_),
    .C(_03783_),
    .A(_03737_),
    .Y(_03804_),
    .D(_03800_));
 sg13g2_nand3b_1 _25791_ (.B(_03783_),
    .C(_03768_),
    .Y(_03805_),
    .A_N(_03769_));
 sg13g2_o21ai_1 _25792_ (.B1(net3461),
    .Y(_03806_),
    .A1(_03766_),
    .A2(_03782_));
 sg13g2_nand3_1 _25793_ (.B(_03805_),
    .C(_03806_),
    .A(_03804_),
    .Y(_03807_));
 sg13g2_a221oi_1 _25794_ (.B2(_03539_),
    .C1(_03807_),
    .B1(_03803_),
    .A1(_03673_),
    .Y(_03808_),
    .A2(_03802_));
 sg13g2_or3_1 _25795_ (.A(_03540_),
    .B(_03674_),
    .C(_03801_),
    .X(_03809_));
 sg13g2_a21oi_1 _25796_ (.A1(_03259_),
    .A2(_03265_),
    .Y(_03810_),
    .B1(_03809_));
 sg13g2_nand2b_2 _25797_ (.Y(_03811_),
    .B(_03808_),
    .A_N(_03810_));
 sg13g2_nand2b_1 _25798_ (.Y(_03812_),
    .B(_03811_),
    .A_N(_03799_));
 sg13g2_xor2_1 _25799_ (.B(_03811_),
    .A(_03799_),
    .X(_03813_));
 sg13g2_a21oi_1 _25800_ (.A1(net4363),
    .A2(_03813_),
    .Y(_03814_),
    .B1(net4238));
 sg13g2_o21ai_1 _25801_ (.B1(_03814_),
    .Y(_03815_),
    .A1(net4363),
    .A2(_03797_));
 sg13g2_o21ai_1 _25802_ (.B1(_03815_),
    .Y(_00436_),
    .A1(_10597_),
    .A2(net4038));
 sg13g2_nand2_1 _25803_ (.Y(_03816_),
    .A(net2685),
    .B(net3977));
 sg13g2_nand2_1 _25804_ (.Y(_03817_),
    .A(_03798_),
    .B(_03812_));
 sg13g2_a21oi_1 _25805_ (.A1(_15232_),
    .A2(_03793_),
    .Y(_03818_),
    .B1(_15202_));
 sg13g2_nand2_1 _25806_ (.Y(_03819_),
    .A(_14760_),
    .B(_14761_));
 sg13g2_a21oi_1 _25807_ (.A1(_14762_),
    .A2(_03793_),
    .Y(_03820_),
    .B1(_03819_));
 sg13g2_nand3b_1 _25808_ (.B(_03818_),
    .C(net4700),
    .Y(_03821_),
    .A_N(_03820_));
 sg13g2_a21oi_1 _25809_ (.A1(net4587),
    .A2(\u_inv.d_next[161] ),
    .Y(_03822_),
    .B1(net3810));
 sg13g2_or2_1 _25810_ (.X(_03823_),
    .B(_03790_),
    .A(_14994_));
 sg13g2_xnor2_1 _25811_ (.Y(_03824_),
    .A(_14760_),
    .B(_03823_));
 sg13g2_a22oi_1 _25812_ (.Y(_03825_),
    .B1(_03824_),
    .B2(net3809),
    .A2(_03822_),
    .A1(_03821_));
 sg13g2_xnor2_1 _25813_ (.Y(_03826_),
    .A(net3452),
    .B(_03825_));
 sg13g2_o21ai_1 _25814_ (.B1(net4363),
    .Y(_03827_),
    .A1(_03817_),
    .A2(_03826_));
 sg13g2_a21oi_1 _25815_ (.A1(_03817_),
    .A2(_03826_),
    .Y(_03828_),
    .B1(_03827_));
 sg13g2_o21ai_1 _25816_ (.B1(net3904),
    .Y(_03829_),
    .A1(net4363),
    .A2(_03825_));
 sg13g2_o21ai_1 _25817_ (.B1(_03816_),
    .Y(_00437_),
    .A1(_03828_),
    .A2(_03829_));
 sg13g2_o21ai_1 _25818_ (.B1(_14764_),
    .Y(_03830_),
    .A1(_14962_),
    .A2(_03788_));
 sg13g2_a21oi_1 _25819_ (.A1(_14995_),
    .A2(_03830_),
    .Y(_03831_),
    .B1(_14755_));
 sg13g2_nand3_1 _25820_ (.B(_14995_),
    .C(_03830_),
    .A(_14755_),
    .Y(_03832_));
 sg13g2_nand2b_1 _25821_ (.Y(_03833_),
    .B(_03832_),
    .A_N(_03831_));
 sg13g2_a221oi_1 _25822_ (.B2(_03793_),
    .C1(_15202_),
    .B1(_15232_),
    .A1(\u_inv.d_next[161] ),
    .Y(_03834_),
    .A2(\u_inv.d_reg[161] ));
 sg13g2_a21oi_1 _25823_ (.A1(_14756_),
    .A2(_03834_),
    .Y(_03835_),
    .B1(net4586));
 sg13g2_o21ai_1 _25824_ (.B1(_03835_),
    .Y(_03836_),
    .A1(_14756_),
    .A2(_03834_));
 sg13g2_a21oi_1 _25825_ (.A1(net4586),
    .A2(\u_inv.d_next[162] ),
    .Y(_03837_),
    .B1(net3806));
 sg13g2_a22oi_1 _25826_ (.Y(_03838_),
    .B1(_03836_),
    .B2(_03837_),
    .A2(_03833_),
    .A1(net3806));
 sg13g2_nand2_1 _25827_ (.Y(_03839_),
    .A(net3452),
    .B(_03838_));
 sg13g2_xnor2_1 _25828_ (.Y(_03840_),
    .A(net3453),
    .B(_03838_));
 sg13g2_o21ai_1 _25829_ (.B1(net3452),
    .Y(_03841_),
    .A1(_03797_),
    .A2(_03825_));
 sg13g2_nand2_1 _25830_ (.Y(_03842_),
    .A(_03812_),
    .B(_03841_));
 sg13g2_o21ai_1 _25831_ (.B1(_03842_),
    .Y(_03843_),
    .A1(net3453),
    .A2(_03825_));
 sg13g2_xnor2_1 _25832_ (.Y(_03844_),
    .A(_03840_),
    .B(_03843_));
 sg13g2_o21ai_1 _25833_ (.B1(net3904),
    .Y(_03845_),
    .A1(net4363),
    .A2(_03838_));
 sg13g2_a21oi_1 _25834_ (.A1(net4363),
    .A2(_03844_),
    .Y(_03846_),
    .B1(_03845_));
 sg13g2_a21o_1 _25835_ (.A2(net3978),
    .A1(net2855),
    .B1(_03846_),
    .X(_00438_));
 sg13g2_a21oi_1 _25836_ (.A1(net4586),
    .A2(\u_inv.d_next[163] ),
    .Y(_03847_),
    .B1(net3806));
 sg13g2_o21ai_1 _25837_ (.B1(_14753_),
    .Y(_03848_),
    .A1(_14756_),
    .A2(_03834_));
 sg13g2_xnor2_1 _25838_ (.Y(_03849_),
    .A(_14752_),
    .B(_03848_));
 sg13g2_o21ai_1 _25839_ (.B1(_03847_),
    .Y(_03850_),
    .A1(net4586),
    .A2(_03849_));
 sg13g2_o21ai_1 _25840_ (.B1(_14752_),
    .Y(_03851_),
    .A1(_14996_),
    .A2(_03831_));
 sg13g2_or3_1 _25841_ (.A(_14752_),
    .B(_14996_),
    .C(_03831_),
    .X(_03852_));
 sg13g2_nand3_1 _25842_ (.B(_03851_),
    .C(_03852_),
    .A(net3806),
    .Y(_03853_));
 sg13g2_and2_1 _25843_ (.A(_03850_),
    .B(_03853_),
    .X(_03854_));
 sg13g2_and3_1 _25844_ (.X(_03855_),
    .A(net3452),
    .B(_03850_),
    .C(_03853_));
 sg13g2_a21oi_1 _25845_ (.A1(_03850_),
    .A2(_03853_),
    .Y(_03856_),
    .B1(net3452));
 sg13g2_nor2_1 _25846_ (.A(_03855_),
    .B(_03856_),
    .Y(_03857_));
 sg13g2_o21ai_1 _25847_ (.B1(_03839_),
    .Y(_03858_),
    .A1(_03840_),
    .A2(_03843_));
 sg13g2_xnor2_1 _25848_ (.Y(_03859_),
    .A(_03857_),
    .B(_03858_));
 sg13g2_o21ai_1 _25849_ (.B1(net3904),
    .Y(_03860_),
    .A1(net4363),
    .A2(_03854_));
 sg13g2_a21oi_1 _25850_ (.A1(net4364),
    .A2(_03859_),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_a21o_1 _25851_ (.A2(net3977),
    .A1(net4801),
    .B1(_03861_),
    .X(_00439_));
 sg13g2_o21ai_1 _25852_ (.B1(_14999_),
    .Y(_03862_),
    .A1(_14757_),
    .A2(_03830_));
 sg13g2_xnor2_1 _25853_ (.Y(_03863_),
    .A(_14746_),
    .B(_03862_));
 sg13g2_o21ai_1 _25854_ (.B1(_15206_),
    .Y(_03864_),
    .A1(_15233_),
    .A2(_03792_));
 sg13g2_xnor2_1 _25855_ (.Y(_03865_),
    .A(_14746_),
    .B(_03864_));
 sg13g2_nand2_1 _25856_ (.Y(_03866_),
    .A(net4701),
    .B(_03865_));
 sg13g2_a21oi_1 _25857_ (.A1(net4589),
    .A2(\u_inv.d_next[164] ),
    .Y(_03867_),
    .B1(net3810));
 sg13g2_a22oi_1 _25858_ (.Y(_03868_),
    .B1(_03866_),
    .B2(_03867_),
    .A2(_03863_),
    .A1(net3810));
 sg13g2_nand2_1 _25859_ (.Y(_03869_),
    .A(net3456),
    .B(_03868_));
 sg13g2_xnor2_1 _25860_ (.Y(_03870_),
    .A(net3456),
    .B(_03868_));
 sg13g2_or3_1 _25861_ (.A(_03840_),
    .B(_03855_),
    .C(_03856_),
    .X(_03871_));
 sg13g2_a21oi_1 _25862_ (.A1(net3452),
    .A2(_03838_),
    .Y(_03872_),
    .B1(_03855_));
 sg13g2_o21ai_1 _25863_ (.B1(_03872_),
    .Y(_03873_),
    .A1(_03841_),
    .A2(_03871_));
 sg13g2_nor3_1 _25864_ (.A(_03799_),
    .B(_03826_),
    .C(_03871_),
    .Y(_03874_));
 sg13g2_a21oi_1 _25865_ (.A1(_03811_),
    .A2(_03874_),
    .Y(_03875_),
    .B1(_03873_));
 sg13g2_nor2_1 _25866_ (.A(_03870_),
    .B(_03875_),
    .Y(_03876_));
 sg13g2_xnor2_1 _25867_ (.Y(_03877_),
    .A(_03870_),
    .B(_03875_));
 sg13g2_o21ai_1 _25868_ (.B1(net3906),
    .Y(_03878_),
    .A1(net4368),
    .A2(_03868_));
 sg13g2_a21oi_1 _25869_ (.A1(net4368),
    .A2(_03877_),
    .Y(_03879_),
    .B1(_03878_));
 sg13g2_a21o_1 _25870_ (.A2(net3977),
    .A1(net3255),
    .B1(_03879_),
    .X(_00440_));
 sg13g2_a21oi_1 _25871_ (.A1(net4589),
    .A2(\u_inv.d_next[165] ),
    .Y(_03880_),
    .B1(net3810));
 sg13g2_a21o_1 _25872_ (.A2(_03864_),
    .A1(_14745_),
    .B1(_14744_),
    .X(_03881_));
 sg13g2_xnor2_1 _25873_ (.Y(_03882_),
    .A(_14743_),
    .B(_03881_));
 sg13g2_nand2_1 _25874_ (.Y(_03883_),
    .A(net4701),
    .B(_03882_));
 sg13g2_a21oi_1 _25875_ (.A1(_14746_),
    .A2(_03862_),
    .Y(_03884_),
    .B1(_15003_));
 sg13g2_or2_1 _25876_ (.X(_03885_),
    .B(_03884_),
    .A(_14743_));
 sg13g2_a21oi_1 _25877_ (.A1(_14743_),
    .A2(_03884_),
    .Y(_03886_),
    .B1(net3864));
 sg13g2_a22oi_1 _25878_ (.Y(_03887_),
    .B1(_03885_),
    .B2(_03886_),
    .A2(_03883_),
    .A1(_03880_));
 sg13g2_nand2_1 _25879_ (.Y(_03888_),
    .A(net3456),
    .B(_03887_));
 sg13g2_nor2_1 _25880_ (.A(net3456),
    .B(_03887_),
    .Y(_03889_));
 sg13g2_xnor2_1 _25881_ (.Y(_03890_),
    .A(net3485),
    .B(_03887_));
 sg13g2_a21oi_1 _25882_ (.A1(net3458),
    .A2(_03868_),
    .Y(_03891_),
    .B1(_03876_));
 sg13g2_xnor2_1 _25883_ (.Y(_03892_),
    .A(_03890_),
    .B(_03891_));
 sg13g2_nor2_1 _25884_ (.A(net4368),
    .B(_03887_),
    .Y(_03893_));
 sg13g2_nor2_1 _25885_ (.A(net4238),
    .B(_03893_),
    .Y(_03894_));
 sg13g2_o21ai_1 _25886_ (.B1(_03894_),
    .Y(_03895_),
    .A1(net4297),
    .A2(_03892_));
 sg13g2_o21ai_1 _25887_ (.B1(_03895_),
    .Y(_00441_),
    .A1(_10596_),
    .A2(net4038));
 sg13g2_a21oi_1 _25888_ (.A1(_14747_),
    .A2(_03862_),
    .Y(_03896_),
    .B1(_15004_));
 sg13g2_xnor2_1 _25889_ (.Y(_03897_),
    .A(_14740_),
    .B(_03896_));
 sg13g2_a21oi_1 _25890_ (.A1(_15200_),
    .A2(_03864_),
    .Y(_03898_),
    .B1(_15208_));
 sg13g2_xnor2_1 _25891_ (.Y(_03899_),
    .A(_14740_),
    .B(_03898_));
 sg13g2_nand2_1 _25892_ (.Y(_03900_),
    .A(net4702),
    .B(_03899_));
 sg13g2_a21oi_1 _25893_ (.A1(net4586),
    .A2(\u_inv.d_next[166] ),
    .Y(_03901_),
    .B1(net3806));
 sg13g2_a22oi_1 _25894_ (.Y(_03902_),
    .B1(_03900_),
    .B2(_03901_),
    .A2(_03897_),
    .A1(net3811));
 sg13g2_nand2_1 _25895_ (.Y(_03903_),
    .A(net3456),
    .B(_03902_));
 sg13g2_xnor2_1 _25896_ (.Y(_03904_),
    .A(net3485),
    .B(_03902_));
 sg13g2_nand2_1 _25897_ (.Y(_03905_),
    .A(_03869_),
    .B(_03888_));
 sg13g2_o21ai_1 _25898_ (.B1(_03888_),
    .Y(_03906_),
    .A1(_03889_),
    .A2(_03891_));
 sg13g2_nand2_1 _25899_ (.Y(_03907_),
    .A(_03904_),
    .B(_03906_));
 sg13g2_xnor2_1 _25900_ (.Y(_03908_),
    .A(_03904_),
    .B(_03906_));
 sg13g2_o21ai_1 _25901_ (.B1(net3906),
    .Y(_03909_),
    .A1(net4370),
    .A2(_03902_));
 sg13g2_a21oi_1 _25902_ (.A1(net4370),
    .A2(_03908_),
    .Y(_03910_),
    .B1(_03909_));
 sg13g2_a21o_1 _25903_ (.A2(net3979),
    .A1(net2935),
    .B1(_03910_),
    .X(_00442_));
 sg13g2_a21oi_1 _25904_ (.A1(net4589),
    .A2(\u_inv.d_next[167] ),
    .Y(_03911_),
    .B1(net3810));
 sg13g2_o21ai_1 _25905_ (.B1(_14738_),
    .Y(_03912_),
    .A1(_14739_),
    .A2(_03898_));
 sg13g2_o21ai_1 _25906_ (.B1(net4701),
    .Y(_03913_),
    .A1(_14737_),
    .A2(_03912_));
 sg13g2_a21o_1 _25907_ (.A2(_03912_),
    .A1(_14737_),
    .B1(_03913_),
    .X(_03914_));
 sg13g2_o21ai_1 _25908_ (.B1(_15000_),
    .Y(_03915_),
    .A1(_14740_),
    .A2(_03896_));
 sg13g2_or2_1 _25909_ (.X(_03916_),
    .B(_03915_),
    .A(_14737_));
 sg13g2_a21oi_1 _25910_ (.A1(_14737_),
    .A2(_03915_),
    .Y(_03917_),
    .B1(net3864));
 sg13g2_a22oi_1 _25911_ (.Y(_03918_),
    .B1(_03916_),
    .B2(_03917_),
    .A2(_03914_),
    .A1(_03911_));
 sg13g2_xnor2_1 _25912_ (.Y(_03919_),
    .A(net3485),
    .B(_03918_));
 sg13g2_nand2_1 _25913_ (.Y(_03920_),
    .A(_03903_),
    .B(_03907_));
 sg13g2_xnor2_1 _25914_ (.Y(_03921_),
    .A(_03919_),
    .B(_03920_));
 sg13g2_o21ai_1 _25915_ (.B1(net3906),
    .Y(_03922_),
    .A1(net4368),
    .A2(_03918_));
 sg13g2_a21oi_1 _25916_ (.A1(net4368),
    .A2(_03921_),
    .Y(_03923_),
    .B1(_03922_));
 sg13g2_a21o_1 _25917_ (.A2(net3977),
    .A1(net3158),
    .B1(_03923_),
    .X(_00443_));
 sg13g2_o21ai_1 _25918_ (.B1(_14766_),
    .Y(_03924_),
    .A1(_14962_),
    .A2(_03788_));
 sg13g2_nand2_1 _25919_ (.Y(_03925_),
    .A(_15005_),
    .B(_03924_));
 sg13g2_xnor2_1 _25920_ (.Y(_03926_),
    .A(_14733_),
    .B(_03925_));
 sg13g2_o21ai_1 _25921_ (.B1(_15213_),
    .Y(_03927_),
    .A1(_15234_),
    .A2(_03792_));
 sg13g2_nand2b_1 _25922_ (.Y(_03928_),
    .B(_03927_),
    .A_N(_14733_));
 sg13g2_nand2b_1 _25923_ (.Y(_03929_),
    .B(_14733_),
    .A_N(_03927_));
 sg13g2_nand3_1 _25924_ (.B(_03928_),
    .C(_03929_),
    .A(net4701),
    .Y(_03930_));
 sg13g2_a21oi_1 _25925_ (.A1(net4589),
    .A2(\u_inv.d_next[168] ),
    .Y(_03931_),
    .B1(net3810));
 sg13g2_a22oi_1 _25926_ (.Y(_03932_),
    .B1(_03930_),
    .B2(_03931_),
    .A2(_03926_),
    .A1(net3810));
 sg13g2_and2_1 _25927_ (.A(net3456),
    .B(_03932_),
    .X(_03933_));
 sg13g2_xnor2_1 _25928_ (.Y(_03934_),
    .A(net3456),
    .B(_03932_));
 sg13g2_nor2b_1 _25929_ (.A(_03870_),
    .B_N(_03890_),
    .Y(_03935_));
 sg13g2_nand4_1 _25930_ (.B(_03904_),
    .C(_03919_),
    .A(_03873_),
    .Y(_03936_),
    .D(_03935_));
 sg13g2_nand3_1 _25931_ (.B(_03905_),
    .C(_03919_),
    .A(_03904_),
    .Y(_03937_));
 sg13g2_o21ai_1 _25932_ (.B1(net3456),
    .Y(_03938_),
    .A1(_03902_),
    .A2(_03918_));
 sg13g2_nand3_1 _25933_ (.B(_03937_),
    .C(_03938_),
    .A(_03936_),
    .Y(_03939_));
 sg13g2_and4_1 _25934_ (.A(_03874_),
    .B(_03904_),
    .C(_03919_),
    .D(_03935_),
    .X(_03940_));
 sg13g2_a21oi_1 _25935_ (.A1(_03811_),
    .A2(_03940_),
    .Y(_03941_),
    .B1(_03939_));
 sg13g2_nor2_1 _25936_ (.A(_03934_),
    .B(_03941_),
    .Y(_03942_));
 sg13g2_xnor2_1 _25937_ (.Y(_03943_),
    .A(_03934_),
    .B(_03941_));
 sg13g2_o21ai_1 _25938_ (.B1(net3906),
    .Y(_03944_),
    .A1(net4368),
    .A2(_03932_));
 sg13g2_a21oi_1 _25939_ (.A1(net4368),
    .A2(_03943_),
    .Y(_03945_),
    .B1(_03944_));
 sg13g2_a21o_1 _25940_ (.A2(net3979),
    .A1(net2794),
    .B1(_03945_),
    .X(_00444_));
 sg13g2_nand2_1 _25941_ (.Y(_03946_),
    .A(net2133),
    .B(net3977));
 sg13g2_nor2_1 _25942_ (.A(_03933_),
    .B(_03942_),
    .Y(_03947_));
 sg13g2_nand3_1 _25943_ (.B(_14732_),
    .C(_03928_),
    .A(_14731_),
    .Y(_03948_));
 sg13g2_a21oi_1 _25944_ (.A1(_15219_),
    .A2(_03927_),
    .Y(_03949_),
    .B1(net4589));
 sg13g2_nand3b_1 _25945_ (.B(_03948_),
    .C(_03949_),
    .Y(_03950_),
    .A_N(_15221_));
 sg13g2_a21oi_1 _25946_ (.A1(net4589),
    .A2(\u_inv.d_next[169] ),
    .Y(_03951_),
    .B1(net3811));
 sg13g2_a21oi_1 _25947_ (.A1(_14733_),
    .A2(_03925_),
    .Y(_03952_),
    .B1(_15007_));
 sg13g2_xor2_1 _25948_ (.B(_03952_),
    .A(_14731_),
    .X(_03953_));
 sg13g2_a22oi_1 _25949_ (.Y(_03954_),
    .B1(_03953_),
    .B2(net3810),
    .A2(_03951_),
    .A1(_03950_));
 sg13g2_xnor2_1 _25950_ (.Y(_03955_),
    .A(net3485),
    .B(_03954_));
 sg13g2_o21ai_1 _25951_ (.B1(net4368),
    .Y(_03956_),
    .A1(_03947_),
    .A2(_03955_));
 sg13g2_a21oi_1 _25952_ (.A1(_03947_),
    .A2(_03955_),
    .Y(_03957_),
    .B1(_03956_));
 sg13g2_o21ai_1 _25953_ (.B1(net3906),
    .Y(_03958_),
    .A1(net4370),
    .A2(_03954_));
 sg13g2_o21ai_1 _25954_ (.B1(_03946_),
    .Y(_00445_),
    .A1(_03957_),
    .A2(_03958_));
 sg13g2_a21oi_2 _25955_ (.B1(_14734_),
    .Y(_03959_),
    .A2(_03924_),
    .A1(_15005_));
 sg13g2_o21ai_1 _25956_ (.B1(_14728_),
    .Y(_03960_),
    .A1(_15009_),
    .A2(_03959_));
 sg13g2_or3_1 _25957_ (.A(_14728_),
    .B(_15009_),
    .C(_03959_),
    .X(_03961_));
 sg13g2_nand2_1 _25958_ (.Y(_03962_),
    .A(_03960_),
    .B(_03961_));
 sg13g2_a221oi_1 _25959_ (.B2(_03927_),
    .C1(_15221_),
    .B1(_15219_),
    .A1(\u_inv.d_next[169] ),
    .Y(_03963_),
    .A2(\u_inv.d_reg[169] ));
 sg13g2_a21oi_1 _25960_ (.A1(_14728_),
    .A2(_03963_),
    .Y(_03964_),
    .B1(net4592));
 sg13g2_o21ai_1 _25961_ (.B1(_03964_),
    .Y(_03965_),
    .A1(_14728_),
    .A2(_03963_));
 sg13g2_a21oi_1 _25962_ (.A1(net4592),
    .A2(\u_inv.d_next[170] ),
    .Y(_03966_),
    .B1(net3814));
 sg13g2_a22oi_1 _25963_ (.Y(_03967_),
    .B1(_03965_),
    .B2(_03966_),
    .A2(_03962_),
    .A1(net3814));
 sg13g2_and2_1 _25964_ (.A(net3457),
    .B(_03967_),
    .X(_03968_));
 sg13g2_nand2b_1 _25965_ (.Y(_03969_),
    .B(net3485),
    .A_N(_03967_));
 sg13g2_xnor2_1 _25966_ (.Y(_03970_),
    .A(net3457),
    .B(_03967_));
 sg13g2_a21oi_1 _25967_ (.A1(net3457),
    .A2(_03954_),
    .Y(_03971_),
    .B1(_03933_));
 sg13g2_inv_1 _25968_ (.Y(_03972_),
    .A(_03971_));
 sg13g2_nand2b_1 _25969_ (.Y(_03973_),
    .B(_03955_),
    .A_N(_03934_));
 sg13g2_o21ai_1 _25970_ (.B1(_03971_),
    .Y(_03974_),
    .A1(_03941_),
    .A2(_03973_));
 sg13g2_xor2_1 _25971_ (.B(_03974_),
    .A(_03970_),
    .X(_03975_));
 sg13g2_a21oi_1 _25972_ (.A1(net4369),
    .A2(_03975_),
    .Y(_03976_),
    .B1(net4238));
 sg13g2_o21ai_1 _25973_ (.B1(_03976_),
    .Y(_03977_),
    .A1(net4369),
    .A2(_03967_));
 sg13g2_o21ai_1 _25974_ (.B1(_03977_),
    .Y(_00446_),
    .A1(_10595_),
    .A2(net4038));
 sg13g2_nand2_1 _25975_ (.Y(_03978_),
    .A(_10594_),
    .B(net3862));
 sg13g2_o21ai_1 _25976_ (.B1(net3862),
    .Y(_03979_),
    .A1(net4708),
    .A2(_10594_));
 sg13g2_o21ai_1 _25977_ (.B1(_14727_),
    .Y(_03980_),
    .A1(_14728_),
    .A2(_03963_));
 sg13g2_xnor2_1 _25978_ (.Y(_03981_),
    .A(_14725_),
    .B(_03980_));
 sg13g2_a22oi_1 _25979_ (.Y(_03982_),
    .B1(_03981_),
    .B2(net4708),
    .A2(_03978_),
    .A1(net3735));
 sg13g2_a21o_1 _25980_ (.A2(_03981_),
    .A1(net4708),
    .B1(_03979_),
    .X(_03983_));
 sg13g2_a21o_1 _25981_ (.A2(_03960_),
    .A1(_15010_),
    .B1(_14725_),
    .X(_03984_));
 sg13g2_nand3_1 _25982_ (.B(_15010_),
    .C(_03960_),
    .A(_14725_),
    .Y(_03985_));
 sg13g2_and3_1 _25983_ (.X(_03986_),
    .A(net3814),
    .B(_03984_),
    .C(_03985_));
 sg13g2_nand3_1 _25984_ (.B(_03984_),
    .C(_03985_),
    .A(net3814),
    .Y(_03987_));
 sg13g2_nor3_1 _25985_ (.A(net3486),
    .B(_03982_),
    .C(_03986_),
    .Y(_03988_));
 sg13g2_a21oi_1 _25986_ (.A1(_03983_),
    .A2(_03987_),
    .Y(_03989_),
    .B1(net3457));
 sg13g2_nor2_1 _25987_ (.A(_03988_),
    .B(_03989_),
    .Y(_03990_));
 sg13g2_a21oi_1 _25988_ (.A1(_03969_),
    .A2(_03974_),
    .Y(_03991_),
    .B1(_03968_));
 sg13g2_xor2_1 _25989_ (.B(_03991_),
    .A(_03990_),
    .X(_03992_));
 sg13g2_o21ai_1 _25990_ (.B1(net4297),
    .Y(_03993_),
    .A1(_03982_),
    .A2(_03986_));
 sg13g2_nand2_1 _25991_ (.Y(_03994_),
    .A(net3910),
    .B(_03993_));
 sg13g2_a21oi_1 _25992_ (.A1(net4369),
    .A2(_03992_),
    .Y(_03995_),
    .B1(_03994_));
 sg13g2_a21o_1 _25993_ (.A2(net3984),
    .A1(net2873),
    .B1(_03995_),
    .X(_00447_));
 sg13g2_a21oi_2 _25994_ (.B1(_15014_),
    .Y(_03996_),
    .A2(_03959_),
    .A1(_14729_));
 sg13g2_xnor2_1 _25995_ (.Y(_03997_),
    .A(_14721_),
    .B(_03996_));
 sg13g2_and3_2 _25996_ (.X(_03998_),
    .A(_15218_),
    .B(_15219_),
    .C(_03927_));
 sg13g2_o21ai_1 _25997_ (.B1(_14721_),
    .Y(_03999_),
    .A1(_15224_),
    .A2(_03998_));
 sg13g2_or3_1 _25998_ (.A(_14721_),
    .B(_15224_),
    .C(_03998_),
    .X(_04000_));
 sg13g2_nand3_1 _25999_ (.B(_03999_),
    .C(_04000_),
    .A(net4708),
    .Y(_04001_));
 sg13g2_a21oi_1 _26000_ (.A1(net4592),
    .A2(\u_inv.d_next[172] ),
    .Y(_04002_),
    .B1(net3814));
 sg13g2_a22oi_1 _26001_ (.Y(_04003_),
    .B1(_04001_),
    .B2(_04002_),
    .A2(_03997_),
    .A1(net3814));
 sg13g2_nand2_1 _26002_ (.Y(_04004_),
    .A(net3457),
    .B(_04003_));
 sg13g2_xnor2_1 _26003_ (.Y(_04005_),
    .A(net3457),
    .B(_04003_));
 sg13g2_or2_1 _26004_ (.X(_04006_),
    .B(_03988_),
    .A(_03968_));
 sg13g2_nor3_1 _26005_ (.A(_03970_),
    .B(_03988_),
    .C(_03989_),
    .Y(_04007_));
 sg13g2_a21o_1 _26006_ (.A2(_04007_),
    .A1(_03974_),
    .B1(_04006_),
    .X(_04008_));
 sg13g2_nand2b_1 _26007_ (.Y(_04009_),
    .B(_04008_),
    .A_N(_04005_));
 sg13g2_xor2_1 _26008_ (.B(_04008_),
    .A(_04005_),
    .X(_04010_));
 sg13g2_a21oi_1 _26009_ (.A1(net4369),
    .A2(_04010_),
    .Y(_04011_),
    .B1(net4239));
 sg13g2_o21ai_1 _26010_ (.B1(_04011_),
    .Y(_04012_),
    .A1(net4370),
    .A2(_04003_));
 sg13g2_o21ai_1 _26011_ (.B1(_04012_),
    .Y(_00448_),
    .A1(_10594_),
    .A2(net4037));
 sg13g2_nand2_1 _26012_ (.Y(_04013_),
    .A(net2987),
    .B(net3984));
 sg13g2_nand3_1 _26013_ (.B(_14720_),
    .C(_03999_),
    .A(_14719_),
    .Y(_04014_));
 sg13g2_o21ai_1 _26014_ (.B1(_15215_),
    .Y(_04015_),
    .A1(_15224_),
    .A2(_03998_));
 sg13g2_nor2_1 _26015_ (.A(net4592),
    .B(_15225_),
    .Y(_04016_));
 sg13g2_nand3_1 _26016_ (.B(_04015_),
    .C(_04016_),
    .A(_04014_),
    .Y(_04017_));
 sg13g2_a21oi_1 _26017_ (.A1(net4592),
    .A2(\u_inv.d_next[173] ),
    .Y(_04018_),
    .B1(net3814));
 sg13g2_o21ai_1 _26018_ (.B1(_15015_),
    .Y(_04019_),
    .A1(_14721_),
    .A2(_03996_));
 sg13g2_xnor2_1 _26019_ (.Y(_04020_),
    .A(_14719_),
    .B(_04019_));
 sg13g2_a22oi_1 _26020_ (.Y(_04021_),
    .B1(_04020_),
    .B2(net3814),
    .A2(_04018_),
    .A1(_04017_));
 sg13g2_nand2_1 _26021_ (.Y(_04022_),
    .A(net3458),
    .B(_04021_));
 sg13g2_xnor2_1 _26022_ (.Y(_04023_),
    .A(net3458),
    .B(_04021_));
 sg13g2_nand2_1 _26023_ (.Y(_04024_),
    .A(_04004_),
    .B(_04009_));
 sg13g2_o21ai_1 _26024_ (.B1(net4370),
    .Y(_04025_),
    .A1(_04023_),
    .A2(_04024_));
 sg13g2_a21oi_1 _26025_ (.A1(_04023_),
    .A2(_04024_),
    .Y(_04026_),
    .B1(_04025_));
 sg13g2_o21ai_1 _26026_ (.B1(net3906),
    .Y(_04027_),
    .A1(net4370),
    .A2(_04021_));
 sg13g2_o21ai_1 _26027_ (.B1(_04013_),
    .Y(_00449_),
    .A1(_04026_),
    .A2(_04027_));
 sg13g2_o21ai_1 _26028_ (.B1(_15018_),
    .Y(_04028_),
    .A1(_14723_),
    .A2(_03996_));
 sg13g2_xnor2_1 _26029_ (.Y(_04029_),
    .A(_14716_),
    .B(_04028_));
 sg13g2_a21o_1 _26030_ (.A2(_04015_),
    .A1(_15226_),
    .B1(_14716_),
    .X(_04030_));
 sg13g2_nand3_1 _26031_ (.B(_15226_),
    .C(_04015_),
    .A(_14716_),
    .Y(_04031_));
 sg13g2_nand3_1 _26032_ (.B(_04030_),
    .C(_04031_),
    .A(net4705),
    .Y(_04032_));
 sg13g2_a21oi_1 _26033_ (.A1(net4590),
    .A2(\u_inv.d_next[174] ),
    .Y(_04033_),
    .B1(net3813));
 sg13g2_a22oi_1 _26034_ (.Y(_04034_),
    .B1(_04032_),
    .B2(_04033_),
    .A2(_04029_),
    .A1(net3813));
 sg13g2_nand2_1 _26035_ (.Y(_04035_),
    .A(net3457),
    .B(_04034_));
 sg13g2_xnor2_1 _26036_ (.Y(_04036_),
    .A(net3486),
    .B(_04034_));
 sg13g2_nand2_1 _26037_ (.Y(_04037_),
    .A(_04004_),
    .B(_04022_));
 sg13g2_nor2_1 _26038_ (.A(_04005_),
    .B(_04023_),
    .Y(_04038_));
 sg13g2_a21o_1 _26039_ (.A2(_04038_),
    .A1(_04008_),
    .B1(_04037_),
    .X(_04039_));
 sg13g2_nand2_1 _26040_ (.Y(_04040_),
    .A(_04036_),
    .B(_04039_));
 sg13g2_xnor2_1 _26041_ (.Y(_04041_),
    .A(_04036_),
    .B(_04039_));
 sg13g2_a21oi_1 _26042_ (.A1(net4369),
    .A2(_04041_),
    .Y(_04042_),
    .B1(net4238));
 sg13g2_o21ai_1 _26043_ (.B1(_04042_),
    .Y(_04043_),
    .A1(net4369),
    .A2(_04034_));
 sg13g2_o21ai_1 _26044_ (.B1(_04043_),
    .Y(_00450_),
    .A1(_10593_),
    .A2(net4035));
 sg13g2_a21oi_1 _26045_ (.A1(net4590),
    .A2(\u_inv.d_next[175] ),
    .Y(_04044_),
    .B1(net3813));
 sg13g2_a21o_1 _26046_ (.A2(_04030_),
    .A1(_14715_),
    .B1(_14714_),
    .X(_04045_));
 sg13g2_nand3_1 _26047_ (.B(_14715_),
    .C(_04030_),
    .A(_14714_),
    .Y(_04046_));
 sg13g2_nand3_1 _26048_ (.B(_04045_),
    .C(_04046_),
    .A(net4705),
    .Y(_04047_));
 sg13g2_a21oi_1 _26049_ (.A1(_14716_),
    .A2(_04028_),
    .Y(_04048_),
    .B1(_15020_));
 sg13g2_or2_1 _26050_ (.X(_04049_),
    .B(_04048_),
    .A(_14714_));
 sg13g2_a21oi_1 _26051_ (.A1(_14714_),
    .A2(_04048_),
    .Y(_04050_),
    .B1(net3860));
 sg13g2_a22oi_1 _26052_ (.Y(_04051_),
    .B1(_04049_),
    .B2(_04050_),
    .A2(_04047_),
    .A1(_04044_));
 sg13g2_nand2_1 _26053_ (.Y(_04052_),
    .A(net3457),
    .B(_04051_));
 sg13g2_xnor2_1 _26054_ (.Y(_04053_),
    .A(net3486),
    .B(_04051_));
 sg13g2_nand2_1 _26055_ (.Y(_04054_),
    .A(_04035_),
    .B(_04040_));
 sg13g2_xnor2_1 _26056_ (.Y(_04055_),
    .A(_04053_),
    .B(_04054_));
 sg13g2_o21ai_1 _26057_ (.B1(net3906),
    .Y(_04056_),
    .A1(net4369),
    .A2(_04051_));
 sg13g2_a21oi_1 _26058_ (.A1(net4369),
    .A2(_04055_),
    .Y(_04057_),
    .B1(_04056_));
 sg13g2_a21o_1 _26059_ (.A2(net3981),
    .A1(net2436),
    .B1(_04057_),
    .X(_00451_));
 sg13g2_o21ai_1 _26060_ (.B1(_14768_),
    .Y(_04058_),
    .A1(_14962_),
    .A2(_03788_));
 sg13g2_nand2_1 _26061_ (.Y(_04059_),
    .A(_15023_),
    .B(_04058_));
 sg13g2_xnor2_1 _26062_ (.Y(_04060_),
    .A(_14708_),
    .B(_04059_));
 sg13g2_a21oi_2 _26063_ (.B1(_15231_),
    .Y(_04061_),
    .A2(_03793_),
    .A1(_15235_));
 sg13g2_a21o_2 _26064_ (.A2(_03793_),
    .A1(_15235_),
    .B1(_15231_),
    .X(_04062_));
 sg13g2_nor2_1 _26065_ (.A(_14708_),
    .B(_04061_),
    .Y(_04063_));
 sg13g2_a21oi_1 _26066_ (.A1(_14708_),
    .A2(_04061_),
    .Y(_04064_),
    .B1(net4590));
 sg13g2_nand2b_1 _26067_ (.Y(_04065_),
    .B(_04064_),
    .A_N(_04063_));
 sg13g2_a21oi_1 _26068_ (.A1(net4590),
    .A2(\u_inv.d_next[176] ),
    .Y(_04066_),
    .B1(net3812));
 sg13g2_a22oi_1 _26069_ (.Y(_04067_),
    .B1(_04065_),
    .B2(_04066_),
    .A2(_04060_),
    .A1(net3812));
 sg13g2_and2_1 _26070_ (.A(net3454),
    .B(_04067_),
    .X(_04068_));
 sg13g2_xnor2_1 _26071_ (.Y(_04069_),
    .A(net3454),
    .B(_04067_));
 sg13g2_nor2b_1 _26072_ (.A(_03973_),
    .B_N(_04007_),
    .Y(_04070_));
 sg13g2_and4_1 _26073_ (.A(_04036_),
    .B(_04038_),
    .C(_04053_),
    .D(_04070_),
    .X(_04071_));
 sg13g2_and2_1 _26074_ (.A(_03939_),
    .B(_04071_),
    .X(_04072_));
 sg13g2_a21o_1 _26075_ (.A2(_04007_),
    .A1(_03972_),
    .B1(_04006_),
    .X(_04073_));
 sg13g2_nand4_1 _26076_ (.B(_04038_),
    .C(_04053_),
    .A(_04036_),
    .Y(_04074_),
    .D(_04073_));
 sg13g2_nand3_1 _26077_ (.B(_04037_),
    .C(_04053_),
    .A(_04036_),
    .Y(_04075_));
 sg13g2_nand4_1 _26078_ (.B(_04052_),
    .C(_04074_),
    .A(_04035_),
    .Y(_04076_),
    .D(_04075_));
 sg13g2_and2_1 _26079_ (.A(_03940_),
    .B(_04071_),
    .X(_04077_));
 sg13g2_a221oi_1 _26080_ (.B2(_03811_),
    .C1(_04076_),
    .B1(_04077_),
    .A1(_03939_),
    .Y(_04078_),
    .A2(_04071_));
 sg13g2_nor2_1 _26081_ (.A(_04069_),
    .B(_04078_),
    .Y(_04079_));
 sg13g2_xnor2_1 _26082_ (.Y(_04080_),
    .A(_04069_),
    .B(_04078_));
 sg13g2_o21ai_1 _26083_ (.B1(net3900),
    .Y(_04081_),
    .A1(net4366),
    .A2(_04067_));
 sg13g2_a21oi_1 _26084_ (.A1(net4366),
    .A2(_04080_),
    .Y(_04082_),
    .B1(_04081_));
 sg13g2_a21o_1 _26085_ (.A2(net3981),
    .A1(net2846),
    .B1(_04082_),
    .X(_00452_));
 sg13g2_nand2_1 _26086_ (.Y(_04083_),
    .A(net2674),
    .B(net3981));
 sg13g2_nor2_1 _26087_ (.A(_04068_),
    .B(_04079_),
    .Y(_04084_));
 sg13g2_nand2_1 _26088_ (.Y(_04085_),
    .A(_14706_),
    .B(_14707_));
 sg13g2_o21ai_1 _26089_ (.B1(net4705),
    .Y(_04086_),
    .A1(_14706_),
    .A2(_14707_));
 sg13g2_a21oi_1 _26090_ (.A1(_15197_),
    .A2(_04062_),
    .Y(_04087_),
    .B1(_04086_));
 sg13g2_o21ai_1 _26091_ (.B1(_04087_),
    .Y(_04088_),
    .A1(_04063_),
    .A2(_04085_));
 sg13g2_a21oi_1 _26092_ (.A1(net4590),
    .A2(\u_inv.d_next[177] ),
    .Y(_04089_),
    .B1(net3812));
 sg13g2_a21oi_1 _26093_ (.A1(_14708_),
    .A2(_04059_),
    .Y(_04090_),
    .B1(_14964_));
 sg13g2_xor2_1 _26094_ (.B(_04090_),
    .A(_14706_),
    .X(_04091_));
 sg13g2_a22oi_1 _26095_ (.Y(_04092_),
    .B1(_04091_),
    .B2(net3812),
    .A2(_04089_),
    .A1(_04088_));
 sg13g2_xnor2_1 _26096_ (.Y(_04093_),
    .A(net3454),
    .B(_04092_));
 sg13g2_inv_1 _26097_ (.Y(_04094_),
    .A(_04093_));
 sg13g2_o21ai_1 _26098_ (.B1(net4366),
    .Y(_04095_),
    .A1(_04084_),
    .A2(_04094_));
 sg13g2_a21oi_1 _26099_ (.A1(_04084_),
    .A2(_04094_),
    .Y(_04096_),
    .B1(_04095_));
 sg13g2_o21ai_1 _26100_ (.B1(net3906),
    .Y(_04097_),
    .A1(net4366),
    .A2(_04092_));
 sg13g2_o21ai_1 _26101_ (.B1(_04083_),
    .Y(_00453_),
    .A1(_04096_),
    .A2(_04097_));
 sg13g2_a21oi_2 _26102_ (.B1(_14709_),
    .Y(_04098_),
    .A2(_04058_),
    .A1(_15023_));
 sg13g2_nor2_1 _26103_ (.A(_14965_),
    .B(_04098_),
    .Y(_04099_));
 sg13g2_o21ai_1 _26104_ (.B1(_14702_),
    .Y(_04100_),
    .A1(_14965_),
    .A2(_04098_));
 sg13g2_xnor2_1 _26105_ (.Y(_04101_),
    .A(_14701_),
    .B(_04099_));
 sg13g2_a21oi_1 _26106_ (.A1(_15197_),
    .A2(_04062_),
    .Y(_04102_),
    .B1(_15311_));
 sg13g2_a21oi_1 _26107_ (.A1(_14702_),
    .A2(_04102_),
    .Y(_04103_),
    .B1(net4590));
 sg13g2_o21ai_1 _26108_ (.B1(_04103_),
    .Y(_04104_),
    .A1(_14702_),
    .A2(_04102_));
 sg13g2_a21oi_1 _26109_ (.A1(net4590),
    .A2(\u_inv.d_next[178] ),
    .Y(_04105_),
    .B1(net3812));
 sg13g2_a22oi_1 _26110_ (.Y(_04106_),
    .B1(_04104_),
    .B2(_04105_),
    .A2(_04101_),
    .A1(net3812));
 sg13g2_and2_1 _26111_ (.A(net3454),
    .B(_04106_),
    .X(_04107_));
 sg13g2_xnor2_1 _26112_ (.Y(_04108_),
    .A(net3455),
    .B(_04106_));
 sg13g2_a21oi_1 _26113_ (.A1(net3454),
    .A2(_04092_),
    .Y(_04109_),
    .B1(_04068_));
 sg13g2_inv_1 _26114_ (.Y(_04110_),
    .A(_04109_));
 sg13g2_nor3_1 _26115_ (.A(_04069_),
    .B(_04078_),
    .C(_04093_),
    .Y(_04111_));
 sg13g2_nor2_1 _26116_ (.A(_04110_),
    .B(_04111_),
    .Y(_04112_));
 sg13g2_nor2_1 _26117_ (.A(_04108_),
    .B(_04112_),
    .Y(_04113_));
 sg13g2_xor2_1 _26118_ (.B(_04112_),
    .A(_04108_),
    .X(_04114_));
 sg13g2_nor2_1 _26119_ (.A(net4366),
    .B(_04106_),
    .Y(_04115_));
 sg13g2_o21ai_1 _26120_ (.B1(net3900),
    .Y(_04116_),
    .A1(net4297),
    .A2(_04114_));
 sg13g2_nand2_1 _26121_ (.Y(_04117_),
    .A(net2635),
    .B(net3981));
 sg13g2_o21ai_1 _26122_ (.B1(_04117_),
    .Y(_00454_),
    .A1(_04115_),
    .A2(_04116_));
 sg13g2_a21oi_1 _26123_ (.A1(net4590),
    .A2(\u_inv.d_next[179] ),
    .Y(_04118_),
    .B1(net3812));
 sg13g2_o21ai_1 _26124_ (.B1(_14700_),
    .Y(_04119_),
    .A1(_14702_),
    .A2(_04102_));
 sg13g2_o21ai_1 _26125_ (.B1(net4705),
    .Y(_04120_),
    .A1(_14699_),
    .A2(_04119_));
 sg13g2_a21o_1 _26126_ (.A2(_04119_),
    .A1(_14699_),
    .B1(_04120_),
    .X(_04121_));
 sg13g2_a21oi_1 _26127_ (.A1(_14966_),
    .A2(_04100_),
    .Y(_04122_),
    .B1(_14698_));
 sg13g2_nand3_1 _26128_ (.B(_14966_),
    .C(_04100_),
    .A(_14698_),
    .Y(_04123_));
 sg13g2_nor2_1 _26129_ (.A(net3860),
    .B(_04122_),
    .Y(_04124_));
 sg13g2_a22oi_1 _26130_ (.Y(_04125_),
    .B1(_04123_),
    .B2(_04124_),
    .A2(_04121_),
    .A1(_04118_));
 sg13g2_xnor2_1 _26131_ (.Y(_04126_),
    .A(net3454),
    .B(_04125_));
 sg13g2_nor2_1 _26132_ (.A(_04107_),
    .B(_04113_),
    .Y(_04127_));
 sg13g2_xnor2_1 _26133_ (.Y(_04128_),
    .A(_04126_),
    .B(_04127_));
 sg13g2_o21ai_1 _26134_ (.B1(net3900),
    .Y(_04129_),
    .A1(net4366),
    .A2(_04125_));
 sg13g2_a21oi_1 _26135_ (.A1(net4366),
    .A2(_04128_),
    .Y(_04130_),
    .B1(_04129_));
 sg13g2_a21o_1 _26136_ (.A2(net3981),
    .A1(net2893),
    .B1(_04130_),
    .X(_00455_));
 sg13g2_a21oi_2 _26137_ (.B1(_14968_),
    .Y(_04131_),
    .A2(_04098_),
    .A1(_14703_));
 sg13g2_xnor2_1 _26138_ (.Y(_04132_),
    .A(_14689_),
    .B(_04131_));
 sg13g2_and4_1 _26139_ (.A(_14699_),
    .B(_14701_),
    .C(_15197_),
    .D(_04062_),
    .X(_04133_));
 sg13g2_nor3_1 _26140_ (.A(_14689_),
    .B(_15314_),
    .C(_04133_),
    .Y(_04134_));
 sg13g2_o21ai_1 _26141_ (.B1(_14689_),
    .Y(_04135_),
    .A1(_15314_),
    .A2(_04133_));
 sg13g2_nand3b_1 _26142_ (.B(_04135_),
    .C(net4698),
    .Y(_04136_),
    .A_N(_04134_));
 sg13g2_a21oi_1 _26143_ (.A1(net4580),
    .A2(\u_inv.d_next[180] ),
    .Y(_04137_),
    .B1(net3812));
 sg13g2_a22oi_1 _26144_ (.Y(_04138_),
    .B1(_04136_),
    .B2(_04137_),
    .A2(_04132_),
    .A1(net3813));
 sg13g2_nand2_1 _26145_ (.Y(_04139_),
    .A(net3455),
    .B(_04138_));
 sg13g2_xnor2_1 _26146_ (.Y(_04140_),
    .A(net3455),
    .B(_04138_));
 sg13g2_a21oi_1 _26147_ (.A1(net3454),
    .A2(_04125_),
    .Y(_04141_),
    .B1(_04107_));
 sg13g2_nor2_1 _26148_ (.A(_04108_),
    .B(_04126_),
    .Y(_04142_));
 sg13g2_o21ai_1 _26149_ (.B1(_04142_),
    .Y(_04143_),
    .A1(_04110_),
    .A2(_04111_));
 sg13g2_a21o_1 _26150_ (.A2(_04143_),
    .A1(_04141_),
    .B1(_04140_),
    .X(_04144_));
 sg13g2_nand3_1 _26151_ (.B(_04141_),
    .C(_04143_),
    .A(_04140_),
    .Y(_04145_));
 sg13g2_nand2_1 _26152_ (.Y(_04146_),
    .A(_04144_),
    .B(_04145_));
 sg13g2_o21ai_1 _26153_ (.B1(net3901),
    .Y(_04147_),
    .A1(net4365),
    .A2(_04138_));
 sg13g2_a21oi_1 _26154_ (.A1(net4365),
    .A2(_04146_),
    .Y(_04148_),
    .B1(_04147_));
 sg13g2_a21o_1 _26155_ (.A2(net3974),
    .A1(net3216),
    .B1(_04148_),
    .X(_00456_));
 sg13g2_nand2_1 _26156_ (.Y(_04149_),
    .A(net3047),
    .B(net3974));
 sg13g2_nand3_1 _26157_ (.B(_14688_),
    .C(_04135_),
    .A(_14687_),
    .Y(_04150_));
 sg13g2_o21ai_1 _26158_ (.B1(_15195_),
    .Y(_04151_),
    .A1(_15314_),
    .A2(_04133_));
 sg13g2_nor2_1 _26159_ (.A(net4581),
    .B(_15315_),
    .Y(_04152_));
 sg13g2_nand3_1 _26160_ (.B(_04151_),
    .C(_04152_),
    .A(_04150_),
    .Y(_04153_));
 sg13g2_a21oi_1 _26161_ (.A1(net4580),
    .A2(\u_inv.d_next[181] ),
    .Y(_04154_),
    .B1(net3801));
 sg13g2_o21ai_1 _26162_ (.B1(_14969_),
    .Y(_04155_),
    .A1(_14689_),
    .A2(_04131_));
 sg13g2_xnor2_1 _26163_ (.Y(_04156_),
    .A(_14687_),
    .B(_04155_));
 sg13g2_a22oi_1 _26164_ (.Y(_04157_),
    .B1(_04156_),
    .B2(net3801),
    .A2(_04154_),
    .A1(_04153_));
 sg13g2_xnor2_1 _26165_ (.Y(_04158_),
    .A(net3455),
    .B(_04157_));
 sg13g2_nand2_1 _26166_ (.Y(_04159_),
    .A(_04139_),
    .B(_04144_));
 sg13g2_o21ai_1 _26167_ (.B1(net4365),
    .Y(_04160_),
    .A1(_04158_),
    .A2(_04159_));
 sg13g2_a21oi_1 _26168_ (.A1(_04158_),
    .A2(_04159_),
    .Y(_04161_),
    .B1(_04160_));
 sg13g2_o21ai_1 _26169_ (.B1(net3901),
    .Y(_04162_),
    .A1(net4365),
    .A2(_04157_));
 sg13g2_o21ai_1 _26170_ (.B1(_04149_),
    .Y(_00457_),
    .A1(_04161_),
    .A2(_04162_));
 sg13g2_o21ai_1 _26171_ (.B1(_14971_),
    .Y(_04163_),
    .A1(_14691_),
    .A2(_04131_));
 sg13g2_xnor2_1 _26172_ (.Y(_04164_),
    .A(_14695_),
    .B(_04163_));
 sg13g2_nand3_1 _26173_ (.B(_15316_),
    .C(_04151_),
    .A(_14695_),
    .Y(_04165_));
 sg13g2_a21o_1 _26174_ (.A2(_04151_),
    .A1(_15316_),
    .B1(_14695_),
    .X(_04166_));
 sg13g2_nand3_1 _26175_ (.B(_04165_),
    .C(_04166_),
    .A(net4698),
    .Y(_04167_));
 sg13g2_a21oi_1 _26176_ (.A1(net4580),
    .A2(\u_inv.d_next[182] ),
    .Y(_04168_),
    .B1(net3801));
 sg13g2_a22oi_1 _26177_ (.Y(_04169_),
    .B1(_04167_),
    .B2(_04168_),
    .A2(_04164_),
    .A1(net3801));
 sg13g2_nand2_1 _26178_ (.Y(_04170_),
    .A(net3455),
    .B(_04169_));
 sg13g2_inv_1 _26179_ (.Y(_04171_),
    .A(_04170_));
 sg13g2_xnor2_1 _26180_ (.Y(_04172_),
    .A(net3485),
    .B(_04169_));
 sg13g2_o21ai_1 _26181_ (.B1(net3455),
    .Y(_04173_),
    .A1(_04138_),
    .A2(_04157_));
 sg13g2_o21ai_1 _26182_ (.B1(_04173_),
    .Y(_04174_),
    .A1(_04144_),
    .A2(_04158_));
 sg13g2_xnor2_1 _26183_ (.Y(_04175_),
    .A(_04172_),
    .B(_04174_));
 sg13g2_a21oi_1 _26184_ (.A1(net4365),
    .A2(_04175_),
    .Y(_04176_),
    .B1(net4236));
 sg13g2_o21ai_1 _26185_ (.B1(_04176_),
    .Y(_04177_),
    .A1(net4365),
    .A2(_04169_));
 sg13g2_o21ai_1 _26186_ (.B1(_04177_),
    .Y(_00458_),
    .A1(_10592_),
    .A2(net4032));
 sg13g2_a21oi_1 _26187_ (.A1(net4581),
    .A2(\u_inv.d_next[183] ),
    .Y(_04178_),
    .B1(net3801));
 sg13g2_nand3_1 _26188_ (.B(_14694_),
    .C(_04166_),
    .A(_14693_),
    .Y(_04179_));
 sg13g2_a21o_1 _26189_ (.A2(_04166_),
    .A1(_14694_),
    .B1(_14693_),
    .X(_04180_));
 sg13g2_nand3_1 _26190_ (.B(_04179_),
    .C(_04180_),
    .A(net4698),
    .Y(_04181_));
 sg13g2_a21oi_1 _26191_ (.A1(_14695_),
    .A2(_04163_),
    .Y(_04182_),
    .B1(_14972_));
 sg13g2_or2_1 _26192_ (.X(_04183_),
    .B(_04182_),
    .A(_14693_));
 sg13g2_a21oi_1 _26193_ (.A1(_14693_),
    .A2(_04182_),
    .Y(_04184_),
    .B1(net3856));
 sg13g2_a22oi_1 _26194_ (.Y(_04185_),
    .B1(_04183_),
    .B2(_04184_),
    .A2(_04181_),
    .A1(_04178_));
 sg13g2_xnor2_1 _26195_ (.Y(_04186_),
    .A(net3485),
    .B(_04185_));
 sg13g2_a21oi_1 _26196_ (.A1(_04172_),
    .A2(_04174_),
    .Y(_04187_),
    .B1(_04171_));
 sg13g2_xor2_1 _26197_ (.B(_04187_),
    .A(_04186_),
    .X(_04188_));
 sg13g2_o21ai_1 _26198_ (.B1(net3901),
    .Y(_04189_),
    .A1(net4365),
    .A2(_04185_));
 sg13g2_a21oi_1 _26199_ (.A1(net4365),
    .A2(_04188_),
    .Y(_04190_),
    .B1(_04189_));
 sg13g2_a21o_1 _26200_ (.A2(net3974),
    .A1(net2507),
    .B1(_04190_),
    .X(_00459_));
 sg13g2_a21oi_2 _26201_ (.B1(_14711_),
    .Y(_04191_),
    .A2(_04058_),
    .A1(_15023_));
 sg13g2_nor2_1 _26202_ (.A(_14976_),
    .B(_04191_),
    .Y(_04192_));
 sg13g2_xnor2_1 _26203_ (.Y(_04193_),
    .A(_14675_),
    .B(_04192_));
 sg13g2_a21oi_1 _26204_ (.A1(_15323_),
    .A2(_04062_),
    .Y(_04194_),
    .B1(_15320_));
 sg13g2_o21ai_1 _26205_ (.B1(_15319_),
    .Y(_04195_),
    .A1(_15198_),
    .A2(_04061_));
 sg13g2_nand2_1 _26206_ (.Y(_04196_),
    .A(_14675_),
    .B(_04195_));
 sg13g2_o21ai_1 _26207_ (.B1(net4698),
    .Y(_04197_),
    .A1(_14675_),
    .A2(_04195_));
 sg13g2_nand2b_1 _26208_ (.Y(_04198_),
    .B(_04196_),
    .A_N(_04197_));
 sg13g2_a21oi_1 _26209_ (.A1(net4580),
    .A2(\u_inv.d_next[184] ),
    .Y(_04199_),
    .B1(net3800));
 sg13g2_a22oi_1 _26210_ (.Y(_04200_),
    .B1(_04198_),
    .B2(_04199_),
    .A2(_04193_),
    .A1(net3800));
 sg13g2_and2_1 _26211_ (.A(net3443),
    .B(_04200_),
    .X(_04201_));
 sg13g2_xnor2_1 _26212_ (.Y(_04202_),
    .A(net3443),
    .B(_04200_));
 sg13g2_nand2_1 _26213_ (.Y(_04203_),
    .A(_04172_),
    .B(_04186_));
 sg13g2_nor2_1 _26214_ (.A(_04140_),
    .B(_04158_),
    .Y(_04204_));
 sg13g2_a221oi_1 _26215_ (.B2(_04110_),
    .C1(_04107_),
    .B1(_04142_),
    .A1(net3454),
    .Y(_04205_),
    .A2(_04125_));
 sg13g2_nor4_1 _26216_ (.A(_04140_),
    .B(_04158_),
    .C(_04203_),
    .D(_04205_),
    .Y(_04206_));
 sg13g2_o21ai_1 _26217_ (.B1(net3455),
    .Y(_04207_),
    .A1(_04169_),
    .A2(_04185_));
 sg13g2_o21ai_1 _26218_ (.B1(_04207_),
    .Y(_04208_),
    .A1(_04173_),
    .A2(_04203_));
 sg13g2_nor2_1 _26219_ (.A(_04206_),
    .B(_04208_),
    .Y(_04209_));
 sg13g2_nor4_1 _26220_ (.A(_04069_),
    .B(_04093_),
    .C(_04108_),
    .D(_04126_),
    .Y(_04210_));
 sg13g2_nand4_1 _26221_ (.B(_04186_),
    .C(_04204_),
    .A(_04172_),
    .Y(_04211_),
    .D(_04210_));
 sg13g2_o21ai_1 _26222_ (.B1(_04209_),
    .Y(_04212_),
    .A1(_04078_),
    .A2(_04211_));
 sg13g2_nor2b_1 _26223_ (.A(_04202_),
    .B_N(_04212_),
    .Y(_04213_));
 sg13g2_xor2_1 _26224_ (.B(_04212_),
    .A(_04202_),
    .X(_04214_));
 sg13g2_o21ai_1 _26225_ (.B1(net3901),
    .Y(_04215_),
    .A1(net4355),
    .A2(_04200_));
 sg13g2_a21oi_1 _26226_ (.A1(net4355),
    .A2(_04214_),
    .Y(_04216_),
    .B1(_04215_));
 sg13g2_a21o_1 _26227_ (.A2(net3974),
    .A1(net2908),
    .B1(_04216_),
    .X(_00460_));
 sg13g2_nand2_1 _26228_ (.Y(_04217_),
    .A(net1065),
    .B(net3974));
 sg13g2_nand2_1 _26229_ (.Y(_04218_),
    .A(_15192_),
    .B(_04195_));
 sg13g2_nand3_1 _26230_ (.B(_14674_),
    .C(_04196_),
    .A(_14673_),
    .Y(_04219_));
 sg13g2_nand4_1 _26231_ (.B(_15300_),
    .C(_04218_),
    .A(net4698),
    .Y(_04220_),
    .D(_04219_));
 sg13g2_a21oi_1 _26232_ (.A1(net4580),
    .A2(\u_inv.d_next[185] ),
    .Y(_04221_),
    .B1(net3800));
 sg13g2_o21ai_1 _26233_ (.B1(_14986_),
    .Y(_04222_),
    .A1(_14675_),
    .A2(_04192_));
 sg13g2_xnor2_1 _26234_ (.Y(_04223_),
    .A(_14673_),
    .B(_04222_));
 sg13g2_a22oi_1 _26235_ (.Y(_04224_),
    .B1(_04223_),
    .B2(net3800),
    .A2(_04221_),
    .A1(_04220_));
 sg13g2_and2_1 _26236_ (.A(net3443),
    .B(_04224_),
    .X(_04225_));
 sg13g2_nand2b_1 _26237_ (.Y(_04226_),
    .B(net3483),
    .A_N(_04224_));
 sg13g2_nand2b_1 _26238_ (.Y(_04227_),
    .B(_04226_),
    .A_N(_04225_));
 sg13g2_inv_1 _26239_ (.Y(_04228_),
    .A(_04227_));
 sg13g2_nor2_1 _26240_ (.A(_04201_),
    .B(_04213_),
    .Y(_04229_));
 sg13g2_o21ai_1 _26241_ (.B1(net4355),
    .Y(_04230_),
    .A1(_04228_),
    .A2(_04229_));
 sg13g2_a21oi_1 _26242_ (.A1(_04228_),
    .A2(_04229_),
    .Y(_04231_),
    .B1(_04230_));
 sg13g2_o21ai_1 _26243_ (.B1(net3902),
    .Y(_04232_),
    .A1(net4355),
    .A2(_04224_));
 sg13g2_o21ai_1 _26244_ (.B1(_04217_),
    .Y(_00461_),
    .A1(_04231_),
    .A2(_04232_));
 sg13g2_o21ai_1 _26245_ (.B1(_14676_),
    .Y(_04233_),
    .A1(_14976_),
    .A2(_04191_));
 sg13g2_a21oi_1 _26246_ (.A1(_14989_),
    .A2(_04233_),
    .Y(_04234_),
    .B1(_14678_));
 sg13g2_nand3_1 _26247_ (.B(_14989_),
    .C(_04233_),
    .A(_14678_),
    .Y(_04235_));
 sg13g2_nand2b_1 _26248_ (.Y(_04236_),
    .B(_04235_),
    .A_N(_04234_));
 sg13g2_a21oi_1 _26249_ (.A1(_15192_),
    .A2(_04195_),
    .Y(_04237_),
    .B1(_15301_));
 sg13g2_a21oi_1 _26250_ (.A1(_14679_),
    .A2(_04237_),
    .Y(_04238_),
    .B1(net4580));
 sg13g2_o21ai_1 _26251_ (.B1(_04238_),
    .Y(_04239_),
    .A1(_14679_),
    .A2(_04237_));
 sg13g2_a21oi_1 _26252_ (.A1(net4580),
    .A2(\u_inv.d_next[186] ),
    .Y(_04240_),
    .B1(net3800));
 sg13g2_a22oi_1 _26253_ (.Y(_04241_),
    .B1(_04239_),
    .B2(_04240_),
    .A2(_04236_),
    .A1(net3800));
 sg13g2_nand2_1 _26254_ (.Y(_04242_),
    .A(net3443),
    .B(_04241_));
 sg13g2_xnor2_1 _26255_ (.Y(_04243_),
    .A(net3443),
    .B(_04241_));
 sg13g2_nor2_1 _26256_ (.A(_04201_),
    .B(_04225_),
    .Y(_04244_));
 sg13g2_or2_1 _26257_ (.X(_04245_),
    .B(_04225_),
    .A(_04201_));
 sg13g2_o21ai_1 _26258_ (.B1(_04226_),
    .Y(_04246_),
    .A1(_04213_),
    .A2(_04245_));
 sg13g2_xnor2_1 _26259_ (.Y(_04247_),
    .A(_04243_),
    .B(_04246_));
 sg13g2_a21oi_1 _26260_ (.A1(net4355),
    .A2(_04247_),
    .Y(_04248_),
    .B1(net4236));
 sg13g2_o21ai_1 _26261_ (.B1(_04248_),
    .Y(_04249_),
    .A1(net4355),
    .A2(_04241_));
 sg13g2_o21ai_1 _26262_ (.B1(_04249_),
    .Y(_00462_),
    .A1(_10591_),
    .A2(net4030));
 sg13g2_a21oi_1 _26263_ (.A1(net4582),
    .A2(\u_inv.d_next[187] ),
    .Y(_04250_),
    .B1(net3799));
 sg13g2_o21ai_1 _26264_ (.B1(_14677_),
    .Y(_04251_),
    .A1(_14679_),
    .A2(_04237_));
 sg13g2_xnor2_1 _26265_ (.Y(_04252_),
    .A(_14681_),
    .B(_04251_));
 sg13g2_o21ai_1 _26266_ (.B1(_04250_),
    .Y(_04253_),
    .A1(net4582),
    .A2(_04252_));
 sg13g2_o21ai_1 _26267_ (.B1(_14681_),
    .Y(_04254_),
    .A1(_14990_),
    .A2(_04234_));
 sg13g2_or3_1 _26268_ (.A(_14681_),
    .B(_14990_),
    .C(_04234_),
    .X(_04255_));
 sg13g2_nand3_1 _26269_ (.B(_04254_),
    .C(_04255_),
    .A(net3800),
    .Y(_04256_));
 sg13g2_nand3_1 _26270_ (.B(_04253_),
    .C(_04256_),
    .A(net3443),
    .Y(_04257_));
 sg13g2_a21o_1 _26271_ (.A2(_04256_),
    .A1(_04253_),
    .B1(net3443),
    .X(_04258_));
 sg13g2_nand2_1 _26272_ (.Y(_04259_),
    .A(_04257_),
    .B(_04258_));
 sg13g2_o21ai_1 _26273_ (.B1(_04242_),
    .Y(_04260_),
    .A1(_04243_),
    .A2(_04246_));
 sg13g2_xnor2_1 _26274_ (.Y(_04261_),
    .A(_04259_),
    .B(_04260_));
 sg13g2_a21oi_1 _26275_ (.A1(_04253_),
    .A2(_04256_),
    .Y(_04262_),
    .B1(net4355));
 sg13g2_nor2_1 _26276_ (.A(net4236),
    .B(_04262_),
    .Y(_04263_));
 sg13g2_o21ai_1 _26277_ (.B1(_04263_),
    .Y(_04264_),
    .A1(net4297),
    .A2(_04261_));
 sg13g2_o21ai_1 _26278_ (.B1(_04264_),
    .Y(_00463_),
    .A1(_10590_),
    .A2(net4030));
 sg13g2_o21ai_1 _26279_ (.B1(_14685_),
    .Y(_04265_),
    .A1(_14976_),
    .A2(_04191_));
 sg13g2_a21oi_1 _26280_ (.A1(_14992_),
    .A2(_04265_),
    .Y(_04266_),
    .B1(_14668_));
 sg13g2_nand3_1 _26281_ (.B(_14992_),
    .C(_04265_),
    .A(_14668_),
    .Y(_04267_));
 sg13g2_nand2b_1 _26282_ (.Y(_04268_),
    .B(_04267_),
    .A_N(_04266_));
 sg13g2_o21ai_1 _26283_ (.B1(_15303_),
    .Y(_04269_),
    .A1(_15193_),
    .A2(_04194_));
 sg13g2_o21ai_1 _26284_ (.B1(net4690),
    .Y(_04270_),
    .A1(_14668_),
    .A2(_04269_));
 sg13g2_a21o_1 _26285_ (.A2(_04269_),
    .A1(_14668_),
    .B1(_04270_),
    .X(_04271_));
 sg13g2_a21oi_1 _26286_ (.A1(net4580),
    .A2(\u_inv.d_next[188] ),
    .Y(_04272_),
    .B1(net3800));
 sg13g2_a22oi_1 _26287_ (.Y(_04273_),
    .B1(_04271_),
    .B2(_04272_),
    .A2(_04268_),
    .A1(net3796));
 sg13g2_and2_1 _26288_ (.A(net3444),
    .B(_04273_),
    .X(_04274_));
 sg13g2_xnor2_1 _26289_ (.Y(_04275_),
    .A(net3443),
    .B(_04273_));
 sg13g2_nand3b_1 _26290_ (.B(_04257_),
    .C(_04258_),
    .Y(_04276_),
    .A_N(_04243_));
 sg13g2_and2_1 _26291_ (.A(_04242_),
    .B(_04257_),
    .X(_04277_));
 sg13g2_o21ai_1 _26292_ (.B1(_04277_),
    .Y(_04278_),
    .A1(_04244_),
    .A2(_04276_));
 sg13g2_or3_1 _26293_ (.A(_04202_),
    .B(_04227_),
    .C(_04276_),
    .X(_04279_));
 sg13g2_inv_1 _26294_ (.Y(_04280_),
    .A(_04279_));
 sg13g2_a21oi_1 _26295_ (.A1(_04212_),
    .A2(_04280_),
    .Y(_04281_),
    .B1(_04278_));
 sg13g2_nor2_1 _26296_ (.A(_04275_),
    .B(_04281_),
    .Y(_04282_));
 sg13g2_xnor2_1 _26297_ (.Y(_04283_),
    .A(_04275_),
    .B(_04281_));
 sg13g2_o21ai_1 _26298_ (.B1(net3902),
    .Y(_04284_),
    .A1(net4355),
    .A2(_04273_));
 sg13g2_a21oi_1 _26299_ (.A1(net4357),
    .A2(_04283_),
    .Y(_04285_),
    .B1(_04284_));
 sg13g2_a21o_1 _26300_ (.A2(net3975),
    .A1(net3138),
    .B1(_04285_),
    .X(_00464_));
 sg13g2_a21oi_1 _26301_ (.A1(net4576),
    .A2(\u_inv.d_next[189] ),
    .Y(_04286_),
    .B1(net3795));
 sg13g2_a21oi_1 _26302_ (.A1(_14668_),
    .A2(_04269_),
    .Y(_04287_),
    .B1(_14667_));
 sg13g2_xnor2_1 _26303_ (.Y(_04288_),
    .A(_14666_),
    .B(_04287_));
 sg13g2_nand2_1 _26304_ (.Y(_04289_),
    .A(net4690),
    .B(_04288_));
 sg13g2_o21ai_1 _26305_ (.B1(_14666_),
    .Y(_04290_),
    .A1(_14978_),
    .A2(_04266_));
 sg13g2_nor3_1 _26306_ (.A(_14666_),
    .B(_14978_),
    .C(_04266_),
    .Y(_04291_));
 sg13g2_nor2_1 _26307_ (.A(net3857),
    .B(_04291_),
    .Y(_04292_));
 sg13g2_a22oi_1 _26308_ (.Y(_04293_),
    .B1(_04290_),
    .B2(_04292_),
    .A2(_04289_),
    .A1(_04286_));
 sg13g2_nor2_1 _26309_ (.A(net3444),
    .B(_04293_),
    .Y(_04294_));
 sg13g2_xnor2_1 _26310_ (.Y(_04295_),
    .A(net3444),
    .B(_04293_));
 sg13g2_nor2_1 _26311_ (.A(_04274_),
    .B(_04282_),
    .Y(_04296_));
 sg13g2_xnor2_1 _26312_ (.Y(_04297_),
    .A(_04295_),
    .B(_04296_));
 sg13g2_o21ai_1 _26313_ (.B1(net3901),
    .Y(_04298_),
    .A1(net4357),
    .A2(_04293_));
 sg13g2_a21oi_1 _26314_ (.A1(net4357),
    .A2(_04297_),
    .Y(_04299_),
    .B1(_04298_));
 sg13g2_a21o_1 _26315_ (.A2(net3974),
    .A1(net2823),
    .B1(_04299_),
    .X(_00465_));
 sg13g2_a21o_1 _26316_ (.A2(_04265_),
    .A1(_14992_),
    .B1(_14670_),
    .X(_04300_));
 sg13g2_a21oi_1 _26317_ (.A1(_14981_),
    .A2(_04300_),
    .Y(_04301_),
    .B1(_14664_));
 sg13g2_nand3_1 _26318_ (.B(_14981_),
    .C(_04300_),
    .A(_14664_),
    .Y(_04302_));
 sg13g2_nand2b_1 _26319_ (.Y(_04303_),
    .B(_04302_),
    .A_N(_04301_));
 sg13g2_a21oi_1 _26320_ (.A1(_15189_),
    .A2(_04269_),
    .Y(_04304_),
    .B1(_15306_));
 sg13g2_xnor2_1 _26321_ (.Y(_04305_),
    .A(_14664_),
    .B(_04304_));
 sg13g2_nand2_1 _26322_ (.Y(_04306_),
    .A(net4691),
    .B(_04305_));
 sg13g2_a21oi_1 _26323_ (.A1(net4576),
    .A2(\u_inv.d_next[190] ),
    .Y(_04307_),
    .B1(net3795));
 sg13g2_a22oi_1 _26324_ (.Y(_04308_),
    .B1(_04306_),
    .B2(_04307_),
    .A2(_04303_),
    .A1(net3795));
 sg13g2_nand2_1 _26325_ (.Y(_04309_),
    .A(net3445),
    .B(_04308_));
 sg13g2_xnor2_1 _26326_ (.Y(_04310_),
    .A(net3483),
    .B(_04308_));
 sg13g2_a21oi_1 _26327_ (.A1(net3444),
    .A2(_04293_),
    .Y(_04311_),
    .B1(_04274_));
 sg13g2_o21ai_1 _26328_ (.B1(_04311_),
    .Y(_04312_),
    .A1(_04275_),
    .A2(_04281_));
 sg13g2_nor2b_1 _26329_ (.A(_04294_),
    .B_N(_04312_),
    .Y(_04313_));
 sg13g2_nand3b_1 _26330_ (.B(_04310_),
    .C(_04312_),
    .Y(_04314_),
    .A_N(_04294_));
 sg13g2_xnor2_1 _26331_ (.Y(_04315_),
    .A(_04310_),
    .B(_04313_));
 sg13g2_a21oi_1 _26332_ (.A1(net4356),
    .A2(_04315_),
    .Y(_04316_),
    .B1(net4237));
 sg13g2_o21ai_1 _26333_ (.B1(_04316_),
    .Y(_04317_),
    .A1(net4356),
    .A2(_04308_));
 sg13g2_o21ai_1 _26334_ (.B1(_04317_),
    .Y(_00466_),
    .A1(_10589_),
    .A2(net4034));
 sg13g2_a21oi_1 _26335_ (.A1(net4576),
    .A2(\u_inv.d_next[191] ),
    .Y(_04318_),
    .B1(net3795));
 sg13g2_o21ai_1 _26336_ (.B1(_14662_),
    .Y(_04319_),
    .A1(_14663_),
    .A2(_04304_));
 sg13g2_xnor2_1 _26337_ (.Y(_04320_),
    .A(_14661_),
    .B(_04319_));
 sg13g2_o21ai_1 _26338_ (.B1(_04318_),
    .Y(_04321_),
    .A1(net4576),
    .A2(_04320_));
 sg13g2_o21ai_1 _26339_ (.B1(_14661_),
    .Y(_04322_),
    .A1(_14982_),
    .A2(_04301_));
 sg13g2_or3_1 _26340_ (.A(_14661_),
    .B(_14982_),
    .C(_04301_),
    .X(_04323_));
 sg13g2_nand3_1 _26341_ (.B(_04322_),
    .C(_04323_),
    .A(net3797),
    .Y(_04324_));
 sg13g2_and2_1 _26342_ (.A(_04321_),
    .B(_04324_),
    .X(_04325_));
 sg13g2_nand3_1 _26343_ (.B(_04321_),
    .C(_04324_),
    .A(net3445),
    .Y(_04326_));
 sg13g2_a21o_1 _26344_ (.A2(_04324_),
    .A1(_04321_),
    .B1(net3445),
    .X(_04327_));
 sg13g2_and2_1 _26345_ (.A(_04326_),
    .B(_04327_),
    .X(_04328_));
 sg13g2_nand2_1 _26346_ (.Y(_04329_),
    .A(_04309_),
    .B(_04314_));
 sg13g2_xnor2_1 _26347_ (.Y(_04330_),
    .A(_04328_),
    .B(_04329_));
 sg13g2_o21ai_1 _26348_ (.B1(net3900),
    .Y(_04331_),
    .A1(net4356),
    .A2(_04325_));
 sg13g2_a21oi_1 _26349_ (.A1(net4356),
    .A2(_04330_),
    .Y(_04332_),
    .B1(_04331_));
 sg13g2_a21o_1 _26350_ (.A2(net3969),
    .A1(net3007),
    .B1(_04332_),
    .X(_00467_));
 sg13g2_nor2_1 _26351_ (.A(_14901_),
    .B(_15026_),
    .Y(_04333_));
 sg13g2_nand2_1 _26352_ (.Y(_04334_),
    .A(_14902_),
    .B(_15025_));
 sg13g2_xnor2_1 _26353_ (.Y(_04335_),
    .A(_13772_),
    .B(_04334_));
 sg13g2_a21oi_1 _26354_ (.A1(_13772_),
    .A2(_15637_),
    .Y(_04336_),
    .B1(net4560));
 sg13g2_o21ai_1 _26355_ (.B1(_04336_),
    .Y(_04337_),
    .A1(_13772_),
    .A2(_15637_));
 sg13g2_a21oi_1 _26356_ (.A1(net4560),
    .A2(\u_inv.d_next[192] ),
    .Y(_04338_),
    .B1(net3778));
 sg13g2_a22oi_1 _26357_ (.Y(_04339_),
    .B1(_04337_),
    .B2(_04338_),
    .A2(_04335_),
    .A1(net3778));
 sg13g2_nand2_1 _26358_ (.Y(_04340_),
    .A(net3425),
    .B(_04339_));
 sg13g2_xnor2_1 _26359_ (.Y(_04341_),
    .A(net3426),
    .B(_04339_));
 sg13g2_nand3_1 _26360_ (.B(_04326_),
    .C(_04327_),
    .A(_04310_),
    .Y(_04342_));
 sg13g2_nor2_1 _26361_ (.A(_04275_),
    .B(_04295_),
    .Y(_04343_));
 sg13g2_or2_1 _26362_ (.X(_04344_),
    .B(_04295_),
    .A(_04275_));
 sg13g2_nand4_1 _26363_ (.B(_04310_),
    .C(_04328_),
    .A(_04280_),
    .Y(_04345_),
    .D(_04343_));
 sg13g2_nor4_2 _26364_ (.A(_04211_),
    .B(_04279_),
    .C(_04342_),
    .Y(_04346_),
    .D(_04344_));
 sg13g2_nand2_1 _26365_ (.Y(_04347_),
    .A(_04077_),
    .B(_04346_));
 sg13g2_nand3b_1 _26366_ (.B(_04077_),
    .C(_04346_),
    .Y(_04348_),
    .A_N(_03809_));
 sg13g2_a21oi_1 _26367_ (.A1(_03259_),
    .A2(_03265_),
    .Y(_04349_),
    .B1(_04348_));
 sg13g2_nor2_1 _26368_ (.A(_03808_),
    .B(_04347_),
    .Y(_04350_));
 sg13g2_o21ai_1 _26369_ (.B1(_04346_),
    .Y(_04351_),
    .A1(_04072_),
    .A2(_04076_));
 sg13g2_nand4_1 _26370_ (.B(_04310_),
    .C(_04328_),
    .A(_04278_),
    .Y(_04352_),
    .D(_04343_));
 sg13g2_or2_1 _26371_ (.X(_04353_),
    .B(_04342_),
    .A(_04311_));
 sg13g2_nand4_1 _26372_ (.B(_04326_),
    .C(_04352_),
    .A(_04309_),
    .Y(_04354_),
    .D(_04353_));
 sg13g2_o21ai_1 _26373_ (.B1(_04351_),
    .Y(_04355_),
    .A1(_04209_),
    .A2(_04345_));
 sg13g2_or4_1 _26374_ (.A(_04349_),
    .B(_04350_),
    .C(_04354_),
    .D(_04355_),
    .X(_04356_));
 sg13g2_nand2b_1 _26375_ (.Y(_04357_),
    .B(_04356_),
    .A_N(_04341_));
 sg13g2_xor2_1 _26376_ (.B(_04356_),
    .A(_04341_),
    .X(_04358_));
 sg13g2_o21ai_1 _26377_ (.B1(net3891),
    .Y(_04359_),
    .A1(net4336),
    .A2(_04339_));
 sg13g2_a21oi_2 _26378_ (.B1(_04359_),
    .Y(_04360_),
    .A2(_04358_),
    .A1(net4336));
 sg13g2_a21o_1 _26379_ (.A2(net3969),
    .A1(net3167),
    .B1(_04360_),
    .X(_00468_));
 sg13g2_o21ai_1 _26380_ (.B1(_13771_),
    .Y(_04361_),
    .A1(_13772_),
    .A2(_15637_));
 sg13g2_a21oi_1 _26381_ (.A1(_13770_),
    .A2(_04361_),
    .Y(_04362_),
    .B1(net4560));
 sg13g2_o21ai_1 _26382_ (.B1(_04362_),
    .Y(_04363_),
    .A1(_13770_),
    .A2(_04361_));
 sg13g2_a21oi_1 _26383_ (.A1(net4560),
    .A2(\u_inv.d_next[193] ),
    .Y(_04364_),
    .B1(net3778));
 sg13g2_a21oi_1 _26384_ (.A1(_13772_),
    .A2(_04334_),
    .Y(_04365_),
    .B1(_13895_));
 sg13g2_o21ai_1 _26385_ (.B1(net3778),
    .Y(_04366_),
    .A1(_13769_),
    .A2(_04365_));
 sg13g2_a21oi_1 _26386_ (.A1(_13769_),
    .A2(_04365_),
    .Y(_04367_),
    .B1(_04366_));
 sg13g2_a21oi_2 _26387_ (.B1(_04367_),
    .Y(_04368_),
    .A2(_04364_),
    .A1(_04363_));
 sg13g2_nand2_1 _26388_ (.Y(_04369_),
    .A(net3425),
    .B(_04368_));
 sg13g2_xnor2_1 _26389_ (.Y(_04370_),
    .A(net3425),
    .B(_04368_));
 sg13g2_nand2_1 _26390_ (.Y(_04371_),
    .A(_04340_),
    .B(_04357_));
 sg13g2_xor2_1 _26391_ (.B(_04371_),
    .A(_04370_),
    .X(_04372_));
 sg13g2_o21ai_1 _26392_ (.B1(net3891),
    .Y(_04373_),
    .A1(net4337),
    .A2(_04368_));
 sg13g2_a21oi_1 _26393_ (.A1(net4336),
    .A2(_04372_),
    .Y(_04374_),
    .B1(_04373_));
 sg13g2_a21o_1 _26394_ (.A2(net3953),
    .A1(net2627),
    .B1(_04374_),
    .X(_00469_));
 sg13g2_o21ai_1 _26395_ (.B1(net3425),
    .Y(_04375_),
    .A1(_04339_),
    .A2(_04368_));
 sg13g2_nand2_1 _26396_ (.Y(_04376_),
    .A(_04340_),
    .B(_04369_));
 sg13g2_o21ai_1 _26397_ (.B1(_04375_),
    .Y(_04377_),
    .A1(_04357_),
    .A2(_04370_));
 sg13g2_a21oi_1 _26398_ (.A1(_14902_),
    .A2(_15025_),
    .Y(_04378_),
    .B1(_13773_));
 sg13g2_or2_1 _26399_ (.X(_04379_),
    .B(_04378_),
    .A(_13897_));
 sg13g2_xnor2_1 _26400_ (.Y(_04380_),
    .A(_13764_),
    .B(_04379_));
 sg13g2_a21oi_1 _26401_ (.A1(_13770_),
    .A2(_04361_),
    .Y(_04381_),
    .B1(_15106_));
 sg13g2_xor2_1 _26402_ (.B(_04381_),
    .A(_13764_),
    .X(_04382_));
 sg13g2_o21ai_1 _26403_ (.B1(net3849),
    .Y(_04383_),
    .A1(net4680),
    .A2(_10587_));
 sg13g2_a21oi_1 _26404_ (.A1(net4680),
    .A2(_04382_),
    .Y(_04384_),
    .B1(_04383_));
 sg13g2_a21oi_1 _26405_ (.A1(net3778),
    .A2(_04380_),
    .Y(_04385_),
    .B1(_04384_));
 sg13g2_and2_1 _26406_ (.A(net3427),
    .B(_04385_),
    .X(_04386_));
 sg13g2_xnor2_1 _26407_ (.Y(_04387_),
    .A(net3427),
    .B(_04385_));
 sg13g2_nor2b_1 _26408_ (.A(_04387_),
    .B_N(_04377_),
    .Y(_04388_));
 sg13g2_xor2_1 _26409_ (.B(_04387_),
    .A(_04377_),
    .X(_04389_));
 sg13g2_o21ai_1 _26410_ (.B1(net3890),
    .Y(_04390_),
    .A1(net4335),
    .A2(_04385_));
 sg13g2_a21oi_1 _26411_ (.A1(net4335),
    .A2(_04389_),
    .Y(_04391_),
    .B1(_04390_));
 sg13g2_a21o_1 _26412_ (.A2(net3953),
    .A1(net2745),
    .B1(_04391_),
    .X(_00470_));
 sg13g2_nor2_1 _26413_ (.A(_04386_),
    .B(_04388_),
    .Y(_04392_));
 sg13g2_a21oi_1 _26414_ (.A1(net4559),
    .A2(\u_inv.d_next[195] ),
    .Y(_04393_),
    .B1(net3777));
 sg13g2_o21ai_1 _26415_ (.B1(_13763_),
    .Y(_04394_),
    .A1(_13764_),
    .A2(_04381_));
 sg13g2_xor2_1 _26416_ (.B(_04394_),
    .A(_13762_),
    .X(_04395_));
 sg13g2_o21ai_1 _26417_ (.B1(_04393_),
    .Y(_04396_),
    .A1(net4559),
    .A2(_04395_));
 sg13g2_a21oi_1 _26418_ (.A1(_13764_),
    .A2(_04379_),
    .Y(_04397_),
    .B1(_13898_));
 sg13g2_a21oi_1 _26419_ (.A1(_13762_),
    .A2(_04397_),
    .Y(_04398_),
    .B1(net3849));
 sg13g2_o21ai_1 _26420_ (.B1(_04398_),
    .Y(_04399_),
    .A1(_13762_),
    .A2(_04397_));
 sg13g2_and3_2 _26421_ (.X(_04400_),
    .A(net3427),
    .B(_04396_),
    .C(_04399_));
 sg13g2_a21oi_1 _26422_ (.A1(_04396_),
    .A2(_04399_),
    .Y(_04401_),
    .B1(net3427));
 sg13g2_nor2_1 _26423_ (.A(_04400_),
    .B(_04401_),
    .Y(_04402_));
 sg13g2_xnor2_1 _26424_ (.Y(_04403_),
    .A(_04392_),
    .B(_04402_));
 sg13g2_a21oi_1 _26425_ (.A1(_04396_),
    .A2(_04399_),
    .Y(_04404_),
    .B1(net4340));
 sg13g2_nor2_1 _26426_ (.A(net4237),
    .B(_04404_),
    .Y(_04405_));
 sg13g2_o21ai_1 _26427_ (.B1(_04405_),
    .Y(_04406_),
    .A1(net4295),
    .A2(_04403_));
 sg13g2_o21ai_1 _26428_ (.B1(_04406_),
    .Y(_00471_),
    .A1(_10587_),
    .A2(net4029));
 sg13g2_o21ai_1 _26429_ (.B1(_13765_),
    .Y(_04407_),
    .A1(_13897_),
    .A2(_04378_));
 sg13g2_a21oi_1 _26430_ (.A1(_13899_),
    .A2(_04407_),
    .Y(_04408_),
    .B1(_13756_));
 sg13g2_nand3_1 _26431_ (.B(_13899_),
    .C(_04407_),
    .A(_13756_),
    .Y(_04409_));
 sg13g2_nand2b_1 _26432_ (.Y(_04410_),
    .B(_04409_),
    .A_N(_04408_));
 sg13g2_a21oi_2 _26433_ (.B1(_15111_),
    .Y(_04411_),
    .A2(_15638_),
    .A1(_15184_));
 sg13g2_a21oi_1 _26434_ (.A1(_13757_),
    .A2(_04411_),
    .Y(_04412_),
    .B1(net4559));
 sg13g2_o21ai_1 _26435_ (.B1(_04412_),
    .Y(_04413_),
    .A1(_13757_),
    .A2(_04411_));
 sg13g2_a21oi_1 _26436_ (.A1(net4559),
    .A2(\u_inv.d_next[196] ),
    .Y(_04414_),
    .B1(net3777));
 sg13g2_a22oi_1 _26437_ (.Y(_04415_),
    .B1(_04413_),
    .B2(_04414_),
    .A2(_04410_),
    .A1(net3777));
 sg13g2_and2_1 _26438_ (.A(net3427),
    .B(_04415_),
    .X(_04416_));
 sg13g2_xnor2_1 _26439_ (.Y(_04417_),
    .A(net3478),
    .B(_04415_));
 sg13g2_or2_1 _26440_ (.X(_04418_),
    .B(_04400_),
    .A(_04386_));
 sg13g2_nor3_2 _26441_ (.A(_04387_),
    .B(_04400_),
    .C(_04401_),
    .Y(_04419_));
 sg13g2_a21o_2 _26442_ (.A2(_04419_),
    .A1(_04377_),
    .B1(_04418_),
    .X(_04420_));
 sg13g2_xnor2_1 _26443_ (.Y(_04421_),
    .A(_04417_),
    .B(_04420_));
 sg13g2_a21oi_1 _26444_ (.A1(net4340),
    .A2(_04421_),
    .Y(_04422_),
    .B1(net4237));
 sg13g2_o21ai_1 _26445_ (.B1(_04422_),
    .Y(_04423_),
    .A1(net4340),
    .A2(_04415_));
 sg13g2_o21ai_1 _26446_ (.B1(_04423_),
    .Y(_00472_),
    .A1(_10586_),
    .A2(net4029));
 sg13g2_a21oi_1 _26447_ (.A1(net4559),
    .A2(\u_inv.d_next[197] ),
    .Y(_04424_),
    .B1(net3777));
 sg13g2_o21ai_1 _26448_ (.B1(_13755_),
    .Y(_04425_),
    .A1(_13757_),
    .A2(_04411_));
 sg13g2_xnor2_1 _26449_ (.Y(_04426_),
    .A(_13753_),
    .B(_04425_));
 sg13g2_o21ai_1 _26450_ (.B1(_04424_),
    .Y(_04427_),
    .A1(net4559),
    .A2(_04426_));
 sg13g2_o21ai_1 _26451_ (.B1(_13753_),
    .Y(_04428_),
    .A1(_13904_),
    .A2(_04408_));
 sg13g2_or3_1 _26452_ (.A(_13753_),
    .B(_13904_),
    .C(_04408_),
    .X(_04429_));
 sg13g2_nand3_1 _26453_ (.B(_04428_),
    .C(_04429_),
    .A(net3777),
    .Y(_04430_));
 sg13g2_and2_1 _26454_ (.A(_04427_),
    .B(_04430_),
    .X(_04431_));
 sg13g2_nand3_1 _26455_ (.B(_04427_),
    .C(_04430_),
    .A(net3427),
    .Y(_04432_));
 sg13g2_a21o_1 _26456_ (.A2(_04430_),
    .A1(_04427_),
    .B1(net3427),
    .X(_04433_));
 sg13g2_nand2_1 _26457_ (.Y(_04434_),
    .A(_04432_),
    .B(_04433_));
 sg13g2_a21oi_1 _26458_ (.A1(_04417_),
    .A2(_04420_),
    .Y(_04435_),
    .B1(_04416_));
 sg13g2_xnor2_1 _26459_ (.Y(_04436_),
    .A(_04434_),
    .B(_04435_));
 sg13g2_o21ai_1 _26460_ (.B1(net3890),
    .Y(_04437_),
    .A1(net4335),
    .A2(_04431_));
 sg13g2_a21oi_1 _26461_ (.A1(net4335),
    .A2(_04436_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_a21o_1 _26462_ (.A2(net3953),
    .A1(net2766),
    .B1(_04438_),
    .X(_00473_));
 sg13g2_a21o_1 _26463_ (.A2(_04407_),
    .A1(_13899_),
    .B1(_13758_),
    .X(_04439_));
 sg13g2_a21oi_1 _26464_ (.A1(_13905_),
    .A2(_04439_),
    .Y(_04440_),
    .B1(_13749_));
 sg13g2_nand3_1 _26465_ (.B(_13905_),
    .C(_04439_),
    .A(_13749_),
    .Y(_04441_));
 sg13g2_nand2b_1 _26466_ (.Y(_04442_),
    .B(_04441_),
    .A_N(_04440_));
 sg13g2_nor2b_1 _26467_ (.A(_04411_),
    .B_N(_15104_),
    .Y(_04443_));
 sg13g2_nor2_1 _26468_ (.A(_15113_),
    .B(_04443_),
    .Y(_04444_));
 sg13g2_a21oi_1 _26469_ (.A1(_13750_),
    .A2(_04444_),
    .Y(_04445_),
    .B1(net4559));
 sg13g2_o21ai_1 _26470_ (.B1(_04445_),
    .Y(_04446_),
    .A1(_13750_),
    .A2(_04444_));
 sg13g2_a21oi_1 _26471_ (.A1(net4559),
    .A2(\u_inv.d_next[198] ),
    .Y(_04447_),
    .B1(net3777));
 sg13g2_a22oi_1 _26472_ (.Y(_04448_),
    .B1(_04446_),
    .B2(_04447_),
    .A2(_04442_),
    .A1(net3777));
 sg13g2_and2_1 _26473_ (.A(net3425),
    .B(_04448_),
    .X(_04449_));
 sg13g2_nand2b_1 _26474_ (.Y(_04450_),
    .B(net3477),
    .A_N(_04448_));
 sg13g2_xnor2_1 _26475_ (.Y(_04451_),
    .A(net3425),
    .B(_04448_));
 sg13g2_nand2b_2 _26476_ (.Y(_04452_),
    .B(_04432_),
    .A_N(_04416_));
 sg13g2_a21o_1 _26477_ (.A2(_04420_),
    .A1(_04417_),
    .B1(_04452_),
    .X(_04453_));
 sg13g2_and2_1 _26478_ (.A(_04433_),
    .B(_04453_),
    .X(_04454_));
 sg13g2_xor2_1 _26479_ (.B(_04454_),
    .A(_04451_),
    .X(_04455_));
 sg13g2_o21ai_1 _26480_ (.B1(net3890),
    .Y(_04456_),
    .A1(net4335),
    .A2(_04448_));
 sg13g2_a21oi_1 _26481_ (.A1(net4335),
    .A2(_04455_),
    .Y(_04457_),
    .B1(_04456_));
 sg13g2_a21o_1 _26482_ (.A2(net3953),
    .A1(net3205),
    .B1(_04457_),
    .X(_00474_));
 sg13g2_nand2_1 _26483_ (.Y(_04458_),
    .A(net2721),
    .B(net3953));
 sg13g2_a21oi_1 _26484_ (.A1(net4561),
    .A2(\u_inv.d_next[199] ),
    .Y(_04459_),
    .B1(net3779));
 sg13g2_o21ai_1 _26485_ (.B1(_13747_),
    .Y(_04460_),
    .A1(_13750_),
    .A2(_04444_));
 sg13g2_xnor2_1 _26486_ (.Y(_04461_),
    .A(_13746_),
    .B(_04460_));
 sg13g2_o21ai_1 _26487_ (.B1(_04459_),
    .Y(_04462_),
    .A1(net4561),
    .A2(_04461_));
 sg13g2_o21ai_1 _26488_ (.B1(_13746_),
    .Y(_04463_),
    .A1(_13901_),
    .A2(_04440_));
 sg13g2_or3_1 _26489_ (.A(_13746_),
    .B(_13901_),
    .C(_04440_),
    .X(_04464_));
 sg13g2_nand3_1 _26490_ (.B(_04463_),
    .C(_04464_),
    .A(net3777),
    .Y(_04465_));
 sg13g2_and2_1 _26491_ (.A(_04462_),
    .B(_04465_),
    .X(_04466_));
 sg13g2_and3_2 _26492_ (.X(_04467_),
    .A(net3426),
    .B(_04462_),
    .C(_04465_));
 sg13g2_a21oi_1 _26493_ (.A1(_04462_),
    .A2(_04465_),
    .Y(_04468_),
    .B1(net3426));
 sg13g2_nor2_1 _26494_ (.A(_04467_),
    .B(_04468_),
    .Y(_04469_));
 sg13g2_a21oi_1 _26495_ (.A1(_04450_),
    .A2(_04454_),
    .Y(_04470_),
    .B1(_04449_));
 sg13g2_o21ai_1 _26496_ (.B1(net4335),
    .Y(_04471_),
    .A1(_04469_),
    .A2(_04470_));
 sg13g2_a21oi_1 _26497_ (.A1(_04469_),
    .A2(_04470_),
    .Y(_04472_),
    .B1(_04471_));
 sg13g2_o21ai_1 _26498_ (.B1(net3890),
    .Y(_04473_),
    .A1(net4335),
    .A2(_04466_));
 sg13g2_o21ai_1 _26499_ (.B1(_04458_),
    .Y(_00475_),
    .A1(_04472_),
    .A2(_04473_));
 sg13g2_a21o_1 _26500_ (.A2(_15025_),
    .A1(_14902_),
    .B1(_13774_),
    .X(_04474_));
 sg13g2_nand2_1 _26501_ (.Y(_04475_),
    .A(_13907_),
    .B(_04474_));
 sg13g2_xnor2_1 _26502_ (.Y(_04476_),
    .A(_13731_),
    .B(_04475_));
 sg13g2_a21oi_2 _26503_ (.B1(_15117_),
    .Y(_04477_),
    .A2(_15638_),
    .A1(_15185_));
 sg13g2_a21oi_1 _26504_ (.A1(_13731_),
    .A2(_04477_),
    .Y(_04478_),
    .B1(net4550));
 sg13g2_o21ai_1 _26505_ (.B1(_04478_),
    .Y(_04479_),
    .A1(_13731_),
    .A2(_04477_));
 sg13g2_a21oi_1 _26506_ (.A1(net4561),
    .A2(\u_inv.d_next[200] ),
    .Y(_04480_),
    .B1(net3779));
 sg13g2_a22oi_1 _26507_ (.Y(_04481_),
    .B1(_04479_),
    .B2(_04480_),
    .A2(_04476_),
    .A1(net3779));
 sg13g2_and2_1 _26508_ (.A(net3424),
    .B(_04481_),
    .X(_04482_));
 sg13g2_xnor2_1 _26509_ (.Y(_04483_),
    .A(net3424),
    .B(_04481_));
 sg13g2_nor3_1 _26510_ (.A(_04451_),
    .B(_04467_),
    .C(_04468_),
    .Y(_04484_));
 sg13g2_nand3_1 _26511_ (.B(_04432_),
    .C(_04433_),
    .A(_04417_),
    .Y(_04485_));
 sg13g2_nor4_1 _26512_ (.A(_04451_),
    .B(_04467_),
    .C(_04468_),
    .D(_04485_),
    .Y(_04486_));
 sg13g2_a21o_1 _26513_ (.A2(_04419_),
    .A1(_04376_),
    .B1(_04418_),
    .X(_04487_));
 sg13g2_or2_1 _26514_ (.X(_04488_),
    .B(_04467_),
    .A(_04449_));
 sg13g2_a21o_1 _26515_ (.A2(_04484_),
    .A1(_04452_),
    .B1(_04488_),
    .X(_04489_));
 sg13g2_a221oi_1 _26516_ (.B2(_04487_),
    .C1(_04488_),
    .B1(_04486_),
    .A1(_04452_),
    .Y(_04490_),
    .A2(_04484_));
 sg13g2_nor2_1 _26517_ (.A(_04341_),
    .B(_04370_),
    .Y(_04491_));
 sg13g2_and3_1 _26518_ (.X(_04492_),
    .A(_04419_),
    .B(_04486_),
    .C(_04491_));
 sg13g2_a221oi_1 _26519_ (.B2(_04356_),
    .C1(_04489_),
    .B1(_04492_),
    .A1(_04486_),
    .Y(_04493_),
    .A2(_04487_));
 sg13g2_nor2_1 _26520_ (.A(_04483_),
    .B(_04493_),
    .Y(_04494_));
 sg13g2_xnor2_1 _26521_ (.Y(_04495_),
    .A(_04483_),
    .B(_04493_));
 sg13g2_o21ai_1 _26522_ (.B1(net3887),
    .Y(_04496_),
    .A1(net4334),
    .A2(_04481_));
 sg13g2_a21oi_1 _26523_ (.A1(net4334),
    .A2(_04495_),
    .Y(_04497_),
    .B1(_04496_));
 sg13g2_a21o_1 _26524_ (.A2(net3953),
    .A1(net2993),
    .B1(_04497_),
    .X(_00476_));
 sg13g2_or2_1 _26525_ (.X(_04498_),
    .B(_04477_),
    .A(_15102_));
 sg13g2_and2_1 _26526_ (.A(_13728_),
    .B(_13730_),
    .X(_04499_));
 sg13g2_o21ai_1 _26527_ (.B1(_04499_),
    .Y(_04500_),
    .A1(_13731_),
    .A2(_04477_));
 sg13g2_nand4_1 _26528_ (.B(_15119_),
    .C(_04498_),
    .A(net4671),
    .Y(_04501_),
    .D(_04500_));
 sg13g2_a21oi_1 _26529_ (.A1(net4551),
    .A2(\u_inv.d_next[201] ),
    .Y(_04502_),
    .B1(net3769));
 sg13g2_a21o_1 _26530_ (.A2(_04475_),
    .A1(_13731_),
    .B1(_13918_),
    .X(_04503_));
 sg13g2_o21ai_1 _26531_ (.B1(net3769),
    .Y(_04504_),
    .A1(_13729_),
    .A2(_04503_));
 sg13g2_a21oi_1 _26532_ (.A1(_13729_),
    .A2(_04503_),
    .Y(_04505_),
    .B1(_04504_));
 sg13g2_a21oi_2 _26533_ (.B1(_04505_),
    .Y(_04506_),
    .A2(_04502_),
    .A1(_04501_));
 sg13g2_and2_1 _26534_ (.A(net3423),
    .B(_04506_),
    .X(_04507_));
 sg13g2_xnor2_1 _26535_ (.Y(_04508_),
    .A(net3424),
    .B(_04506_));
 sg13g2_nor2_1 _26536_ (.A(_04482_),
    .B(_04494_),
    .Y(_04509_));
 sg13g2_xnor2_1 _26537_ (.Y(_04510_),
    .A(_04508_),
    .B(_04509_));
 sg13g2_o21ai_1 _26538_ (.B1(net3886),
    .Y(_04511_),
    .A1(net4336),
    .A2(_04506_));
 sg13g2_a21oi_1 _26539_ (.A1(net4336),
    .A2(_04510_),
    .Y(_04512_),
    .B1(_04511_));
 sg13g2_a21o_1 _26540_ (.A2(net3953),
    .A1(net2897),
    .B1(_04512_),
    .X(_00477_));
 sg13g2_a21oi_1 _26541_ (.A1(_13907_),
    .A2(_04474_),
    .Y(_04513_),
    .B1(_13733_));
 sg13g2_nor2_1 _26542_ (.A(_13920_),
    .B(_04513_),
    .Y(_04514_));
 sg13g2_xnor2_1 _26543_ (.Y(_04515_),
    .A(_13736_),
    .B(_04514_));
 sg13g2_a21oi_1 _26544_ (.A1(_15121_),
    .A2(_04498_),
    .Y(_04516_),
    .B1(_13737_));
 sg13g2_nand3_1 _26545_ (.B(_15121_),
    .C(_04498_),
    .A(_13737_),
    .Y(_04517_));
 sg13g2_nand3b_1 _26546_ (.B(_04517_),
    .C(net4671),
    .Y(_04518_),
    .A_N(_04516_));
 sg13g2_a21oi_1 _26547_ (.A1(net4554),
    .A2(\u_inv.d_next[202] ),
    .Y(_04519_),
    .B1(net3769));
 sg13g2_a22oi_1 _26548_ (.Y(_04520_),
    .B1(_04518_),
    .B2(_04519_),
    .A2(_04515_),
    .A1(net3769));
 sg13g2_nand2_1 _26549_ (.Y(_04521_),
    .A(net3424),
    .B(_04520_));
 sg13g2_xnor2_1 _26550_ (.Y(_04522_),
    .A(net3424),
    .B(_04520_));
 sg13g2_nor2_1 _26551_ (.A(_04482_),
    .B(_04507_),
    .Y(_04523_));
 sg13g2_or2_1 _26552_ (.X(_04524_),
    .B(_04507_),
    .A(_04482_));
 sg13g2_nor3_1 _26553_ (.A(_04483_),
    .B(_04493_),
    .C(_04508_),
    .Y(_04525_));
 sg13g2_nor2_1 _26554_ (.A(_04524_),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_xnor2_1 _26555_ (.Y(_04527_),
    .A(_04522_),
    .B(_04526_));
 sg13g2_a21oi_1 _26556_ (.A1(net4334),
    .A2(_04527_),
    .Y(_04528_),
    .B1(net4235));
 sg13g2_o21ai_1 _26557_ (.B1(_04528_),
    .Y(_04529_),
    .A1(net4334),
    .A2(_04520_));
 sg13g2_o21ai_1 _26558_ (.B1(_04529_),
    .Y(_00478_),
    .A1(_10585_),
    .A2(net4025));
 sg13g2_a21oi_1 _26559_ (.A1(net4554),
    .A2(\u_inv.d_next[203] ),
    .Y(_04530_),
    .B1(net3769));
 sg13g2_o21ai_1 _26560_ (.B1(_13740_),
    .Y(_04531_),
    .A1(_13735_),
    .A2(_04516_));
 sg13g2_or3_1 _26561_ (.A(_13735_),
    .B(_13740_),
    .C(_04516_),
    .X(_04532_));
 sg13g2_nand3_1 _26562_ (.B(_04531_),
    .C(_04532_),
    .A(net4671),
    .Y(_04533_));
 sg13g2_o21ai_1 _26563_ (.B1(_13922_),
    .Y(_04534_),
    .A1(_13736_),
    .A2(_04514_));
 sg13g2_or2_1 _26564_ (.X(_04535_),
    .B(_04534_),
    .A(_13740_));
 sg13g2_a21oi_1 _26565_ (.A1(_13740_),
    .A2(_04534_),
    .Y(_04536_),
    .B1(net3842));
 sg13g2_a22oi_1 _26566_ (.Y(_04537_),
    .B1(_04535_),
    .B2(_04536_),
    .A2(_04533_),
    .A1(_04530_));
 sg13g2_xnor2_1 _26567_ (.Y(_04538_),
    .A(net3477),
    .B(_04537_));
 sg13g2_o21ai_1 _26568_ (.B1(_04521_),
    .Y(_04539_),
    .A1(_04522_),
    .A2(_04526_));
 sg13g2_xnor2_1 _26569_ (.Y(_04540_),
    .A(_04538_),
    .B(_04539_));
 sg13g2_o21ai_1 _26570_ (.B1(net3886),
    .Y(_04541_),
    .A1(net4334),
    .A2(_04537_));
 sg13g2_a21oi_1 _26571_ (.A1(net4334),
    .A2(_04540_),
    .Y(_04542_),
    .B1(_04541_));
 sg13g2_a21o_1 _26572_ (.A2(net3944),
    .A1(net2538),
    .B1(_04542_),
    .X(_00479_));
 sg13g2_o21ai_1 _26573_ (.B1(_13741_),
    .Y(_04543_),
    .A1(_13920_),
    .A2(_04513_));
 sg13g2_a21oi_1 _26574_ (.A1(_13923_),
    .A2(_04543_),
    .Y(_04544_),
    .B1(_13724_));
 sg13g2_nand3_1 _26575_ (.B(_13923_),
    .C(_04543_),
    .A(_13724_),
    .Y(_04545_));
 sg13g2_nand2b_1 _26576_ (.Y(_04546_),
    .B(_04545_),
    .A_N(_04544_));
 sg13g2_nor3_1 _26577_ (.A(_15101_),
    .B(_15102_),
    .C(_04477_),
    .Y(_04547_));
 sg13g2_o21ai_1 _26578_ (.B1(_13724_),
    .Y(_04548_),
    .A1(_15124_),
    .A2(_04547_));
 sg13g2_or3_1 _26579_ (.A(_13724_),
    .B(_15124_),
    .C(_04547_),
    .X(_04549_));
 sg13g2_nand3_1 _26580_ (.B(_04548_),
    .C(_04549_),
    .A(net4671),
    .Y(_04550_));
 sg13g2_a21oi_1 _26581_ (.A1(net4550),
    .A2(\u_inv.d_next[204] ),
    .Y(_04551_),
    .B1(net3768));
 sg13g2_a22oi_1 _26582_ (.Y(_04552_),
    .B1(_04550_),
    .B2(_04551_),
    .A2(_04546_),
    .A1(net3768));
 sg13g2_and2_1 _26583_ (.A(net3423),
    .B(_04552_),
    .X(_04553_));
 sg13g2_xnor2_1 _26584_ (.Y(_04554_),
    .A(net3423),
    .B(_04552_));
 sg13g2_o21ai_1 _26585_ (.B1(net3424),
    .Y(_04555_),
    .A1(_04520_),
    .A2(_04537_));
 sg13g2_nand2b_1 _26586_ (.Y(_04556_),
    .B(_04538_),
    .A_N(_04522_));
 sg13g2_inv_1 _26587_ (.Y(_04557_),
    .A(_04556_));
 sg13g2_o21ai_1 _26588_ (.B1(_04557_),
    .Y(_04558_),
    .A1(_04524_),
    .A2(_04525_));
 sg13g2_a21oi_1 _26589_ (.A1(_04555_),
    .A2(_04558_),
    .Y(_04559_),
    .B1(_04554_));
 sg13g2_and3_1 _26590_ (.X(_04560_),
    .A(_04554_),
    .B(_04555_),
    .C(_04558_));
 sg13g2_o21ai_1 _26591_ (.B1(net4334),
    .Y(_04561_),
    .A1(_04559_),
    .A2(_04560_));
 sg13g2_o21ai_1 _26592_ (.B1(net3886),
    .Y(_04562_),
    .A1(net4334),
    .A2(_04552_));
 sg13g2_nor2b_1 _26593_ (.A(_04562_),
    .B_N(_04561_),
    .Y(_04563_));
 sg13g2_a21o_1 _26594_ (.A2(net3944),
    .A1(net2657),
    .B1(_04563_),
    .X(_00480_));
 sg13g2_nand3_1 _26595_ (.B(_13723_),
    .C(_04548_),
    .A(_13721_),
    .Y(_04564_));
 sg13g2_nor2_1 _26596_ (.A(_13721_),
    .B(_04548_),
    .Y(_04565_));
 sg13g2_o21ai_1 _26597_ (.B1(_15099_),
    .Y(_04566_),
    .A1(_15124_),
    .A2(_04547_));
 sg13g2_nor3_1 _26598_ (.A(net4550),
    .B(_15127_),
    .C(_04565_),
    .Y(_04567_));
 sg13g2_a221oi_1 _26599_ (.B2(_04567_),
    .C1(net3768),
    .B1(_04564_),
    .A1(net4550),
    .Y(_04568_),
    .A2(\u_inv.d_next[205] ));
 sg13g2_nand3b_1 _26600_ (.B(_13721_),
    .C(_13910_),
    .Y(_04569_),
    .A_N(_04544_));
 sg13g2_o21ai_1 _26601_ (.B1(_13722_),
    .Y(_04570_),
    .A1(_13909_),
    .A2(_04544_));
 sg13g2_and3_1 _26602_ (.X(_04571_),
    .A(net3768),
    .B(_04569_),
    .C(_04570_));
 sg13g2_nor2_1 _26603_ (.A(_04568_),
    .B(_04571_),
    .Y(_04572_));
 sg13g2_or3_1 _26604_ (.A(net3477),
    .B(_04568_),
    .C(_04571_),
    .X(_04573_));
 sg13g2_o21ai_1 _26605_ (.B1(net3477),
    .Y(_04574_),
    .A1(_04568_),
    .A2(_04571_));
 sg13g2_nand2_1 _26606_ (.Y(_04575_),
    .A(_04573_),
    .B(_04574_));
 sg13g2_nor2_1 _26607_ (.A(_04553_),
    .B(_04559_),
    .Y(_04576_));
 sg13g2_xnor2_1 _26608_ (.Y(_04577_),
    .A(_04575_),
    .B(_04576_));
 sg13g2_o21ai_1 _26609_ (.B1(net3886),
    .Y(_04578_),
    .A1(net4328),
    .A2(_04572_));
 sg13g2_a21oi_1 _26610_ (.A1(net4328),
    .A2(_04577_),
    .Y(_04579_),
    .B1(_04578_));
 sg13g2_a21o_1 _26611_ (.A2(net3944),
    .A1(net2905),
    .B1(_04579_),
    .X(_00481_));
 sg13g2_a21oi_1 _26612_ (.A1(_13923_),
    .A2(_04543_),
    .Y(_04580_),
    .B1(_13726_));
 sg13g2_o21ai_1 _26613_ (.B1(_13717_),
    .Y(_04581_),
    .A1(_13911_),
    .A2(_04580_));
 sg13g2_or3_1 _26614_ (.A(_13717_),
    .B(_13911_),
    .C(_04580_),
    .X(_04582_));
 sg13g2_nand2_1 _26615_ (.Y(_04583_),
    .A(_04581_),
    .B(_04582_));
 sg13g2_and2_1 _26616_ (.A(_15128_),
    .B(_04566_),
    .X(_04584_));
 sg13g2_a21oi_1 _26617_ (.A1(_13717_),
    .A2(_04584_),
    .Y(_04585_),
    .B1(net4550));
 sg13g2_o21ai_1 _26618_ (.B1(_04585_),
    .Y(_04586_),
    .A1(_13717_),
    .A2(_04584_));
 sg13g2_a21oi_1 _26619_ (.A1(net4550),
    .A2(\u_inv.d_next[206] ),
    .Y(_04587_),
    .B1(net3768));
 sg13g2_a22oi_1 _26620_ (.Y(_04588_),
    .B1(_04586_),
    .B2(_04587_),
    .A2(_04583_),
    .A1(net3768));
 sg13g2_nand2_1 _26621_ (.Y(_04589_),
    .A(net3423),
    .B(_04588_));
 sg13g2_xnor2_1 _26622_ (.Y(_04590_),
    .A(net3423),
    .B(_04588_));
 sg13g2_nand2b_1 _26623_ (.Y(_04591_),
    .B(_04573_),
    .A_N(_04553_));
 sg13g2_nand3b_1 _26624_ (.B(_04573_),
    .C(_04574_),
    .Y(_04592_),
    .A_N(_04554_));
 sg13g2_a21oi_1 _26625_ (.A1(_04555_),
    .A2(_04558_),
    .Y(_04593_),
    .B1(_04592_));
 sg13g2_nor2_1 _26626_ (.A(_04591_),
    .B(_04593_),
    .Y(_04594_));
 sg13g2_xnor2_1 _26627_ (.Y(_04595_),
    .A(_04590_),
    .B(_04594_));
 sg13g2_o21ai_1 _26628_ (.B1(net3887),
    .Y(_04596_),
    .A1(net4328),
    .A2(_04588_));
 sg13g2_a21oi_1 _26629_ (.A1(net4330),
    .A2(_04595_),
    .Y(_04597_),
    .B1(_04596_));
 sg13g2_a21o_1 _26630_ (.A2(net3944),
    .A1(net3244),
    .B1(_04597_),
    .X(_00482_));
 sg13g2_a21oi_1 _26631_ (.A1(net4550),
    .A2(\u_inv.d_next[207] ),
    .Y(_04598_),
    .B1(net3768));
 sg13g2_o21ai_1 _26632_ (.B1(_13716_),
    .Y(_04599_),
    .A1(_13717_),
    .A2(_04584_));
 sg13g2_xor2_1 _26633_ (.B(_04599_),
    .A(_13715_),
    .X(_04600_));
 sg13g2_o21ai_1 _26634_ (.B1(_04598_),
    .Y(_04601_),
    .A1(net4550),
    .A2(_04600_));
 sg13g2_a21o_1 _26635_ (.A2(_04581_),
    .A1(_13915_),
    .B1(_13715_),
    .X(_04602_));
 sg13g2_nand3_1 _26636_ (.B(_13915_),
    .C(_04581_),
    .A(_13715_),
    .Y(_04603_));
 sg13g2_nand3_1 _26637_ (.B(_04602_),
    .C(_04603_),
    .A(net3768),
    .Y(_04604_));
 sg13g2_and2_1 _26638_ (.A(_04601_),
    .B(_04604_),
    .X(_04605_));
 sg13g2_and3_2 _26639_ (.X(_04606_),
    .A(net3423),
    .B(_04601_),
    .C(_04604_));
 sg13g2_a21oi_1 _26640_ (.A1(_04601_),
    .A2(_04604_),
    .Y(_04607_),
    .B1(net3423));
 sg13g2_nor2_1 _26641_ (.A(_04606_),
    .B(_04607_),
    .Y(_04608_));
 sg13g2_o21ai_1 _26642_ (.B1(_04589_),
    .Y(_04609_),
    .A1(_04590_),
    .A2(_04594_));
 sg13g2_xnor2_1 _26643_ (.Y(_04610_),
    .A(_04608_),
    .B(_04609_));
 sg13g2_o21ai_1 _26644_ (.B1(net3887),
    .Y(_04611_),
    .A1(net4330),
    .A2(_04605_));
 sg13g2_a21oi_1 _26645_ (.A1(net4328),
    .A2(_04610_),
    .Y(_04612_),
    .B1(_04611_));
 sg13g2_a21o_1 _26646_ (.A2(net3944),
    .A1(net3001),
    .B1(_04612_),
    .X(_00483_));
 sg13g2_o21ai_1 _26647_ (.B1(_13775_),
    .Y(_04613_),
    .A1(_14901_),
    .A2(_15026_));
 sg13g2_nand2_1 _26648_ (.Y(_04614_),
    .A(_13925_),
    .B(_04613_));
 sg13g2_xnor2_1 _26649_ (.Y(_04615_),
    .A(net4431),
    .B(_04614_));
 sg13g2_a21oi_2 _26650_ (.B1(_15131_),
    .Y(_04616_),
    .A2(_15638_),
    .A1(_15186_));
 sg13g2_a21o_1 _26651_ (.A2(_15638_),
    .A1(_15186_),
    .B1(_15131_),
    .X(_04617_));
 sg13g2_a21oi_1 _26652_ (.A1(net4431),
    .A2(_04616_),
    .Y(_04618_),
    .B1(net4551));
 sg13g2_o21ai_1 _26653_ (.B1(_04618_),
    .Y(_04619_),
    .A1(net4431),
    .A2(_04616_));
 sg13g2_a21oi_1 _26654_ (.A1(net4551),
    .A2(\u_inv.d_next[208] ),
    .Y(_04620_),
    .B1(net3770));
 sg13g2_a22oi_1 _26655_ (.Y(_04621_),
    .B1(_04619_),
    .B2(_04620_),
    .A2(_04615_),
    .A1(net3770));
 sg13g2_and2_1 _26656_ (.A(net3419),
    .B(_04621_),
    .X(_04622_));
 sg13g2_xnor2_1 _26657_ (.Y(_04623_),
    .A(net3419),
    .B(_04621_));
 sg13g2_nor3_1 _26658_ (.A(_04590_),
    .B(_04606_),
    .C(_04607_),
    .Y(_04624_));
 sg13g2_nor4_1 _26659_ (.A(_04590_),
    .B(_04592_),
    .C(_04606_),
    .D(_04607_),
    .Y(_04625_));
 sg13g2_nor3_1 _26660_ (.A(_04483_),
    .B(_04508_),
    .C(_04556_),
    .Y(_04626_));
 sg13g2_nand3b_1 _26661_ (.B(_04625_),
    .C(_04626_),
    .Y(_04627_),
    .A_N(_04490_));
 sg13g2_a221oi_1 _26662_ (.B2(_04624_),
    .C1(_04606_),
    .B1(_04591_),
    .A1(net3423),
    .Y(_04628_),
    .A2(_04588_));
 sg13g2_o21ai_1 _26663_ (.B1(_04555_),
    .Y(_04629_),
    .A1(_04523_),
    .A2(_04556_));
 sg13g2_nand2_1 _26664_ (.Y(_04630_),
    .A(_04625_),
    .B(_04629_));
 sg13g2_nand3_1 _26665_ (.B(_04628_),
    .C(_04630_),
    .A(_04627_),
    .Y(_04631_));
 sg13g2_and3_2 _26666_ (.X(_04632_),
    .A(_04492_),
    .B(_04625_),
    .C(_04626_));
 sg13g2_a21oi_2 _26667_ (.B1(_04631_),
    .Y(_04633_),
    .A2(_04632_),
    .A1(_04356_));
 sg13g2_nor2_1 _26668_ (.A(_04623_),
    .B(_04633_),
    .Y(_04634_));
 sg13g2_xnor2_1 _26669_ (.Y(_04635_),
    .A(_04623_),
    .B(_04633_));
 sg13g2_o21ai_1 _26670_ (.B1(net3885),
    .Y(_04636_),
    .A1(net4328),
    .A2(_04621_));
 sg13g2_a21oi_1 _26671_ (.A1(net4328),
    .A2(_04635_),
    .Y(_04637_),
    .B1(_04636_));
 sg13g2_a21o_1 _26672_ (.A2(net3944),
    .A1(net2730),
    .B1(_04637_),
    .X(_00484_));
 sg13g2_nor2_1 _26673_ (.A(_13823_),
    .B(_13824_),
    .Y(_04638_));
 sg13g2_o21ai_1 _26674_ (.B1(_04638_),
    .Y(_04639_),
    .A1(net4431),
    .A2(_04616_));
 sg13g2_nor3_1 _26675_ (.A(_13822_),
    .B(_13825_),
    .C(_04616_),
    .Y(_04640_));
 sg13g2_a21oi_1 _26676_ (.A1(_13823_),
    .A2(_13824_),
    .Y(_04641_),
    .B1(net4551));
 sg13g2_nor2b_1 _26677_ (.A(_04640_),
    .B_N(_04641_),
    .Y(_04642_));
 sg13g2_a22oi_1 _26678_ (.Y(_04643_),
    .B1(_04639_),
    .B2(_04642_),
    .A2(\u_inv.d_next[209] ),
    .A1(net4551));
 sg13g2_a21oi_1 _26679_ (.A1(_13825_),
    .A2(_04614_),
    .Y(_04644_),
    .B1(_13939_));
 sg13g2_or2_1 _26680_ (.X(_04645_),
    .B(_04644_),
    .A(_13822_));
 sg13g2_a21oi_1 _26681_ (.A1(_13822_),
    .A2(_04644_),
    .Y(_04646_),
    .B1(net3847));
 sg13g2_a22oi_1 _26682_ (.Y(_04647_),
    .B1(_04645_),
    .B2(_04646_),
    .A2(_04643_),
    .A1(net3847));
 sg13g2_and2_1 _26683_ (.A(net3419),
    .B(_04647_),
    .X(_04648_));
 sg13g2_nor2_1 _26684_ (.A(net3419),
    .B(_04647_),
    .Y(_04649_));
 sg13g2_nor2_1 _26685_ (.A(_04648_),
    .B(_04649_),
    .Y(_04650_));
 sg13g2_nor2_1 _26686_ (.A(_04622_),
    .B(_04634_),
    .Y(_04651_));
 sg13g2_xor2_1 _26687_ (.B(_04651_),
    .A(_04650_),
    .X(_04652_));
 sg13g2_o21ai_1 _26688_ (.B1(net3885),
    .Y(_04653_),
    .A1(net4328),
    .A2(_04647_));
 sg13g2_a21oi_1 _26689_ (.A1(net4328),
    .A2(_04652_),
    .Y(_04654_),
    .B1(_04653_));
 sg13g2_a21o_1 _26690_ (.A2(net3944),
    .A1(net2962),
    .B1(_04654_),
    .X(_00485_));
 sg13g2_a21o_1 _26691_ (.A2(_04613_),
    .A1(_13925_),
    .B1(_13826_),
    .X(_04655_));
 sg13g2_a21o_2 _26692_ (.A2(_04655_),
    .A1(_13941_),
    .B1(_13818_),
    .X(_04656_));
 sg13g2_nand3_1 _26693_ (.B(_13941_),
    .C(_04655_),
    .A(_13818_),
    .Y(_04657_));
 sg13g2_a21oi_1 _26694_ (.A1(_04656_),
    .A2(_04657_),
    .Y(_04658_),
    .B1(net3847));
 sg13g2_o21ai_1 _26695_ (.B1(_13818_),
    .Y(_04659_),
    .A1(_15073_),
    .A2(_04640_));
 sg13g2_nor3_1 _26696_ (.A(_13818_),
    .B(_15073_),
    .C(_04640_),
    .Y(_04660_));
 sg13g2_nor2_1 _26697_ (.A(net4551),
    .B(_04660_),
    .Y(_04661_));
 sg13g2_a221oi_1 _26698_ (.B2(_04661_),
    .C1(net3770),
    .B1(_04659_),
    .A1(net4551),
    .Y(_04662_),
    .A2(\u_inv.d_next[210] ));
 sg13g2_or2_1 _26699_ (.X(_04663_),
    .B(_04662_),
    .A(_04658_));
 sg13g2_nor2_1 _26700_ (.A(net3474),
    .B(_04663_),
    .Y(_04664_));
 sg13g2_inv_1 _26701_ (.Y(_04665_),
    .A(_04664_));
 sg13g2_xnor2_1 _26702_ (.Y(_04666_),
    .A(net3475),
    .B(_04663_));
 sg13g2_or2_1 _26703_ (.X(_04667_),
    .B(_04648_),
    .A(_04622_));
 sg13g2_nor2_1 _26704_ (.A(_04649_),
    .B(_04651_),
    .Y(_04668_));
 sg13g2_nor2_1 _26705_ (.A(_04648_),
    .B(_04668_),
    .Y(_04669_));
 sg13g2_xor2_1 _26706_ (.B(_04669_),
    .A(_04666_),
    .X(_04670_));
 sg13g2_o21ai_1 _26707_ (.B1(net3885),
    .Y(_04671_),
    .A1(net4293),
    .A2(_04670_));
 sg13g2_a21oi_1 _26708_ (.A1(net4293),
    .A2(_04663_),
    .Y(_04672_),
    .B1(_04671_));
 sg13g2_a21o_1 _26709_ (.A2(net3944),
    .A1(net2804),
    .B1(_04672_),
    .X(_00486_));
 sg13g2_a21oi_1 _26710_ (.A1(net4548),
    .A2(\u_inv.d_next[211] ),
    .Y(_04673_),
    .B1(net3765));
 sg13g2_a21o_1 _26711_ (.A2(_04659_),
    .A1(_13817_),
    .B1(_13815_),
    .X(_04674_));
 sg13g2_nand3_1 _26712_ (.B(_13817_),
    .C(_04659_),
    .A(_13815_),
    .Y(_04675_));
 sg13g2_nand3_1 _26713_ (.B(_04674_),
    .C(_04675_),
    .A(net4670),
    .Y(_04676_));
 sg13g2_a21oi_1 _26714_ (.A1(_13942_),
    .A2(_04656_),
    .Y(_04677_),
    .B1(_13815_));
 sg13g2_nand3_1 _26715_ (.B(_13942_),
    .C(_04656_),
    .A(_13815_),
    .Y(_04678_));
 sg13g2_nor2_1 _26716_ (.A(net3841),
    .B(_04677_),
    .Y(_04679_));
 sg13g2_a22oi_1 _26717_ (.Y(_04680_),
    .B1(_04678_),
    .B2(_04679_),
    .A2(_04676_),
    .A1(_04673_));
 sg13g2_xnor2_1 _26718_ (.Y(_04681_),
    .A(net3474),
    .B(_04680_));
 sg13g2_o21ai_1 _26719_ (.B1(_04665_),
    .Y(_04682_),
    .A1(_04666_),
    .A2(_04669_));
 sg13g2_xnor2_1 _26720_ (.Y(_04683_),
    .A(_04681_),
    .B(_04682_));
 sg13g2_o21ai_1 _26721_ (.B1(net3885),
    .Y(_04684_),
    .A1(net4326),
    .A2(_04680_));
 sg13g2_a21oi_1 _26722_ (.A1(net4326),
    .A2(_04683_),
    .Y(_04685_),
    .B1(_04684_));
 sg13g2_a21o_1 _26723_ (.A2(net3943),
    .A1(net2623),
    .B1(_04685_),
    .X(_00487_));
 sg13g2_a21oi_1 _26724_ (.A1(_13943_),
    .A2(_04656_),
    .Y(_04686_),
    .B1(_13814_));
 sg13g2_xnor2_1 _26725_ (.Y(_04687_),
    .A(_13810_),
    .B(_04686_));
 sg13g2_nor4_1 _26726_ (.A(_13822_),
    .B(net4431),
    .C(_15094_),
    .D(_04616_),
    .Y(_04688_));
 sg13g2_o21ai_1 _26727_ (.B1(_13809_),
    .Y(_04689_),
    .A1(_15075_),
    .A2(_04688_));
 sg13g2_nor3_1 _26728_ (.A(_13809_),
    .B(_15075_),
    .C(_04688_),
    .Y(_04690_));
 sg13g2_nand3b_1 _26729_ (.B(net4670),
    .C(_04689_),
    .Y(_04691_),
    .A_N(_04690_));
 sg13g2_a21oi_1 _26730_ (.A1(net4548),
    .A2(\u_inv.d_next[212] ),
    .Y(_04692_),
    .B1(net3766));
 sg13g2_a22oi_1 _26731_ (.Y(_04693_),
    .B1(_04691_),
    .B2(_04692_),
    .A2(_04687_),
    .A1(net3766));
 sg13g2_and2_1 _26732_ (.A(net3417),
    .B(_04693_),
    .X(_04694_));
 sg13g2_xnor2_1 _26733_ (.Y(_04695_),
    .A(net3418),
    .B(_04693_));
 sg13g2_nor2b_1 _26734_ (.A(_04666_),
    .B_N(_04681_),
    .Y(_04696_));
 sg13g2_a221oi_1 _26735_ (.B2(_04667_),
    .C1(_04664_),
    .B1(_04696_),
    .A1(net3417),
    .Y(_04697_),
    .A2(_04680_));
 sg13g2_nand3b_1 _26736_ (.B(_04650_),
    .C(_04696_),
    .Y(_04698_),
    .A_N(_04623_));
 sg13g2_o21ai_1 _26737_ (.B1(_04697_),
    .Y(_04699_),
    .A1(_04633_),
    .A2(_04698_));
 sg13g2_nand2b_1 _26738_ (.Y(_04700_),
    .B(_04699_),
    .A_N(_04695_));
 sg13g2_xor2_1 _26739_ (.B(_04699_),
    .A(_04695_),
    .X(_04701_));
 sg13g2_a21oi_1 _26740_ (.A1(net4326),
    .A2(_04701_),
    .Y(_04702_),
    .B1(net4235));
 sg13g2_o21ai_1 _26741_ (.B1(_04702_),
    .Y(_04703_),
    .A1(net4326),
    .A2(_04693_));
 sg13g2_o21ai_1 _26742_ (.B1(_04703_),
    .Y(_00488_),
    .A1(_10584_),
    .A2(net4025));
 sg13g2_nand3_1 _26743_ (.B(_13808_),
    .C(_04689_),
    .A(_13807_),
    .Y(_04704_));
 sg13g2_o21ai_1 _26744_ (.B1(_15068_),
    .Y(_04705_),
    .A1(_15075_),
    .A2(_04688_));
 sg13g2_o21ai_1 _26745_ (.B1(net4670),
    .Y(_04706_),
    .A1(_13807_),
    .A2(_13808_));
 sg13g2_nand3b_1 _26746_ (.B(_04705_),
    .C(_04704_),
    .Y(_04707_),
    .A_N(_04706_));
 sg13g2_a21oi_1 _26747_ (.A1(net4548),
    .A2(\u_inv.d_next[213] ),
    .Y(_04708_),
    .B1(net3766));
 sg13g2_a21oi_1 _26748_ (.A1(_13810_),
    .A2(_04686_),
    .Y(_04709_),
    .B1(_13949_));
 sg13g2_or2_1 _26749_ (.X(_04710_),
    .B(_04709_),
    .A(_13807_));
 sg13g2_a21oi_1 _26750_ (.A1(_13807_),
    .A2(_04709_),
    .Y(_04711_),
    .B1(net3841));
 sg13g2_a22oi_1 _26751_ (.Y(_04712_),
    .B1(_04710_),
    .B2(_04711_),
    .A2(_04708_),
    .A1(_04707_));
 sg13g2_nor2_1 _26752_ (.A(net3417),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_xnor2_1 _26753_ (.Y(_04714_),
    .A(net3417),
    .B(_04712_));
 sg13g2_nor2b_1 _26754_ (.A(_04694_),
    .B_N(_04700_),
    .Y(_04715_));
 sg13g2_xnor2_1 _26755_ (.Y(_04716_),
    .A(_04714_),
    .B(_04715_));
 sg13g2_o21ai_1 _26756_ (.B1(net3885),
    .Y(_04717_),
    .A1(net4326),
    .A2(_04712_));
 sg13g2_a21oi_1 _26757_ (.A1(net4326),
    .A2(_04716_),
    .Y(_04718_),
    .B1(_04717_));
 sg13g2_a21o_1 _26758_ (.A2(net3943),
    .A1(net3112),
    .B1(_04718_),
    .X(_00489_));
 sg13g2_a221oi_1 _26759_ (.B2(_04656_),
    .C1(_13812_),
    .B1(_13943_),
    .A1(_10584_),
    .Y(_04719_),
    .A2(\u_inv.d_reg[211] ));
 sg13g2_o21ai_1 _26760_ (.B1(_13803_),
    .Y(_04720_),
    .A1(_13950_),
    .A2(_04719_));
 sg13g2_or3_1 _26761_ (.A(_13803_),
    .B(_13950_),
    .C(_04719_),
    .X(_04721_));
 sg13g2_nand2_1 _26762_ (.Y(_04722_),
    .A(_04720_),
    .B(_04721_));
 sg13g2_a21o_1 _26763_ (.A2(_04705_),
    .A1(_15078_),
    .B1(_13803_),
    .X(_04723_));
 sg13g2_nand3_1 _26764_ (.B(_15078_),
    .C(_04705_),
    .A(_13803_),
    .Y(_04724_));
 sg13g2_nand3_1 _26765_ (.B(_04723_),
    .C(_04724_),
    .A(net4670),
    .Y(_04725_));
 sg13g2_a21oi_1 _26766_ (.A1(net4549),
    .A2(\u_inv.d_next[214] ),
    .Y(_04726_),
    .B1(net3766));
 sg13g2_a22oi_1 _26767_ (.Y(_04727_),
    .B1(_04725_),
    .B2(_04726_),
    .A2(_04722_),
    .A1(net3766));
 sg13g2_and2_1 _26768_ (.A(net3416),
    .B(_04727_),
    .X(_04728_));
 sg13g2_xnor2_1 _26769_ (.Y(_04729_),
    .A(net3417),
    .B(_04727_));
 sg13g2_a21oi_1 _26770_ (.A1(net3417),
    .A2(_04712_),
    .Y(_04730_),
    .B1(_04694_));
 sg13g2_a21oi_1 _26771_ (.A1(_04700_),
    .A2(_04730_),
    .Y(_04731_),
    .B1(_04713_));
 sg13g2_nor2b_1 _26772_ (.A(_04729_),
    .B_N(_04731_),
    .Y(_04732_));
 sg13g2_xor2_1 _26773_ (.B(_04731_),
    .A(_04729_),
    .X(_04733_));
 sg13g2_o21ai_1 _26774_ (.B1(net3885),
    .Y(_04734_),
    .A1(net4325),
    .A2(_04727_));
 sg13g2_a21oi_1 _26775_ (.A1(net4327),
    .A2(_04733_),
    .Y(_04735_),
    .B1(_04734_));
 sg13g2_a21o_1 _26776_ (.A2(net3943),
    .A1(net2703),
    .B1(_04735_),
    .X(_00490_));
 sg13g2_nand3_1 _26777_ (.B(_13802_),
    .C(_04723_),
    .A(_13801_),
    .Y(_04736_));
 sg13g2_a21oi_1 _26778_ (.A1(_13802_),
    .A2(_04723_),
    .Y(_04737_),
    .B1(_13801_));
 sg13g2_nor2_1 _26779_ (.A(net4549),
    .B(_04737_),
    .Y(_04738_));
 sg13g2_a221oi_1 _26780_ (.B2(_04738_),
    .C1(net3766),
    .B1(_04736_),
    .A1(net4549),
    .Y(_04739_),
    .A2(\u_inv.d_next[215] ));
 sg13g2_a21oi_1 _26781_ (.A1(_13948_),
    .A2(_04720_),
    .Y(_04740_),
    .B1(_13801_));
 sg13g2_and3_1 _26782_ (.X(_04741_),
    .A(_13801_),
    .B(_13948_),
    .C(_04720_));
 sg13g2_nor3_1 _26783_ (.A(net3841),
    .B(_04740_),
    .C(_04741_),
    .Y(_04742_));
 sg13g2_nor2_1 _26784_ (.A(_04739_),
    .B(_04742_),
    .Y(_04743_));
 sg13g2_nor3_1 _26785_ (.A(net3474),
    .B(_04739_),
    .C(_04742_),
    .Y(_04744_));
 sg13g2_xnor2_1 _26786_ (.Y(_04745_),
    .A(net3416),
    .B(_04743_));
 sg13g2_nor2_1 _26787_ (.A(_04728_),
    .B(_04732_),
    .Y(_04746_));
 sg13g2_xnor2_1 _26788_ (.Y(_04747_),
    .A(_04745_),
    .B(_04746_));
 sg13g2_o21ai_1 _26789_ (.B1(net3885),
    .Y(_04748_),
    .A1(net4325),
    .A2(_04743_));
 sg13g2_a21oi_1 _26790_ (.A1(net4325),
    .A2(_04747_),
    .Y(_04749_),
    .B1(_04748_));
 sg13g2_a21o_1 _26791_ (.A2(net3943),
    .A1(net2773),
    .B1(_04749_),
    .X(_00491_));
 sg13g2_a21oi_1 _26792_ (.A1(_13925_),
    .A2(_04613_),
    .Y(_04750_),
    .B1(_13829_));
 sg13g2_o21ai_1 _26793_ (.B1(_13790_),
    .Y(_04751_),
    .A1(_13952_),
    .A2(_04750_));
 sg13g2_nand3b_1 _26794_ (.B(_13953_),
    .C(_13789_),
    .Y(_04752_),
    .A_N(_04750_));
 sg13g2_nand2_1 _26795_ (.Y(_04753_),
    .A(_04751_),
    .B(_04752_));
 sg13g2_a21oi_2 _26796_ (.B1(_15082_),
    .Y(_04754_),
    .A2(_04617_),
    .A1(_15095_));
 sg13g2_a21oi_1 _26797_ (.A1(_13790_),
    .A2(_04754_),
    .Y(_04755_),
    .B1(net4548));
 sg13g2_o21ai_1 _26798_ (.B1(_04755_),
    .Y(_04756_),
    .A1(_13790_),
    .A2(_04754_));
 sg13g2_a21oi_1 _26799_ (.A1(net4548),
    .A2(\u_inv.d_next[216] ),
    .Y(_04757_),
    .B1(net3765));
 sg13g2_a22oi_1 _26800_ (.Y(_04758_),
    .B1(_04756_),
    .B2(_04757_),
    .A2(_04753_),
    .A1(net3765));
 sg13g2_and2_1 _26801_ (.A(net3417),
    .B(_04758_),
    .X(_04759_));
 sg13g2_nand2b_1 _26802_ (.Y(_04760_),
    .B(net3474),
    .A_N(_04758_));
 sg13g2_nand2b_1 _26803_ (.Y(_04761_),
    .B(_04760_),
    .A_N(_04759_));
 sg13g2_or2_1 _26804_ (.X(_04762_),
    .B(_04714_),
    .A(_04695_));
 sg13g2_nor4_1 _26805_ (.A(_04697_),
    .B(_04729_),
    .C(_04745_),
    .D(_04762_),
    .Y(_04763_));
 sg13g2_nor3_1 _26806_ (.A(_04729_),
    .B(_04730_),
    .C(_04745_),
    .Y(_04764_));
 sg13g2_nor4_1 _26807_ (.A(_04728_),
    .B(_04744_),
    .C(_04763_),
    .D(_04764_),
    .Y(_04765_));
 sg13g2_or4_1 _26808_ (.A(_04698_),
    .B(_04729_),
    .C(_04745_),
    .D(_04762_),
    .X(_04766_));
 sg13g2_o21ai_1 _26809_ (.B1(_04765_),
    .Y(_04767_),
    .A1(_04633_),
    .A2(_04766_));
 sg13g2_xor2_1 _26810_ (.B(_04767_),
    .A(_04761_),
    .X(_04768_));
 sg13g2_o21ai_1 _26811_ (.B1(net3883),
    .Y(_04769_),
    .A1(net4325),
    .A2(_04758_));
 sg13g2_a21oi_1 _26812_ (.A1(net4325),
    .A2(_04768_),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_a21o_1 _26813_ (.A2(net3943),
    .A1(net2929),
    .B1(_04770_),
    .X(_00492_));
 sg13g2_a21oi_1 _26814_ (.A1(_04760_),
    .A2(_04767_),
    .Y(_04771_),
    .B1(_04759_));
 sg13g2_a21oi_1 _26815_ (.A1(net4543),
    .A2(\u_inv.d_next[217] ),
    .Y(_04772_),
    .B1(net3759));
 sg13g2_o21ai_1 _26816_ (.B1(_13788_),
    .Y(_04773_),
    .A1(_13790_),
    .A2(_04754_));
 sg13g2_a21oi_1 _26817_ (.A1(_13795_),
    .A2(_04773_),
    .Y(_04774_),
    .B1(net4544));
 sg13g2_o21ai_1 _26818_ (.B1(_04774_),
    .Y(_04775_),
    .A1(_13795_),
    .A2(_04773_));
 sg13g2_o21ai_1 _26819_ (.B1(_04751_),
    .Y(_04776_),
    .A1(_10583_),
    .A2(\u_inv.d_reg[216] ));
 sg13g2_o21ai_1 _26820_ (.B1(net3760),
    .Y(_04777_),
    .A1(_13795_),
    .A2(_04776_));
 sg13g2_a21oi_1 _26821_ (.A1(_13795_),
    .A2(_04776_),
    .Y(_04778_),
    .B1(_04777_));
 sg13g2_a21oi_2 _26822_ (.B1(_04778_),
    .Y(_04779_),
    .A2(_04775_),
    .A1(_04772_));
 sg13g2_xnor2_1 _26823_ (.Y(_04780_),
    .A(net3415),
    .B(_04779_));
 sg13g2_xnor2_1 _26824_ (.Y(_04781_),
    .A(_04771_),
    .B(_04780_));
 sg13g2_o21ai_1 _26825_ (.B1(net3884),
    .Y(_04782_),
    .A1(net4321),
    .A2(_04779_));
 sg13g2_a21o_1 _26826_ (.A2(_04781_),
    .A1(net4321),
    .B1(_04782_),
    .X(_04783_));
 sg13g2_o21ai_1 _26827_ (.B1(_04783_),
    .Y(_00493_),
    .A1(_10583_),
    .A2(net4019));
 sg13g2_a21o_1 _26828_ (.A2(_04751_),
    .A1(_13928_),
    .B1(_13794_),
    .X(_04784_));
 sg13g2_a221oi_1 _26829_ (.B2(_04751_),
    .C1(_13792_),
    .B1(_13928_),
    .A1(_10582_),
    .Y(_04785_),
    .A2(\u_inv.d_reg[217] ));
 sg13g2_xnor2_1 _26830_ (.Y(_04786_),
    .A(_13792_),
    .B(_04784_));
 sg13g2_o21ai_1 _26831_ (.B1(_15084_),
    .Y(_04787_),
    .A1(_15065_),
    .A2(_04754_));
 sg13g2_xnor2_1 _26832_ (.Y(_04788_),
    .A(_13793_),
    .B(_04787_));
 sg13g2_nand2b_1 _26833_ (.Y(_04789_),
    .B(net3836),
    .A_N(\u_inv.d_next[218] ));
 sg13g2_a22oi_1 _26834_ (.Y(_04790_),
    .B1(_04789_),
    .B2(net3726),
    .A2(_04788_),
    .A1(net4659));
 sg13g2_a21o_2 _26835_ (.A2(_04786_),
    .A1(net3759),
    .B1(_04790_),
    .X(_04791_));
 sg13g2_nor2_1 _26836_ (.A(net3473),
    .B(_04791_),
    .Y(_04792_));
 sg13g2_nand2b_1 _26837_ (.Y(_04793_),
    .B(net3415),
    .A_N(_04791_));
 sg13g2_xnor2_1 _26838_ (.Y(_04794_),
    .A(net3473),
    .B(_04791_));
 sg13g2_a21o_1 _26839_ (.A2(_04779_),
    .A1(net3415),
    .B1(_04759_),
    .X(_04795_));
 sg13g2_or2_1 _26840_ (.X(_04796_),
    .B(_04780_),
    .A(_04761_));
 sg13g2_inv_1 _26841_ (.Y(_04797_),
    .A(_04796_));
 sg13g2_a21oi_1 _26842_ (.A1(_04767_),
    .A2(_04797_),
    .Y(_04798_),
    .B1(_04795_));
 sg13g2_xnor2_1 _26843_ (.Y(_04799_),
    .A(_04794_),
    .B(_04798_));
 sg13g2_nand2_1 _26844_ (.Y(_04800_),
    .A(net4293),
    .B(_04791_));
 sg13g2_a21oi_1 _26845_ (.A1(net4322),
    .A2(_04799_),
    .Y(_04801_),
    .B1(net4234));
 sg13g2_nand2_1 _26846_ (.Y(_04802_),
    .A(_04800_),
    .B(_04801_));
 sg13g2_o21ai_1 _26847_ (.B1(_04802_),
    .Y(_00494_),
    .A1(_10582_),
    .A2(net4019));
 sg13g2_a21oi_1 _26848_ (.A1(net4544),
    .A2(\u_inv.d_next[219] ),
    .Y(_04803_),
    .B1(net3760));
 sg13g2_a21oi_1 _26849_ (.A1(_13792_),
    .A2(_04787_),
    .Y(_04804_),
    .B1(_13791_));
 sg13g2_xnor2_1 _26850_ (.Y(_04805_),
    .A(_13797_),
    .B(_04804_));
 sg13g2_nand2_1 _26851_ (.Y(_04806_),
    .A(net4659),
    .B(_04805_));
 sg13g2_o21ai_1 _26852_ (.B1(_13797_),
    .Y(_04807_),
    .A1(_13927_),
    .A2(_04785_));
 sg13g2_nor3_1 _26853_ (.A(_13797_),
    .B(_13927_),
    .C(_04785_),
    .Y(_04808_));
 sg13g2_nor2_1 _26854_ (.A(net3836),
    .B(_04808_),
    .Y(_04809_));
 sg13g2_a22oi_1 _26855_ (.Y(_04810_),
    .B1(_04807_),
    .B2(_04809_),
    .A2(_04806_),
    .A1(_04803_));
 sg13g2_xnor2_1 _26856_ (.Y(_04811_),
    .A(net3415),
    .B(_04810_));
 sg13g2_o21ai_1 _26857_ (.B1(_04793_),
    .Y(_04812_),
    .A1(_04794_),
    .A2(_04798_));
 sg13g2_xor2_1 _26858_ (.B(_04812_),
    .A(_04811_),
    .X(_04813_));
 sg13g2_o21ai_1 _26859_ (.B1(net3883),
    .Y(_04814_),
    .A1(net4322),
    .A2(_04810_));
 sg13g2_a21oi_1 _26860_ (.A1(net4322),
    .A2(_04813_),
    .Y(_04815_),
    .B1(_04814_));
 sg13g2_a21o_1 _26861_ (.A2(net3934),
    .A1(net2789),
    .B1(_04815_),
    .X(_00495_));
 sg13g2_o21ai_1 _26862_ (.B1(_13798_),
    .Y(_04816_),
    .A1(_13952_),
    .A2(_04750_));
 sg13g2_nand2b_2 _26863_ (.Y(_04817_),
    .B(_04816_),
    .A_N(_13931_));
 sg13g2_xnor2_1 _26864_ (.Y(_04818_),
    .A(_13780_),
    .B(_04817_));
 sg13g2_a21oi_1 _26865_ (.A1(_15063_),
    .A2(_04787_),
    .Y(_04819_),
    .B1(_15087_));
 sg13g2_a21o_1 _26866_ (.A2(_04787_),
    .A1(_15063_),
    .B1(_15087_),
    .X(_04820_));
 sg13g2_a21oi_1 _26867_ (.A1(_13780_),
    .A2(_04819_),
    .Y(_04821_),
    .B1(net4548));
 sg13g2_o21ai_1 _26868_ (.B1(_04821_),
    .Y(_04822_),
    .A1(_13780_),
    .A2(_04819_));
 sg13g2_a21oi_1 _26869_ (.A1(net4548),
    .A2(\u_inv.d_next[220] ),
    .Y(_04823_),
    .B1(net3765));
 sg13g2_a22oi_1 _26870_ (.Y(_04824_),
    .B1(_04822_),
    .B2(_04823_),
    .A2(_04818_),
    .A1(net3765));
 sg13g2_and2_1 _26871_ (.A(net3416),
    .B(_04824_),
    .X(_04825_));
 sg13g2_xnor2_1 _26872_ (.Y(_04826_),
    .A(net3416),
    .B(_04824_));
 sg13g2_nor2_1 _26873_ (.A(_04794_),
    .B(_04811_),
    .Y(_04827_));
 sg13g2_a221oi_1 _26874_ (.B2(_04795_),
    .C1(_04792_),
    .B1(_04827_),
    .A1(net3415),
    .Y(_04828_),
    .A2(_04810_));
 sg13g2_nand3_1 _26875_ (.B(_04797_),
    .C(_04827_),
    .A(_04767_),
    .Y(_04829_));
 sg13g2_a21oi_1 _26876_ (.A1(_04828_),
    .A2(_04829_),
    .Y(_04830_),
    .B1(_04826_));
 sg13g2_nand3_1 _26877_ (.B(_04828_),
    .C(_04829_),
    .A(_04826_),
    .Y(_04831_));
 sg13g2_nand2b_1 _26878_ (.Y(_04832_),
    .B(_04831_),
    .A_N(_04830_));
 sg13g2_o21ai_1 _26879_ (.B1(net3883),
    .Y(_04833_),
    .A1(net4324),
    .A2(_04824_));
 sg13g2_a21oi_1 _26880_ (.A1(net4324),
    .A2(_04832_),
    .Y(_04834_),
    .B1(_04833_));
 sg13g2_a21o_1 _26881_ (.A2(net3934),
    .A1(net2938),
    .B1(_04834_),
    .X(_00496_));
 sg13g2_nor2_1 _26882_ (.A(_04825_),
    .B(_04830_),
    .Y(_04835_));
 sg13g2_nand2_1 _26883_ (.Y(_04836_),
    .A(_10581_),
    .B(net3841));
 sg13g2_o21ai_1 _26884_ (.B1(_13779_),
    .Y(_04837_),
    .A1(_13780_),
    .A2(_04819_));
 sg13g2_xnor2_1 _26885_ (.Y(_04838_),
    .A(_13778_),
    .B(_04837_));
 sg13g2_a22oi_1 _26886_ (.Y(_04839_),
    .B1(_04838_),
    .B2(net4670),
    .A2(_04836_),
    .A1(net3728));
 sg13g2_a21oi_1 _26887_ (.A1(_13780_),
    .A2(_04817_),
    .Y(_04840_),
    .B1(_13933_));
 sg13g2_o21ai_1 _26888_ (.B1(net3765),
    .Y(_04841_),
    .A1(_13778_),
    .A2(_04840_));
 sg13g2_a21oi_1 _26889_ (.A1(_13778_),
    .A2(_04840_),
    .Y(_04842_),
    .B1(_04841_));
 sg13g2_nor2_1 _26890_ (.A(_04839_),
    .B(_04842_),
    .Y(_04843_));
 sg13g2_xnor2_1 _26891_ (.Y(_04844_),
    .A(net3474),
    .B(_04843_));
 sg13g2_xor2_1 _26892_ (.B(_04844_),
    .A(_04835_),
    .X(_04845_));
 sg13g2_o21ai_1 _26893_ (.B1(net3883),
    .Y(_04846_),
    .A1(net4324),
    .A2(_04843_));
 sg13g2_a21oi_1 _26894_ (.A1(net4324),
    .A2(_04845_),
    .Y(_04847_),
    .B1(_04846_));
 sg13g2_a21o_1 _26895_ (.A2(net3943),
    .A1(net2810),
    .B1(_04847_),
    .X(_00497_));
 sg13g2_a21oi_1 _26896_ (.A1(_13781_),
    .A2(_04817_),
    .Y(_04848_),
    .B1(_13935_));
 sg13g2_xnor2_1 _26897_ (.Y(_04849_),
    .A(_13785_),
    .B(_04848_));
 sg13g2_a21oi_1 _26898_ (.A1(_15061_),
    .A2(_04820_),
    .Y(_04850_),
    .B1(_15090_));
 sg13g2_xnor2_1 _26899_ (.Y(_04851_),
    .A(_13785_),
    .B(_04850_));
 sg13g2_nand2_1 _26900_ (.Y(_04852_),
    .A(net4670),
    .B(_04851_));
 sg13g2_a21oi_1 _26901_ (.A1(net4548),
    .A2(\u_inv.d_next[222] ),
    .Y(_04853_),
    .B1(net3765));
 sg13g2_a22oi_1 _26902_ (.Y(_04854_),
    .B1(_04852_),
    .B2(_04853_),
    .A2(_04849_),
    .A1(net3765));
 sg13g2_nand2_1 _26903_ (.Y(_04855_),
    .A(net3416),
    .B(_04854_));
 sg13g2_xnor2_1 _26904_ (.Y(_04856_),
    .A(net3474),
    .B(_04854_));
 sg13g2_inv_1 _26905_ (.Y(_04857_),
    .A(_04856_));
 sg13g2_a21o_1 _26906_ (.A2(_04843_),
    .A1(net3416),
    .B1(_04825_),
    .X(_04858_));
 sg13g2_nand2b_1 _26907_ (.Y(_04859_),
    .B(_04844_),
    .A_N(_04826_));
 sg13g2_a21oi_1 _26908_ (.A1(_04830_),
    .A2(_04844_),
    .Y(_04860_),
    .B1(_04858_));
 sg13g2_xnor2_1 _26909_ (.Y(_04861_),
    .A(_04857_),
    .B(_04860_));
 sg13g2_a21oi_1 _26910_ (.A1(net4324),
    .A2(_04861_),
    .Y(_04862_),
    .B1(net4234));
 sg13g2_o21ai_1 _26911_ (.B1(_04862_),
    .Y(_04863_),
    .A1(net4324),
    .A2(_04854_));
 sg13g2_o21ai_1 _26912_ (.B1(_04863_),
    .Y(_00498_),
    .A1(_10581_),
    .A2(net4025));
 sg13g2_a21oi_1 _26913_ (.A1(net4544),
    .A2(\u_inv.d_next[223] ),
    .Y(_04864_),
    .B1(net3760));
 sg13g2_o21ai_1 _26914_ (.B1(_13783_),
    .Y(_04865_),
    .A1(_13784_),
    .A2(_04850_));
 sg13g2_xnor2_1 _26915_ (.Y(_04866_),
    .A(_13782_),
    .B(_04865_));
 sg13g2_o21ai_1 _26916_ (.B1(_04864_),
    .Y(_04867_),
    .A1(net4544),
    .A2(_04866_));
 sg13g2_o21ai_1 _26917_ (.B1(_13932_),
    .Y(_04868_),
    .A1(_13785_),
    .A2(_04848_));
 sg13g2_a21oi_1 _26918_ (.A1(_13782_),
    .A2(_04868_),
    .Y(_04869_),
    .B1(net3841));
 sg13g2_o21ai_1 _26919_ (.B1(_04869_),
    .Y(_04870_),
    .A1(_13782_),
    .A2(_04868_));
 sg13g2_and2_1 _26920_ (.A(_04867_),
    .B(_04870_),
    .X(_04871_));
 sg13g2_nand3_1 _26921_ (.B(_04867_),
    .C(_04870_),
    .A(net3416),
    .Y(_04872_));
 sg13g2_a21o_1 _26922_ (.A2(_04870_),
    .A1(_04867_),
    .B1(net3416),
    .X(_04873_));
 sg13g2_and2_1 _26923_ (.A(_04872_),
    .B(_04873_),
    .X(_04874_));
 sg13g2_o21ai_1 _26924_ (.B1(_04855_),
    .Y(_04875_),
    .A1(_04857_),
    .A2(_04860_));
 sg13g2_xnor2_1 _26925_ (.Y(_04876_),
    .A(_04874_),
    .B(_04875_));
 sg13g2_o21ai_1 _26926_ (.B1(net3883),
    .Y(_04877_),
    .A1(net4324),
    .A2(_04871_));
 sg13g2_a21oi_1 _26927_ (.A1(net4324),
    .A2(_04876_),
    .Y(_04878_),
    .B1(_04877_));
 sg13g2_a21o_1 _26928_ (.A2(net3943),
    .A1(net3240),
    .B1(_04878_),
    .X(_00499_));
 sg13g2_o21ai_1 _26929_ (.B1(_13955_),
    .Y(_04879_),
    .A1(_13830_),
    .A2(_04333_));
 sg13g2_xnor2_1 _26930_ (.Y(_04880_),
    .A(_13708_),
    .B(_04879_));
 sg13g2_a21oi_2 _26931_ (.B1(_15133_),
    .Y(_04881_),
    .A2(_15638_),
    .A1(_15187_));
 sg13g2_or2_1 _26932_ (.X(_04882_),
    .B(_04881_),
    .A(_13708_));
 sg13g2_a21oi_1 _26933_ (.A1(_13708_),
    .A2(_04881_),
    .Y(_04883_),
    .B1(net4541));
 sg13g2_nand2_1 _26934_ (.Y(_04884_),
    .A(_04882_),
    .B(_04883_));
 sg13g2_a21oi_1 _26935_ (.A1(net4541),
    .A2(\u_inv.d_next[224] ),
    .Y(_04885_),
    .B1(net3756));
 sg13g2_a22oi_1 _26936_ (.Y(_04886_),
    .B1(_04884_),
    .B2(_04885_),
    .A2(_04880_),
    .A1(net3756));
 sg13g2_and2_1 _26937_ (.A(net3411),
    .B(_04886_),
    .X(_04887_));
 sg13g2_xnor2_1 _26938_ (.Y(_04888_),
    .A(net3472),
    .B(_04886_));
 sg13g2_nand3_1 _26939_ (.B(_04872_),
    .C(_04873_),
    .A(_04856_),
    .Y(_04889_));
 sg13g2_or2_1 _26940_ (.X(_04890_),
    .B(_04889_),
    .A(_04859_));
 sg13g2_nand2b_1 _26941_ (.Y(_04891_),
    .B(_04827_),
    .A_N(_04796_));
 sg13g2_nor4_1 _26942_ (.A(_04766_),
    .B(_04859_),
    .C(_04889_),
    .D(_04891_),
    .Y(_04892_));
 sg13g2_and2_1 _26943_ (.A(_04632_),
    .B(_04892_),
    .X(_04893_));
 sg13g2_and2_1 _26944_ (.A(_04631_),
    .B(_04892_),
    .X(_04894_));
 sg13g2_nand2b_1 _26945_ (.Y(_04895_),
    .B(_04858_),
    .A_N(_04889_));
 sg13g2_nand2_1 _26946_ (.Y(_04896_),
    .A(_04855_),
    .B(_04895_));
 sg13g2_o21ai_1 _26947_ (.B1(_04872_),
    .Y(_04897_),
    .A1(_04828_),
    .A2(_04890_));
 sg13g2_nor3_1 _26948_ (.A(_04765_),
    .B(_04890_),
    .C(_04891_),
    .Y(_04898_));
 sg13g2_or4_1 _26949_ (.A(_04894_),
    .B(_04896_),
    .C(_04897_),
    .D(_04898_),
    .X(_04899_));
 sg13g2_a21oi_2 _26950_ (.B1(_04899_),
    .Y(_04900_),
    .A2(_04893_),
    .A1(_04356_));
 sg13g2_a21o_2 _26951_ (.A2(_04893_),
    .A1(_04356_),
    .B1(_04899_),
    .X(_04901_));
 sg13g2_xnor2_1 _26952_ (.Y(_04902_),
    .A(_04888_),
    .B(_04900_));
 sg13g2_nor2_1 _26953_ (.A(net4322),
    .B(_04886_),
    .Y(_04903_));
 sg13g2_o21ai_1 _26954_ (.B1(net3882),
    .Y(_04904_),
    .A1(net4292),
    .A2(_04902_));
 sg13g2_nand2_1 _26955_ (.Y(_04905_),
    .A(net2413),
    .B(net3934));
 sg13g2_o21ai_1 _26956_ (.B1(_04905_),
    .Y(_00500_),
    .A1(_04903_),
    .A2(_04904_));
 sg13g2_nand3_1 _26957_ (.B(_13707_),
    .C(_04882_),
    .A(_13706_),
    .Y(_04906_));
 sg13g2_a21o_1 _26958_ (.A2(_04882_),
    .A1(_13707_),
    .B1(_13706_),
    .X(_04907_));
 sg13g2_nand3_1 _26959_ (.B(_04906_),
    .C(_04907_),
    .A(net4657),
    .Y(_04908_));
 sg13g2_a21oi_1 _26960_ (.A1(net4541),
    .A2(\u_inv.d_next[225] ),
    .Y(_04909_),
    .B1(net3756));
 sg13g2_a21oi_1 _26961_ (.A1(_13708_),
    .A2(_04879_),
    .Y(_04910_),
    .B1(_13839_));
 sg13g2_o21ai_1 _26962_ (.B1(net3756),
    .Y(_04911_),
    .A1(_13706_),
    .A2(_04910_));
 sg13g2_a21oi_1 _26963_ (.A1(_13706_),
    .A2(_04910_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_a21oi_2 _26964_ (.B1(_04912_),
    .Y(_04913_),
    .A2(_04909_),
    .A1(_04908_));
 sg13g2_xnor2_1 _26965_ (.Y(_04914_),
    .A(net3472),
    .B(_04913_));
 sg13g2_a21oi_1 _26966_ (.A1(_04888_),
    .A2(_04901_),
    .Y(_04915_),
    .B1(_04887_));
 sg13g2_xor2_1 _26967_ (.B(_04915_),
    .A(_04914_),
    .X(_04916_));
 sg13g2_o21ai_1 _26968_ (.B1(net3882),
    .Y(_04917_),
    .A1(net4319),
    .A2(_04913_));
 sg13g2_a21oi_1 _26969_ (.A1(net4318),
    .A2(_04916_),
    .Y(_04918_),
    .B1(_04917_));
 sg13g2_a21o_1 _26970_ (.A2(net3932),
    .A1(net2449),
    .B1(_04918_),
    .X(_00501_));
 sg13g2_a21oi_1 _26971_ (.A1(_13709_),
    .A2(_04879_),
    .Y(_04919_),
    .B1(_13840_));
 sg13g2_nor2_1 _26972_ (.A(_13701_),
    .B(_04919_),
    .Y(_04920_));
 sg13g2_xnor2_1 _26973_ (.Y(_04921_),
    .A(_13701_),
    .B(_04919_));
 sg13g2_nand2_1 _26974_ (.Y(_04922_),
    .A(_15149_),
    .B(_04907_));
 sg13g2_xnor2_1 _26975_ (.Y(_04923_),
    .A(_13702_),
    .B(_04922_));
 sg13g2_nand2_1 _26976_ (.Y(_04924_),
    .A(net4657),
    .B(_04923_));
 sg13g2_a21oi_1 _26977_ (.A1(net4541),
    .A2(\u_inv.d_next[226] ),
    .Y(_04925_),
    .B1(net3756));
 sg13g2_a22oi_1 _26978_ (.Y(_04926_),
    .B1(_04924_),
    .B2(_04925_),
    .A2(_04921_),
    .A1(net3756));
 sg13g2_and2_1 _26979_ (.A(net3410),
    .B(_04926_),
    .X(_04927_));
 sg13g2_xnor2_1 _26980_ (.Y(_04928_),
    .A(net3410),
    .B(_04926_));
 sg13g2_a21oi_2 _26981_ (.B1(_04887_),
    .Y(_04929_),
    .A2(_04913_),
    .A1(net3410));
 sg13g2_nand3_1 _26982_ (.B(_04901_),
    .C(_04914_),
    .A(_04888_),
    .Y(_04930_));
 sg13g2_a21oi_1 _26983_ (.A1(_04929_),
    .A2(_04930_),
    .Y(_04931_),
    .B1(_04928_));
 sg13g2_nand3_1 _26984_ (.B(_04929_),
    .C(_04930_),
    .A(_04928_),
    .Y(_04932_));
 sg13g2_nand2b_1 _26985_ (.Y(_04933_),
    .B(_04932_),
    .A_N(_04931_));
 sg13g2_o21ai_1 _26986_ (.B1(net3882),
    .Y(_04934_),
    .A1(net4318),
    .A2(_04926_));
 sg13g2_a21oi_1 _26987_ (.A1(net4318),
    .A2(_04933_),
    .Y(_04935_),
    .B1(_04934_));
 sg13g2_a21o_1 _26988_ (.A2(net3932),
    .A1(net2895),
    .B1(_04935_),
    .X(_00502_));
 sg13g2_a21oi_1 _26989_ (.A1(net4540),
    .A2(\u_inv.d_next[227] ),
    .Y(_04936_),
    .B1(net3757));
 sg13g2_a21o_1 _26990_ (.A2(_04922_),
    .A1(_13701_),
    .B1(_13699_),
    .X(_04937_));
 sg13g2_xnor2_1 _26991_ (.Y(_04938_),
    .A(_13698_),
    .B(_04937_));
 sg13g2_nand2_1 _26992_ (.Y(_04939_),
    .A(net4657),
    .B(_04938_));
 sg13g2_nor2_1 _26993_ (.A(_13842_),
    .B(_04920_),
    .Y(_04940_));
 sg13g2_or2_1 _26994_ (.X(_04941_),
    .B(_04940_),
    .A(_13698_));
 sg13g2_a21oi_1 _26995_ (.A1(_13698_),
    .A2(_04940_),
    .Y(_04942_),
    .B1(net3835));
 sg13g2_a22oi_1 _26996_ (.Y(_04943_),
    .B1(_04941_),
    .B2(_04942_),
    .A2(_04939_),
    .A1(_04936_));
 sg13g2_xnor2_1 _26997_ (.Y(_04944_),
    .A(net3410),
    .B(_04943_));
 sg13g2_nor2_1 _26998_ (.A(_04927_),
    .B(_04931_),
    .Y(_04945_));
 sg13g2_xnor2_1 _26999_ (.Y(_04946_),
    .A(_04944_),
    .B(_04945_));
 sg13g2_o21ai_1 _27000_ (.B1(net3879),
    .Y(_04947_),
    .A1(net4318),
    .A2(_04943_));
 sg13g2_a21oi_1 _27001_ (.A1(net4318),
    .A2(_04946_),
    .Y(_04948_),
    .B1(_04947_));
 sg13g2_a21o_1 _27002_ (.A2(net3933),
    .A1(net3009),
    .B1(_04948_),
    .X(_00503_));
 sg13g2_o21ai_1 _27003_ (.B1(_13843_),
    .Y(_04949_),
    .A1(_13703_),
    .A2(_04919_));
 sg13g2_nand2_1 _27004_ (.Y(_04950_),
    .A(_13693_),
    .B(_04949_));
 sg13g2_xnor2_1 _27005_ (.Y(_04951_),
    .A(_13693_),
    .B(_04949_));
 sg13g2_o21ai_1 _27006_ (.B1(_15153_),
    .Y(_04952_),
    .A1(_15057_),
    .A2(_04881_));
 sg13g2_nand2_1 _27007_ (.Y(_04953_),
    .A(_13692_),
    .B(_04952_));
 sg13g2_o21ai_1 _27008_ (.B1(net4656),
    .Y(_04954_),
    .A1(_13692_),
    .A2(_04952_));
 sg13g2_nand2b_1 _27009_ (.Y(_04955_),
    .B(_04953_),
    .A_N(_04954_));
 sg13g2_a21oi_1 _27010_ (.A1(net4540),
    .A2(\u_inv.d_next[228] ),
    .Y(_04956_),
    .B1(net3757));
 sg13g2_a22oi_1 _27011_ (.Y(_04957_),
    .B1(_04955_),
    .B2(_04956_),
    .A2(_04951_),
    .A1(net3757));
 sg13g2_and2_1 _27012_ (.A(net3403),
    .B(_04957_),
    .X(_04958_));
 sg13g2_xnor2_1 _27013_ (.Y(_04959_),
    .A(net3403),
    .B(_04957_));
 sg13g2_inv_1 _27014_ (.Y(_04960_),
    .A(_04959_));
 sg13g2_a21o_1 _27015_ (.A2(_04943_),
    .A1(net3410),
    .B1(_04927_),
    .X(_04961_));
 sg13g2_nor2_1 _27016_ (.A(_04928_),
    .B(_04944_),
    .Y(_04962_));
 sg13g2_inv_1 _27017_ (.Y(_04963_),
    .A(_04962_));
 sg13g2_a21oi_1 _27018_ (.A1(_04929_),
    .A2(_04930_),
    .Y(_04964_),
    .B1(_04963_));
 sg13g2_o21ai_1 _27019_ (.B1(_04960_),
    .Y(_04965_),
    .A1(_04961_),
    .A2(_04964_));
 sg13g2_or3_1 _27020_ (.A(_04960_),
    .B(_04961_),
    .C(_04964_),
    .X(_04966_));
 sg13g2_nand2_1 _27021_ (.Y(_04967_),
    .A(_04965_),
    .B(_04966_));
 sg13g2_o21ai_1 _27022_ (.B1(net3880),
    .Y(_04968_),
    .A1(net4313),
    .A2(_04957_));
 sg13g2_a21oi_1 _27023_ (.A1(net4318),
    .A2(_04967_),
    .Y(_04969_),
    .B1(_04968_));
 sg13g2_a21o_1 _27024_ (.A2(net3932),
    .A1(net2752),
    .B1(_04969_),
    .X(_00504_));
 sg13g2_nand2_1 _27025_ (.Y(_04970_),
    .A(net2822),
    .B(net3932));
 sg13g2_nand3_1 _27026_ (.B(_13691_),
    .C(_04953_),
    .A(_13690_),
    .Y(_04971_));
 sg13g2_nand2_1 _27027_ (.Y(_04972_),
    .A(_15055_),
    .B(_04952_));
 sg13g2_nand4_1 _27028_ (.B(_15154_),
    .C(_04971_),
    .A(net4656),
    .Y(_04973_),
    .D(_04972_));
 sg13g2_a21oi_1 _27029_ (.A1(net4540),
    .A2(\u_inv.d_next[229] ),
    .Y(_04974_),
    .B1(net3757));
 sg13g2_and2_1 _27030_ (.A(_13847_),
    .B(_04950_),
    .X(_04975_));
 sg13g2_xor2_1 _27031_ (.B(_04975_),
    .A(_13690_),
    .X(_04976_));
 sg13g2_a22oi_1 _27032_ (.Y(_04977_),
    .B1(_04976_),
    .B2(net3757),
    .A2(_04974_),
    .A1(_04973_));
 sg13g2_inv_1 _27033_ (.Y(_04978_),
    .A(_04977_));
 sg13g2_xnor2_1 _27034_ (.Y(_04979_),
    .A(net3403),
    .B(_04977_));
 sg13g2_nand2b_1 _27035_ (.Y(_04980_),
    .B(_04965_),
    .A_N(_04958_));
 sg13g2_o21ai_1 _27036_ (.B1(net4313),
    .Y(_04981_),
    .A1(_04979_),
    .A2(_04980_));
 sg13g2_a21oi_1 _27037_ (.A1(_04979_),
    .A2(_04980_),
    .Y(_04982_),
    .B1(_04981_));
 sg13g2_o21ai_1 _27038_ (.B1(net3879),
    .Y(_04983_),
    .A1(net4313),
    .A2(_04977_));
 sg13g2_o21ai_1 _27039_ (.B1(_04970_),
    .Y(_00505_),
    .A1(_04982_),
    .A2(_04983_));
 sg13g2_a21oi_1 _27040_ (.A1(_13694_),
    .A2(_04949_),
    .Y(_04984_),
    .B1(_13848_));
 sg13g2_xnor2_1 _27041_ (.Y(_04985_),
    .A(_13685_),
    .B(_04984_));
 sg13g2_nand3_1 _27042_ (.B(_15156_),
    .C(_04972_),
    .A(_13686_),
    .Y(_04986_));
 sg13g2_a21o_1 _27043_ (.A2(_04972_),
    .A1(_15156_),
    .B1(_13686_),
    .X(_04987_));
 sg13g2_nand3_1 _27044_ (.B(_04986_),
    .C(_04987_),
    .A(net4656),
    .Y(_04988_));
 sg13g2_a21oi_1 _27045_ (.A1(net4540),
    .A2(\u_inv.d_next[230] ),
    .Y(_04989_),
    .B1(net3757));
 sg13g2_a22oi_1 _27046_ (.Y(_04990_),
    .B1(_04988_),
    .B2(_04989_),
    .A2(_04985_),
    .A1(net3757));
 sg13g2_and2_1 _27047_ (.A(net3404),
    .B(_04990_),
    .X(_04991_));
 sg13g2_nand2b_1 _27048_ (.Y(_04992_),
    .B(net3471),
    .A_N(_04990_));
 sg13g2_nand2b_1 _27049_ (.Y(_04993_),
    .B(_04992_),
    .A_N(_04991_));
 sg13g2_a21oi_1 _27050_ (.A1(net3403),
    .A2(_04977_),
    .Y(_04994_),
    .B1(_04958_));
 sg13g2_a22oi_1 _27051_ (.Y(_04995_),
    .B1(_04994_),
    .B2(_04965_),
    .A2(_04978_),
    .A1(net3471));
 sg13g2_xnor2_1 _27052_ (.Y(_04996_),
    .A(_04993_),
    .B(_04995_));
 sg13g2_nor2_1 _27053_ (.A(net4313),
    .B(_04990_),
    .Y(_04997_));
 sg13g2_o21ai_1 _27054_ (.B1(net3880),
    .Y(_04998_),
    .A1(net4292),
    .A2(_04996_));
 sg13g2_nand2_1 _27055_ (.Y(_04999_),
    .A(net2515),
    .B(net3932));
 sg13g2_o21ai_1 _27056_ (.B1(_04999_),
    .Y(_00506_),
    .A1(_04997_),
    .A2(_04998_));
 sg13g2_a21oi_1 _27057_ (.A1(net4540),
    .A2(\u_inv.d_next[231] ),
    .Y(_05000_),
    .B1(net3757));
 sg13g2_nand2_1 _27058_ (.Y(_05001_),
    .A(_13684_),
    .B(_04987_));
 sg13g2_xor2_1 _27059_ (.B(_05001_),
    .A(_13683_),
    .X(_05002_));
 sg13g2_nand2_1 _27060_ (.Y(_05003_),
    .A(net4656),
    .B(_05002_));
 sg13g2_o21ai_1 _27061_ (.B1(_13845_),
    .Y(_05004_),
    .A1(_13685_),
    .A2(_04984_));
 sg13g2_or2_1 _27062_ (.X(_05005_),
    .B(_05004_),
    .A(_13683_));
 sg13g2_a21oi_1 _27063_ (.A1(_13683_),
    .A2(_05004_),
    .Y(_05006_),
    .B1(net3835));
 sg13g2_a22oi_1 _27064_ (.Y(_05007_),
    .B1(_05005_),
    .B2(_05006_),
    .A2(_05003_),
    .A1(_05000_));
 sg13g2_xnor2_1 _27065_ (.Y(_05008_),
    .A(net3403),
    .B(_05007_));
 sg13g2_a21oi_1 _27066_ (.A1(_04992_),
    .A2(_04995_),
    .Y(_05009_),
    .B1(_04991_));
 sg13g2_xnor2_1 _27067_ (.Y(_05010_),
    .A(_05008_),
    .B(_05009_));
 sg13g2_o21ai_1 _27068_ (.B1(net3879),
    .Y(_05011_),
    .A1(net4313),
    .A2(_05007_));
 sg13g2_a21oi_1 _27069_ (.A1(net4313),
    .A2(_05010_),
    .Y(_05012_),
    .B1(_05011_));
 sg13g2_a21o_1 _27070_ (.A2(net3932),
    .A1(net3051),
    .B1(_05012_),
    .X(_00507_));
 sg13g2_a21oi_2 _27071_ (.B1(_13850_),
    .Y(_05013_),
    .A2(_04879_),
    .A1(_13710_));
 sg13g2_inv_1 _27072_ (.Y(_05014_),
    .A(_05013_));
 sg13g2_xor2_1 _27073_ (.B(_05013_),
    .A(_13661_),
    .X(_05015_));
 sg13g2_o21ai_1 _27074_ (.B1(_15161_),
    .Y(_05016_),
    .A1(_15058_),
    .A2(_04881_));
 sg13g2_nand2b_1 _27075_ (.Y(_05017_),
    .B(_05016_),
    .A_N(_13661_));
 sg13g2_nand2b_1 _27076_ (.Y(_05018_),
    .B(_13661_),
    .A_N(_05016_));
 sg13g2_nand3_1 _27077_ (.B(_05017_),
    .C(_05018_),
    .A(net4645),
    .Y(_05019_));
 sg13g2_a21oi_1 _27078_ (.A1(net4535),
    .A2(\u_inv.d_next[232] ),
    .Y(_05020_),
    .B1(net3748));
 sg13g2_a22oi_1 _27079_ (.Y(_05021_),
    .B1(_05019_),
    .B2(_05020_),
    .A2(_05015_),
    .A1(net3748));
 sg13g2_and2_1 _27080_ (.A(net3402),
    .B(_05021_),
    .X(_05022_));
 sg13g2_xnor2_1 _27081_ (.Y(_05023_),
    .A(net3402),
    .B(_05021_));
 sg13g2_or2_1 _27082_ (.X(_05024_),
    .B(_05008_),
    .A(_04993_));
 sg13g2_nor3_1 _27083_ (.A(_04959_),
    .B(_04979_),
    .C(_05024_),
    .Y(_05025_));
 sg13g2_nor3_1 _27084_ (.A(_04928_),
    .B(_04929_),
    .C(_04944_),
    .Y(_05026_));
 sg13g2_o21ai_1 _27085_ (.B1(_05025_),
    .Y(_05027_),
    .A1(_04961_),
    .A2(_05026_));
 sg13g2_a21oi_1 _27086_ (.A1(net3403),
    .A2(_05007_),
    .Y(_05028_),
    .B1(_04991_));
 sg13g2_o21ai_1 _27087_ (.B1(_05028_),
    .Y(_05029_),
    .A1(_04994_),
    .A2(_05024_));
 sg13g2_nand2b_2 _27088_ (.Y(_05030_),
    .B(_05027_),
    .A_N(_05029_));
 sg13g2_nand4_1 _27089_ (.B(_04914_),
    .C(_04962_),
    .A(_04888_),
    .Y(_05031_),
    .D(_05025_));
 sg13g2_inv_1 _27090_ (.Y(_05032_),
    .A(_05031_));
 sg13g2_a21oi_1 _27091_ (.A1(_04901_),
    .A2(_05032_),
    .Y(_05033_),
    .B1(_05030_));
 sg13g2_nor2_1 _27092_ (.A(_05023_),
    .B(_05033_),
    .Y(_05034_));
 sg13g2_xnor2_1 _27093_ (.Y(_05035_),
    .A(_05023_),
    .B(_05033_));
 sg13g2_o21ai_1 _27094_ (.B1(net3880),
    .Y(_05036_),
    .A1(net4312),
    .A2(_05021_));
 sg13g2_a21oi_1 _27095_ (.A1(net4312),
    .A2(_05035_),
    .Y(_05037_),
    .B1(_05036_));
 sg13g2_a21o_1 _27096_ (.A2(net3923),
    .A1(net3032),
    .B1(_05037_),
    .X(_00508_));
 sg13g2_nor2_1 _27097_ (.A(_05022_),
    .B(_05034_),
    .Y(_05038_));
 sg13g2_nand3_1 _27098_ (.B(_13664_),
    .C(_05017_),
    .A(_13660_),
    .Y(_05039_));
 sg13g2_nand2_1 _27099_ (.Y(_05040_),
    .A(_15052_),
    .B(_05016_));
 sg13g2_nor2_1 _27100_ (.A(net4532),
    .B(_15167_),
    .Y(_05041_));
 sg13g2_nand3_1 _27101_ (.B(_05040_),
    .C(_05041_),
    .A(_05039_),
    .Y(_05042_));
 sg13g2_a21oi_1 _27102_ (.A1(net4535),
    .A2(\u_inv.d_next[233] ),
    .Y(_05043_),
    .B1(net3748));
 sg13g2_a21o_1 _27103_ (.A2(_05014_),
    .A1(_13661_),
    .B1(_13834_),
    .X(_05044_));
 sg13g2_xnor2_1 _27104_ (.Y(_05045_),
    .A(_13664_),
    .B(_05044_));
 sg13g2_a22oi_1 _27105_ (.Y(_05046_),
    .B1(_05045_),
    .B2(net3748),
    .A2(_05043_),
    .A1(_05042_));
 sg13g2_xnor2_1 _27106_ (.Y(_05047_),
    .A(net3471),
    .B(_05046_));
 sg13g2_a21oi_1 _27107_ (.A1(_05038_),
    .A2(_05047_),
    .Y(_05048_),
    .B1(net4291));
 sg13g2_o21ai_1 _27108_ (.B1(_05048_),
    .Y(_05049_),
    .A1(_05038_),
    .A2(_05047_));
 sg13g2_nor2_1 _27109_ (.A(net4312),
    .B(_05046_),
    .Y(_05050_));
 sg13g2_nor2_1 _27110_ (.A(net4233),
    .B(_05050_),
    .Y(_05051_));
 sg13g2_a22oi_1 _27111_ (.Y(_05052_),
    .B1(_05049_),
    .B2(_05051_),
    .A2(net3924),
    .A1(net2519));
 sg13g2_inv_1 _27112_ (.Y(_00509_),
    .A(_05052_));
 sg13g2_and3_1 _27113_ (.X(_05053_),
    .A(_13661_),
    .B(_13662_),
    .C(_05014_));
 sg13g2_nor2_1 _27114_ (.A(_13836_),
    .B(_05053_),
    .Y(_05054_));
 sg13g2_o21ai_1 _27115_ (.B1(_13659_),
    .Y(_05055_),
    .A1(_13836_),
    .A2(_05053_));
 sg13g2_xnor2_1 _27116_ (.Y(_05056_),
    .A(_13659_),
    .B(_05054_));
 sg13g2_nand2_1 _27117_ (.Y(_05057_),
    .A(_15168_),
    .B(_05040_));
 sg13g2_nand2_1 _27118_ (.Y(_05058_),
    .A(_13658_),
    .B(_05057_));
 sg13g2_nand3_1 _27119_ (.B(_15168_),
    .C(_05040_),
    .A(_13659_),
    .Y(_05059_));
 sg13g2_and3_1 _27120_ (.X(_05060_),
    .A(net4645),
    .B(_05058_),
    .C(_05059_));
 sg13g2_a21oi_1 _27121_ (.A1(net4532),
    .A2(\u_inv.d_next[234] ),
    .Y(_05061_),
    .B1(net3747));
 sg13g2_nand2b_1 _27122_ (.Y(_05062_),
    .B(_05061_),
    .A_N(_05060_));
 sg13g2_o21ai_1 _27123_ (.B1(_05062_),
    .Y(_05063_),
    .A1(net3830),
    .A2(_05056_));
 sg13g2_nand2b_1 _27124_ (.Y(_05064_),
    .B(net3402),
    .A_N(_05063_));
 sg13g2_xnor2_1 _27125_ (.Y(_05065_),
    .A(net3471),
    .B(_05063_));
 sg13g2_a21o_1 _27126_ (.A2(_05046_),
    .A1(net3402),
    .B1(_05022_),
    .X(_05066_));
 sg13g2_nor2b_1 _27127_ (.A(_05023_),
    .B_N(_05047_),
    .Y(_05067_));
 sg13g2_inv_1 _27128_ (.Y(_05068_),
    .A(_05067_));
 sg13g2_a21oi_1 _27129_ (.A1(_05034_),
    .A2(_05047_),
    .Y(_05069_),
    .B1(_05066_));
 sg13g2_xnor2_1 _27130_ (.Y(_05070_),
    .A(_05065_),
    .B(_05069_));
 sg13g2_nand2_1 _27131_ (.Y(_05071_),
    .A(net4291),
    .B(_05063_));
 sg13g2_a21oi_1 _27132_ (.A1(net4314),
    .A2(_05070_),
    .Y(_05072_),
    .B1(net4233));
 sg13g2_a22oi_1 _27133_ (.Y(_05073_),
    .B1(_05071_),
    .B2(_05072_),
    .A2(net3924),
    .A1(net2918));
 sg13g2_inv_1 _27134_ (.Y(_00510_),
    .A(_05073_));
 sg13g2_a21oi_1 _27135_ (.A1(net4532),
    .A2(\u_inv.d_next[235] ),
    .Y(_05074_),
    .B1(net3748));
 sg13g2_nand2_1 _27136_ (.Y(_05075_),
    .A(_13657_),
    .B(_05058_));
 sg13g2_xnor2_1 _27137_ (.Y(_05076_),
    .A(_13667_),
    .B(_05075_));
 sg13g2_nand2_1 _27138_ (.Y(_05077_),
    .A(net4645),
    .B(_05076_));
 sg13g2_a21oi_1 _27139_ (.A1(_13833_),
    .A2(_05055_),
    .Y(_05078_),
    .B1(_13667_));
 sg13g2_nand3_1 _27140_ (.B(_13833_),
    .C(_05055_),
    .A(_13667_),
    .Y(_05079_));
 sg13g2_nor2_1 _27141_ (.A(net3830),
    .B(_05078_),
    .Y(_05080_));
 sg13g2_a22oi_1 _27142_ (.Y(_05081_),
    .B1(_05079_),
    .B2(_05080_),
    .A2(_05077_),
    .A1(_05074_));
 sg13g2_nand2_1 _27143_ (.Y(_05082_),
    .A(net3402),
    .B(_05081_));
 sg13g2_xnor2_1 _27144_ (.Y(_05083_),
    .A(net3403),
    .B(_05081_));
 sg13g2_o21ai_1 _27145_ (.B1(_05064_),
    .Y(_05084_),
    .A1(_05065_),
    .A2(_05069_));
 sg13g2_xor2_1 _27146_ (.B(_05084_),
    .A(_05083_),
    .X(_05085_));
 sg13g2_o21ai_1 _27147_ (.B1(net3878),
    .Y(_05086_),
    .A1(net4312),
    .A2(_05081_));
 sg13g2_a21oi_1 _27148_ (.A1(net4312),
    .A2(_05085_),
    .Y(_05087_),
    .B1(_05086_));
 sg13g2_a21o_1 _27149_ (.A2(net3923),
    .A1(net3035),
    .B1(_05087_),
    .X(_00511_));
 sg13g2_o21ai_1 _27150_ (.B1(_13838_),
    .Y(_05088_),
    .A1(_13668_),
    .A2(_05013_));
 sg13g2_xnor2_1 _27151_ (.Y(_05089_),
    .A(_13673_),
    .B(_05088_));
 sg13g2_a21oi_2 _27152_ (.B1(_15170_),
    .Y(_05090_),
    .A2(_05057_),
    .A1(_15051_));
 sg13g2_xor2_1 _27153_ (.B(_05090_),
    .A(_13673_),
    .X(_05091_));
 sg13g2_nand2_1 _27154_ (.Y(_05092_),
    .A(net4645),
    .B(_05091_));
 sg13g2_a21oi_1 _27155_ (.A1(net4532),
    .A2(\u_inv.d_next[236] ),
    .Y(_05093_),
    .B1(net3747));
 sg13g2_a22oi_1 _27156_ (.Y(_05094_),
    .B1(_05092_),
    .B2(_05093_),
    .A2(_05089_),
    .A1(net3747));
 sg13g2_and2_1 _27157_ (.A(net3402),
    .B(_05094_),
    .X(_05095_));
 sg13g2_xnor2_1 _27158_ (.Y(_05096_),
    .A(net3476),
    .B(_05094_));
 sg13g2_inv_1 _27159_ (.Y(_05097_),
    .A(_05096_));
 sg13g2_nor2_1 _27160_ (.A(_05065_),
    .B(_05083_),
    .Y(_05098_));
 sg13g2_nand2_1 _27161_ (.Y(_05099_),
    .A(_05066_),
    .B(_05098_));
 sg13g2_nand3_1 _27162_ (.B(_05082_),
    .C(_05099_),
    .A(_05064_),
    .Y(_05100_));
 sg13g2_nor4_1 _27163_ (.A(_05033_),
    .B(_05065_),
    .C(_05068_),
    .D(_05083_),
    .Y(_05101_));
 sg13g2_o21ai_1 _27164_ (.B1(_05096_),
    .Y(_05102_),
    .A1(_05100_),
    .A2(_05101_));
 sg13g2_or3_1 _27165_ (.A(_05096_),
    .B(_05100_),
    .C(_05101_),
    .X(_05103_));
 sg13g2_nand2_1 _27166_ (.Y(_05104_),
    .A(_05102_),
    .B(_05103_));
 sg13g2_o21ai_1 _27167_ (.B1(net3878),
    .Y(_05105_),
    .A1(net4312),
    .A2(_05094_));
 sg13g2_a21oi_1 _27168_ (.A1(net4312),
    .A2(_05104_),
    .Y(_05106_),
    .B1(_05105_));
 sg13g2_a21o_1 _27169_ (.A2(net3923),
    .A1(net2644),
    .B1(_05106_),
    .X(_00512_));
 sg13g2_nand2_1 _27170_ (.Y(_05107_),
    .A(net2194),
    .B(net3923));
 sg13g2_a21oi_1 _27171_ (.A1(net4532),
    .A2(\u_inv.d_next[237] ),
    .Y(_05108_),
    .B1(net3747));
 sg13g2_o21ai_1 _27172_ (.B1(_13672_),
    .Y(_05109_),
    .A1(_13673_),
    .A2(_05090_));
 sg13g2_xnor2_1 _27173_ (.Y(_05110_),
    .A(_13671_),
    .B(_05109_));
 sg13g2_nand2_1 _27174_ (.Y(_05111_),
    .A(net4645),
    .B(_05110_));
 sg13g2_a21oi_1 _27175_ (.A1(_13673_),
    .A2(_05088_),
    .Y(_05112_),
    .B1(_13855_));
 sg13g2_o21ai_1 _27176_ (.B1(net3747),
    .Y(_05113_),
    .A1(_13671_),
    .A2(_05112_));
 sg13g2_a21oi_1 _27177_ (.A1(_13671_),
    .A2(_05112_),
    .Y(_05114_),
    .B1(_05113_));
 sg13g2_a21oi_2 _27178_ (.B1(_05114_),
    .Y(_05115_),
    .A2(_05111_),
    .A1(_05108_));
 sg13g2_xnor2_1 _27179_ (.Y(_05116_),
    .A(net3402),
    .B(_05115_));
 sg13g2_nand2b_1 _27180_ (.Y(_05117_),
    .B(_05102_),
    .A_N(_05095_));
 sg13g2_o21ai_1 _27181_ (.B1(net4312),
    .Y(_05118_),
    .A1(_05116_),
    .A2(_05117_));
 sg13g2_a21oi_1 _27182_ (.A1(_05116_),
    .A2(_05117_),
    .Y(_05119_),
    .B1(_05118_));
 sg13g2_o21ai_1 _27183_ (.B1(net3878),
    .Y(_05120_),
    .A1(net4310),
    .A2(_05115_));
 sg13g2_o21ai_1 _27184_ (.B1(_05107_),
    .Y(_00513_),
    .A1(_05119_),
    .A2(_05120_));
 sg13g2_a21oi_1 _27185_ (.A1(_13674_),
    .A2(_05088_),
    .Y(_05121_),
    .B1(_13856_));
 sg13g2_xnor2_1 _27186_ (.Y(_05122_),
    .A(_13679_),
    .B(_05121_));
 sg13g2_o21ai_1 _27187_ (.B1(_15163_),
    .Y(_05123_),
    .A1(_15049_),
    .A2(_05090_));
 sg13g2_xor2_1 _27188_ (.B(_05123_),
    .A(_13679_),
    .X(_05124_));
 sg13g2_nand2_1 _27189_ (.Y(_05125_),
    .A(net4645),
    .B(_05124_));
 sg13g2_a21oi_1 _27190_ (.A1(net4532),
    .A2(\u_inv.d_next[238] ),
    .Y(_05126_),
    .B1(net3747));
 sg13g2_a22oi_1 _27191_ (.Y(_05127_),
    .B1(_05125_),
    .B2(_05126_),
    .A2(_05122_),
    .A1(net3747));
 sg13g2_and2_1 _27192_ (.A(net3401),
    .B(_05127_),
    .X(_05128_));
 sg13g2_xnor2_1 _27193_ (.Y(_05129_),
    .A(net3400),
    .B(_05127_));
 sg13g2_inv_1 _27194_ (.Y(_05130_),
    .A(_05129_));
 sg13g2_a21oi_1 _27195_ (.A1(net3402),
    .A2(_05115_),
    .Y(_05131_),
    .B1(_05095_));
 sg13g2_o21ai_1 _27196_ (.B1(_05131_),
    .Y(_05132_),
    .A1(_05102_),
    .A2(_05116_));
 sg13g2_xnor2_1 _27197_ (.Y(_05133_),
    .A(_05130_),
    .B(_05132_));
 sg13g2_o21ai_1 _27198_ (.B1(net3878),
    .Y(_05134_),
    .A1(net4309),
    .A2(_05127_));
 sg13g2_a21oi_1 _27199_ (.A1(net4310),
    .A2(_05133_),
    .Y(_05135_),
    .B1(_05134_));
 sg13g2_a21o_1 _27200_ (.A2(net3923),
    .A1(net2390),
    .B1(_05135_),
    .X(_00514_));
 sg13g2_a21oi_1 _27201_ (.A1(net4532),
    .A2(\u_inv.d_next[239] ),
    .Y(_05136_),
    .B1(net3747));
 sg13g2_a21oi_1 _27202_ (.A1(_13679_),
    .A2(_05123_),
    .Y(_05137_),
    .B1(_13678_));
 sg13g2_xor2_1 _27203_ (.B(_05137_),
    .A(_13677_),
    .X(_05138_));
 sg13g2_o21ai_1 _27204_ (.B1(_05136_),
    .Y(_05139_),
    .A1(net4532),
    .A2(_05138_));
 sg13g2_o21ai_1 _27205_ (.B1(_13851_),
    .Y(_05140_),
    .A1(_13679_),
    .A2(_05121_));
 sg13g2_a21oi_1 _27206_ (.A1(_13677_),
    .A2(_05140_),
    .Y(_05141_),
    .B1(net3830));
 sg13g2_o21ai_1 _27207_ (.B1(_05141_),
    .Y(_05142_),
    .A1(_13677_),
    .A2(_05140_));
 sg13g2_and2_1 _27208_ (.A(_05139_),
    .B(_05142_),
    .X(_05143_));
 sg13g2_xnor2_1 _27209_ (.Y(_05144_),
    .A(net3400),
    .B(_05143_));
 sg13g2_a21oi_1 _27210_ (.A1(_05130_),
    .A2(_05132_),
    .Y(_05145_),
    .B1(_05128_));
 sg13g2_xnor2_1 _27211_ (.Y(_05146_),
    .A(_05144_),
    .B(_05145_));
 sg13g2_o21ai_1 _27212_ (.B1(net3878),
    .Y(_05147_),
    .A1(net4310),
    .A2(_05143_));
 sg13g2_a21oi_1 _27213_ (.A1(net4310),
    .A2(_05146_),
    .Y(_05148_),
    .B1(_05147_));
 sg13g2_a21o_1 _27214_ (.A2(net3923),
    .A1(net2669),
    .B1(_05148_),
    .X(_00515_));
 sg13g2_a21oi_2 _27215_ (.B1(_13860_),
    .Y(_05149_),
    .A2(_04879_),
    .A1(_13712_));
 sg13g2_or2_1 _27216_ (.X(_05150_),
    .B(_05149_),
    .A(_13654_));
 sg13g2_xnor2_1 _27217_ (.Y(_05151_),
    .A(_13654_),
    .B(_05149_));
 sg13g2_o21ai_1 _27218_ (.B1(_15173_),
    .Y(_05152_),
    .A1(_15059_),
    .A2(_04881_));
 sg13g2_o21ai_1 _27219_ (.B1(net4643),
    .Y(_05153_),
    .A1(_13654_),
    .A2(_05152_));
 sg13g2_a21o_1 _27220_ (.A2(_05152_),
    .A1(_13654_),
    .B1(_05153_),
    .X(_05154_));
 sg13g2_a21oi_1 _27221_ (.A1(net4531),
    .A2(\u_inv.d_next[240] ),
    .Y(_05155_),
    .B1(net3745));
 sg13g2_a22oi_1 _27222_ (.Y(_05156_),
    .B1(_05154_),
    .B2(_05155_),
    .A2(_05151_),
    .A1(net3745));
 sg13g2_and2_1 _27223_ (.A(net3400),
    .B(_05156_),
    .X(_05157_));
 sg13g2_xnor2_1 _27224_ (.Y(_05158_),
    .A(net3400),
    .B(_05156_));
 sg13g2_or4_1 _27225_ (.A(_05097_),
    .B(_05116_),
    .C(_05129_),
    .D(_05144_),
    .X(_05159_));
 sg13g2_inv_1 _27226_ (.Y(_05160_),
    .A(_05159_));
 sg13g2_nand2_1 _27227_ (.Y(_05161_),
    .A(_05067_),
    .B(_05098_));
 sg13g2_nor2_1 _27228_ (.A(_05159_),
    .B(_05161_),
    .Y(_05162_));
 sg13g2_nor3_1 _27229_ (.A(_05031_),
    .B(_05159_),
    .C(_05161_),
    .Y(_05163_));
 sg13g2_nand2_1 _27230_ (.Y(_05164_),
    .A(_05032_),
    .B(_05162_));
 sg13g2_nor3_1 _27231_ (.A(_05129_),
    .B(_05131_),
    .C(_05144_),
    .Y(_05165_));
 sg13g2_a21oi_1 _27232_ (.A1(net3401),
    .A2(_05143_),
    .Y(_05166_),
    .B1(_05128_));
 sg13g2_nand2b_1 _27233_ (.Y(_05167_),
    .B(_05166_),
    .A_N(_05165_));
 sg13g2_a21o_1 _27234_ (.A2(_05160_),
    .A1(_05100_),
    .B1(_05167_),
    .X(_05168_));
 sg13g2_a221oi_1 _27235_ (.B2(_05030_),
    .C1(_05167_),
    .B1(_05162_),
    .A1(_05100_),
    .Y(_05169_),
    .A2(_05160_));
 sg13g2_a221oi_1 _27236_ (.B2(_04901_),
    .C1(_05168_),
    .B1(_05163_),
    .A1(_05030_),
    .Y(_05170_),
    .A2(_05162_));
 sg13g2_o21ai_1 _27237_ (.B1(_05169_),
    .Y(_05171_),
    .A1(_04900_),
    .A2(_05164_));
 sg13g2_nor2_1 _27238_ (.A(_05158_),
    .B(_05170_),
    .Y(_05172_));
 sg13g2_xnor2_1 _27239_ (.Y(_05173_),
    .A(_05158_),
    .B(_05170_));
 sg13g2_o21ai_1 _27240_ (.B1(net3878),
    .Y(_05174_),
    .A1(net4309),
    .A2(_05156_));
 sg13g2_a21oi_1 _27241_ (.A1(net4309),
    .A2(_05173_),
    .Y(_05175_),
    .B1(_05174_));
 sg13g2_a21o_1 _27242_ (.A2(net3923),
    .A1(net3045),
    .B1(_05175_),
    .X(_00516_));
 sg13g2_nand2_1 _27243_ (.Y(_05176_),
    .A(net2230),
    .B(net3921));
 sg13g2_a21oi_1 _27244_ (.A1(_13654_),
    .A2(_05152_),
    .Y(_05177_),
    .B1(_13636_));
 sg13g2_nand2_1 _27245_ (.Y(_05178_),
    .A(_13653_),
    .B(_05177_));
 sg13g2_nand3_1 _27246_ (.B(_13654_),
    .C(_05152_),
    .A(_13636_),
    .Y(_05179_));
 sg13g2_nand4_1 _27247_ (.B(_15139_),
    .C(_05178_),
    .A(net4643),
    .Y(_05180_),
    .D(_05179_));
 sg13g2_a21oi_1 _27248_ (.A1(net4530),
    .A2(\u_inv.d_next[241] ),
    .Y(_05181_),
    .B1(net3745));
 sg13g2_nand2b_1 _27249_ (.Y(_05182_),
    .B(_05150_),
    .A_N(_13865_));
 sg13g2_xnor2_1 _27250_ (.Y(_05183_),
    .A(_13635_),
    .B(_05182_));
 sg13g2_a22oi_1 _27251_ (.Y(_05184_),
    .B1(_05183_),
    .B2(net3745),
    .A2(_05181_),
    .A1(_05180_));
 sg13g2_xnor2_1 _27252_ (.Y(_05185_),
    .A(net3471),
    .B(_05184_));
 sg13g2_nor2_1 _27253_ (.A(_05157_),
    .B(_05172_),
    .Y(_05186_));
 sg13g2_o21ai_1 _27254_ (.B1(net4309),
    .Y(_05187_),
    .A1(_05185_),
    .A2(_05186_));
 sg13g2_a21oi_1 _27255_ (.A1(_05185_),
    .A2(_05186_),
    .Y(_05188_),
    .B1(_05187_));
 sg13g2_o21ai_1 _27256_ (.B1(net3878),
    .Y(_05189_),
    .A1(net4309),
    .A2(_05184_));
 sg13g2_o21ai_1 _27257_ (.B1(_05176_),
    .Y(_00517_),
    .A1(_05188_),
    .A2(_05189_));
 sg13g2_o21ai_1 _27258_ (.B1(_13632_),
    .Y(_05190_),
    .A1(_13633_),
    .A2(_05182_));
 sg13g2_xnor2_1 _27259_ (.Y(_05191_),
    .A(_13631_),
    .B(_05190_));
 sg13g2_nand2_1 _27260_ (.Y(_05192_),
    .A(_15140_),
    .B(_05179_));
 sg13g2_nand2_1 _27261_ (.Y(_05193_),
    .A(_13631_),
    .B(_05192_));
 sg13g2_nand3_1 _27262_ (.B(_15140_),
    .C(_05179_),
    .A(_13630_),
    .Y(_05194_));
 sg13g2_nand3_1 _27263_ (.B(_05193_),
    .C(_05194_),
    .A(net4643),
    .Y(_05195_));
 sg13g2_a21oi_1 _27264_ (.A1(net4531),
    .A2(\u_inv.d_next[242] ),
    .Y(_05196_),
    .B1(net3745));
 sg13g2_a22oi_1 _27265_ (.Y(_05197_),
    .B1(_05195_),
    .B2(_05196_),
    .A2(_05191_),
    .A1(net3745));
 sg13g2_nand2_1 _27266_ (.Y(_05198_),
    .A(net3400),
    .B(_05197_));
 sg13g2_xnor2_1 _27267_ (.Y(_05199_),
    .A(net3471),
    .B(_05197_));
 sg13g2_inv_1 _27268_ (.Y(_05200_),
    .A(_05199_));
 sg13g2_a21o_1 _27269_ (.A2(_05184_),
    .A1(net3400),
    .B1(_05157_),
    .X(_05201_));
 sg13g2_nand2b_1 _27270_ (.Y(_05202_),
    .B(_05185_),
    .A_N(_05158_));
 sg13g2_a21oi_1 _27271_ (.A1(_05172_),
    .A2(_05185_),
    .Y(_05203_),
    .B1(_05201_));
 sg13g2_xnor2_1 _27272_ (.Y(_05204_),
    .A(_05199_),
    .B(_05203_));
 sg13g2_nor2_1 _27273_ (.A(net4309),
    .B(_05197_),
    .Y(_05205_));
 sg13g2_o21ai_1 _27274_ (.B1(net3878),
    .Y(_05206_),
    .A1(net4291),
    .A2(_05204_));
 sg13g2_nand2_1 _27275_ (.Y(_05207_),
    .A(net2088),
    .B(net3921));
 sg13g2_o21ai_1 _27276_ (.B1(_05207_),
    .Y(_00518_),
    .A1(_05205_),
    .A2(_05206_));
 sg13g2_a21oi_1 _27277_ (.A1(net4530),
    .A2(\u_inv.d_next[243] ),
    .Y(_05208_),
    .B1(net3744));
 sg13g2_nand2_1 _27278_ (.Y(_05209_),
    .A(_13629_),
    .B(_05193_));
 sg13g2_xnor2_1 _27279_ (.Y(_05210_),
    .A(_13639_),
    .B(_05209_));
 sg13g2_nand2_1 _27280_ (.Y(_05211_),
    .A(net4643),
    .B(_05210_));
 sg13g2_o21ai_1 _27281_ (.B1(_13864_),
    .Y(_05212_),
    .A1(_13631_),
    .A2(_05190_));
 sg13g2_nand2b_1 _27282_ (.Y(_05213_),
    .B(_13639_),
    .A_N(_05212_));
 sg13g2_a21oi_1 _27283_ (.A1(_13640_),
    .A2(_05212_),
    .Y(_05214_),
    .B1(net3829));
 sg13g2_a22oi_1 _27284_ (.Y(_05215_),
    .B1(_05213_),
    .B2(_05214_),
    .A2(_05211_),
    .A1(_05208_));
 sg13g2_xnor2_1 _27285_ (.Y(_05216_),
    .A(net3400),
    .B(_05215_));
 sg13g2_o21ai_1 _27286_ (.B1(_05198_),
    .Y(_05217_),
    .A1(_05200_),
    .A2(_05203_));
 sg13g2_xor2_1 _27287_ (.B(_05217_),
    .A(_05216_),
    .X(_05218_));
 sg13g2_o21ai_1 _27288_ (.B1(net3875),
    .Y(_05219_),
    .A1(net4309),
    .A2(_05215_));
 sg13g2_a21oi_1 _27289_ (.A1(net4309),
    .A2(_05218_),
    .Y(_05220_),
    .B1(_05219_));
 sg13g2_a21o_1 _27290_ (.A2(net3921),
    .A1(net2758),
    .B1(_05220_),
    .X(_00519_));
 sg13g2_or2_1 _27291_ (.X(_05221_),
    .B(_05150_),
    .A(_13641_));
 sg13g2_nand2_1 _27292_ (.Y(_05222_),
    .A(_13868_),
    .B(_05221_));
 sg13g2_xnor2_1 _27293_ (.Y(_05223_),
    .A(_13644_),
    .B(_05222_));
 sg13g2_a21oi_2 _27294_ (.B1(_15137_),
    .Y(_05224_),
    .A2(_05192_),
    .A1(_15043_));
 sg13g2_a21oi_1 _27295_ (.A1(_13644_),
    .A2(_05224_),
    .Y(_05225_),
    .B1(net4530));
 sg13g2_o21ai_1 _27296_ (.B1(_05225_),
    .Y(_05226_),
    .A1(_13644_),
    .A2(_05224_));
 sg13g2_a21oi_1 _27297_ (.A1(net4530),
    .A2(\u_inv.d_next[244] ),
    .Y(_05227_),
    .B1(net3744));
 sg13g2_a22oi_1 _27298_ (.Y(_05228_),
    .B1(_05226_),
    .B2(_05227_),
    .A2(_05223_),
    .A1(net3745));
 sg13g2_and2_1 _27299_ (.A(net3396),
    .B(_05228_),
    .X(_05229_));
 sg13g2_xnor2_1 _27300_ (.Y(_05230_),
    .A(net3396),
    .B(_05228_));
 sg13g2_inv_1 _27301_ (.Y(_05231_),
    .A(_05230_));
 sg13g2_or2_1 _27302_ (.X(_05232_),
    .B(_05216_),
    .A(_05200_));
 sg13g2_nand2b_1 _27303_ (.Y(_05233_),
    .B(_05201_),
    .A_N(_05232_));
 sg13g2_o21ai_1 _27304_ (.B1(net3400),
    .Y(_05234_),
    .A1(_05197_),
    .A2(_05215_));
 sg13g2_nand2_1 _27305_ (.Y(_05235_),
    .A(_05233_),
    .B(_05234_));
 sg13g2_nor3_1 _27306_ (.A(_05170_),
    .B(_05202_),
    .C(_05232_),
    .Y(_05236_));
 sg13g2_o21ai_1 _27307_ (.B1(_05231_),
    .Y(_05237_),
    .A1(_05235_),
    .A2(_05236_));
 sg13g2_or3_1 _27308_ (.A(_05231_),
    .B(_05235_),
    .C(_05236_),
    .X(_05238_));
 sg13g2_nand2_1 _27309_ (.Y(_05239_),
    .A(_05237_),
    .B(_05238_));
 sg13g2_o21ai_1 _27310_ (.B1(net3875),
    .Y(_05240_),
    .A1(net4302),
    .A2(_05228_));
 sg13g2_a21oi_1 _27311_ (.A1(net4303),
    .A2(_05239_),
    .Y(_05241_),
    .B1(_05240_));
 sg13g2_a21o_1 _27312_ (.A2(net3921),
    .A1(net2850),
    .B1(_05241_),
    .X(_00520_));
 sg13g2_nand2_1 _27313_ (.Y(_05242_),
    .A(net2127),
    .B(net3921));
 sg13g2_a21oi_1 _27314_ (.A1(net4530),
    .A2(\u_inv.d_next[245] ),
    .Y(_05243_),
    .B1(net3744));
 sg13g2_o21ai_1 _27315_ (.B1(_13643_),
    .Y(_05244_),
    .A1(_13644_),
    .A2(_05224_));
 sg13g2_xnor2_1 _27316_ (.Y(_05245_),
    .A(_13642_),
    .B(_05244_));
 sg13g2_nand2_1 _27317_ (.Y(_05246_),
    .A(net4643),
    .B(_05245_));
 sg13g2_a21oi_1 _27318_ (.A1(_13644_),
    .A2(_05222_),
    .Y(_05247_),
    .B1(_13872_));
 sg13g2_o21ai_1 _27319_ (.B1(net3744),
    .Y(_05248_),
    .A1(_13642_),
    .A2(_05247_));
 sg13g2_a21oi_1 _27320_ (.A1(_13642_),
    .A2(_05247_),
    .Y(_05249_),
    .B1(_05248_));
 sg13g2_a21oi_1 _27321_ (.A1(_05243_),
    .A2(_05246_),
    .Y(_05250_),
    .B1(_05249_));
 sg13g2_xnor2_1 _27322_ (.Y(_05251_),
    .A(net3395),
    .B(_05250_));
 sg13g2_nand2b_1 _27323_ (.Y(_05252_),
    .B(_05237_),
    .A_N(_05229_));
 sg13g2_o21ai_1 _27324_ (.B1(net4303),
    .Y(_05253_),
    .A1(_05251_),
    .A2(_05252_));
 sg13g2_a21oi_1 _27325_ (.A1(_05251_),
    .A2(_05252_),
    .Y(_05254_),
    .B1(_05253_));
 sg13g2_o21ai_1 _27326_ (.B1(net3875),
    .Y(_05255_),
    .A1(net4302),
    .A2(_05250_));
 sg13g2_o21ai_1 _27327_ (.B1(_05242_),
    .Y(_00521_),
    .A1(_05254_),
    .A2(_05255_));
 sg13g2_a21oi_1 _27328_ (.A1(_13645_),
    .A2(_05222_),
    .Y(_05256_),
    .B1(_13874_));
 sg13g2_xnor2_1 _27329_ (.Y(_05257_),
    .A(_13650_),
    .B(_05256_));
 sg13g2_o21ai_1 _27330_ (.B1(_15136_),
    .Y(_05258_),
    .A1(_15042_),
    .A2(_05224_));
 sg13g2_o21ai_1 _27331_ (.B1(net4643),
    .Y(_05259_),
    .A1(_13650_),
    .A2(_05258_));
 sg13g2_a21o_1 _27332_ (.A2(_05258_),
    .A1(_13650_),
    .B1(_05259_),
    .X(_05260_));
 sg13g2_a21oi_1 _27333_ (.A1(net4530),
    .A2(\u_inv.d_next[246] ),
    .Y(_05261_),
    .B1(net3744));
 sg13g2_a22oi_1 _27334_ (.Y(_05262_),
    .B1(_05260_),
    .B2(_05261_),
    .A2(_05257_),
    .A1(net3744));
 sg13g2_and2_1 _27335_ (.A(net3395),
    .B(_05262_),
    .X(_05263_));
 sg13g2_xnor2_1 _27336_ (.Y(_05264_),
    .A(net3396),
    .B(_05262_));
 sg13g2_inv_1 _27337_ (.Y(_05265_),
    .A(_05264_));
 sg13g2_a21oi_1 _27338_ (.A1(net3396),
    .A2(_05250_),
    .Y(_05266_),
    .B1(_05229_));
 sg13g2_o21ai_1 _27339_ (.B1(_05266_),
    .Y(_05267_),
    .A1(_05237_),
    .A2(_05251_));
 sg13g2_xnor2_1 _27340_ (.Y(_05268_),
    .A(_05265_),
    .B(_05267_));
 sg13g2_a21oi_1 _27341_ (.A1(net4302),
    .A2(_05268_),
    .Y(_05269_),
    .B1(net4232));
 sg13g2_o21ai_1 _27342_ (.B1(_05269_),
    .Y(_05270_),
    .A1(net4303),
    .A2(_05262_));
 sg13g2_o21ai_1 _27343_ (.B1(_05270_),
    .Y(_00522_),
    .A1(_10578_),
    .A2(net4013));
 sg13g2_a21oi_1 _27344_ (.A1(net4530),
    .A2(\u_inv.d_next[247] ),
    .Y(_05271_),
    .B1(net3744));
 sg13g2_a21oi_1 _27345_ (.A1(_13650_),
    .A2(_05258_),
    .Y(_05272_),
    .B1(_13649_));
 sg13g2_a21oi_1 _27346_ (.A1(_13648_),
    .A2(_05272_),
    .Y(_05273_),
    .B1(net4530));
 sg13g2_o21ai_1 _27347_ (.B1(_05273_),
    .Y(_05274_),
    .A1(_13648_),
    .A2(_05272_));
 sg13g2_o21ai_1 _27348_ (.B1(_13871_),
    .Y(_05275_),
    .A1(_13650_),
    .A2(_05256_));
 sg13g2_o21ai_1 _27349_ (.B1(net3744),
    .Y(_05276_),
    .A1(_13647_),
    .A2(_05275_));
 sg13g2_a21oi_1 _27350_ (.A1(_13647_),
    .A2(_05275_),
    .Y(_05277_),
    .B1(_05276_));
 sg13g2_a21oi_1 _27351_ (.A1(_05271_),
    .A2(_05274_),
    .Y(_05278_),
    .B1(_05277_));
 sg13g2_xnor2_1 _27352_ (.Y(_05279_),
    .A(net3395),
    .B(_05278_));
 sg13g2_a21oi_1 _27353_ (.A1(_05265_),
    .A2(_05267_),
    .Y(_05280_),
    .B1(_05263_));
 sg13g2_xnor2_1 _27354_ (.Y(_05281_),
    .A(_05279_),
    .B(_05280_));
 sg13g2_o21ai_1 _27355_ (.B1(net3875),
    .Y(_05282_),
    .A1(net4302),
    .A2(_05278_));
 sg13g2_a21oi_1 _27356_ (.A1(net4303),
    .A2(_05281_),
    .Y(_05283_),
    .B1(_05282_));
 sg13g2_a21o_1 _27357_ (.A2(net3921),
    .A1(net3073),
    .B1(_05283_),
    .X(_00523_));
 sg13g2_o21ai_1 _27358_ (.B1(_13877_),
    .Y(_05284_),
    .A1(_13652_),
    .A2(_05221_));
 sg13g2_xnor2_1 _27359_ (.Y(_05285_),
    .A(_13625_),
    .B(_05284_));
 sg13g2_a21oi_2 _27360_ (.B1(_15147_),
    .Y(_05286_),
    .A2(_05152_),
    .A1(_15046_));
 sg13g2_a21oi_1 _27361_ (.A1(_13625_),
    .A2(_05286_),
    .Y(_05287_),
    .B1(net4523));
 sg13g2_o21ai_1 _27362_ (.B1(_05287_),
    .Y(_05288_),
    .A1(_13625_),
    .A2(_05286_));
 sg13g2_a21oi_1 _27363_ (.A1(net4523),
    .A2(\u_inv.d_next[248] ),
    .Y(_05289_),
    .B1(net3738));
 sg13g2_a22oi_1 _27364_ (.Y(_05290_),
    .B1(_05288_),
    .B2(_05289_),
    .A2(_05285_),
    .A1(net3738));
 sg13g2_nand2_1 _27365_ (.Y(_05291_),
    .A(net3395),
    .B(_05290_));
 sg13g2_xnor2_1 _27366_ (.Y(_05292_),
    .A(net3395),
    .B(_05290_));
 sg13g2_nor2_1 _27367_ (.A(_05264_),
    .B(_05279_),
    .Y(_05293_));
 sg13g2_or4_1 _27368_ (.A(_05230_),
    .B(_05251_),
    .C(_05264_),
    .D(_05279_),
    .X(_05294_));
 sg13g2_nor3_1 _27369_ (.A(_05202_),
    .B(_05232_),
    .C(_05294_),
    .Y(_05295_));
 sg13g2_nand2b_1 _27370_ (.Y(_05296_),
    .B(_05235_),
    .A_N(_05294_));
 sg13g2_a21oi_1 _27371_ (.A1(net3395),
    .A2(_05278_),
    .Y(_05297_),
    .B1(_05263_));
 sg13g2_nand2b_1 _27372_ (.Y(_05298_),
    .B(_05293_),
    .A_N(_05266_));
 sg13g2_nand3_1 _27373_ (.B(_05297_),
    .C(_05298_),
    .A(_05296_),
    .Y(_05299_));
 sg13g2_a21oi_2 _27374_ (.B1(_05299_),
    .Y(_05300_),
    .A2(_05295_),
    .A1(_05171_));
 sg13g2_nor2_1 _27375_ (.A(_05292_),
    .B(_05300_),
    .Y(_05301_));
 sg13g2_xnor2_1 _27376_ (.Y(_05302_),
    .A(_05292_),
    .B(_05300_));
 sg13g2_o21ai_1 _27377_ (.B1(net3875),
    .Y(_05303_),
    .A1(net4302),
    .A2(_05290_));
 sg13g2_a21oi_1 _27378_ (.A1(net4302),
    .A2(_05302_),
    .Y(_05304_),
    .B1(_05303_));
 sg13g2_a21o_1 _27379_ (.A2(net3912),
    .A1(net3131),
    .B1(_05304_),
    .X(_00524_));
 sg13g2_nand2b_1 _27380_ (.Y(_05305_),
    .B(net3823),
    .A_N(\u_inv.d_next[249] ));
 sg13g2_o21ai_1 _27381_ (.B1(_13624_),
    .Y(_05306_),
    .A1(_13625_),
    .A2(_05286_));
 sg13g2_xnor2_1 _27382_ (.Y(_05307_),
    .A(_13623_),
    .B(_05306_));
 sg13g2_a22oi_1 _27383_ (.Y(_05308_),
    .B1(_05307_),
    .B2(net4634),
    .A2(_05305_),
    .A1(net3723));
 sg13g2_a21oi_1 _27384_ (.A1(_13625_),
    .A2(_05284_),
    .Y(_05309_),
    .B1(_13890_));
 sg13g2_o21ai_1 _27385_ (.B1(net3738),
    .Y(_05310_),
    .A1(_13623_),
    .A2(_05309_));
 sg13g2_a21oi_1 _27386_ (.A1(_13623_),
    .A2(_05309_),
    .Y(_05311_),
    .B1(_05310_));
 sg13g2_nor2_1 _27387_ (.A(_05308_),
    .B(_05311_),
    .Y(_05312_));
 sg13g2_nand2_1 _27388_ (.Y(_05313_),
    .A(net3395),
    .B(_05312_));
 sg13g2_nand2b_1 _27389_ (.Y(_05314_),
    .B(net3470),
    .A_N(_05312_));
 sg13g2_nand2_1 _27390_ (.Y(_05315_),
    .A(_05313_),
    .B(_05314_));
 sg13g2_o21ai_1 _27391_ (.B1(_05291_),
    .Y(_05316_),
    .A1(_05292_),
    .A2(_05300_));
 sg13g2_xor2_1 _27392_ (.B(_05316_),
    .A(_05315_),
    .X(_05317_));
 sg13g2_o21ai_1 _27393_ (.B1(net3875),
    .Y(_05318_),
    .A1(net4302),
    .A2(_05312_));
 sg13g2_a21oi_1 _27394_ (.A1(net4302),
    .A2(_05317_),
    .Y(_05319_),
    .B1(_05318_));
 sg13g2_a21o_1 _27395_ (.A2(net3912),
    .A1(net2388),
    .B1(_05319_),
    .X(_00525_));
 sg13g2_a21oi_1 _27396_ (.A1(_13626_),
    .A2(_05284_),
    .Y(_05320_),
    .B1(_13891_));
 sg13g2_nor2_1 _27397_ (.A(_13618_),
    .B(_05320_),
    .Y(_05321_));
 sg13g2_xnor2_1 _27398_ (.Y(_05322_),
    .A(_13618_),
    .B(_05320_));
 sg13g2_nor2_1 _27399_ (.A(_15040_),
    .B(_05286_),
    .Y(_05323_));
 sg13g2_nor2_2 _27400_ (.A(_15178_),
    .B(_05323_),
    .Y(_05324_));
 sg13g2_inv_1 _27401_ (.Y(_05325_),
    .A(_05324_));
 sg13g2_a21oi_1 _27402_ (.A1(_13619_),
    .A2(_05324_),
    .Y(_05326_),
    .B1(net4522));
 sg13g2_o21ai_1 _27403_ (.B1(_05326_),
    .Y(_05327_),
    .A1(_13619_),
    .A2(_05324_));
 sg13g2_a21oi_1 _27404_ (.A1(net4523),
    .A2(\u_inv.d_next[250] ),
    .Y(_05328_),
    .B1(net3737));
 sg13g2_a22oi_1 _27405_ (.Y(_05329_),
    .B1(_05327_),
    .B2(_05328_),
    .A2(_05322_),
    .A1(net3738));
 sg13g2_nand2_1 _27406_ (.Y(_05330_),
    .A(net3393),
    .B(_05329_));
 sg13g2_inv_1 _27407_ (.Y(_05331_),
    .A(_05330_));
 sg13g2_xnor2_1 _27408_ (.Y(_05332_),
    .A(net3393),
    .B(_05329_));
 sg13g2_nand2_1 _27409_ (.Y(_05333_),
    .A(_05291_),
    .B(_05313_));
 sg13g2_o21ai_1 _27410_ (.B1(_05314_),
    .Y(_05334_),
    .A1(_05301_),
    .A2(_05333_));
 sg13g2_xor2_1 _27411_ (.B(_05334_),
    .A(_05332_),
    .X(_05335_));
 sg13g2_nor2_1 _27412_ (.A(net4300),
    .B(_05329_),
    .Y(_05336_));
 sg13g2_o21ai_1 _27413_ (.B1(net3874),
    .Y(_05337_),
    .A1(net4290),
    .A2(_05335_));
 sg13g2_nand2_1 _27414_ (.Y(_05338_),
    .A(net1870),
    .B(net3912));
 sg13g2_o21ai_1 _27415_ (.B1(_05338_),
    .Y(_00526_),
    .A1(_05336_),
    .A2(_05337_));
 sg13g2_a21oi_1 _27416_ (.A1(net4522),
    .A2(\u_inv.d_next[251] ),
    .Y(_05339_),
    .B1(net3737));
 sg13g2_o21ai_1 _27417_ (.B1(_13617_),
    .Y(_05340_),
    .A1(_13619_),
    .A2(_05324_));
 sg13g2_xor2_1 _27418_ (.B(_05340_),
    .A(_13616_),
    .X(_05341_));
 sg13g2_o21ai_1 _27419_ (.B1(_05339_),
    .Y(_05342_),
    .A1(net4522),
    .A2(_05341_));
 sg13g2_nor2_1 _27420_ (.A(_13887_),
    .B(_05321_),
    .Y(_05343_));
 sg13g2_a21oi_1 _27421_ (.A1(_13616_),
    .A2(_05343_),
    .Y(_05344_),
    .B1(net3823));
 sg13g2_o21ai_1 _27422_ (.B1(_05344_),
    .Y(_05345_),
    .A1(_13616_),
    .A2(_05343_));
 sg13g2_and2_1 _27423_ (.A(_05342_),
    .B(_05345_),
    .X(_05346_));
 sg13g2_xnor2_1 _27424_ (.Y(_05347_),
    .A(net3470),
    .B(_05346_));
 sg13g2_o21ai_1 _27425_ (.B1(_05330_),
    .Y(_05348_),
    .A1(_05332_),
    .A2(_05334_));
 sg13g2_xnor2_1 _27426_ (.Y(_05349_),
    .A(_05347_),
    .B(_05348_));
 sg13g2_o21ai_1 _27427_ (.B1(net3874),
    .Y(_05350_),
    .A1(net4300),
    .A2(_05346_));
 sg13g2_a21oi_1 _27428_ (.A1(net4300),
    .A2(_05349_),
    .Y(_05351_),
    .B1(_05350_));
 sg13g2_a21o_1 _27429_ (.A2(net3913),
    .A1(net2776),
    .B1(_05351_),
    .X(_00527_));
 sg13g2_o21ai_1 _27430_ (.B1(_13888_),
    .Y(_05352_),
    .A1(_13620_),
    .A2(_05320_));
 sg13g2_xnor2_1 _27431_ (.Y(_05353_),
    .A(_13611_),
    .B(_05352_));
 sg13g2_a21oi_2 _27432_ (.B1(_15179_),
    .Y(_05354_),
    .A2(_05325_),
    .A1(_15039_));
 sg13g2_inv_1 _27433_ (.Y(_05355_),
    .A(_05354_));
 sg13g2_a21oi_1 _27434_ (.A1(_13611_),
    .A2(_05354_),
    .Y(_05356_),
    .B1(net4522));
 sg13g2_o21ai_1 _27435_ (.B1(_05356_),
    .Y(_05357_),
    .A1(_13611_),
    .A2(_05354_));
 sg13g2_a21oi_1 _27436_ (.A1(net4522),
    .A2(\u_inv.d_next[252] ),
    .Y(_05358_),
    .B1(net3737));
 sg13g2_a22oi_1 _27437_ (.Y(_05359_),
    .B1(_05357_),
    .B2(_05358_),
    .A2(_05353_),
    .A1(net3737));
 sg13g2_nand2_1 _27438_ (.Y(_05360_),
    .A(net3393),
    .B(_05359_));
 sg13g2_inv_1 _27439_ (.Y(_05361_),
    .A(_05360_));
 sg13g2_xnor2_1 _27440_ (.Y(_05362_),
    .A(net3393),
    .B(_05359_));
 sg13g2_nor2b_1 _27441_ (.A(_05332_),
    .B_N(_05347_),
    .Y(_05363_));
 sg13g2_nor2_1 _27442_ (.A(_05292_),
    .B(_05315_),
    .Y(_05364_));
 sg13g2_nand2_1 _27443_ (.Y(_05365_),
    .A(_05363_),
    .B(_05364_));
 sg13g2_a221oi_1 _27444_ (.B2(_05333_),
    .C1(_05331_),
    .B1(_05363_),
    .A1(net3395),
    .Y(_05366_),
    .A2(_05346_));
 sg13g2_o21ai_1 _27445_ (.B1(_05366_),
    .Y(_05367_),
    .A1(_05300_),
    .A2(_05365_));
 sg13g2_nand2b_1 _27446_ (.Y(_05368_),
    .B(_05367_),
    .A_N(_05362_));
 sg13g2_xor2_1 _27447_ (.B(_05367_),
    .A(_05362_),
    .X(_05369_));
 sg13g2_o21ai_1 _27448_ (.B1(net3874),
    .Y(_05370_),
    .A1(net4300),
    .A2(_05359_));
 sg13g2_a21oi_1 _27449_ (.A1(net4300),
    .A2(_05369_),
    .Y(_05371_),
    .B1(_05370_));
 sg13g2_a21o_1 _27450_ (.A2(net3912),
    .A1(net3056),
    .B1(_05371_),
    .X(_00528_));
 sg13g2_a21oi_1 _27451_ (.A1(net4522),
    .A2(\u_inv.d_next[253] ),
    .Y(_05372_),
    .B1(net3737));
 sg13g2_o21ai_1 _27452_ (.B1(_13610_),
    .Y(_05373_),
    .A1(_13611_),
    .A2(_05354_));
 sg13g2_xnor2_1 _27453_ (.Y(_05374_),
    .A(_13609_),
    .B(_05373_));
 sg13g2_nand2_1 _27454_ (.Y(_05375_),
    .A(net4634),
    .B(_05374_));
 sg13g2_a21oi_1 _27455_ (.A1(_13611_),
    .A2(_05352_),
    .Y(_05376_),
    .B1(_13880_));
 sg13g2_o21ai_1 _27456_ (.B1(net3737),
    .Y(_05377_),
    .A1(_13609_),
    .A2(_05376_));
 sg13g2_a21oi_1 _27457_ (.A1(_13609_),
    .A2(_05376_),
    .Y(_05378_),
    .B1(_05377_));
 sg13g2_a21oi_2 _27458_ (.B1(_05378_),
    .Y(_05379_),
    .A2(_05375_),
    .A1(_05372_));
 sg13g2_xnor2_1 _27459_ (.Y(_05380_),
    .A(net3393),
    .B(_05379_));
 sg13g2_nand2_1 _27460_ (.Y(_05381_),
    .A(_05360_),
    .B(_05368_));
 sg13g2_xor2_1 _27461_ (.B(_05381_),
    .A(_05380_),
    .X(_05382_));
 sg13g2_o21ai_1 _27462_ (.B1(net3874),
    .Y(_05383_),
    .A1(net4300),
    .A2(_05379_));
 sg13g2_a21oi_1 _27463_ (.A1(net4300),
    .A2(_05382_),
    .Y(_05384_),
    .B1(_05383_));
 sg13g2_a21o_1 _27464_ (.A2(net3912),
    .A1(net2743),
    .B1(_05384_),
    .X(_00529_));
 sg13g2_a221oi_1 _27465_ (.B2(_13612_),
    .C1(_13879_),
    .B1(_05352_),
    .A1(_13609_),
    .Y(_05385_),
    .A2(_13880_));
 sg13g2_nor2_1 _27466_ (.A(_13604_),
    .B(_05385_),
    .Y(_05386_));
 sg13g2_xnor2_1 _27467_ (.Y(_05387_),
    .A(_13604_),
    .B(_05385_));
 sg13g2_a21oi_1 _27468_ (.A1(_15037_),
    .A2(_05355_),
    .Y(_05388_),
    .B1(_15175_));
 sg13g2_a21oi_1 _27469_ (.A1(_13605_),
    .A2(_05388_),
    .Y(_05389_),
    .B1(net4522));
 sg13g2_o21ai_1 _27470_ (.B1(_05389_),
    .Y(_05390_),
    .A1(_13605_),
    .A2(_05388_));
 sg13g2_a21oi_1 _27471_ (.A1(net4523),
    .A2(\u_inv.d_next[254] ),
    .Y(_05391_),
    .B1(net3738));
 sg13g2_a22oi_1 _27472_ (.Y(_05392_),
    .B1(_05390_),
    .B2(_05391_),
    .A2(_05387_),
    .A1(net3738));
 sg13g2_nand2_1 _27473_ (.Y(_05393_),
    .A(net3394),
    .B(_05392_));
 sg13g2_xnor2_1 _27474_ (.Y(_05394_),
    .A(net3394),
    .B(_05392_));
 sg13g2_nor2_1 _27475_ (.A(_05362_),
    .B(_05380_),
    .Y(_05395_));
 sg13g2_a221oi_1 _27476_ (.B2(_05367_),
    .C1(_05361_),
    .B1(_05395_),
    .A1(net3393),
    .Y(_05396_),
    .A2(_05379_));
 sg13g2_xnor2_1 _27477_ (.Y(_05397_),
    .A(_05394_),
    .B(_05396_));
 sg13g2_o21ai_1 _27478_ (.B1(net3875),
    .Y(_05398_),
    .A1(net4301),
    .A2(_05392_));
 sg13g2_a21oi_1 _27479_ (.A1(net4301),
    .A2(_05397_),
    .Y(_05399_),
    .B1(_05398_));
 sg13g2_a21o_1 _27480_ (.A2(net3912),
    .A1(net2637),
    .B1(_05399_),
    .X(_00530_));
 sg13g2_a21oi_1 _27481_ (.A1(net4522),
    .A2(\u_inv.d_next[255] ),
    .Y(_05400_),
    .B1(net3737));
 sg13g2_o21ai_1 _27482_ (.B1(_13603_),
    .Y(_05401_),
    .A1(_13605_),
    .A2(_05388_));
 sg13g2_xnor2_1 _27483_ (.Y(_05402_),
    .A(_13602_),
    .B(_05401_));
 sg13g2_nand2_1 _27484_ (.Y(_05403_),
    .A(net4634),
    .B(_05402_));
 sg13g2_nor2_1 _27485_ (.A(_13882_),
    .B(_05386_),
    .Y(_05404_));
 sg13g2_o21ai_1 _27486_ (.B1(net3737),
    .Y(_05405_),
    .A1(_13602_),
    .A2(_05404_));
 sg13g2_a21oi_1 _27487_ (.A1(_13602_),
    .A2(_05404_),
    .Y(_05406_),
    .B1(_05405_));
 sg13g2_a21oi_2 _27488_ (.B1(_05406_),
    .Y(_05407_),
    .A2(_05403_),
    .A1(_05400_));
 sg13g2_xnor2_1 _27489_ (.Y(_05408_),
    .A(net3470),
    .B(_05407_));
 sg13g2_o21ai_1 _27490_ (.B1(_05393_),
    .Y(_05409_),
    .A1(_05394_),
    .A2(_05396_));
 sg13g2_xnor2_1 _27491_ (.Y(_05410_),
    .A(_05408_),
    .B(_05409_));
 sg13g2_o21ai_1 _27492_ (.B1(net3874),
    .Y(_05411_),
    .A1(net4301),
    .A2(_05407_));
 sg13g2_a21oi_1 _27493_ (.A1(net4301),
    .A2(_05410_),
    .Y(_05412_),
    .B1(_05411_));
 sg13g2_a21o_1 _27494_ (.A2(net3912),
    .A1(net2714),
    .B1(_05412_),
    .X(_00531_));
 sg13g2_or3_1 _27495_ (.A(_13600_),
    .B(_15028_),
    .C(_15031_),
    .X(_05413_));
 sg13g2_and3_1 _27496_ (.X(_05414_),
    .A(net4656),
    .B(_13600_),
    .C(_15639_));
 sg13g2_nor2_1 _27497_ (.A(_15643_),
    .B(_05414_),
    .Y(_05415_));
 sg13g2_a22oi_1 _27498_ (.Y(_05416_),
    .B1(_05415_),
    .B2(_15642_),
    .A2(_05413_),
    .A1(_15033_));
 sg13g2_nor2_1 _27499_ (.A(net4304),
    .B(_05416_),
    .Y(_05417_));
 sg13g2_xnor2_1 _27500_ (.Y(_05418_),
    .A(net3470),
    .B(_05416_));
 sg13g2_nand2b_1 _27501_ (.Y(_05419_),
    .B(_05408_),
    .A_N(_05394_));
 sg13g2_o21ai_1 _27502_ (.B1(net3394),
    .Y(_05420_),
    .A1(_05392_),
    .A2(_05407_));
 sg13g2_o21ai_1 _27503_ (.B1(_05420_),
    .Y(_05421_),
    .A1(_05396_),
    .A2(_05419_));
 sg13g2_or2_1 _27504_ (.X(_05422_),
    .B(_05421_),
    .A(_05418_));
 sg13g2_a21oi_1 _27505_ (.A1(_05418_),
    .A2(_05421_),
    .Y(_05423_),
    .B1(net4290));
 sg13g2_a21oi_1 _27506_ (.A1(_05422_),
    .A2(_05423_),
    .Y(_05424_),
    .B1(_05417_));
 sg13g2_nand2_1 _27507_ (.Y(_05425_),
    .A(net2452),
    .B(net3912));
 sg13g2_o21ai_1 _27508_ (.B1(_05425_),
    .Y(_00532_),
    .A1(net4233),
    .A2(_05424_));
 sg13g2_nand2_1 _27509_ (.Y(_05426_),
    .A(net2570),
    .B(net3923));
 sg13g2_a21oi_1 _27510_ (.A1(net3397),
    .A2(net4290),
    .Y(_05427_),
    .B1(_05423_));
 sg13g2_o21ai_1 _27511_ (.B1(net3879),
    .Y(_05428_),
    .A1(net3401),
    .A2(_05416_));
 sg13g2_o21ai_1 _27512_ (.B1(_05426_),
    .Y(_00533_),
    .A1(_05427_),
    .A2(_05428_));
 sg13g2_nor2_2 _27513_ (.A(net4445),
    .B(net3780),
    .Y(_05429_));
 sg13g2_nand2_1 _27514_ (.Y(_05430_),
    .A(net4382),
    .B(net3841));
 sg13g2_nand2_1 _27515_ (.Y(_05431_),
    .A(net4027),
    .B(net3704));
 sg13g2_nor2_1 _27516_ (.A(net4443),
    .B(net3845),
    .Y(_05432_));
 sg13g2_nand2_1 _27517_ (.Y(_05433_),
    .A(net4381),
    .B(net3767));
 sg13g2_nor2_1 _27518_ (.A(net3841),
    .B(net4234),
    .Y(_05434_));
 sg13g2_a22oi_1 _27519_ (.Y(_05435_),
    .B1(net3589),
    .B2(net2479),
    .A2(net3496),
    .A1(net4799));
 sg13g2_inv_1 _27520_ (.Y(_00534_),
    .A(net2480));
 sg13g2_a22oi_1 _27521_ (.Y(_05436_),
    .B1(net3589),
    .B2(net2558),
    .A2(net3496),
    .A1(net4797));
 sg13g2_inv_1 _27522_ (.Y(_00535_),
    .A(net2559));
 sg13g2_a22oi_1 _27523_ (.Y(_05437_),
    .B1(net3589),
    .B2(net3030),
    .A2(net3496),
    .A1(net4796));
 sg13g2_inv_1 _27524_ (.Y(_00536_),
    .A(_05437_));
 sg13g2_a22oi_1 _27525_ (.Y(_05438_),
    .B1(net3589),
    .B2(net2797),
    .A2(net3496),
    .A1(\u_inv.d_reg[3] ));
 sg13g2_inv_1 _27526_ (.Y(_00537_),
    .A(net2798));
 sg13g2_a22oi_1 _27527_ (.Y(_05439_),
    .B1(net3589),
    .B2(net2155),
    .A2(net3496),
    .A1(net2982));
 sg13g2_inv_1 _27528_ (.Y(_00538_),
    .A(_05439_));
 sg13g2_a22oi_1 _27529_ (.Y(_05440_),
    .B1(net3589),
    .B2(net2816),
    .A2(net3496),
    .A1(\u_inv.d_reg[5] ));
 sg13g2_inv_1 _27530_ (.Y(_00539_),
    .A(net2817));
 sg13g2_a22oi_1 _27531_ (.Y(_05441_),
    .B1(net3589),
    .B2(net2170),
    .A2(net3496),
    .A1(net4795));
 sg13g2_inv_1 _27532_ (.Y(_00540_),
    .A(_05441_));
 sg13g2_a22oi_1 _27533_ (.Y(_05442_),
    .B1(net3587),
    .B2(net2547),
    .A2(net3494),
    .A1(net4794));
 sg13g2_inv_1 _27534_ (.Y(_00541_),
    .A(net2548));
 sg13g2_a22oi_1 _27535_ (.Y(_05443_),
    .B1(net3587),
    .B2(net2516),
    .A2(net3494),
    .A1(net3053));
 sg13g2_inv_1 _27536_ (.Y(_00542_),
    .A(_05443_));
 sg13g2_a22oi_1 _27537_ (.Y(_05444_),
    .B1(net3587),
    .B2(net2901),
    .A2(net3494),
    .A1(\u_inv.d_reg[9] ));
 sg13g2_inv_1 _27538_ (.Y(_00543_),
    .A(net2902));
 sg13g2_a22oi_1 _27539_ (.Y(_05445_),
    .B1(net3587),
    .B2(net2066),
    .A2(net3494),
    .A1(net2331));
 sg13g2_inv_1 _27540_ (.Y(_00544_),
    .A(_05445_));
 sg13g2_a22oi_1 _27541_ (.Y(_05446_),
    .B1(net3587),
    .B2(net2492),
    .A2(net3494),
    .A1(net4792));
 sg13g2_inv_1 _27542_ (.Y(_00545_),
    .A(net2493));
 sg13g2_a22oi_1 _27543_ (.Y(_05447_),
    .B1(net3587),
    .B2(net2511),
    .A2(net3494),
    .A1(\u_inv.d_reg[12] ));
 sg13g2_inv_1 _27544_ (.Y(_00546_),
    .A(net2512));
 sg13g2_a22oi_1 _27545_ (.Y(_05448_),
    .B1(net3587),
    .B2(net2727),
    .A2(net3494),
    .A1(\u_inv.d_reg[13] ));
 sg13g2_inv_1 _27546_ (.Y(_00547_),
    .A(net2728));
 sg13g2_a22oi_1 _27547_ (.Y(_05449_),
    .B1(net3587),
    .B2(net2945),
    .A2(net3494),
    .A1(\u_inv.d_reg[14] ));
 sg13g2_inv_1 _27548_ (.Y(_00548_),
    .A(net2946));
 sg13g2_a22oi_1 _27549_ (.Y(_05450_),
    .B1(net3595),
    .B2(net3215),
    .A2(net3502),
    .A1(net3243));
 sg13g2_inv_1 _27550_ (.Y(_00549_),
    .A(_05450_));
 sg13g2_a22oi_1 _27551_ (.Y(_05451_),
    .B1(net3597),
    .B2(net2028),
    .A2(net3504),
    .A1(net2761));
 sg13g2_inv_1 _27552_ (.Y(_00550_),
    .A(_05451_));
 sg13g2_a22oi_1 _27553_ (.Y(_05452_),
    .B1(net3597),
    .B2(net4805),
    .A2(net3504),
    .A1(net4791));
 sg13g2_inv_1 _27554_ (.Y(_00551_),
    .A(net4961));
 sg13g2_a22oi_1 _27555_ (.Y(_05453_),
    .B1(net3597),
    .B2(net3191),
    .A2(net3504),
    .A1(net4790));
 sg13g2_inv_1 _27556_ (.Y(_00552_),
    .A(net3192));
 sg13g2_a22oi_1 _27557_ (.Y(_05454_),
    .B1(net3597),
    .B2(net2134),
    .A2(net3504),
    .A1(net2867));
 sg13g2_inv_1 _27558_ (.Y(_00553_),
    .A(_05454_));
 sg13g2_a22oi_1 _27559_ (.Y(_05455_),
    .B1(net3597),
    .B2(net2911),
    .A2(net3504),
    .A1(\u_inv.d_reg[20] ));
 sg13g2_inv_1 _27560_ (.Y(_00554_),
    .A(net2912));
 sg13g2_a22oi_1 _27561_ (.Y(_05456_),
    .B1(net3599),
    .B2(net3085),
    .A2(net3506),
    .A1(\u_inv.d_reg[21] ));
 sg13g2_inv_1 _27562_ (.Y(_00555_),
    .A(net3086));
 sg13g2_a22oi_1 _27563_ (.Y(_05457_),
    .B1(net3599),
    .B2(net2840),
    .A2(net3506),
    .A1(net4789));
 sg13g2_inv_1 _27564_ (.Y(_00556_),
    .A(_05457_));
 sg13g2_a22oi_1 _27565_ (.Y(_05458_),
    .B1(net3599),
    .B2(\u_inv.d_next[23] ),
    .A2(net3506),
    .A1(net3223));
 sg13g2_inv_1 _27566_ (.Y(_00557_),
    .A(net3224));
 sg13g2_a22oi_1 _27567_ (.Y(_05459_),
    .B1(net3599),
    .B2(\u_inv.d_next[24] ),
    .A2(net3506),
    .A1(net2693));
 sg13g2_inv_1 _27568_ (.Y(_00558_),
    .A(net2694));
 sg13g2_a22oi_1 _27569_ (.Y(_05460_),
    .B1(net3599),
    .B2(net2465),
    .A2(net3506),
    .A1(net4788));
 sg13g2_inv_1 _27570_ (.Y(_00559_),
    .A(_05460_));
 sg13g2_a22oi_1 _27571_ (.Y(_05461_),
    .B1(net3599),
    .B2(net3143),
    .A2(net3506),
    .A1(net4787));
 sg13g2_inv_1 _27572_ (.Y(_00560_),
    .A(net3144));
 sg13g2_a22oi_1 _27573_ (.Y(_05462_),
    .B1(net3600),
    .B2(net2780),
    .A2(net3507),
    .A1(\u_inv.d_reg[27] ));
 sg13g2_inv_1 _27574_ (.Y(_00561_),
    .A(net2781));
 sg13g2_a22oi_1 _27575_ (.Y(_05463_),
    .B1(net3599),
    .B2(net2605),
    .A2(net3506),
    .A1(\u_inv.d_reg[28] ));
 sg13g2_inv_1 _27576_ (.Y(_00562_),
    .A(net2606));
 sg13g2_a22oi_1 _27577_ (.Y(_05464_),
    .B1(net3609),
    .B2(net2649),
    .A2(net3516),
    .A1(\u_inv.d_reg[29] ));
 sg13g2_inv_1 _27578_ (.Y(_00563_),
    .A(net2650));
 sg13g2_a22oi_1 _27579_ (.Y(_05465_),
    .B1(net3599),
    .B2(net3281),
    .A2(net3506),
    .A1(net3287));
 sg13g2_inv_1 _27580_ (.Y(_00564_),
    .A(_05465_));
 sg13g2_a22oi_1 _27581_ (.Y(_05466_),
    .B1(net3609),
    .B2(\u_inv.d_next[31] ),
    .A2(net3516),
    .A1(net3213));
 sg13g2_inv_1 _27582_ (.Y(_00565_),
    .A(net3214));
 sg13g2_a22oi_1 _27583_ (.Y(_05467_),
    .B1(net3609),
    .B2(net3104),
    .A2(net3516),
    .A1(\u_inv.d_reg[32] ));
 sg13g2_inv_1 _27584_ (.Y(_00566_),
    .A(net3105));
 sg13g2_a22oi_1 _27585_ (.Y(_05468_),
    .B1(net3609),
    .B2(net2864),
    .A2(net3516),
    .A1(net3266));
 sg13g2_inv_1 _27586_ (.Y(_00567_),
    .A(_05468_));
 sg13g2_a22oi_1 _27587_ (.Y(_05469_),
    .B1(net3609),
    .B2(net2889),
    .A2(net3516),
    .A1(net3203));
 sg13g2_inv_1 _27588_ (.Y(_00568_),
    .A(_05469_));
 sg13g2_a22oi_1 _27589_ (.Y(_05470_),
    .B1(net3612),
    .B2(net2844),
    .A2(net3519),
    .A1(\u_inv.d_reg[35] ));
 sg13g2_inv_1 _27590_ (.Y(_00569_),
    .A(net2845));
 sg13g2_a22oi_1 _27591_ (.Y(_05471_),
    .B1(net3609),
    .B2(net3122),
    .A2(net3516),
    .A1(\u_inv.d_reg[36] ));
 sg13g2_inv_1 _27592_ (.Y(_00570_),
    .A(net3123));
 sg13g2_a22oi_1 _27593_ (.Y(_05472_),
    .B1(net3609),
    .B2(net2922),
    .A2(net3516),
    .A1(\u_inv.d_reg[37] ));
 sg13g2_inv_1 _27594_ (.Y(_00571_),
    .A(net2923));
 sg13g2_a22oi_1 _27595_ (.Y(_05473_),
    .B1(net3610),
    .B2(net2957),
    .A2(net3517),
    .A1(\u_inv.d_reg[38] ));
 sg13g2_inv_1 _27596_ (.Y(_00572_),
    .A(net2958));
 sg13g2_a22oi_1 _27597_ (.Y(_05474_),
    .B1(net3608),
    .B2(net3168),
    .A2(net3515),
    .A1(net3302));
 sg13g2_inv_1 _27598_ (.Y(_00573_),
    .A(_05474_));
 sg13g2_a22oi_1 _27599_ (.Y(_05475_),
    .B1(net3610),
    .B2(net3117),
    .A2(net3517),
    .A1(\u_inv.d_reg[40] ));
 sg13g2_inv_1 _27600_ (.Y(_00574_),
    .A(net3118));
 sg13g2_a22oi_1 _27601_ (.Y(_05476_),
    .B1(net3612),
    .B2(net2970),
    .A2(net3519),
    .A1(\u_inv.d_reg[41] ));
 sg13g2_inv_1 _27602_ (.Y(_00575_),
    .A(net2971));
 sg13g2_a22oi_1 _27603_ (.Y(_05477_),
    .B1(net3611),
    .B2(net3094),
    .A2(net3518),
    .A1(net4786));
 sg13g2_inv_1 _27604_ (.Y(_00576_),
    .A(net3095));
 sg13g2_a22oi_1 _27605_ (.Y(_05478_),
    .B1(net3611),
    .B2(net3273),
    .A2(net3518),
    .A1(net3288));
 sg13g2_inv_1 _27606_ (.Y(_00577_),
    .A(_05478_));
 sg13g2_a22oi_1 _27607_ (.Y(_05479_),
    .B1(net3611),
    .B2(net3146),
    .A2(net3518),
    .A1(\u_inv.d_reg[44] ));
 sg13g2_inv_1 _27608_ (.Y(_00578_),
    .A(net3147));
 sg13g2_a22oi_1 _27609_ (.Y(_05480_),
    .B1(net3611),
    .B2(net3023),
    .A2(net3518),
    .A1(\u_inv.d_reg[45] ));
 sg13g2_inv_1 _27610_ (.Y(_00579_),
    .A(net3024));
 sg13g2_a22oi_1 _27611_ (.Y(_05481_),
    .B1(net3611),
    .B2(net3182),
    .A2(net3518),
    .A1(net3237));
 sg13g2_inv_1 _27612_ (.Y(_00580_),
    .A(_05481_));
 sg13g2_a22oi_1 _27613_ (.Y(_05482_),
    .B1(net3612),
    .B2(net3225),
    .A2(net3519),
    .A1(\u_inv.d_reg[47] ));
 sg13g2_inv_1 _27614_ (.Y(_00581_),
    .A(net3226));
 sg13g2_a22oi_1 _27615_ (.Y(_05483_),
    .B1(net3621),
    .B2(net2215),
    .A2(net3528),
    .A1(net2537));
 sg13g2_inv_1 _27616_ (.Y(_00582_),
    .A(_05483_));
 sg13g2_a22oi_1 _27617_ (.Y(_05484_),
    .B1(net3625),
    .B2(net3038),
    .A2(net3532),
    .A1(\u_inv.d_reg[49] ));
 sg13g2_inv_1 _27618_ (.Y(_00583_),
    .A(net3039));
 sg13g2_a22oi_1 _27619_ (.Y(_05485_),
    .B1(net3625),
    .B2(net2064),
    .A2(net3532),
    .A1(net2879));
 sg13g2_inv_1 _27620_ (.Y(_00584_),
    .A(_05485_));
 sg13g2_a22oi_1 _27621_ (.Y(_05486_),
    .B1(net3625),
    .B2(net2625),
    .A2(net3532),
    .A1(\u_inv.d_reg[51] ));
 sg13g2_inv_1 _27622_ (.Y(_00585_),
    .A(net2626));
 sg13g2_a22oi_1 _27623_ (.Y(_05487_),
    .B1(net3623),
    .B2(net2447),
    .A2(net3530),
    .A1(net3049));
 sg13g2_inv_1 _27624_ (.Y(_00586_),
    .A(_05487_));
 sg13g2_a22oi_1 _27625_ (.Y(_05488_),
    .B1(net3623),
    .B2(net3079),
    .A2(net3530),
    .A1(\u_inv.d_reg[53] ));
 sg13g2_inv_1 _27626_ (.Y(_00587_),
    .A(net3080));
 sg13g2_a22oi_1 _27627_ (.Y(_05489_),
    .B1(net3623),
    .B2(net3026),
    .A2(net3530),
    .A1(\u_inv.d_reg[54] ));
 sg13g2_inv_1 _27628_ (.Y(_00588_),
    .A(net3027));
 sg13g2_a22oi_1 _27629_ (.Y(_05490_),
    .B1(net3623),
    .B2(net2458),
    .A2(net3530),
    .A1(\u_inv.d_reg[55] ));
 sg13g2_inv_1 _27630_ (.Y(_00589_),
    .A(net2459));
 sg13g2_a22oi_1 _27631_ (.Y(_05491_),
    .B1(net3623),
    .B2(net2112),
    .A2(net3530),
    .A1(net2510));
 sg13g2_inv_1 _27632_ (.Y(_00590_),
    .A(_05491_));
 sg13g2_a22oi_1 _27633_ (.Y(_05492_),
    .B1(net3623),
    .B2(net2991),
    .A2(net3530),
    .A1(\u_inv.d_reg[57] ));
 sg13g2_inv_1 _27634_ (.Y(_00591_),
    .A(net2992));
 sg13g2_a22oi_1 _27635_ (.Y(_05493_),
    .B1(net3623),
    .B2(net4804),
    .A2(net3530),
    .A1(net2422));
 sg13g2_inv_1 _27636_ (.Y(_00592_),
    .A(net2423));
 sg13g2_a22oi_1 _27637_ (.Y(_05494_),
    .B1(net3623),
    .B2(net3219),
    .A2(net3530),
    .A1(\u_inv.d_reg[59] ));
 sg13g2_inv_1 _27638_ (.Y(_00593_),
    .A(net3220));
 sg13g2_a22oi_1 _27639_ (.Y(_05495_),
    .B1(net3631),
    .B2(net2094),
    .A2(net3538),
    .A1(net2803));
 sg13g2_inv_1 _27640_ (.Y(_00594_),
    .A(_05495_));
 sg13g2_a22oi_1 _27641_ (.Y(_05496_),
    .B1(net3624),
    .B2(net2647),
    .A2(net3531),
    .A1(\u_inv.d_reg[61] ));
 sg13g2_inv_1 _27642_ (.Y(_00595_),
    .A(net2648));
 sg13g2_a22oi_1 _27643_ (.Y(_05497_),
    .B1(net3624),
    .B2(net2665),
    .A2(net3531),
    .A1(\u_inv.d_reg[62] ));
 sg13g2_inv_1 _27644_ (.Y(_00596_),
    .A(net2666));
 sg13g2_a22oi_1 _27645_ (.Y(_05498_),
    .B1(net3622),
    .B2(net3114),
    .A2(net3529),
    .A1(net3210));
 sg13g2_inv_1 _27646_ (.Y(_00597_),
    .A(_05498_));
 sg13g2_a22oi_1 _27647_ (.Y(_05499_),
    .B1(net3631),
    .B2(net3241),
    .A2(net3538),
    .A1(net4784));
 sg13g2_inv_1 _27648_ (.Y(_00598_),
    .A(_05499_));
 sg13g2_a22oi_1 _27649_ (.Y(_05500_),
    .B1(net3631),
    .B2(net2607),
    .A2(net3538),
    .A1(\u_inv.d_reg[65] ));
 sg13g2_inv_1 _27650_ (.Y(_00599_),
    .A(net2608));
 sg13g2_a22oi_1 _27651_ (.Y(_05501_),
    .B1(net3631),
    .B2(net2948),
    .A2(net3538),
    .A1(\u_inv.d_reg[66] ));
 sg13g2_inv_1 _27652_ (.Y(_00600_),
    .A(net2949));
 sg13g2_a22oi_1 _27653_ (.Y(_05502_),
    .B1(net3631),
    .B2(net2524),
    .A2(net3538),
    .A1(\u_inv.d_reg[67] ));
 sg13g2_inv_1 _27654_ (.Y(_00601_),
    .A(net2525));
 sg13g2_a22oi_1 _27655_ (.Y(_05503_),
    .B1(net3631),
    .B2(net3150),
    .A2(net3538),
    .A1(\u_inv.d_reg[68] ));
 sg13g2_inv_1 _27656_ (.Y(_00602_),
    .A(net3151));
 sg13g2_a22oi_1 _27657_ (.Y(_05504_),
    .B1(net3636),
    .B2(net1949),
    .A2(net3543),
    .A1(\u_inv.d_reg[69] ));
 sg13g2_inv_1 _27658_ (.Y(_00603_),
    .A(net1950));
 sg13g2_a22oi_1 _27659_ (.Y(_05505_),
    .B1(net3636),
    .B2(net2374),
    .A2(net3543),
    .A1(net2652));
 sg13g2_inv_1 _27660_ (.Y(_00604_),
    .A(_05505_));
 sg13g2_a22oi_1 _27661_ (.Y(_05506_),
    .B1(net3631),
    .B2(net2787),
    .A2(net3538),
    .A1(\u_inv.d_reg[71] ));
 sg13g2_inv_1 _27662_ (.Y(_00605_),
    .A(net2788));
 sg13g2_a22oi_1 _27663_ (.Y(_05507_),
    .B1(net3631),
    .B2(net3058),
    .A2(net3538),
    .A1(net4783));
 sg13g2_inv_1 _27664_ (.Y(_00606_),
    .A(_05507_));
 sg13g2_a22oi_1 _27665_ (.Y(_05508_),
    .B1(net3634),
    .B2(net2315),
    .A2(net3541),
    .A1(net3127));
 sg13g2_inv_1 _27666_ (.Y(_00607_),
    .A(_05508_));
 sg13g2_a22oi_1 _27667_ (.Y(_05509_),
    .B1(net3634),
    .B2(net3211),
    .A2(net3541),
    .A1(\u_inv.d_reg[74] ));
 sg13g2_inv_1 _27668_ (.Y(_00608_),
    .A(net3212));
 sg13g2_a22oi_1 _27669_ (.Y(_05510_),
    .B1(net3648),
    .B2(net3020),
    .A2(net3555),
    .A1(\u_inv.d_reg[75] ));
 sg13g2_inv_1 _27670_ (.Y(_00609_),
    .A(net3021));
 sg13g2_a22oi_1 _27671_ (.Y(_05511_),
    .B1(net3634),
    .B2(net2716),
    .A2(net3541),
    .A1(net4782));
 sg13g2_inv_1 _27672_ (.Y(_00610_),
    .A(_05511_));
 sg13g2_a22oi_1 _27673_ (.Y(_05512_),
    .B1(net3634),
    .B2(net3267),
    .A2(net3541),
    .A1(net4781));
 sg13g2_inv_1 _27674_ (.Y(_00611_),
    .A(net3268));
 sg13g2_a22oi_1 _27675_ (.Y(_05513_),
    .B1(net3634),
    .B2(net2829),
    .A2(net3541),
    .A1(\u_inv.d_reg[78] ));
 sg13g2_inv_1 _27676_ (.Y(_00612_),
    .A(net2830));
 sg13g2_a22oi_1 _27677_ (.Y(_05514_),
    .B1(net3634),
    .B2(net2848),
    .A2(net3541),
    .A1(\u_inv.d_reg[79] ));
 sg13g2_inv_1 _27678_ (.Y(_00613_),
    .A(net2849));
 sg13g2_a22oi_1 _27679_ (.Y(_05515_),
    .B1(net3634),
    .B2(net1997),
    .A2(net3541),
    .A1(net2582));
 sg13g2_inv_1 _27680_ (.Y(_00614_),
    .A(_05515_));
 sg13g2_a22oi_1 _27681_ (.Y(_05516_),
    .B1(net3634),
    .B2(net2241),
    .A2(net3541),
    .A1(net2775));
 sg13g2_inv_1 _27682_ (.Y(_00615_),
    .A(_05516_));
 sg13g2_a22oi_1 _27683_ (.Y(_05517_),
    .B1(net3635),
    .B2(net2862),
    .A2(net3542),
    .A1(\u_inv.d_reg[82] ));
 sg13g2_inv_1 _27684_ (.Y(_00616_),
    .A(net2863));
 sg13g2_a22oi_1 _27685_ (.Y(_05518_),
    .B1(net3633),
    .B2(net2662),
    .A2(net3540),
    .A1(\u_inv.d_reg[83] ));
 sg13g2_inv_1 _27686_ (.Y(_00617_),
    .A(net2663));
 sg13g2_a22oi_1 _27687_ (.Y(_05519_),
    .B1(net3633),
    .B2(net2615),
    .A2(net3540),
    .A1(net2981));
 sg13g2_inv_1 _27688_ (.Y(_00618_),
    .A(_05519_));
 sg13g2_a22oi_1 _27689_ (.Y(_05520_),
    .B1(net3635),
    .B2(net2695),
    .A2(net3542),
    .A1(net3040));
 sg13g2_inv_1 _27690_ (.Y(_00619_),
    .A(_05520_));
 sg13g2_a22oi_1 _27691_ (.Y(_05521_),
    .B1(net3633),
    .B2(net3174),
    .A2(net3540),
    .A1(\u_inv.d_reg[86] ));
 sg13g2_inv_1 _27692_ (.Y(_00620_),
    .A(net3175));
 sg13g2_a22oi_1 _27693_ (.Y(_05522_),
    .B1(net3633),
    .B2(net2815),
    .A2(net3540),
    .A1(net3161));
 sg13g2_inv_1 _27694_ (.Y(_00621_),
    .A(_05522_));
 sg13g2_a22oi_1 _27695_ (.Y(_05523_),
    .B1(net3642),
    .B2(net3098),
    .A2(net3549),
    .A1(net3269));
 sg13g2_inv_1 _27696_ (.Y(_00622_),
    .A(_05523_));
 sg13g2_a22oi_1 _27697_ (.Y(_05524_),
    .B1(net3633),
    .B2(net2351),
    .A2(net3540),
    .A1(\u_inv.d_reg[89] ));
 sg13g2_inv_1 _27698_ (.Y(_00623_),
    .A(net2352));
 sg13g2_a22oi_1 _27699_ (.Y(_05525_),
    .B1(net3633),
    .B2(net2708),
    .A2(net3540),
    .A1(net3173));
 sg13g2_inv_1 _27700_ (.Y(_00624_),
    .A(_05525_));
 sg13g2_a22oi_1 _27701_ (.Y(_05526_),
    .B1(net3633),
    .B2(net2732),
    .A2(net3540),
    .A1(\u_inv.d_reg[91] ));
 sg13g2_inv_1 _27702_ (.Y(_00625_),
    .A(net2733));
 sg13g2_a22oi_1 _27703_ (.Y(_05527_),
    .B1(net3633),
    .B2(net2198),
    .A2(net3540),
    .A1(net2360));
 sg13g2_inv_1 _27704_ (.Y(_00626_),
    .A(_05527_));
 sg13g2_a22oi_1 _27705_ (.Y(_05528_),
    .B1(net3642),
    .B2(net2631),
    .A2(net3549),
    .A1(\u_inv.d_reg[93] ));
 sg13g2_inv_1 _27706_ (.Y(_00627_),
    .A(net2632));
 sg13g2_a22oi_1 _27707_ (.Y(_05529_),
    .B1(net3635),
    .B2(net2210),
    .A2(net3542),
    .A1(net2599));
 sg13g2_inv_1 _27708_ (.Y(_00628_),
    .A(_05529_));
 sg13g2_a22oi_1 _27709_ (.Y(_05530_),
    .B1(net3642),
    .B2(net4955),
    .A2(net3549),
    .A1(\u_inv.d_reg[95] ));
 sg13g2_inv_1 _27710_ (.Y(_00629_),
    .A(net4956));
 sg13g2_a22oi_1 _27711_ (.Y(_05531_),
    .B1(net3643),
    .B2(net2139),
    .A2(net3550),
    .A1(net2859));
 sg13g2_inv_1 _27712_ (.Y(_00630_),
    .A(_05531_));
 sg13g2_a22oi_1 _27713_ (.Y(_05532_),
    .B1(net3643),
    .B2(net2782),
    .A2(net3550),
    .A1(\u_inv.d_reg[97] ));
 sg13g2_inv_1 _27714_ (.Y(_00631_),
    .A(net2783));
 sg13g2_a22oi_1 _27715_ (.Y(_05533_),
    .B1(net3642),
    .B2(net2724),
    .A2(net3549),
    .A1(\u_inv.d_reg[98] ));
 sg13g2_inv_1 _27716_ (.Y(_00632_),
    .A(net2725));
 sg13g2_a22oi_1 _27717_ (.Y(_05534_),
    .B1(net3642),
    .B2(net2612),
    .A2(net3549),
    .A1(net3097));
 sg13g2_inv_1 _27718_ (.Y(_00633_),
    .A(_05534_));
 sg13g2_a22oi_1 _27719_ (.Y(_05535_),
    .B1(net3642),
    .B2(net3066),
    .A2(net3549),
    .A1(\u_inv.d_reg[100] ));
 sg13g2_inv_1 _27720_ (.Y(_00634_),
    .A(net3067));
 sg13g2_a22oi_1 _27721_ (.Y(_05536_),
    .B1(net3642),
    .B2(net2263),
    .A2(net3549),
    .A1(\u_inv.d_reg[101] ));
 sg13g2_inv_1 _27722_ (.Y(_00635_),
    .A(net2264));
 sg13g2_a22oi_1 _27723_ (.Y(_05537_),
    .B1(net3642),
    .B2(net3068),
    .A2(net3549),
    .A1(\u_inv.d_reg[102] ));
 sg13g2_inv_1 _27724_ (.Y(_00636_),
    .A(net3069));
 sg13g2_a22oi_1 _27725_ (.Y(_05538_),
    .B1(net3643),
    .B2(net2834),
    .A2(net3550),
    .A1(\u_inv.d_reg[103] ));
 sg13g2_inv_1 _27726_ (.Y(_00637_),
    .A(net2835));
 sg13g2_a22oi_1 _27727_ (.Y(_05539_),
    .B1(net3644),
    .B2(net2796),
    .A2(net3551),
    .A1(net4780));
 sg13g2_inv_1 _27728_ (.Y(_00638_),
    .A(_05539_));
 sg13g2_a22oi_1 _27729_ (.Y(_05540_),
    .B1(net3644),
    .B2(net2806),
    .A2(net3551),
    .A1(\u_inv.d_reg[105] ));
 sg13g2_inv_1 _27730_ (.Y(_00639_),
    .A(net2807));
 sg13g2_a22oi_1 _27731_ (.Y(_05541_),
    .B1(net3644),
    .B2(net2445),
    .A2(net3551),
    .A1(net2872));
 sg13g2_inv_1 _27732_ (.Y(_00640_),
    .A(_05541_));
 sg13g2_a22oi_1 _27733_ (.Y(_05542_),
    .B1(net3644),
    .B2(net2292),
    .A2(net3551),
    .A1(net2875));
 sg13g2_inv_1 _27734_ (.Y(_00641_),
    .A(_05542_));
 sg13g2_a22oi_1 _27735_ (.Y(_05543_),
    .B1(net3644),
    .B2(net2237),
    .A2(net3551),
    .A1(net2737));
 sg13g2_inv_1 _27736_ (.Y(_00642_),
    .A(_05543_));
 sg13g2_a22oi_1 _27737_ (.Y(_05544_),
    .B1(net3647),
    .B2(net3293),
    .A2(net3554),
    .A1(net3294));
 sg13g2_inv_1 _27738_ (.Y(_00643_),
    .A(_05544_));
 sg13g2_a22oi_1 _27739_ (.Y(_05545_),
    .B1(net3647),
    .B2(net3217),
    .A2(net3554),
    .A1(\u_inv.d_reg[110] ));
 sg13g2_inv_1 _27740_ (.Y(_00644_),
    .A(net3218));
 sg13g2_a22oi_1 _27741_ (.Y(_05546_),
    .B1(net3643),
    .B2(net2976),
    .A2(net3550),
    .A1(\u_inv.d_reg[111] ));
 sg13g2_inv_1 _27742_ (.Y(_00645_),
    .A(net2977));
 sg13g2_a22oi_1 _27743_ (.Y(_05547_),
    .B1(net3646),
    .B2(net2876),
    .A2(net3553),
    .A1(\u_inv.d_reg[112] ));
 sg13g2_inv_1 _27744_ (.Y(_00646_),
    .A(net2877));
 sg13g2_a22oi_1 _27745_ (.Y(_05548_),
    .B1(net3645),
    .B2(net2917),
    .A2(net3552),
    .A1(net3289));
 sg13g2_inv_1 _27746_ (.Y(_00647_),
    .A(_05548_));
 sg13g2_a22oi_1 _27747_ (.Y(_05549_),
    .B1(net3645),
    .B2(net2540),
    .A2(net3552),
    .A1(net3196));
 sg13g2_inv_1 _27748_ (.Y(_00648_),
    .A(_05549_));
 sg13g2_a22oi_1 _27749_ (.Y(_05550_),
    .B1(net3645),
    .B2(net3201),
    .A2(net3552),
    .A1(\u_inv.d_reg[115] ));
 sg13g2_inv_1 _27750_ (.Y(_00649_),
    .A(net3202));
 sg13g2_a22oi_1 _27751_ (.Y(_05551_),
    .B1(net3645),
    .B2(net2344),
    .A2(net3552),
    .A1(net3000));
 sg13g2_inv_1 _27752_ (.Y(_00650_),
    .A(_05551_));
 sg13g2_a22oi_1 _27753_ (.Y(_05552_),
    .B1(net3645),
    .B2(net3081),
    .A2(net3552),
    .A1(\u_inv.d_reg[117] ));
 sg13g2_inv_1 _27754_ (.Y(_00651_),
    .A(net3082));
 sg13g2_a22oi_1 _27755_ (.Y(_05553_),
    .B1(net3645),
    .B2(net2598),
    .A2(net3552),
    .A1(net3238));
 sg13g2_inv_1 _27756_ (.Y(_00652_),
    .A(_05553_));
 sg13g2_a22oi_1 _27757_ (.Y(_05554_),
    .B1(net3645),
    .B2(net2926),
    .A2(net3552),
    .A1(\u_inv.d_reg[119] ));
 sg13g2_inv_1 _27758_ (.Y(_00653_),
    .A(net2927));
 sg13g2_a22oi_1 _27759_ (.Y(_05555_),
    .B1(net3647),
    .B2(net3060),
    .A2(net3554),
    .A1(\u_inv.d_reg[120] ));
 sg13g2_inv_1 _27760_ (.Y(_00654_),
    .A(net3061));
 sg13g2_a22oi_1 _27761_ (.Y(_05556_),
    .B1(net3646),
    .B2(net2756),
    .A2(net3553),
    .A1(\u_inv.d_reg[121] ));
 sg13g2_inv_1 _27762_ (.Y(_00655_),
    .A(net2757));
 sg13g2_a22oi_1 _27763_ (.Y(_05557_),
    .B1(net3646),
    .B2(net3230),
    .A2(net3553),
    .A1(\u_inv.d_reg[122] ));
 sg13g2_inv_1 _27764_ (.Y(_00656_),
    .A(net3231));
 sg13g2_a22oi_1 _27765_ (.Y(_05558_),
    .B1(net3647),
    .B2(net3235),
    .A2(net3554),
    .A1(\u_inv.d_reg[123] ));
 sg13g2_inv_1 _27766_ (.Y(_00657_),
    .A(net3236));
 sg13g2_a22oi_1 _27767_ (.Y(_05559_),
    .B1(net3655),
    .B2(net2955),
    .A2(net3562),
    .A1(\u_inv.d_reg[124] ));
 sg13g2_inv_1 _27768_ (.Y(_00658_),
    .A(net2956));
 sg13g2_a22oi_1 _27769_ (.Y(_05560_),
    .B1(net3647),
    .B2(net3126),
    .A2(net3554),
    .A1(net3195));
 sg13g2_inv_1 _27770_ (.Y(_00659_),
    .A(_05560_));
 sg13g2_a22oi_1 _27771_ (.Y(_05561_),
    .B1(net3647),
    .B2(net2030),
    .A2(net3554),
    .A1(net2369));
 sg13g2_inv_1 _27772_ (.Y(_00660_),
    .A(_05561_));
 sg13g2_a22oi_1 _27773_ (.Y(_05562_),
    .B1(net3655),
    .B2(net2489),
    .A2(net3562),
    .A1(\u_inv.d_reg[127] ));
 sg13g2_inv_1 _27774_ (.Y(_00661_),
    .A(net2490));
 sg13g2_a22oi_1 _27775_ (.Y(_05563_),
    .B1(net3654),
    .B2(net2580),
    .A2(net3561),
    .A1(\u_inv.d_reg[128] ));
 sg13g2_inv_1 _27776_ (.Y(_00662_),
    .A(net2581));
 sg13g2_a22oi_1 _27777_ (.Y(_05564_),
    .B1(net3654),
    .B2(net2934),
    .A2(net3561),
    .A1(net4779));
 sg13g2_inv_1 _27778_ (.Y(_00663_),
    .A(_05564_));
 sg13g2_a22oi_1 _27779_ (.Y(_05565_),
    .B1(net3645),
    .B2(net4802),
    .A2(net3552),
    .A1(net4778));
 sg13g2_inv_1 _27780_ (.Y(_00664_),
    .A(_05565_));
 sg13g2_a22oi_1 _27781_ (.Y(_05566_),
    .B1(net3654),
    .B2(net3274),
    .A2(net3561),
    .A1(\u_inv.d_reg[131] ));
 sg13g2_inv_1 _27782_ (.Y(_00665_),
    .A(net3275));
 sg13g2_a22oi_1 _27783_ (.Y(_05567_),
    .B1(net3654),
    .B2(net2825),
    .A2(net3561),
    .A1(\u_inv.d_reg[132] ));
 sg13g2_inv_1 _27784_ (.Y(_00666_),
    .A(net2826));
 sg13g2_a22oi_1 _27785_ (.Y(_05568_),
    .B1(net3654),
    .B2(net2909),
    .A2(net3561),
    .A1(\u_inv.d_reg[133] ));
 sg13g2_inv_1 _27786_ (.Y(_00667_),
    .A(net2910));
 sg13g2_a22oi_1 _27787_ (.Y(_05569_),
    .B1(net3654),
    .B2(net2924),
    .A2(net3561),
    .A1(\u_inv.d_reg[134] ));
 sg13g2_inv_1 _27788_ (.Y(_00668_),
    .A(net2925));
 sg13g2_a22oi_1 _27789_ (.Y(_05570_),
    .B1(net3654),
    .B2(net3090),
    .A2(net3561),
    .A1(net3149));
 sg13g2_inv_1 _27790_ (.Y(_00669_),
    .A(_05570_));
 sg13g2_a22oi_1 _27791_ (.Y(_05571_),
    .B1(net3654),
    .B2(net2565),
    .A2(net3561),
    .A1(net3166));
 sg13g2_inv_1 _27792_ (.Y(_00670_),
    .A(_05571_));
 sg13g2_a22oi_1 _27793_ (.Y(_05572_),
    .B1(net3655),
    .B2(net3292),
    .A2(net3562),
    .A1(net4952));
 sg13g2_inv_1 _27794_ (.Y(_00671_),
    .A(_05572_));
 sg13g2_a22oi_1 _27795_ (.Y(_05573_),
    .B1(net3657),
    .B2(net3291),
    .A2(net3564),
    .A1(net4777));
 sg13g2_inv_1 _27796_ (.Y(_00672_),
    .A(_05573_));
 sg13g2_a22oi_1 _27797_ (.Y(_05574_),
    .B1(net3656),
    .B2(net3207),
    .A2(net3563),
    .A1(\u_inv.d_reg[139] ));
 sg13g2_inv_1 _27798_ (.Y(_00673_),
    .A(net3208));
 sg13g2_a22oi_1 _27799_ (.Y(_05575_),
    .B1(net3656),
    .B2(net2852),
    .A2(net3563),
    .A1(\u_inv.d_reg[140] ));
 sg13g2_inv_1 _27800_ (.Y(_00674_),
    .A(net2853));
 sg13g2_a22oi_1 _27801_ (.Y(_05576_),
    .B1(net3656),
    .B2(net2899),
    .A2(net3563),
    .A1(\u_inv.d_reg[141] ));
 sg13g2_inv_1 _27802_ (.Y(_00675_),
    .A(net2900));
 sg13g2_a22oi_1 _27803_ (.Y(_05577_),
    .B1(net3656),
    .B2(net2641),
    .A2(net3563),
    .A1(\u_inv.d_reg[142] ));
 sg13g2_inv_1 _27804_ (.Y(_00676_),
    .A(net2642));
 sg13g2_a22oi_1 _27805_ (.Y(_05578_),
    .B1(net3656),
    .B2(net2567),
    .A2(net3563),
    .A1(net3055));
 sg13g2_inv_1 _27806_ (.Y(_00677_),
    .A(_05578_));
 sg13g2_a22oi_1 _27807_ (.Y(_05579_),
    .B1(net3668),
    .B2(net2150),
    .A2(net3575),
    .A1(net2476));
 sg13g2_inv_1 _27808_ (.Y(_00678_),
    .A(_05579_));
 sg13g2_a22oi_1 _27809_ (.Y(_05580_),
    .B1(net3668),
    .B2(net2959),
    .A2(net3575),
    .A1(\u_inv.d_reg[145] ));
 sg13g2_inv_1 _27810_ (.Y(_00679_),
    .A(net2960));
 sg13g2_a22oi_1 _27811_ (.Y(_05581_),
    .B1(net3668),
    .B2(net2881),
    .A2(net3575),
    .A1(\u_inv.d_reg[146] ));
 sg13g2_inv_1 _27812_ (.Y(_00680_),
    .A(net2882));
 sg13g2_a22oi_1 _27813_ (.Y(_05582_),
    .B1(net3667),
    .B2(net3197),
    .A2(net3574),
    .A1(net3262));
 sg13g2_inv_1 _27814_ (.Y(_00681_),
    .A(_05582_));
 sg13g2_a22oi_1 _27815_ (.Y(_05583_),
    .B1(net3667),
    .B2(net2837),
    .A2(net3574),
    .A1(\u_inv.d_reg[148] ));
 sg13g2_inv_1 _27816_ (.Y(_00682_),
    .A(net2838));
 sg13g2_a22oi_1 _27817_ (.Y(_05584_),
    .B1(net3667),
    .B2(net2972),
    .A2(net3574),
    .A1(\u_inv.d_reg[149] ));
 sg13g2_inv_1 _27818_ (.Y(_00683_),
    .A(net2973));
 sg13g2_a22oi_1 _27819_ (.Y(_05585_),
    .B1(net3668),
    .B2(\u_inv.d_next[150] ),
    .A2(net3575),
    .A1(net2734));
 sg13g2_inv_1 _27820_ (.Y(_00684_),
    .A(net2735));
 sg13g2_a22oi_1 _27821_ (.Y(_05586_),
    .B1(net3668),
    .B2(net2364),
    .A2(net3575),
    .A1(\u_inv.d_reg[151] ));
 sg13g2_inv_1 _27822_ (.Y(_00685_),
    .A(net2365));
 sg13g2_a22oi_1 _27823_ (.Y(_05587_),
    .B1(net3668),
    .B2(net2501),
    .A2(net3575),
    .A1(net2659));
 sg13g2_inv_1 _27824_ (.Y(_00686_),
    .A(_05587_));
 sg13g2_a22oi_1 _27825_ (.Y(_05588_),
    .B1(net3668),
    .B2(net2870),
    .A2(net3575),
    .A1(\u_inv.d_reg[153] ));
 sg13g2_inv_1 _27826_ (.Y(_00687_),
    .A(net2871));
 sg13g2_a22oi_1 _27827_ (.Y(_05589_),
    .B1(net3656),
    .B2(net2747),
    .A2(net3563),
    .A1(\u_inv.d_reg[154] ));
 sg13g2_inv_1 _27828_ (.Y(_00688_),
    .A(net2748));
 sg13g2_a22oi_1 _27829_ (.Y(_05590_),
    .B1(net3656),
    .B2(\u_inv.d_next[155] ),
    .A2(net3563),
    .A1(net2951));
 sg13g2_inv_1 _27830_ (.Y(_00689_),
    .A(net2952));
 sg13g2_a22oi_1 _27831_ (.Y(_05591_),
    .B1(net3657),
    .B2(net3190),
    .A2(net3564),
    .A1(net3300));
 sg13g2_inv_1 _27832_ (.Y(_00690_),
    .A(_05591_));
 sg13g2_a22oi_1 _27833_ (.Y(_05592_),
    .B1(net3657),
    .B2(net3106),
    .A2(net3564),
    .A1(\u_inv.d_reg[157] ));
 sg13g2_inv_1 _27834_ (.Y(_00691_),
    .A(net3107));
 sg13g2_a22oi_1 _27835_ (.Y(_05593_),
    .B1(net3656),
    .B2(net2460),
    .A2(net3563),
    .A1(net3136));
 sg13g2_inv_1 _27836_ (.Y(_00692_),
    .A(_05593_));
 sg13g2_a22oi_1 _27837_ (.Y(_05594_),
    .B1(net3657),
    .B2(net2311),
    .A2(net3564),
    .A1(\u_inv.d_reg[159] ));
 sg13g2_inv_1 _27838_ (.Y(_00693_),
    .A(net2312));
 sg13g2_a22oi_1 _27839_ (.Y(_05595_),
    .B1(net3657),
    .B2(net2685),
    .A2(net3564),
    .A1(net3046));
 sg13g2_inv_1 _27840_ (.Y(_00694_),
    .A(_05595_));
 sg13g2_a22oi_1 _27841_ (.Y(_05596_),
    .B1(net3658),
    .B2(net2855),
    .A2(net3565),
    .A1(\u_inv.d_reg[161] ));
 sg13g2_inv_1 _27842_ (.Y(_00695_),
    .A(net2856));
 sg13g2_a22oi_1 _27843_ (.Y(_05597_),
    .B1(net3655),
    .B2(net4801),
    .A2(net3562),
    .A1(net4775));
 sg13g2_inv_1 _27844_ (.Y(_00696_),
    .A(_05597_));
 sg13g2_a22oi_1 _27845_ (.Y(_05598_),
    .B1(net3658),
    .B2(net3255),
    .A2(net3565),
    .A1(\u_inv.d_reg[163] ));
 sg13g2_inv_1 _27846_ (.Y(_00697_),
    .A(net3256));
 sg13g2_a22oi_1 _27847_ (.Y(_05599_),
    .B1(net3658),
    .B2(net2269),
    .A2(net3565),
    .A1(\u_inv.d_reg[164] ));
 sg13g2_inv_1 _27848_ (.Y(_00698_),
    .A(net2270));
 sg13g2_a22oi_1 _27849_ (.Y(_05600_),
    .B1(net3658),
    .B2(net2935),
    .A2(net3565),
    .A1(\u_inv.d_reg[165] ));
 sg13g2_inv_1 _27850_ (.Y(_00699_),
    .A(net2936));
 sg13g2_a22oi_1 _27851_ (.Y(_05601_),
    .B1(net3655),
    .B2(net3158),
    .A2(net3562),
    .A1(\u_inv.d_reg[166] ));
 sg13g2_inv_1 _27852_ (.Y(_00700_),
    .A(net3159));
 sg13g2_a22oi_1 _27853_ (.Y(_05602_),
    .B1(net3658),
    .B2(net2794),
    .A2(net3565),
    .A1(\u_inv.d_reg[167] ));
 sg13g2_inv_1 _27854_ (.Y(_00701_),
    .A(net2795));
 sg13g2_a22oi_1 _27855_ (.Y(_05603_),
    .B1(net3658),
    .B2(net2133),
    .A2(net3565),
    .A1(net2564));
 sg13g2_inv_1 _27856_ (.Y(_00702_),
    .A(_05603_));
 sg13g2_a22oi_1 _27857_ (.Y(_05604_),
    .B1(net3658),
    .B2(net2906),
    .A2(net3565),
    .A1(\u_inv.d_reg[169] ));
 sg13g2_inv_1 _27858_ (.Y(_00703_),
    .A(net2907));
 sg13g2_a22oi_1 _27859_ (.Y(_05605_),
    .B1(net3663),
    .B2(net2873),
    .A2(net3570),
    .A1(\u_inv.d_reg[170] ));
 sg13g2_inv_1 _27860_ (.Y(_00704_),
    .A(net2874));
 sg13g2_a22oi_1 _27861_ (.Y(_05606_),
    .B1(net3663),
    .B2(net3164),
    .A2(net3570),
    .A1(\u_inv.d_reg[171] ));
 sg13g2_inv_1 _27862_ (.Y(_00705_),
    .A(net3165));
 sg13g2_a22oi_1 _27863_ (.Y(_05607_),
    .B1(net3663),
    .B2(net2987),
    .A2(net3570),
    .A1(\u_inv.d_reg[172] ));
 sg13g2_inv_1 _27864_ (.Y(_00706_),
    .A(net2988));
 sg13g2_a22oi_1 _27865_ (.Y(_05608_),
    .B1(net3660),
    .B2(net2342),
    .A2(net3567),
    .A1(\u_inv.d_reg[173] ));
 sg13g2_inv_1 _27866_ (.Y(_00707_),
    .A(net2343));
 sg13g2_a22oi_1 _27867_ (.Y(_05609_),
    .B1(net3660),
    .B2(net2436),
    .A2(net3567),
    .A1(\u_inv.d_reg[174] ));
 sg13g2_inv_1 _27868_ (.Y(_00708_),
    .A(net2437));
 sg13g2_a22oi_1 _27869_ (.Y(_05610_),
    .B1(net3660),
    .B2(net2846),
    .A2(net3567),
    .A1(\u_inv.d_reg[175] ));
 sg13g2_inv_1 _27870_ (.Y(_00709_),
    .A(net2847));
 sg13g2_a22oi_1 _27871_ (.Y(_05611_),
    .B1(net3660),
    .B2(net2674),
    .A2(net3567),
    .A1(\u_inv.d_reg[176] ));
 sg13g2_inv_1 _27872_ (.Y(_00710_),
    .A(net2675));
 sg13g2_a22oi_1 _27873_ (.Y(_05612_),
    .B1(net3660),
    .B2(net2635),
    .A2(net3567),
    .A1(net2740));
 sg13g2_inv_1 _27874_ (.Y(_00711_),
    .A(_05612_));
 sg13g2_a22oi_1 _27875_ (.Y(_05613_),
    .B1(net3660),
    .B2(net2893),
    .A2(net3567),
    .A1(\u_inv.d_reg[178] ));
 sg13g2_inv_1 _27876_ (.Y(_00712_),
    .A(net2894));
 sg13g2_a22oi_1 _27877_ (.Y(_05614_),
    .B1(net3652),
    .B2(net3216),
    .A2(net3559),
    .A1(net3234));
 sg13g2_inv_1 _27878_ (.Y(_00713_),
    .A(_05614_));
 sg13g2_a22oi_1 _27879_ (.Y(_05615_),
    .B1(net3652),
    .B2(net3047),
    .A2(net3559),
    .A1(\u_inv.d_reg[180] ));
 sg13g2_inv_1 _27880_ (.Y(_00714_),
    .A(net3048));
 sg13g2_a22oi_1 _27881_ (.Y(_05616_),
    .B1(net3652),
    .B2(net2392),
    .A2(net3559),
    .A1(\u_inv.d_reg[181] ));
 sg13g2_inv_1 _27882_ (.Y(_00715_),
    .A(net2393));
 sg13g2_a22oi_1 _27883_ (.Y(_05617_),
    .B1(net3652),
    .B2(net2507),
    .A2(net3559),
    .A1(\u_inv.d_reg[182] ));
 sg13g2_inv_1 _27884_ (.Y(_00716_),
    .A(net2508));
 sg13g2_a22oi_1 _27885_ (.Y(_05618_),
    .B1(net3652),
    .B2(net2908),
    .A2(net3559),
    .A1(net3017));
 sg13g2_inv_1 _27886_ (.Y(_00717_),
    .A(_05618_));
 sg13g2_a22oi_1 _27887_ (.Y(_05619_),
    .B1(net3652),
    .B2(net1065),
    .A2(net3559),
    .A1(\u_inv.d_reg[184] ));
 sg13g2_inv_1 _27888_ (.Y(_00718_),
    .A(net1066));
 sg13g2_a22oi_1 _27889_ (.Y(_05620_),
    .B1(net3649),
    .B2(net2273),
    .A2(net3556),
    .A1(\u_inv.d_reg[185] ));
 sg13g2_inv_1 _27890_ (.Y(_00719_),
    .A(net2274));
 sg13g2_a22oi_1 _27891_ (.Y(_05621_),
    .B1(net3649),
    .B2(net2672),
    .A2(net3556),
    .A1(\u_inv.d_reg[186] ));
 sg13g2_inv_1 _27892_ (.Y(_00720_),
    .A(net2673));
 sg13g2_a22oi_1 _27893_ (.Y(_05622_),
    .B1(net3644),
    .B2(net3138),
    .A2(net3551),
    .A1(net4774));
 sg13g2_inv_1 _27894_ (.Y(_00721_),
    .A(net3139));
 sg13g2_a22oi_1 _27895_ (.Y(_05623_),
    .B1(net3652),
    .B2(net2823),
    .A2(net3559),
    .A1(\u_inv.d_reg[188] ));
 sg13g2_inv_1 _27896_ (.Y(_00722_),
    .A(net2824));
 sg13g2_a22oi_1 _27897_ (.Y(_05624_),
    .B1(net3647),
    .B2(net2297),
    .A2(net3554),
    .A1(\u_inv.d_reg[189] ));
 sg13g2_inv_1 _27898_ (.Y(_00723_),
    .A(net2298));
 sg13g2_a22oi_1 _27899_ (.Y(_05625_),
    .B1(net3647),
    .B2(net3007),
    .A2(net3554),
    .A1(\u_inv.d_reg[190] ));
 sg13g2_inv_1 _27900_ (.Y(_00724_),
    .A(net3008));
 sg13g2_a22oi_1 _27901_ (.Y(_05626_),
    .B1(net3648),
    .B2(net3167),
    .A2(net3555),
    .A1(net3176));
 sg13g2_inv_1 _27902_ (.Y(_00725_),
    .A(_05626_));
 sg13g2_a22oi_1 _27903_ (.Y(_05627_),
    .B1(net3632),
    .B2(net2627),
    .A2(net3539),
    .A1(\u_inv.d_reg[192] ));
 sg13g2_inv_1 _27904_ (.Y(_00726_),
    .A(net2628));
 sg13g2_a22oi_1 _27905_ (.Y(_05628_),
    .B1(net3632),
    .B2(net2745),
    .A2(net3539),
    .A1(\u_inv.d_reg[193] ));
 sg13g2_inv_1 _27906_ (.Y(_00727_),
    .A(net2746));
 sg13g2_a22oi_1 _27907_ (.Y(_05629_),
    .B1(net3632),
    .B2(net2454),
    .A2(net3539),
    .A1(\u_inv.d_reg[194] ));
 sg13g2_inv_1 _27908_ (.Y(_00728_),
    .A(net2455));
 sg13g2_a22oi_1 _27909_ (.Y(_05630_),
    .B1(net3632),
    .B2(net2762),
    .A2(net3539),
    .A1(\u_inv.d_reg[195] ));
 sg13g2_inv_1 _27910_ (.Y(_00729_),
    .A(net2763));
 sg13g2_a22oi_1 _27911_ (.Y(_05631_),
    .B1(net3632),
    .B2(net2766),
    .A2(net3539),
    .A1(net4773));
 sg13g2_inv_1 _27912_ (.Y(_00730_),
    .A(_05631_));
 sg13g2_a22oi_1 _27913_ (.Y(_05632_),
    .B1(net3632),
    .B2(net3205),
    .A2(net3539),
    .A1(net4772));
 sg13g2_inv_1 _27914_ (.Y(_00731_),
    .A(net3206));
 sg13g2_a22oi_1 _27915_ (.Y(_05633_),
    .B1(net3632),
    .B2(net2721),
    .A2(net3539),
    .A1(net4771));
 sg13g2_inv_1 _27916_ (.Y(_00732_),
    .A(_05633_));
 sg13g2_a22oi_1 _27917_ (.Y(_05634_),
    .B1(net3632),
    .B2(net2993),
    .A2(net3539),
    .A1(\u_inv.d_reg[199] ));
 sg13g2_inv_1 _27918_ (.Y(_00733_),
    .A(net2994));
 sg13g2_a22oi_1 _27919_ (.Y(_05635_),
    .B1(net3624),
    .B2(net2897),
    .A2(net3531),
    .A1(net3108));
 sg13g2_inv_1 _27920_ (.Y(_00734_),
    .A(_05635_));
 sg13g2_a22oi_1 _27921_ (.Y(_05636_),
    .B1(net3622),
    .B2(net2998),
    .A2(net3529),
    .A1(\u_inv.d_reg[201] ));
 sg13g2_inv_1 _27922_ (.Y(_00735_),
    .A(net2999));
 sg13g2_a22oi_1 _27923_ (.Y(_05637_),
    .B1(net3622),
    .B2(net2538),
    .A2(net3529),
    .A1(\u_inv.d_reg[202] ));
 sg13g2_inv_1 _27924_ (.Y(_00736_),
    .A(net2539));
 sg13g2_a22oi_1 _27925_ (.Y(_05638_),
    .B1(net3624),
    .B2(net2657),
    .A2(net3531),
    .A1(\u_inv.d_reg[203] ));
 sg13g2_inv_1 _27926_ (.Y(_00737_),
    .A(net2658));
 sg13g2_a22oi_1 _27927_ (.Y(_05639_),
    .B1(net3622),
    .B2(net2905),
    .A2(net3529),
    .A1(net3059));
 sg13g2_inv_1 _27928_ (.Y(_00738_),
    .A(_05639_));
 sg13g2_a22oi_1 _27929_ (.Y(_05640_),
    .B1(net3624),
    .B2(net3244),
    .A2(net3531),
    .A1(net3286));
 sg13g2_inv_1 _27930_ (.Y(_00739_),
    .A(_05640_));
 sg13g2_a22oi_1 _27931_ (.Y(_05641_),
    .B1(net3622),
    .B2(net3001),
    .A2(net3529),
    .A1(\u_inv.d_reg[206] ));
 sg13g2_inv_1 _27932_ (.Y(_00740_),
    .A(net3002));
 sg13g2_a22oi_1 _27933_ (.Y(_05642_),
    .B1(net3622),
    .B2(net2730),
    .A2(net3529),
    .A1(\u_inv.d_reg[207] ));
 sg13g2_inv_1 _27934_ (.Y(_00741_),
    .A(net2731));
 sg13g2_a22oi_1 _27935_ (.Y(_05643_),
    .B1(net3622),
    .B2(net2962),
    .A2(net3529),
    .A1(net4770));
 sg13g2_inv_1 _27936_ (.Y(_00742_),
    .A(net2963));
 sg13g2_a22oi_1 _27937_ (.Y(_05644_),
    .B1(net3622),
    .B2(net2804),
    .A2(net3529),
    .A1(net4769));
 sg13g2_inv_1 _27938_ (.Y(_00743_),
    .A(net2805));
 sg13g2_a22oi_1 _27939_ (.Y(_05645_),
    .B1(net3621),
    .B2(net2623),
    .A2(net3528),
    .A1(\u_inv.d_reg[210] ));
 sg13g2_inv_1 _27940_ (.Y(_00744_),
    .A(net2624));
 sg13g2_a22oi_1 _27941_ (.Y(_05646_),
    .B1(net3621),
    .B2(net2913),
    .A2(net3528),
    .A1(\u_inv.d_reg[211] ));
 sg13g2_inv_1 _27942_ (.Y(_00745_),
    .A(net2914));
 sg13g2_a22oi_1 _27943_ (.Y(_05647_),
    .B1(net3621),
    .B2(net3112),
    .A2(net3528),
    .A1(\u_inv.d_reg[212] ));
 sg13g2_inv_1 _27944_ (.Y(_00746_),
    .A(net3113));
 sg13g2_a22oi_1 _27945_ (.Y(_05648_),
    .B1(net3621),
    .B2(net2703),
    .A2(net3528),
    .A1(\u_inv.d_reg[213] ));
 sg13g2_inv_1 _27946_ (.Y(_00747_),
    .A(net2704));
 sg13g2_a22oi_1 _27947_ (.Y(_05649_),
    .B1(net3621),
    .B2(net2773),
    .A2(net3528),
    .A1(\u_inv.d_reg[214] ));
 sg13g2_inv_1 _27948_ (.Y(_00748_),
    .A(net2774));
 sg13g2_a22oi_1 _27949_ (.Y(_05650_),
    .B1(net3621),
    .B2(net2929),
    .A2(net3528),
    .A1(\u_inv.d_reg[215] ));
 sg13g2_inv_1 _27950_ (.Y(_00749_),
    .A(net2930));
 sg13g2_a22oi_1 _27951_ (.Y(_05651_),
    .B1(net3610),
    .B2(net2967),
    .A2(net3517),
    .A1(\u_inv.d_reg[216] ));
 sg13g2_inv_1 _27952_ (.Y(_00750_),
    .A(net2968));
 sg13g2_a22oi_1 _27953_ (.Y(_05652_),
    .B1(net3610),
    .B2(net2931),
    .A2(net3517),
    .A1(\u_inv.d_reg[217] ));
 sg13g2_inv_1 _27954_ (.Y(_00751_),
    .A(net2932));
 sg13g2_a22oi_1 _27955_ (.Y(_05653_),
    .B1(net3610),
    .B2(net2789),
    .A2(net3517),
    .A1(\u_inv.d_reg[218] ));
 sg13g2_inv_1 _27956_ (.Y(_00752_),
    .A(net2790));
 sg13g2_a22oi_1 _27957_ (.Y(_05654_),
    .B1(net3610),
    .B2(net2938),
    .A2(net3517),
    .A1(\u_inv.d_reg[219] ));
 sg13g2_inv_1 _27958_ (.Y(_00753_),
    .A(net2939));
 sg13g2_a22oi_1 _27959_ (.Y(_05655_),
    .B1(net3621),
    .B2(net2810),
    .A2(net3528),
    .A1(\u_inv.d_reg[220] ));
 sg13g2_inv_1 _27960_ (.Y(_00754_),
    .A(net2811));
 sg13g2_a22oi_1 _27961_ (.Y(_05656_),
    .B1(net3610),
    .B2(net2013),
    .A2(net3517),
    .A1(\u_inv.d_reg[221] ));
 sg13g2_inv_1 _27962_ (.Y(_00755_),
    .A(net2014));
 sg13g2_a22oi_1 _27963_ (.Y(_05657_),
    .B1(net3611),
    .B2(net3240),
    .A2(net3518),
    .A1(net3252));
 sg13g2_inv_1 _27964_ (.Y(_00756_),
    .A(_05657_));
 sg13g2_a22oi_1 _27965_ (.Y(_05658_),
    .B1(net3611),
    .B2(net2413),
    .A2(net3518),
    .A1(net3041));
 sg13g2_inv_1 _27966_ (.Y(_00757_),
    .A(_05658_));
 sg13g2_a22oi_1 _27967_ (.Y(_05659_),
    .B1(net3610),
    .B2(net2449),
    .A2(net3517),
    .A1(\u_inv.d_reg[224] ));
 sg13g2_inv_1 _27968_ (.Y(_00758_),
    .A(net2450));
 sg13g2_a22oi_1 _27969_ (.Y(_05660_),
    .B1(net3608),
    .B2(net2895),
    .A2(net3515),
    .A1(net3004));
 sg13g2_inv_1 _27970_ (.Y(_00759_),
    .A(_05660_));
 sg13g2_a22oi_1 _27971_ (.Y(_05661_),
    .B1(net3608),
    .B2(net3009),
    .A2(net3515),
    .A1(net4768));
 sg13g2_inv_1 _27972_ (.Y(_00760_),
    .A(net3010));
 sg13g2_a22oi_1 _27973_ (.Y(_05662_),
    .B1(net3608),
    .B2(net2752),
    .A2(net3515),
    .A1(\u_inv.d_reg[227] ));
 sg13g2_inv_1 _27974_ (.Y(_00761_),
    .A(net2753));
 sg13g2_a22oi_1 _27975_ (.Y(_05663_),
    .B1(net3608),
    .B2(net2822),
    .A2(net3515),
    .A1(net4767));
 sg13g2_inv_1 _27976_ (.Y(_00762_),
    .A(_05663_));
 sg13g2_a22oi_1 _27977_ (.Y(_05664_),
    .B1(net3608),
    .B2(net2515),
    .A2(net3515),
    .A1(net4766));
 sg13g2_inv_1 _27978_ (.Y(_00763_),
    .A(_05664_));
 sg13g2_a22oi_1 _27979_ (.Y(_05665_),
    .B1(net3608),
    .B2(net3051),
    .A2(net3515),
    .A1(\u_inv.d_reg[230] ));
 sg13g2_inv_1 _27980_ (.Y(_00764_),
    .A(net3052));
 sg13g2_a22oi_1 _27981_ (.Y(_05666_),
    .B1(net3598),
    .B2(net3032),
    .A2(net3505),
    .A1(\u_inv.d_reg[231] ));
 sg13g2_inv_1 _27982_ (.Y(_00765_),
    .A(net3033));
 sg13g2_a22oi_1 _27983_ (.Y(_05667_),
    .B1(net3598),
    .B2(net2519),
    .A2(net3505),
    .A1(\u_inv.d_reg[232] ));
 sg13g2_inv_1 _27984_ (.Y(_00766_),
    .A(net2520));
 sg13g2_a22oi_1 _27985_ (.Y(_05668_),
    .B1(net3600),
    .B2(net2918),
    .A2(net3507),
    .A1(\u_inv.d_reg[233] ));
 sg13g2_inv_1 _27986_ (.Y(_00767_),
    .A(net2919));
 sg13g2_a22oi_1 _27987_ (.Y(_05669_),
    .B1(net3598),
    .B2(net3035),
    .A2(net3505),
    .A1(\u_inv.d_reg[234] ));
 sg13g2_inv_1 _27988_ (.Y(_00768_),
    .A(net3036));
 sg13g2_a22oi_1 _27989_ (.Y(_05670_),
    .B1(net3598),
    .B2(net2644),
    .A2(net3505),
    .A1(\u_inv.d_reg[235] ));
 sg13g2_inv_1 _27990_ (.Y(_00769_),
    .A(net2645));
 sg13g2_a22oi_1 _27991_ (.Y(_05671_),
    .B1(net3598),
    .B2(net2194),
    .A2(net3505),
    .A1(net2800));
 sg13g2_inv_1 _27992_ (.Y(_00770_),
    .A(_05671_));
 sg13g2_a22oi_1 _27993_ (.Y(_05672_),
    .B1(net3598),
    .B2(net2390),
    .A2(net3505),
    .A1(\u_inv.d_reg[237] ));
 sg13g2_inv_1 _27994_ (.Y(_00771_),
    .A(net2391));
 sg13g2_a22oi_1 _27995_ (.Y(_05673_),
    .B1(net3598),
    .B2(net2669),
    .A2(net3505),
    .A1(\u_inv.d_reg[238] ));
 sg13g2_inv_1 _27996_ (.Y(_00772_),
    .A(net2670));
 sg13g2_a22oi_1 _27997_ (.Y(_05674_),
    .B1(net3598),
    .B2(net3045),
    .A2(net3505),
    .A1(net3155));
 sg13g2_inv_1 _27998_ (.Y(_00773_),
    .A(_05674_));
 sg13g2_a22oi_1 _27999_ (.Y(_05675_),
    .B1(net3596),
    .B2(net2230),
    .A2(net3503),
    .A1(net2699));
 sg13g2_inv_1 _28000_ (.Y(_00774_),
    .A(_05675_));
 sg13g2_a22oi_1 _28001_ (.Y(_05676_),
    .B1(net3596),
    .B2(net2088),
    .A2(net3503),
    .A1(net2760));
 sg13g2_inv_1 _28002_ (.Y(_00775_),
    .A(_05676_));
 sg13g2_a22oi_1 _28003_ (.Y(_05677_),
    .B1(net3596),
    .B2(net2758),
    .A2(net3503),
    .A1(\u_inv.d_reg[242] ));
 sg13g2_inv_1 _28004_ (.Y(_00776_),
    .A(net2759));
 sg13g2_a22oi_1 _28005_ (.Y(_05678_),
    .B1(net3596),
    .B2(net2850),
    .A2(net3503),
    .A1(\u_inv.d_reg[243] ));
 sg13g2_inv_1 _28006_ (.Y(_00777_),
    .A(net2851));
 sg13g2_a22oi_1 _28007_ (.Y(_05679_),
    .B1(net3596),
    .B2(net2127),
    .A2(net3503),
    .A1(net2692));
 sg13g2_inv_1 _28008_ (.Y(_00778_),
    .A(_05679_));
 sg13g2_a22oi_1 _28009_ (.Y(_05680_),
    .B1(net3596),
    .B2(net2275),
    .A2(net3503),
    .A1(\u_inv.d_reg[245] ));
 sg13g2_inv_1 _28010_ (.Y(_00779_),
    .A(net2276));
 sg13g2_a22oi_1 _28011_ (.Y(_05681_),
    .B1(net3596),
    .B2(net3073),
    .A2(net3503),
    .A1(\u_inv.d_reg[246] ));
 sg13g2_inv_1 _28012_ (.Y(_00780_),
    .A(net3074));
 sg13g2_a22oi_1 _28013_ (.Y(_05682_),
    .B1(net3596),
    .B2(net3131),
    .A2(net3503),
    .A1(\u_inv.d_reg[247] ));
 sg13g2_inv_1 _28014_ (.Y(_00781_),
    .A(net3132));
 sg13g2_a22oi_1 _28015_ (.Y(_05683_),
    .B1(net3588),
    .B2(net2388),
    .A2(net3495),
    .A1(\u_inv.d_reg[248] ));
 sg13g2_inv_1 _28016_ (.Y(_00782_),
    .A(net2389));
 sg13g2_a22oi_1 _28017_ (.Y(_05684_),
    .B1(net3588),
    .B2(net1870),
    .A2(net3495),
    .A1(net2384));
 sg13g2_inv_1 _28018_ (.Y(_00783_),
    .A(_05684_));
 sg13g2_a22oi_1 _28019_ (.Y(_05685_),
    .B1(net3588),
    .B2(net2776),
    .A2(net3495),
    .A1(\u_inv.d_reg[250] ));
 sg13g2_inv_1 _28020_ (.Y(_00784_),
    .A(net2777));
 sg13g2_a22oi_1 _28021_ (.Y(_05686_),
    .B1(net3588),
    .B2(net3056),
    .A2(net3495),
    .A1(\u_inv.d_reg[251] ));
 sg13g2_inv_1 _28022_ (.Y(_00785_),
    .A(net3057));
 sg13g2_a22oi_1 _28023_ (.Y(_05687_),
    .B1(net3588),
    .B2(net2743),
    .A2(net3495),
    .A1(\u_inv.d_reg[252] ));
 sg13g2_inv_1 _28024_ (.Y(_00786_),
    .A(net2744));
 sg13g2_a22oi_1 _28025_ (.Y(_05688_),
    .B1(net3588),
    .B2(net2637),
    .A2(net3495),
    .A1(\u_inv.d_reg[253] ));
 sg13g2_inv_1 _28026_ (.Y(_00787_),
    .A(net2638));
 sg13g2_a22oi_1 _28027_ (.Y(_05689_),
    .B1(net3588),
    .B2(net2714),
    .A2(net3495),
    .A1(net2892));
 sg13g2_inv_1 _28028_ (.Y(_00788_),
    .A(_05689_));
 sg13g2_a22oi_1 _28029_ (.Y(_05690_),
    .B1(net3588),
    .B2(net2452),
    .A2(net3495),
    .A1(net3022));
 sg13g2_inv_1 _28030_ (.Y(_00789_),
    .A(_05690_));
 sg13g2_a22oi_1 _28031_ (.Y(_05691_),
    .B1(net3608),
    .B2(net2570),
    .A2(net3515),
    .A1(net3034));
 sg13g2_inv_1 _28032_ (.Y(_00790_),
    .A(_05691_));
 sg13g2_nand2b_1 _28033_ (.Y(_00791_),
    .B(net3499),
    .A_N(net1297));
 sg13g2_a22oi_1 _28034_ (.Y(_00792_),
    .B1(net3592),
    .B2(_10576_),
    .A2(net3499),
    .A1(_10883_));
 sg13g2_a22oi_1 _28035_ (.Y(_00793_),
    .B1(net3592),
    .B2(_10575_),
    .A2(net3499),
    .A1(_10882_));
 sg13g2_a22oi_1 _28036_ (.Y(_00794_),
    .B1(net3593),
    .B2(_10574_),
    .A2(net3500),
    .A1(_10881_));
 sg13g2_a22oi_1 _28037_ (.Y(_05692_),
    .B1(net3593),
    .B2(\u_inv.f_next[4] ),
    .A2(net3500),
    .A1(net2424));
 sg13g2_inv_1 _28038_ (.Y(_00795_),
    .A(net2425));
 sg13g2_a22oi_1 _28039_ (.Y(_00796_),
    .B1(net3593),
    .B2(_10573_),
    .A2(net3500),
    .A1(_10880_));
 sg13g2_a22oi_1 _28040_ (.Y(_05693_),
    .B1(net3593),
    .B2(net2143),
    .A2(net3500),
    .A1(\u_inv.f_reg[6] ));
 sg13g2_inv_1 _28041_ (.Y(_00797_),
    .A(net2144));
 sg13g2_a22oi_1 _28042_ (.Y(_05694_),
    .B1(net3593),
    .B2(\u_inv.f_next[7] ),
    .A2(net3500),
    .A1(net2562));
 sg13g2_inv_1 _28043_ (.Y(_00798_),
    .A(net2563));
 sg13g2_a22oi_1 _28044_ (.Y(_05695_),
    .B1(net3594),
    .B2(\u_inv.f_next[8] ),
    .A2(net3501),
    .A1(net2613));
 sg13g2_inv_1 _28045_ (.Y(_00799_),
    .A(net2614));
 sg13g2_a22oi_1 _28046_ (.Y(_05696_),
    .B1(net3594),
    .B2(net2394),
    .A2(net3501),
    .A1(net2786));
 sg13g2_inv_1 _28047_ (.Y(_00800_),
    .A(_05696_));
 sg13g2_a22oi_1 _28048_ (.Y(_00801_),
    .B1(net3593),
    .B2(_10571_),
    .A2(net3500),
    .A1(_10879_));
 sg13g2_a22oi_1 _28049_ (.Y(_00802_),
    .B1(net3593),
    .B2(_10570_),
    .A2(net3500),
    .A1(_10878_));
 sg13g2_a22oi_1 _28050_ (.Y(_00803_),
    .B1(net3593),
    .B2(_10569_),
    .A2(net3500),
    .A1(_10877_));
 sg13g2_a22oi_1 _28051_ (.Y(_00804_),
    .B1(net3603),
    .B2(_10568_),
    .A2(net3510),
    .A1(_10876_));
 sg13g2_a22oi_1 _28052_ (.Y(_00805_),
    .B1(net3603),
    .B2(_10567_),
    .A2(net3510),
    .A1(_10875_));
 sg13g2_a22oi_1 _28053_ (.Y(_00806_),
    .B1(net3603),
    .B2(_10566_),
    .A2(net3510),
    .A1(_10874_));
 sg13g2_a22oi_1 _28054_ (.Y(_00807_),
    .B1(net3603),
    .B2(_10565_),
    .A2(net3510),
    .A1(_10873_));
 sg13g2_a22oi_1 _28055_ (.Y(_00808_),
    .B1(net3603),
    .B2(_10564_),
    .A2(net3510),
    .A1(_10872_));
 sg13g2_a22oi_1 _28056_ (.Y(_00809_),
    .B1(net3604),
    .B2(_10563_),
    .A2(net3511),
    .A1(_10871_));
 sg13g2_a22oi_1 _28057_ (.Y(_00810_),
    .B1(net3604),
    .B2(_10562_),
    .A2(net3511),
    .A1(_10870_));
 sg13g2_a22oi_1 _28058_ (.Y(_00811_),
    .B1(net3603),
    .B2(_10561_),
    .A2(net3510),
    .A1(_10869_));
 sg13g2_a22oi_1 _28059_ (.Y(_00812_),
    .B1(net3605),
    .B2(_10560_),
    .A2(net3512),
    .A1(_10868_));
 sg13g2_a22oi_1 _28060_ (.Y(_00813_),
    .B1(net3603),
    .B2(_10559_),
    .A2(net3510),
    .A1(_10867_));
 sg13g2_a22oi_1 _28061_ (.Y(_00814_),
    .B1(net3603),
    .B2(_10558_),
    .A2(net3510),
    .A1(_10866_));
 sg13g2_a22oi_1 _28062_ (.Y(_00815_),
    .B1(net3605),
    .B2(_10557_),
    .A2(net3512),
    .A1(_10865_));
 sg13g2_a22oi_1 _28063_ (.Y(_00816_),
    .B1(net3605),
    .B2(_10556_),
    .A2(net3512),
    .A1(_10864_));
 sg13g2_a22oi_1 _28064_ (.Y(_00817_),
    .B1(net3605),
    .B2(_10555_),
    .A2(net3512),
    .A1(_10863_));
 sg13g2_a22oi_1 _28065_ (.Y(_00818_),
    .B1(net3605),
    .B2(_10554_),
    .A2(net3512),
    .A1(_10862_));
 sg13g2_a22oi_1 _28066_ (.Y(_00819_),
    .B1(net3605),
    .B2(_10553_),
    .A2(net3512),
    .A1(_10861_));
 sg13g2_a22oi_1 _28067_ (.Y(_00820_),
    .B1(net3605),
    .B2(_10552_),
    .A2(net3512),
    .A1(_10860_));
 sg13g2_a22oi_1 _28068_ (.Y(_00821_),
    .B1(net3605),
    .B2(_10551_),
    .A2(net3512),
    .A1(_10859_));
 sg13g2_a22oi_1 _28069_ (.Y(_00822_),
    .B1(net3606),
    .B2(_10550_),
    .A2(net3513),
    .A1(_10858_));
 sg13g2_a22oi_1 _28070_ (.Y(_05697_),
    .B1(net3614),
    .B2(net2280),
    .A2(net3521),
    .A1(net2326));
 sg13g2_inv_1 _28071_ (.Y(_00823_),
    .A(_05697_));
 sg13g2_a22oi_1 _28072_ (.Y(_00824_),
    .B1(net3614),
    .B2(_10548_),
    .A2(net3521),
    .A1(_10857_));
 sg13g2_a22oi_1 _28073_ (.Y(_00825_),
    .B1(net3614),
    .B2(_10547_),
    .A2(net3521),
    .A1(_10856_));
 sg13g2_a22oi_1 _28074_ (.Y(_00826_),
    .B1(net3614),
    .B2(_10546_),
    .A2(net3521),
    .A1(_10855_));
 sg13g2_a22oi_1 _28075_ (.Y(_00827_),
    .B1(net3614),
    .B2(_10545_),
    .A2(net3521),
    .A1(_10854_));
 sg13g2_a22oi_1 _28076_ (.Y(_00828_),
    .B1(net3614),
    .B2(_10544_),
    .A2(net3521),
    .A1(_10853_));
 sg13g2_a22oi_1 _28077_ (.Y(_00829_),
    .B1(net3614),
    .B2(_10543_),
    .A2(net3521),
    .A1(_10852_));
 sg13g2_a22oi_1 _28078_ (.Y(_00830_),
    .B1(net3614),
    .B2(_10542_),
    .A2(net3521),
    .A1(_10851_));
 sg13g2_a22oi_1 _28079_ (.Y(_00831_),
    .B1(net3615),
    .B2(_10541_),
    .A2(net3522),
    .A1(_10850_));
 sg13g2_a22oi_1 _28080_ (.Y(_00832_),
    .B1(net3615),
    .B2(_10540_),
    .A2(net3522),
    .A1(_10849_));
 sg13g2_a22oi_1 _28081_ (.Y(_00833_),
    .B1(net3615),
    .B2(_10539_),
    .A2(net3522),
    .A1(_10848_));
 sg13g2_a22oi_1 _28082_ (.Y(_00834_),
    .B1(net3615),
    .B2(_10538_),
    .A2(net3522),
    .A1(_10847_));
 sg13g2_a22oi_1 _28083_ (.Y(_00835_),
    .B1(net3618),
    .B2(_10537_),
    .A2(net3525),
    .A1(_10846_));
 sg13g2_a22oi_1 _28084_ (.Y(_00836_),
    .B1(net3618),
    .B2(_10536_),
    .A2(net3525),
    .A1(_10845_));
 sg13g2_a22oi_1 _28085_ (.Y(_00837_),
    .B1(net3618),
    .B2(_10535_),
    .A2(net3525),
    .A1(_10844_));
 sg13g2_a22oi_1 _28086_ (.Y(_00838_),
    .B1(net3618),
    .B2(_10534_),
    .A2(net3525),
    .A1(_10843_));
 sg13g2_a22oi_1 _28087_ (.Y(_00839_),
    .B1(net3618),
    .B2(_10533_),
    .A2(net3525),
    .A1(_10842_));
 sg13g2_a22oi_1 _28088_ (.Y(_00840_),
    .B1(net3618),
    .B2(_10532_),
    .A2(net3525),
    .A1(_10841_));
 sg13g2_a22oi_1 _28089_ (.Y(_00841_),
    .B1(net3618),
    .B2(_10531_),
    .A2(net3525),
    .A1(_10840_));
 sg13g2_a22oi_1 _28090_ (.Y(_00842_),
    .B1(net3619),
    .B2(_10530_),
    .A2(net3526),
    .A1(_10839_));
 sg13g2_a22oi_1 _28091_ (.Y(_00843_),
    .B1(net3619),
    .B2(_10529_),
    .A2(net3526),
    .A1(_10838_));
 sg13g2_a22oi_1 _28092_ (.Y(_00844_),
    .B1(net3618),
    .B2(_10528_),
    .A2(net3525),
    .A1(_10837_));
 sg13g2_a22oi_1 _28093_ (.Y(_00845_),
    .B1(net3619),
    .B2(_10527_),
    .A2(net3526),
    .A1(_10836_));
 sg13g2_a22oi_1 _28094_ (.Y(_00846_),
    .B1(net3626),
    .B2(_10526_),
    .A2(net3533),
    .A1(_10835_));
 sg13g2_a22oi_1 _28095_ (.Y(_00847_),
    .B1(net3626),
    .B2(_10525_),
    .A2(net3533),
    .A1(_10834_));
 sg13g2_a22oi_1 _28096_ (.Y(_00848_),
    .B1(net3626),
    .B2(_10524_),
    .A2(net3533),
    .A1(_10833_));
 sg13g2_a22oi_1 _28097_ (.Y(_00849_),
    .B1(net3626),
    .B2(_10523_),
    .A2(net3533),
    .A1(_10832_));
 sg13g2_a22oi_1 _28098_ (.Y(_00850_),
    .B1(net3626),
    .B2(_10522_),
    .A2(net3533),
    .A1(_10831_));
 sg13g2_a22oi_1 _28099_ (.Y(_00851_),
    .B1(net3626),
    .B2(_10521_),
    .A2(net3533),
    .A1(_10830_));
 sg13g2_a22oi_1 _28100_ (.Y(_00852_),
    .B1(net3626),
    .B2(_10520_),
    .A2(net3533),
    .A1(_10829_));
 sg13g2_a22oi_1 _28101_ (.Y(_00853_),
    .B1(net3626),
    .B2(_10519_),
    .A2(net3533),
    .A1(_10828_));
 sg13g2_a22oi_1 _28102_ (.Y(_00854_),
    .B1(net3627),
    .B2(_10518_),
    .A2(net3534),
    .A1(_10827_));
 sg13g2_a22oi_1 _28103_ (.Y(_00855_),
    .B1(net3628),
    .B2(_10517_),
    .A2(net3535),
    .A1(_10826_));
 sg13g2_a22oi_1 _28104_ (.Y(_00856_),
    .B1(net3628),
    .B2(_10516_),
    .A2(net3535),
    .A1(_10825_));
 sg13g2_a22oi_1 _28105_ (.Y(_00857_),
    .B1(net3628),
    .B2(_10515_),
    .A2(net3535),
    .A1(_10824_));
 sg13g2_a22oi_1 _28106_ (.Y(_00858_),
    .B1(net3628),
    .B2(_10514_),
    .A2(net3535),
    .A1(_10823_));
 sg13g2_a22oi_1 _28107_ (.Y(_00859_),
    .B1(net3629),
    .B2(_10513_),
    .A2(net3536),
    .A1(_10822_));
 sg13g2_a22oi_1 _28108_ (.Y(_00860_),
    .B1(net3628),
    .B2(_10512_),
    .A2(net3535),
    .A1(_10821_));
 sg13g2_a22oi_1 _28109_ (.Y(_00861_),
    .B1(net3628),
    .B2(_10511_),
    .A2(net3535),
    .A1(_10820_));
 sg13g2_a22oi_1 _28110_ (.Y(_00862_),
    .B1(net3628),
    .B2(_10510_),
    .A2(net3535),
    .A1(_10819_));
 sg13g2_a22oi_1 _28111_ (.Y(_00863_),
    .B1(net3637),
    .B2(_10509_),
    .A2(net3544),
    .A1(_10818_));
 sg13g2_a22oi_1 _28112_ (.Y(_00864_),
    .B1(net3637),
    .B2(_10508_),
    .A2(net3544),
    .A1(_10817_));
 sg13g2_a22oi_1 _28113_ (.Y(_00865_),
    .B1(net3637),
    .B2(_10507_),
    .A2(net3544),
    .A1(_10816_));
 sg13g2_a22oi_1 _28114_ (.Y(_00866_),
    .B1(net3637),
    .B2(_10506_),
    .A2(net3544),
    .A1(_10815_));
 sg13g2_a22oi_1 _28115_ (.Y(_00867_),
    .B1(net3637),
    .B2(_10505_),
    .A2(net3544),
    .A1(_10814_));
 sg13g2_a22oi_1 _28116_ (.Y(_00868_),
    .B1(net3637),
    .B2(_10504_),
    .A2(net3544),
    .A1(_10813_));
 sg13g2_a22oi_1 _28117_ (.Y(_00869_),
    .B1(net3637),
    .B2(_10503_),
    .A2(net3544),
    .A1(_10812_));
 sg13g2_a22oi_1 _28118_ (.Y(_00870_),
    .B1(net3638),
    .B2(_10502_),
    .A2(net3545),
    .A1(_10811_));
 sg13g2_a22oi_1 _28119_ (.Y(_00871_),
    .B1(net3638),
    .B2(_10501_),
    .A2(net3545),
    .A1(_10810_));
 sg13g2_a22oi_1 _28120_ (.Y(_00872_),
    .B1(net3638),
    .B2(_10500_),
    .A2(net3545),
    .A1(_10809_));
 sg13g2_a22oi_1 _28121_ (.Y(_00873_),
    .B1(net3639),
    .B2(_10499_),
    .A2(net3546),
    .A1(_10808_));
 sg13g2_a22oi_1 _28122_ (.Y(_00874_),
    .B1(net3638),
    .B2(_10498_),
    .A2(net3545),
    .A1(_10807_));
 sg13g2_a22oi_1 _28123_ (.Y(_00875_),
    .B1(net3639),
    .B2(_10497_),
    .A2(net3546),
    .A1(_10806_));
 sg13g2_a22oi_1 _28124_ (.Y(_00876_),
    .B1(net3639),
    .B2(_10496_),
    .A2(net3546),
    .A1(_10805_));
 sg13g2_a22oi_1 _28125_ (.Y(_00877_),
    .B1(net3637),
    .B2(_10495_),
    .A2(net3544),
    .A1(_10804_));
 sg13g2_a22oi_1 _28126_ (.Y(_00878_),
    .B1(net3638),
    .B2(_10494_),
    .A2(net3545),
    .A1(_10803_));
 sg13g2_a22oi_1 _28127_ (.Y(_00879_),
    .B1(net3639),
    .B2(_10493_),
    .A2(net3546),
    .A1(_10802_));
 sg13g2_a22oi_1 _28128_ (.Y(_00880_),
    .B1(net3639),
    .B2(_10492_),
    .A2(net3546),
    .A1(_10801_));
 sg13g2_a22oi_1 _28129_ (.Y(_00881_),
    .B1(net3639),
    .B2(_10491_),
    .A2(net3546),
    .A1(_10800_));
 sg13g2_a22oi_1 _28130_ (.Y(_00882_),
    .B1(net3639),
    .B2(_10490_),
    .A2(net3546),
    .A1(_10799_));
 sg13g2_a22oi_1 _28131_ (.Y(_00883_),
    .B1(net3640),
    .B2(_10489_),
    .A2(net3547),
    .A1(_10798_));
 sg13g2_a22oi_1 _28132_ (.Y(_00884_),
    .B1(net3640),
    .B2(_10488_),
    .A2(net3547),
    .A1(_10797_));
 sg13g2_a22oi_1 _28133_ (.Y(_00885_),
    .B1(net3639),
    .B2(_10487_),
    .A2(net3546),
    .A1(_10796_));
 sg13g2_a22oi_1 _28134_ (.Y(_00886_),
    .B1(net3640),
    .B2(_10486_),
    .A2(net3547),
    .A1(_10795_));
 sg13g2_a22oi_1 _28135_ (.Y(_00887_),
    .B1(net3651),
    .B2(_10485_),
    .A2(net3558),
    .A1(_10794_));
 sg13g2_a22oi_1 _28136_ (.Y(_00888_),
    .B1(net3651),
    .B2(_10484_),
    .A2(net3558),
    .A1(_10793_));
 sg13g2_a22oi_1 _28137_ (.Y(_00889_),
    .B1(net3651),
    .B2(_10483_),
    .A2(net3558),
    .A1(_10792_));
 sg13g2_a22oi_1 _28138_ (.Y(_00890_),
    .B1(net3651),
    .B2(_10482_),
    .A2(net3558),
    .A1(_10791_));
 sg13g2_a22oi_1 _28139_ (.Y(_00891_),
    .B1(net3659),
    .B2(_10481_),
    .A2(net3566),
    .A1(_10790_));
 sg13g2_a22oi_1 _28140_ (.Y(_00892_),
    .B1(net3659),
    .B2(_10480_),
    .A2(net3566),
    .A1(_10789_));
 sg13g2_a22oi_1 _28141_ (.Y(_00893_),
    .B1(net3659),
    .B2(_10479_),
    .A2(net3566),
    .A1(_10788_));
 sg13g2_a22oi_1 _28142_ (.Y(_00894_),
    .B1(net3659),
    .B2(_10478_),
    .A2(net3566),
    .A1(_10787_));
 sg13g2_a22oi_1 _28143_ (.Y(_00895_),
    .B1(net3661),
    .B2(_10477_),
    .A2(net3568),
    .A1(_10786_));
 sg13g2_a22oi_1 _28144_ (.Y(_00896_),
    .B1(net3661),
    .B2(_10476_),
    .A2(net3568),
    .A1(_10785_));
 sg13g2_a22oi_1 _28145_ (.Y(_00897_),
    .B1(net3659),
    .B2(_10475_),
    .A2(net3566),
    .A1(_10784_));
 sg13g2_a22oi_1 _28146_ (.Y(_00898_),
    .B1(net3661),
    .B2(_10474_),
    .A2(net3568),
    .A1(_10783_));
 sg13g2_a22oi_1 _28147_ (.Y(_00899_),
    .B1(net3662),
    .B2(_10473_),
    .A2(net3569),
    .A1(_10782_));
 sg13g2_a22oi_1 _28148_ (.Y(_00900_),
    .B1(net3662),
    .B2(_10472_),
    .A2(net3569),
    .A1(_10781_));
 sg13g2_a22oi_1 _28149_ (.Y(_00901_),
    .B1(net3662),
    .B2(_10471_),
    .A2(net3569),
    .A1(_10780_));
 sg13g2_a22oi_1 _28150_ (.Y(_00902_),
    .B1(net3662),
    .B2(_10470_),
    .A2(net3569),
    .A1(_10779_));
 sg13g2_a22oi_1 _28151_ (.Y(_00903_),
    .B1(net3670),
    .B2(_10469_),
    .A2(net3577),
    .A1(_10778_));
 sg13g2_a22oi_1 _28152_ (.Y(_00904_),
    .B1(net3670),
    .B2(_10468_),
    .A2(net3577),
    .A1(_10777_));
 sg13g2_a22oi_1 _28153_ (.Y(_00905_),
    .B1(net3670),
    .B2(_10467_),
    .A2(net3577),
    .A1(_10776_));
 sg13g2_a22oi_1 _28154_ (.Y(_00906_),
    .B1(net3669),
    .B2(_10466_),
    .A2(net3576),
    .A1(_10775_));
 sg13g2_a22oi_1 _28155_ (.Y(_00907_),
    .B1(net3674),
    .B2(_10465_),
    .A2(net3581),
    .A1(_10774_));
 sg13g2_a22oi_1 _28156_ (.Y(_00908_),
    .B1(net3674),
    .B2(_10464_),
    .A2(net3581),
    .A1(_10773_));
 sg13g2_a22oi_1 _28157_ (.Y(_00909_),
    .B1(net3674),
    .B2(_10463_),
    .A2(net3581),
    .A1(_10772_));
 sg13g2_a22oi_1 _28158_ (.Y(_00910_),
    .B1(net3674),
    .B2(_10462_),
    .A2(net3581),
    .A1(_10771_));
 sg13g2_a22oi_1 _28159_ (.Y(_00911_),
    .B1(net3675),
    .B2(_10461_),
    .A2(net3582),
    .A1(_10770_));
 sg13g2_a22oi_1 _28160_ (.Y(_00912_),
    .B1(net3675),
    .B2(_10460_),
    .A2(net3582),
    .A1(_10769_));
 sg13g2_a22oi_1 _28161_ (.Y(_00913_),
    .B1(net3674),
    .B2(_10459_),
    .A2(net3581),
    .A1(_10768_));
 sg13g2_a22oi_1 _28162_ (.Y(_00914_),
    .B1(net3674),
    .B2(_10458_),
    .A2(net3581),
    .A1(_10767_));
 sg13g2_a22oi_1 _28163_ (.Y(_00915_),
    .B1(net3674),
    .B2(_10457_),
    .A2(net3581),
    .A1(_10766_));
 sg13g2_a22oi_1 _28164_ (.Y(_00916_),
    .B1(net3674),
    .B2(_10456_),
    .A2(net3581),
    .A1(_10765_));
 sg13g2_a22oi_1 _28165_ (.Y(_00917_),
    .B1(net3669),
    .B2(_10455_),
    .A2(net3576),
    .A1(_10764_));
 sg13g2_a22oi_1 _28166_ (.Y(_00918_),
    .B1(net3670),
    .B2(_10454_),
    .A2(net3577),
    .A1(_10763_));
 sg13g2_a22oi_1 _28167_ (.Y(_00919_),
    .B1(net3671),
    .B2(_10453_),
    .A2(net3578),
    .A1(_10762_));
 sg13g2_a22oi_1 _28168_ (.Y(_00920_),
    .B1(net3672),
    .B2(_10452_),
    .A2(net3579),
    .A1(_10761_));
 sg13g2_a22oi_1 _28169_ (.Y(_00921_),
    .B1(net3671),
    .B2(_10451_),
    .A2(net3578),
    .A1(_10760_));
 sg13g2_a22oi_1 _28170_ (.Y(_00922_),
    .B1(net3672),
    .B2(_10450_),
    .A2(net3579),
    .A1(_10759_));
 sg13g2_a22oi_1 _28171_ (.Y(_00923_),
    .B1(net3667),
    .B2(_10449_),
    .A2(net3574),
    .A1(_10758_));
 sg13g2_a22oi_1 _28172_ (.Y(_00924_),
    .B1(net3667),
    .B2(_10448_),
    .A2(net3574),
    .A1(_10757_));
 sg13g2_a22oi_1 _28173_ (.Y(_00925_),
    .B1(net3667),
    .B2(_10447_),
    .A2(net3574),
    .A1(_10756_));
 sg13g2_a22oi_1 _28174_ (.Y(_00926_),
    .B1(net3665),
    .B2(_10446_),
    .A2(net3572),
    .A1(_10755_));
 sg13g2_a22oi_1 _28175_ (.Y(_00927_),
    .B1(net3665),
    .B2(_10445_),
    .A2(net3572),
    .A1(_10754_));
 sg13g2_a22oi_1 _28176_ (.Y(_00928_),
    .B1(net3665),
    .B2(_10444_),
    .A2(net3572),
    .A1(_10753_));
 sg13g2_a22oi_1 _28177_ (.Y(_00929_),
    .B1(net3667),
    .B2(_10443_),
    .A2(net3574),
    .A1(_10752_));
 sg13g2_a22oi_1 _28178_ (.Y(_00930_),
    .B1(net3665),
    .B2(_10442_),
    .A2(net3572),
    .A1(_10751_));
 sg13g2_a22oi_1 _28179_ (.Y(_00931_),
    .B1(net3665),
    .B2(_10441_),
    .A2(net3572),
    .A1(_10750_));
 sg13g2_a22oi_1 _28180_ (.Y(_00932_),
    .B1(net3665),
    .B2(_10440_),
    .A2(net3572),
    .A1(_10749_));
 sg13g2_a22oi_1 _28181_ (.Y(_00933_),
    .B1(net3666),
    .B2(_10439_),
    .A2(net3573),
    .A1(_10748_));
 sg13g2_a22oi_1 _28182_ (.Y(_00934_),
    .B1(net3666),
    .B2(_10438_),
    .A2(net3573),
    .A1(_10747_));
 sg13g2_a22oi_1 _28183_ (.Y(_00935_),
    .B1(net3665),
    .B2(_10437_),
    .A2(net3572),
    .A1(_10746_));
 sg13g2_a22oi_1 _28184_ (.Y(_00936_),
    .B1(net3666),
    .B2(_10436_),
    .A2(net3573),
    .A1(_10745_));
 sg13g2_a22oi_1 _28185_ (.Y(_00937_),
    .B1(net3666),
    .B2(_10435_),
    .A2(net3573),
    .A1(_10744_));
 sg13g2_a22oi_1 _28186_ (.Y(_00938_),
    .B1(net3665),
    .B2(_10434_),
    .A2(net3572),
    .A1(_10743_));
 sg13g2_a22oi_1 _28187_ (.Y(_00939_),
    .B1(net3672),
    .B2(_10433_),
    .A2(net3579),
    .A1(_10742_));
 sg13g2_a22oi_1 _28188_ (.Y(_00940_),
    .B1(net3672),
    .B2(_10432_),
    .A2(net3579),
    .A1(_10741_));
 sg13g2_a22oi_1 _28189_ (.Y(_00941_),
    .B1(net3673),
    .B2(_10431_),
    .A2(net3580),
    .A1(_10740_));
 sg13g2_a22oi_1 _28190_ (.Y(_00942_),
    .B1(net3673),
    .B2(_10430_),
    .A2(net3580),
    .A1(_10739_));
 sg13g2_a22oi_1 _28191_ (.Y(_00943_),
    .B1(net3673),
    .B2(_10429_),
    .A2(net3580),
    .A1(_10738_));
 sg13g2_a22oi_1 _28192_ (.Y(_00944_),
    .B1(net3673),
    .B2(_10428_),
    .A2(net3580),
    .A1(_10737_));
 sg13g2_a22oi_1 _28193_ (.Y(_00945_),
    .B1(net3673),
    .B2(_10427_),
    .A2(net3580),
    .A1(_10736_));
 sg13g2_a22oi_1 _28194_ (.Y(_00946_),
    .B1(net3672),
    .B2(_10426_),
    .A2(net3579),
    .A1(_10735_));
 sg13g2_a22oi_1 _28195_ (.Y(_00947_),
    .B1(net3672),
    .B2(_10425_),
    .A2(net3579),
    .A1(_10734_));
 sg13g2_a22oi_1 _28196_ (.Y(_00948_),
    .B1(net3672),
    .B2(_10424_),
    .A2(net3579),
    .A1(_10733_));
 sg13g2_a22oi_1 _28197_ (.Y(_00949_),
    .B1(net3672),
    .B2(_10423_),
    .A2(net3579),
    .A1(_10732_));
 sg13g2_a22oi_1 _28198_ (.Y(_00950_),
    .B1(net3671),
    .B2(_10422_),
    .A2(net3578),
    .A1(_10731_));
 sg13g2_a22oi_1 _28199_ (.Y(_00951_),
    .B1(net3669),
    .B2(_10421_),
    .A2(net3576),
    .A1(_10730_));
 sg13g2_a22oi_1 _28200_ (.Y(_00952_),
    .B1(net3669),
    .B2(_10420_),
    .A2(net3576),
    .A1(_10729_));
 sg13g2_a22oi_1 _28201_ (.Y(_00953_),
    .B1(net3669),
    .B2(_10419_),
    .A2(net3576),
    .A1(_10728_));
 sg13g2_a22oi_1 _28202_ (.Y(_00954_),
    .B1(net3669),
    .B2(_10418_),
    .A2(net3576),
    .A1(_10727_));
 sg13g2_a22oi_1 _28203_ (.Y(_00955_),
    .B1(net3669),
    .B2(_10417_),
    .A2(net3576),
    .A1(_10726_));
 sg13g2_a22oi_1 _28204_ (.Y(_00956_),
    .B1(net3669),
    .B2(_10416_),
    .A2(net3576),
    .A1(_10725_));
 sg13g2_a22oi_1 _28205_ (.Y(_00957_),
    .B1(net3662),
    .B2(_10415_),
    .A2(net3569),
    .A1(_10724_));
 sg13g2_a22oi_1 _28206_ (.Y(_00958_),
    .B1(net3661),
    .B2(_10414_),
    .A2(net3568),
    .A1(_10723_));
 sg13g2_a22oi_1 _28207_ (.Y(_00959_),
    .B1(net3661),
    .B2(_10413_),
    .A2(net3568),
    .A1(_10722_));
 sg13g2_a22oi_1 _28208_ (.Y(_00960_),
    .B1(net3661),
    .B2(_10412_),
    .A2(net3568),
    .A1(_10721_));
 sg13g2_a22oi_1 _28209_ (.Y(_00961_),
    .B1(net3661),
    .B2(_10411_),
    .A2(net3568),
    .A1(_10720_));
 sg13g2_a22oi_1 _28210_ (.Y(_00962_),
    .B1(net3661),
    .B2(_10410_),
    .A2(net3568),
    .A1(_10719_));
 sg13g2_a22oi_1 _28211_ (.Y(_00963_),
    .B1(net3659),
    .B2(_10409_),
    .A2(net3566),
    .A1(_10718_));
 sg13g2_a22oi_1 _28212_ (.Y(_00964_),
    .B1(net3659),
    .B2(_10408_),
    .A2(net3566),
    .A1(_10717_));
 sg13g2_a22oi_1 _28213_ (.Y(_00965_),
    .B1(net3659),
    .B2(_10407_),
    .A2(net3566),
    .A1(_10716_));
 sg13g2_a22oi_1 _28214_ (.Y(_00966_),
    .B1(net3660),
    .B2(_10406_),
    .A2(net3567),
    .A1(_10715_));
 sg13g2_a22oi_1 _28215_ (.Y(_00967_),
    .B1(net3650),
    .B2(_10405_),
    .A2(net3557),
    .A1(_10714_));
 sg13g2_a22oi_1 _28216_ (.Y(_00968_),
    .B1(net3650),
    .B2(_10404_),
    .A2(net3557),
    .A1(_10713_));
 sg13g2_a22oi_1 _28217_ (.Y(_00969_),
    .B1(net3650),
    .B2(_10403_),
    .A2(net3557),
    .A1(_10712_));
 sg13g2_a22oi_1 _28218_ (.Y(_00970_),
    .B1(net3650),
    .B2(_10402_),
    .A2(net3557),
    .A1(_10711_));
 sg13g2_a22oi_1 _28219_ (.Y(_00971_),
    .B1(net3650),
    .B2(_10401_),
    .A2(net3557),
    .A1(_10710_));
 sg13g2_a22oi_1 _28220_ (.Y(_00972_),
    .B1(net3650),
    .B2(_10400_),
    .A2(net3557),
    .A1(_10709_));
 sg13g2_a22oi_1 _28221_ (.Y(_00973_),
    .B1(net3650),
    .B2(_10399_),
    .A2(net3557),
    .A1(_10708_));
 sg13g2_a22oi_1 _28222_ (.Y(_00974_),
    .B1(net3650),
    .B2(_10398_),
    .A2(net3557),
    .A1(_10707_));
 sg13g2_a22oi_1 _28223_ (.Y(_00975_),
    .B1(net3649),
    .B2(_10397_),
    .A2(net3556),
    .A1(_10706_));
 sg13g2_a22oi_1 _28224_ (.Y(_00976_),
    .B1(net3649),
    .B2(_10396_),
    .A2(net3556),
    .A1(_10705_));
 sg13g2_a22oi_1 _28225_ (.Y(_00977_),
    .B1(net3649),
    .B2(_10395_),
    .A2(net3556),
    .A1(_10704_));
 sg13g2_a22oi_1 _28226_ (.Y(_00978_),
    .B1(net3649),
    .B2(_10394_),
    .A2(net3556),
    .A1(_10703_));
 sg13g2_a22oi_1 _28227_ (.Y(_00979_),
    .B1(net3653),
    .B2(_10393_),
    .A2(net3560),
    .A1(_10702_));
 sg13g2_a22oi_1 _28228_ (.Y(_00980_),
    .B1(net3649),
    .B2(_10392_),
    .A2(net3556),
    .A1(_10701_));
 sg13g2_a22oi_1 _28229_ (.Y(_00981_),
    .B1(net3649),
    .B2(_10391_),
    .A2(net3556),
    .A1(_10700_));
 sg13g2_a22oi_1 _28230_ (.Y(_00982_),
    .B1(net3653),
    .B2(_10390_),
    .A2(net3560),
    .A1(_10699_));
 sg13g2_a22oi_1 _28231_ (.Y(_00983_),
    .B1(net3628),
    .B2(_10389_),
    .A2(net3535),
    .A1(_10698_));
 sg13g2_a22oi_1 _28232_ (.Y(_00984_),
    .B1(net3629),
    .B2(_10388_),
    .A2(net3536),
    .A1(_10697_));
 sg13g2_a22oi_1 _28233_ (.Y(_00985_),
    .B1(net3629),
    .B2(_10387_),
    .A2(net3536),
    .A1(_10696_));
 sg13g2_a22oi_1 _28234_ (.Y(_00986_),
    .B1(net3629),
    .B2(_10386_),
    .A2(net3536),
    .A1(_10695_));
 sg13g2_a22oi_1 _28235_ (.Y(_00987_),
    .B1(net3627),
    .B2(_10385_),
    .A2(net3534),
    .A1(_10694_));
 sg13g2_a22oi_1 _28236_ (.Y(_00988_),
    .B1(net3627),
    .B2(_10384_),
    .A2(net3534),
    .A1(_10693_));
 sg13g2_a22oi_1 _28237_ (.Y(_00989_),
    .B1(net3627),
    .B2(_10383_),
    .A2(net3534),
    .A1(_10692_));
 sg13g2_a22oi_1 _28238_ (.Y(_00990_),
    .B1(net3627),
    .B2(_10382_),
    .A2(net3534),
    .A1(_10691_));
 sg13g2_a22oi_1 _28239_ (.Y(_00991_),
    .B1(net3627),
    .B2(_10381_),
    .A2(net3534),
    .A1(_10690_));
 sg13g2_a22oi_1 _28240_ (.Y(_00992_),
    .B1(net3627),
    .B2(_10380_),
    .A2(net3534),
    .A1(_10689_));
 sg13g2_a22oi_1 _28241_ (.Y(_00993_),
    .B1(net3617),
    .B2(_10379_),
    .A2(net3524),
    .A1(_10688_));
 sg13g2_a22oi_1 _28242_ (.Y(_00994_),
    .B1(net3620),
    .B2(_10378_),
    .A2(net3527),
    .A1(_10687_));
 sg13g2_a22oi_1 _28243_ (.Y(_00995_),
    .B1(net3619),
    .B2(_10377_),
    .A2(net3526),
    .A1(_10686_));
 sg13g2_a22oi_1 _28244_ (.Y(_00996_),
    .B1(net3620),
    .B2(_10376_),
    .A2(net3527),
    .A1(_10685_));
 sg13g2_a22oi_1 _28245_ (.Y(_00997_),
    .B1(net3617),
    .B2(_10375_),
    .A2(net3524),
    .A1(_10684_));
 sg13g2_a22oi_1 _28246_ (.Y(_00998_),
    .B1(net3620),
    .B2(_10374_),
    .A2(net3527),
    .A1(_10683_));
 sg13g2_a22oi_1 _28247_ (.Y(_00999_),
    .B1(net3617),
    .B2(_10373_),
    .A2(net3524),
    .A1(_10682_));
 sg13g2_a22oi_1 _28248_ (.Y(_01000_),
    .B1(net3617),
    .B2(_10372_),
    .A2(net3524),
    .A1(_10681_));
 sg13g2_a22oi_1 _28249_ (.Y(_01001_),
    .B1(net3617),
    .B2(_10371_),
    .A2(net3524),
    .A1(_10680_));
 sg13g2_a22oi_1 _28250_ (.Y(_01002_),
    .B1(net3617),
    .B2(_10370_),
    .A2(net3524),
    .A1(_10679_));
 sg13g2_a22oi_1 _28251_ (.Y(_01003_),
    .B1(net3617),
    .B2(_10369_),
    .A2(net3524),
    .A1(_10678_));
 sg13g2_a22oi_1 _28252_ (.Y(_01004_),
    .B1(net3617),
    .B2(_10368_),
    .A2(net3524),
    .A1(_10677_));
 sg13g2_a22oi_1 _28253_ (.Y(_01005_),
    .B1(net3613),
    .B2(_10367_),
    .A2(net3520),
    .A1(_10676_));
 sg13g2_a22oi_1 _28254_ (.Y(_01006_),
    .B1(net3616),
    .B2(_10366_),
    .A2(net3523),
    .A1(_10675_));
 sg13g2_a22oi_1 _28255_ (.Y(_01007_),
    .B1(net3613),
    .B2(_10365_),
    .A2(net3520),
    .A1(_10674_));
 sg13g2_a22oi_1 _28256_ (.Y(_01008_),
    .B1(net3613),
    .B2(_10364_),
    .A2(net3520),
    .A1(_10673_));
 sg13g2_a22oi_1 _28257_ (.Y(_01009_),
    .B1(net3613),
    .B2(_10363_),
    .A2(net3520),
    .A1(_10672_));
 sg13g2_a22oi_1 _28258_ (.Y(_01010_),
    .B1(net3613),
    .B2(_10362_),
    .A2(net3520),
    .A1(_10671_));
 sg13g2_a22oi_1 _28259_ (.Y(_01011_),
    .B1(net3606),
    .B2(_10361_),
    .A2(net3513),
    .A1(_10670_));
 sg13g2_a22oi_1 _28260_ (.Y(_01012_),
    .B1(net3613),
    .B2(_10360_),
    .A2(net3520),
    .A1(_10669_));
 sg13g2_a22oi_1 _28261_ (.Y(_01013_),
    .B1(net3613),
    .B2(_10359_),
    .A2(net3520),
    .A1(_10668_));
 sg13g2_a22oi_1 _28262_ (.Y(_01014_),
    .B1(net3613),
    .B2(_10358_),
    .A2(net3520),
    .A1(_10667_));
 sg13g2_a22oi_1 _28263_ (.Y(_01015_),
    .B1(net3606),
    .B2(_10357_),
    .A2(net3513),
    .A1(_10666_));
 sg13g2_a22oi_1 _28264_ (.Y(_01016_),
    .B1(net3606),
    .B2(_10356_),
    .A2(net3513),
    .A1(_10665_));
 sg13g2_a22oi_1 _28265_ (.Y(_01017_),
    .B1(net3602),
    .B2(_10355_),
    .A2(net3509),
    .A1(_10664_));
 sg13g2_a22oi_1 _28266_ (.Y(_01018_),
    .B1(net3601),
    .B2(_10354_),
    .A2(net3508),
    .A1(_10663_));
 sg13g2_a22oi_1 _28267_ (.Y(_01019_),
    .B1(net3602),
    .B2(_10353_),
    .A2(net3509),
    .A1(_10662_));
 sg13g2_a22oi_1 _28268_ (.Y(_01020_),
    .B1(net3604),
    .B2(_10352_),
    .A2(net3511),
    .A1(_10661_));
 sg13g2_a22oi_1 _28269_ (.Y(_01021_),
    .B1(net3601),
    .B2(_10351_),
    .A2(net3508),
    .A1(_10660_));
 sg13g2_a22oi_1 _28270_ (.Y(_01022_),
    .B1(net3602),
    .B2(_10350_),
    .A2(net3509),
    .A1(_10659_));
 sg13g2_a22oi_1 _28271_ (.Y(_01023_),
    .B1(net3602),
    .B2(_10349_),
    .A2(net3509),
    .A1(_10658_));
 sg13g2_a22oi_1 _28272_ (.Y(_01024_),
    .B1(net3602),
    .B2(_10348_),
    .A2(net3509),
    .A1(_10657_));
 sg13g2_a22oi_1 _28273_ (.Y(_01025_),
    .B1(net3601),
    .B2(_10347_),
    .A2(net3508),
    .A1(_10656_));
 sg13g2_a22oi_1 _28274_ (.Y(_01026_),
    .B1(net3601),
    .B2(_10346_),
    .A2(net3508),
    .A1(_10655_));
 sg13g2_a22oi_1 _28275_ (.Y(_01027_),
    .B1(net3601),
    .B2(_10345_),
    .A2(net3508),
    .A1(_10654_));
 sg13g2_a22oi_1 _28276_ (.Y(_01028_),
    .B1(net3601),
    .B2(_10344_),
    .A2(net3508),
    .A1(_10653_));
 sg13g2_a22oi_1 _28277_ (.Y(_01029_),
    .B1(net3601),
    .B2(_10343_),
    .A2(net3508),
    .A1(_10652_));
 sg13g2_a22oi_1 _28278_ (.Y(_01030_),
    .B1(net3601),
    .B2(_10342_),
    .A2(net3508),
    .A1(_10651_));
 sg13g2_a22oi_1 _28279_ (.Y(_01031_),
    .B1(net3590),
    .B2(_10341_),
    .A2(net3497),
    .A1(_10650_));
 sg13g2_a22oi_1 _28280_ (.Y(_01032_),
    .B1(net3591),
    .B2(_10340_),
    .A2(net3498),
    .A1(_10649_));
 sg13g2_a22oi_1 _28281_ (.Y(_01033_),
    .B1(net3591),
    .B2(_10339_),
    .A2(net3498),
    .A1(_10648_));
 sg13g2_a22oi_1 _28282_ (.Y(_01034_),
    .B1(net3590),
    .B2(_10338_),
    .A2(net3497),
    .A1(_10647_));
 sg13g2_a22oi_1 _28283_ (.Y(_01035_),
    .B1(net3590),
    .B2(_10337_),
    .A2(net3497),
    .A1(_10646_));
 sg13g2_a22oi_1 _28284_ (.Y(_01036_),
    .B1(net3590),
    .B2(_10336_),
    .A2(net3497),
    .A1(_10645_));
 sg13g2_a22oi_1 _28285_ (.Y(_01037_),
    .B1(net3590),
    .B2(_10335_),
    .A2(net3497),
    .A1(_10644_));
 sg13g2_a22oi_1 _28286_ (.Y(_01038_),
    .B1(net3590),
    .B2(_10334_),
    .A2(net3497),
    .A1(_10643_));
 sg13g2_a22oi_1 _28287_ (.Y(_01039_),
    .B1(net3590),
    .B2(_10333_),
    .A2(net3497),
    .A1(_10642_));
 sg13g2_a22oi_1 _28288_ (.Y(_01040_),
    .B1(net3591),
    .B2(_10332_),
    .A2(net3498),
    .A1(_10641_));
 sg13g2_a22oi_1 _28289_ (.Y(_01041_),
    .B1(net3591),
    .B2(_10331_),
    .A2(net3498),
    .A1(_10640_));
 sg13g2_a22oi_1 _28290_ (.Y(_01042_),
    .B1(net3592),
    .B2(_10330_),
    .A2(net3499),
    .A1(_10639_));
 sg13g2_a22oi_1 _28291_ (.Y(_01043_),
    .B1(net3592),
    .B2(_10329_),
    .A2(net3499),
    .A1(_10638_));
 sg13g2_a22oi_1 _28292_ (.Y(_01044_),
    .B1(net3592),
    .B2(_10328_),
    .A2(net3499),
    .A1(_10637_));
 sg13g2_a22oi_1 _28293_ (.Y(_01045_),
    .B1(net3592),
    .B2(_10327_),
    .A2(net3499),
    .A1(_10636_));
 sg13g2_a22oi_1 _28294_ (.Y(_01046_),
    .B1(net3591),
    .B2(_10326_),
    .A2(net3498),
    .A1(_10635_));
 sg13g2_a22oi_1 _28295_ (.Y(_05698_),
    .B1(net3590),
    .B2(net4959),
    .A2(net3497),
    .A1(net4725));
 sg13g2_inv_2 _28296_ (.Y(_01047_),
    .A(_05698_));
 sg13g2_a21oi_2 _28297_ (.B1(_11046_),
    .Y(_05699_),
    .A2(net4453),
    .A1(inv_done));
 sg13g2_nand2b_2 _28298_ (.Y(_05700_),
    .B(_11043_),
    .A_N(_11046_));
 sg13g2_or2_1 _28299_ (.X(_05701_),
    .B(\u_inv.d_reg[152] ),
    .A(\u_inv.d_reg[153] ));
 sg13g2_or2_1 _28300_ (.X(_05702_),
    .B(_05701_),
    .A(\u_inv.d_reg[154] ));
 sg13g2_nand2b_1 _28301_ (.Y(_05703_),
    .B(_10915_),
    .A_N(_05702_));
 sg13g2_or2_1 _28302_ (.X(_05704_),
    .B(_05703_),
    .A(\u_inv.d_reg[156] ));
 sg13g2_nor2_1 _28303_ (.A(\u_inv.d_reg[157] ),
    .B(_05704_),
    .Y(_05705_));
 sg13g2_inv_1 _28304_ (.Y(_05706_),
    .A(_05705_));
 sg13g2_or2_1 _28305_ (.X(_05707_),
    .B(\u_inv.d_reg[144] ),
    .A(\u_inv.d_reg[145] ));
 sg13g2_or2_1 _28306_ (.X(_05708_),
    .B(_05707_),
    .A(\u_inv.d_reg[146] ));
 sg13g2_nor2_1 _28307_ (.A(\u_inv.d_reg[147] ),
    .B(_05708_),
    .Y(_05709_));
 sg13g2_or2_1 _28308_ (.X(_05710_),
    .B(\u_inv.d_reg[148] ),
    .A(\u_inv.d_reg[149] ));
 sg13g2_or2_1 _28309_ (.X(_05711_),
    .B(_05710_),
    .A(net4776));
 sg13g2_nor2_1 _28310_ (.A(\u_inv.d_reg[158] ),
    .B(_05706_),
    .Y(_05712_));
 sg13g2_nor2_1 _28311_ (.A(\u_inv.d_reg[151] ),
    .B(_05711_),
    .Y(_05713_));
 sg13g2_nor3_1 _28312_ (.A(\u_inv.d_reg[159] ),
    .B(\u_inv.d_reg[151] ),
    .C(_05711_),
    .Y(_05714_));
 sg13g2_or2_1 _28313_ (.X(_05715_),
    .B(\u_inv.d_reg[120] ),
    .A(\u_inv.d_reg[121] ));
 sg13g2_or2_1 _28314_ (.X(_05716_),
    .B(_05715_),
    .A(\u_inv.d_reg[122] ));
 sg13g2_or2_1 _28315_ (.X(_05717_),
    .B(_05716_),
    .A(\u_inv.d_reg[123] ));
 sg13g2_or3_1 _28316_ (.A(\u_inv.d_reg[125] ),
    .B(\u_inv.d_reg[124] ),
    .C(_05717_),
    .X(_05718_));
 sg13g2_or3_1 _28317_ (.A(net4797),
    .B(net4799),
    .C(net4796),
    .X(_05719_));
 sg13g2_or4_1 _28318_ (.A(net4797),
    .B(net4799),
    .C(\u_inv.d_reg[3] ),
    .D(net4796),
    .X(_05720_));
 sg13g2_or2_1 _28319_ (.X(_05721_),
    .B(_05720_),
    .A(\u_inv.d_reg[4] ));
 sg13g2_or4_1 _28320_ (.A(net4795),
    .B(\u_inv.d_reg[5] ),
    .C(\u_inv.d_reg[4] ),
    .D(_05720_),
    .X(_05722_));
 sg13g2_nor3_1 _28321_ (.A(\u_inv.d_reg[8] ),
    .B(net4794),
    .C(_05722_),
    .Y(_05723_));
 sg13g2_nand2_1 _28322_ (.Y(_05724_),
    .A(_10955_),
    .B(_10956_));
 sg13g2_or4_1 _28323_ (.A(\u_inv.d_reg[10] ),
    .B(\u_inv.d_reg[7] ),
    .C(_05722_),
    .D(_05724_),
    .X(_05725_));
 sg13g2_nor3_1 _28324_ (.A(\u_inv.d_reg[12] ),
    .B(net4792),
    .C(_05725_),
    .Y(_05726_));
 sg13g2_nor4_1 _28325_ (.A(\u_inv.d_reg[13] ),
    .B(\u_inv.d_reg[12] ),
    .C(net4792),
    .D(_05725_),
    .Y(_05727_));
 sg13g2_or4_1 _28326_ (.A(\u_inv.d_reg[13] ),
    .B(\u_inv.d_reg[12] ),
    .C(net4792),
    .D(_05725_),
    .X(_05728_));
 sg13g2_nor3_1 _28327_ (.A(\u_inv.d_reg[15] ),
    .B(\u_inv.d_reg[14] ),
    .C(_05728_),
    .Y(_05729_));
 sg13g2_nor2_1 _28328_ (.A(net4791),
    .B(\u_inv.d_reg[16] ),
    .Y(_05730_));
 sg13g2_nand4_1 _28329_ (.B(_10953_),
    .C(_05727_),
    .A(_10952_),
    .Y(_05731_),
    .D(_05730_));
 sg13g2_or4_1 _28330_ (.A(\u_inv.d_reg[19] ),
    .B(net4790),
    .C(net4791),
    .D(\u_inv.d_reg[16] ),
    .X(_05732_));
 sg13g2_nor4_2 _28331_ (.A(\u_inv.d_reg[15] ),
    .B(\u_inv.d_reg[14] ),
    .C(_05728_),
    .Y(_05733_),
    .D(_05732_));
 sg13g2_or4_1 _28332_ (.A(\u_inv.d_reg[15] ),
    .B(\u_inv.d_reg[14] ),
    .C(_05728_),
    .D(_05732_),
    .X(_05734_));
 sg13g2_nor2_1 _28333_ (.A(\u_inv.d_reg[21] ),
    .B(\u_inv.d_reg[20] ),
    .Y(_05735_));
 sg13g2_nand2_1 _28334_ (.Y(_05736_),
    .A(_05733_),
    .B(_05735_));
 sg13g2_nor2_1 _28335_ (.A(\u_inv.d_reg[23] ),
    .B(\u_inv.d_reg[22] ),
    .Y(_05737_));
 sg13g2_nand3_1 _28336_ (.B(_05735_),
    .C(_05737_),
    .A(_05733_),
    .Y(_05738_));
 sg13g2_nand4_1 _28337_ (.B(_05733_),
    .C(_05735_),
    .A(_10949_),
    .Y(_05739_),
    .D(_05737_));
 sg13g2_nor3_1 _28338_ (.A(\u_inv.d_reg[26] ),
    .B(net4788),
    .C(_05739_),
    .Y(_05740_));
 sg13g2_nor4_2 _28339_ (.A(\u_inv.d_reg[27] ),
    .B(net4787),
    .C(net4788),
    .Y(_05741_),
    .D(_05739_));
 sg13g2_nor2_1 _28340_ (.A(\u_inv.d_reg[29] ),
    .B(\u_inv.d_reg[28] ),
    .Y(_05742_));
 sg13g2_nand2_1 _28341_ (.Y(_05743_),
    .A(_05741_),
    .B(_05742_));
 sg13g2_and4_1 _28342_ (.A(_10946_),
    .B(_10947_),
    .C(_05741_),
    .D(_05742_),
    .X(_05744_));
 sg13g2_nand4_1 _28343_ (.B(_10947_),
    .C(_05741_),
    .A(_10946_),
    .Y(_05745_),
    .D(_05742_));
 sg13g2_or2_1 _28344_ (.X(_05746_),
    .B(\u_inv.d_reg[32] ),
    .A(\u_inv.d_reg[33] ));
 sg13g2_or3_1 _28345_ (.A(\u_inv.d_reg[35] ),
    .B(\u_inv.d_reg[34] ),
    .C(_05746_),
    .X(_05747_));
 sg13g2_or2_1 _28346_ (.X(_05748_),
    .B(_05747_),
    .A(\u_inv.d_reg[36] ));
 sg13g2_nor4_2 _28347_ (.A(\u_inv.d_reg[39] ),
    .B(\u_inv.d_reg[38] ),
    .C(\u_inv.d_reg[37] ),
    .Y(_05749_),
    .D(_05748_));
 sg13g2_nand2_1 _28348_ (.Y(_05750_),
    .A(_05744_),
    .B(_05749_));
 sg13g2_or2_1 _28349_ (.X(_05751_),
    .B(\u_inv.d_reg[40] ),
    .A(\u_inv.d_reg[41] ));
 sg13g2_nor3_1 _28350_ (.A(\u_inv.d_reg[43] ),
    .B(net4786),
    .C(_05751_),
    .Y(_05752_));
 sg13g2_nand3_1 _28351_ (.B(_05749_),
    .C(_05752_),
    .A(_05744_),
    .Y(_05753_));
 sg13g2_or2_1 _28352_ (.X(_05754_),
    .B(\u_inv.d_reg[44] ),
    .A(\u_inv.d_reg[45] ));
 sg13g2_nor3_1 _28353_ (.A(\u_inv.d_reg[47] ),
    .B(\u_inv.d_reg[46] ),
    .C(_05754_),
    .Y(_05755_));
 sg13g2_nand4_1 _28354_ (.B(_05749_),
    .C(_05752_),
    .A(_05744_),
    .Y(_05756_),
    .D(_05755_));
 sg13g2_or2_1 _28355_ (.X(_05757_),
    .B(\u_inv.d_reg[48] ),
    .A(\u_inv.d_reg[49] ));
 sg13g2_nor3_1 _28356_ (.A(\u_inv.d_reg[51] ),
    .B(\u_inv.d_reg[50] ),
    .C(_05757_),
    .Y(_05758_));
 sg13g2_inv_1 _28357_ (.Y(_05759_),
    .A(_05758_));
 sg13g2_nand2_1 _28358_ (.Y(_05760_),
    .A(_10937_),
    .B(_10938_));
 sg13g2_or3_1 _28359_ (.A(_05756_),
    .B(_05759_),
    .C(_05760_),
    .X(_05761_));
 sg13g2_or2_1 _28360_ (.X(_05762_),
    .B(\u_inv.d_reg[54] ),
    .A(\u_inv.d_reg[55] ));
 sg13g2_nor4_2 _28361_ (.A(_05756_),
    .B(_05759_),
    .C(_05760_),
    .Y(_05763_),
    .D(_05762_));
 sg13g2_nor4_2 _28362_ (.A(\u_inv.d_reg[59] ),
    .B(net4785),
    .C(\u_inv.d_reg[57] ),
    .Y(_05764_),
    .D(\u_inv.d_reg[56] ));
 sg13g2_nand2_1 _28363_ (.Y(_05765_),
    .A(net3493),
    .B(_05764_));
 sg13g2_nor4_2 _28364_ (.A(\u_inv.d_reg[63] ),
    .B(\u_inv.d_reg[62] ),
    .C(\u_inv.d_reg[61] ),
    .Y(_05766_),
    .D(\u_inv.d_reg[60] ));
 sg13g2_nand3_1 _28365_ (.B(_05764_),
    .C(_05766_),
    .A(net3493),
    .Y(_05767_));
 sg13g2_or2_1 _28366_ (.X(_05768_),
    .B(net4784),
    .A(\u_inv.d_reg[65] ));
 sg13g2_or2_1 _28367_ (.X(_05769_),
    .B(_05768_),
    .A(\u_inv.d_reg[66] ));
 sg13g2_nor2_1 _28368_ (.A(\u_inv.d_reg[67] ),
    .B(_05769_),
    .Y(_05770_));
 sg13g2_or2_1 _28369_ (.X(_05771_),
    .B(\u_inv.d_reg[68] ),
    .A(\u_inv.d_reg[69] ));
 sg13g2_or2_1 _28370_ (.X(_05772_),
    .B(_05771_),
    .A(\u_inv.d_reg[70] ));
 sg13g2_nor4_1 _28371_ (.A(\u_inv.d_reg[71] ),
    .B(\u_inv.d_reg[67] ),
    .C(_05769_),
    .D(_05772_),
    .Y(_05773_));
 sg13g2_or2_1 _28372_ (.X(_05774_),
    .B(\u_inv.d_reg[72] ),
    .A(\u_inv.d_reg[73] ));
 sg13g2_or2_1 _28373_ (.X(_05775_),
    .B(_05774_),
    .A(\u_inv.d_reg[74] ));
 sg13g2_nor2_1 _28374_ (.A(\u_inv.d_reg[75] ),
    .B(_05775_),
    .Y(_05776_));
 sg13g2_nor4_1 _28375_ (.A(\u_inv.d_reg[79] ),
    .B(\u_inv.d_reg[78] ),
    .C(\u_inv.d_reg[77] ),
    .D(\u_inv.d_reg[76] ),
    .Y(_05777_));
 sg13g2_nand3_1 _28376_ (.B(_05776_),
    .C(_05777_),
    .A(_05773_),
    .Y(_05778_));
 sg13g2_inv_1 _28377_ (.Y(_05779_),
    .A(_05778_));
 sg13g2_or2_1 _28378_ (.X(_05780_),
    .B(\u_inv.d_reg[80] ),
    .A(\u_inv.d_reg[81] ));
 sg13g2_or2_1 _28379_ (.X(_05781_),
    .B(_05780_),
    .A(\u_inv.d_reg[82] ));
 sg13g2_or2_1 _28380_ (.X(_05782_),
    .B(\u_inv.d_reg[84] ),
    .A(\u_inv.d_reg[85] ));
 sg13g2_or2_1 _28381_ (.X(_05783_),
    .B(_05781_),
    .A(\u_inv.d_reg[83] ));
 sg13g2_nor2_1 _28382_ (.A(\u_inv.d_reg[86] ),
    .B(_05782_),
    .Y(_05784_));
 sg13g2_nand2b_1 _28383_ (.Y(_05785_),
    .B(_05784_),
    .A_N(\u_inv.d_reg[87] ));
 sg13g2_nor3_1 _28384_ (.A(_05778_),
    .B(_05783_),
    .C(_05785_),
    .Y(_05786_));
 sg13g2_or2_1 _28385_ (.X(_05787_),
    .B(\u_inv.d_reg[88] ),
    .A(\u_inv.d_reg[89] ));
 sg13g2_nor3_1 _28386_ (.A(\u_inv.d_reg[91] ),
    .B(\u_inv.d_reg[90] ),
    .C(_05787_),
    .Y(_05788_));
 sg13g2_nand2_1 _28387_ (.Y(_05789_),
    .A(_05786_),
    .B(_05788_));
 sg13g2_inv_1 _28388_ (.Y(_05790_),
    .A(_05789_));
 sg13g2_or2_1 _28389_ (.X(_05791_),
    .B(\u_inv.d_reg[92] ),
    .A(\u_inv.d_reg[93] ));
 sg13g2_or2_1 _28390_ (.X(_05792_),
    .B(_05791_),
    .A(\u_inv.d_reg[94] ));
 sg13g2_nor3_1 _28391_ (.A(\u_inv.d_reg[95] ),
    .B(_05789_),
    .C(_05792_),
    .Y(_05793_));
 sg13g2_nand4_1 _28392_ (.B(_05764_),
    .C(_05766_),
    .A(net3493),
    .Y(_05794_),
    .D(_05793_));
 sg13g2_or3_1 _28393_ (.A(\u_inv.d_reg[106] ),
    .B(\u_inv.d_reg[105] ),
    .C(net4780),
    .X(_05795_));
 sg13g2_nor2_1 _28394_ (.A(\u_inv.d_reg[107] ),
    .B(_05795_),
    .Y(_05796_));
 sg13g2_nand2b_1 _28395_ (.Y(_05797_),
    .B(_05796_),
    .A_N(\u_inv.d_reg[108] ));
 sg13g2_nor2_1 _28396_ (.A(\u_inv.d_reg[109] ),
    .B(_05797_),
    .Y(_05798_));
 sg13g2_or2_1 _28397_ (.X(_05799_),
    .B(\u_inv.d_reg[100] ),
    .A(\u_inv.d_reg[101] ));
 sg13g2_or2_1 _28398_ (.X(_05800_),
    .B(_05799_),
    .A(\u_inv.d_reg[102] ));
 sg13g2_nor2_1 _28399_ (.A(\u_inv.d_reg[103] ),
    .B(_05800_),
    .Y(_05801_));
 sg13g2_or2_1 _28400_ (.X(_05802_),
    .B(\u_inv.d_reg[96] ),
    .A(\u_inv.d_reg[97] ));
 sg13g2_nor3_1 _28401_ (.A(\u_inv.d_reg[99] ),
    .B(\u_inv.d_reg[98] ),
    .C(_05802_),
    .Y(_05803_));
 sg13g2_nor2_1 _28402_ (.A(\u_inv.d_reg[111] ),
    .B(\u_inv.d_reg[110] ),
    .Y(_05804_));
 sg13g2_nand4_1 _28403_ (.B(_05801_),
    .C(_05803_),
    .A(_05798_),
    .Y(_05805_),
    .D(_05804_));
 sg13g2_or2_1 _28404_ (.X(_05806_),
    .B(_05805_),
    .A(net3492));
 sg13g2_or2_1 _28405_ (.X(_05807_),
    .B(\u_inv.d_reg[112] ),
    .A(\u_inv.d_reg[113] ));
 sg13g2_or2_1 _28406_ (.X(_05808_),
    .B(_05807_),
    .A(\u_inv.d_reg[114] ));
 sg13g2_or2_1 _28407_ (.X(_05809_),
    .B(\u_inv.d_reg[116] ),
    .A(\u_inv.d_reg[117] ));
 sg13g2_or2_1 _28408_ (.X(_05810_),
    .B(_05809_),
    .A(\u_inv.d_reg[118] ));
 sg13g2_or4_1 _28409_ (.A(\u_inv.d_reg[119] ),
    .B(\u_inv.d_reg[115] ),
    .C(_05808_),
    .D(_05810_),
    .X(_05811_));
 sg13g2_or3_1 _28410_ (.A(net3492),
    .B(_05805_),
    .C(_05811_),
    .X(_05812_));
 sg13g2_or4_1 _28411_ (.A(\u_inv.d_reg[127] ),
    .B(\u_inv.d_reg[126] ),
    .C(_05718_),
    .D(_05811_),
    .X(_05813_));
 sg13g2_nor3_2 _28412_ (.A(net3492),
    .B(_05805_),
    .C(_05813_),
    .Y(_05814_));
 sg13g2_or2_1 _28413_ (.X(_05815_),
    .B(\u_inv.d_reg[136] ),
    .A(\u_inv.d_reg[137] ));
 sg13g2_or3_1 _28414_ (.A(\u_inv.d_reg[139] ),
    .B(net4777),
    .C(_05815_),
    .X(_05816_));
 sg13g2_nor3_1 _28415_ (.A(\u_inv.d_reg[141] ),
    .B(\u_inv.d_reg[140] ),
    .C(_05816_),
    .Y(_05817_));
 sg13g2_inv_1 _28416_ (.Y(_05818_),
    .A(_05817_));
 sg13g2_nor2_1 _28417_ (.A(net4778),
    .B(net4779),
    .Y(_05819_));
 sg13g2_nor4_2 _28418_ (.A(\u_inv.d_reg[131] ),
    .B(\u_inv.d_reg[130] ),
    .C(net4779),
    .Y(_05820_),
    .D(\u_inv.d_reg[128] ));
 sg13g2_or2_1 _28419_ (.X(_05821_),
    .B(\u_inv.d_reg[132] ),
    .A(\u_inv.d_reg[133] ));
 sg13g2_or2_1 _28420_ (.X(_05822_),
    .B(_05821_),
    .A(\u_inv.d_reg[134] ));
 sg13g2_nor2_1 _28421_ (.A(\u_inv.d_reg[135] ),
    .B(_05822_),
    .Y(_05823_));
 sg13g2_nor2_1 _28422_ (.A(\u_inv.d_reg[143] ),
    .B(\u_inv.d_reg[142] ),
    .Y(_05824_));
 sg13g2_and4_1 _28423_ (.A(_05817_),
    .B(_05820_),
    .C(_05823_),
    .D(_05824_),
    .X(_05825_));
 sg13g2_nand2_2 _28424_ (.Y(_05826_),
    .A(net3489),
    .B(_05825_));
 sg13g2_nand4_1 _28425_ (.B(_05712_),
    .C(_05714_),
    .A(_05709_),
    .Y(_05827_),
    .D(_05825_));
 sg13g2_inv_2 _28426_ (.Y(_05828_),
    .A(_05827_));
 sg13g2_nand2_2 _28427_ (.Y(_05829_),
    .A(net3489),
    .B(_05828_));
 sg13g2_or2_1 _28428_ (.X(_05830_),
    .B(\u_inv.d_reg[160] ),
    .A(\u_inv.d_reg[161] ));
 sg13g2_nor2_1 _28429_ (.A(net4775),
    .B(_05830_),
    .Y(_05831_));
 sg13g2_inv_1 _28430_ (.Y(_05832_),
    .A(_05831_));
 sg13g2_or2_1 _28431_ (.X(_05833_),
    .B(\u_inv.d_reg[164] ),
    .A(\u_inv.d_reg[165] ));
 sg13g2_nor3_1 _28432_ (.A(\u_inv.d_reg[167] ),
    .B(\u_inv.d_reg[163] ),
    .C(_05833_),
    .Y(_05834_));
 sg13g2_nand3_1 _28433_ (.B(_05831_),
    .C(_05834_),
    .A(_10911_),
    .Y(_05835_));
 sg13g2_nand2_1 _28434_ (.Y(_05836_),
    .A(_10909_),
    .B(_10910_));
 sg13g2_or4_1 _28435_ (.A(\u_inv.d_reg[171] ),
    .B(\u_inv.d_reg[170] ),
    .C(_05835_),
    .D(_05836_),
    .X(_05837_));
 sg13g2_nand2_1 _28436_ (.Y(_05838_),
    .A(_10906_),
    .B(_10907_));
 sg13g2_or2_1 _28437_ (.X(_05839_),
    .B(_05838_),
    .A(\u_inv.d_reg[174] ));
 sg13g2_nor3_1 _28438_ (.A(\u_inv.d_reg[175] ),
    .B(_05837_),
    .C(_05839_),
    .Y(_05840_));
 sg13g2_nand3_1 _28439_ (.B(_05828_),
    .C(_05840_),
    .A(_05814_),
    .Y(_05841_));
 sg13g2_or2_1 _28440_ (.X(_05842_),
    .B(\u_inv.d_reg[184] ),
    .A(\u_inv.d_reg[185] ));
 sg13g2_or2_1 _28441_ (.X(_05843_),
    .B(_05842_),
    .A(\u_inv.d_reg[186] ));
 sg13g2_nor2_1 _28442_ (.A(net4774),
    .B(_05843_),
    .Y(_05844_));
 sg13g2_inv_1 _28443_ (.Y(_05845_),
    .A(_05844_));
 sg13g2_or4_1 _28444_ (.A(\u_inv.d_reg[190] ),
    .B(\u_inv.d_reg[189] ),
    .C(\u_inv.d_reg[188] ),
    .D(_05845_),
    .X(_05846_));
 sg13g2_or2_1 _28445_ (.X(_05847_),
    .B(\u_inv.d_reg[180] ),
    .A(\u_inv.d_reg[181] ));
 sg13g2_nand3b_1 _28446_ (.B(_10903_),
    .C(_10902_),
    .Y(_05848_),
    .A_N(_05847_));
 sg13g2_or2_1 _28447_ (.X(_05849_),
    .B(\u_inv.d_reg[176] ),
    .A(\u_inv.d_reg[177] ));
 sg13g2_or3_1 _28448_ (.A(\u_inv.d_reg[179] ),
    .B(\u_inv.d_reg[178] ),
    .C(_05849_),
    .X(_05850_));
 sg13g2_nor4_2 _28449_ (.A(\u_inv.d_reg[191] ),
    .B(_05846_),
    .C(_05848_),
    .Y(_05851_),
    .D(_05850_));
 sg13g2_nand2b_2 _28450_ (.Y(_05852_),
    .B(_05851_),
    .A_N(_05841_));
 sg13g2_or2_1 _28451_ (.X(_05853_),
    .B(\u_inv.d_reg[192] ),
    .A(\u_inv.d_reg[193] ));
 sg13g2_nand2b_1 _28452_ (.Y(_05854_),
    .B(_10898_),
    .A_N(_05853_));
 sg13g2_nor2_2 _28453_ (.A(\u_inv.d_reg[195] ),
    .B(_05854_),
    .Y(_05855_));
 sg13g2_nor4_2 _28454_ (.A(\u_inv.d_reg[199] ),
    .B(\u_inv.d_reg[198] ),
    .C(\u_inv.d_reg[197] ),
    .Y(_05856_),
    .D(\u_inv.d_reg[196] ));
 sg13g2_nor2_1 _28455_ (.A(\u_inv.d_reg[205] ),
    .B(\u_inv.d_reg[204] ),
    .Y(_05857_));
 sg13g2_nand2b_1 _28456_ (.Y(_05858_),
    .B(_05857_),
    .A_N(\u_inv.d_reg[206] ));
 sg13g2_nor4_1 _28457_ (.A(\u_inv.d_reg[203] ),
    .B(\u_inv.d_reg[202] ),
    .C(\u_inv.d_reg[201] ),
    .D(\u_inv.d_reg[200] ),
    .Y(_05859_));
 sg13g2_nand3_1 _28458_ (.B(_05856_),
    .C(_05859_),
    .A(_05855_),
    .Y(_05860_));
 sg13g2_nor3_1 _28459_ (.A(\u_inv.d_reg[207] ),
    .B(_05858_),
    .C(_05860_),
    .Y(_05861_));
 sg13g2_nand3b_1 _28460_ (.B(_05851_),
    .C(_05861_),
    .Y(_05862_),
    .A_N(_05841_));
 sg13g2_or4_1 _28461_ (.A(\u_inv.d_reg[211] ),
    .B(\u_inv.d_reg[210] ),
    .C(net4769),
    .D(net4770),
    .X(_05863_));
 sg13g2_or4_1 _28462_ (.A(\u_inv.d_reg[215] ),
    .B(\u_inv.d_reg[214] ),
    .C(\u_inv.d_reg[213] ),
    .D(\u_inv.d_reg[212] ),
    .X(_05864_));
 sg13g2_nor3_2 _28463_ (.A(_05862_),
    .B(_05863_),
    .C(_05864_),
    .Y(_05865_));
 sg13g2_or4_1 _28464_ (.A(\u_inv.d_reg[219] ),
    .B(\u_inv.d_reg[218] ),
    .C(\u_inv.d_reg[217] ),
    .D(\u_inv.d_reg[216] ),
    .X(_05866_));
 sg13g2_nor3_1 _28465_ (.A(\u_inv.d_reg[221] ),
    .B(\u_inv.d_reg[220] ),
    .C(_05866_),
    .Y(_05867_));
 sg13g2_nand4_1 _28466_ (.B(_10889_),
    .C(_05865_),
    .A(_10888_),
    .Y(_05868_),
    .D(_05867_));
 sg13g2_nor4_1 _28467_ (.A(\u_inv.d_reg[235] ),
    .B(\u_inv.d_reg[234] ),
    .C(\u_inv.d_reg[233] ),
    .D(\u_inv.d_reg[232] ),
    .Y(_05869_));
 sg13g2_nor3_1 _28468_ (.A(\u_inv.d_reg[238] ),
    .B(\u_inv.d_reg[237] ),
    .C(\u_inv.d_reg[236] ),
    .Y(_05870_));
 sg13g2_nand2_1 _28469_ (.Y(_05871_),
    .A(_05869_),
    .B(_05870_));
 sg13g2_or2_1 _28470_ (.X(_05872_),
    .B(\u_inv.d_reg[224] ),
    .A(\u_inv.d_reg[225] ));
 sg13g2_nor3_1 _28471_ (.A(\u_inv.d_reg[227] ),
    .B(\u_inv.d_reg[226] ),
    .C(_05872_),
    .Y(_05873_));
 sg13g2_inv_1 _28472_ (.Y(_05874_),
    .A(_05873_));
 sg13g2_nor4_1 _28473_ (.A(\u_inv.d_reg[231] ),
    .B(\u_inv.d_reg[230] ),
    .C(net4766),
    .D(\u_inv.d_reg[228] ),
    .Y(_05875_));
 sg13g2_nand2_2 _28474_ (.Y(_05876_),
    .A(_05873_),
    .B(_05875_));
 sg13g2_or4_1 _28475_ (.A(\u_inv.d_reg[239] ),
    .B(_05868_),
    .C(_05871_),
    .D(_05876_),
    .X(_05877_));
 sg13g2_or2_1 _28476_ (.X(_05878_),
    .B(\u_inv.d_reg[240] ),
    .A(\u_inv.d_reg[241] ));
 sg13g2_or3_1 _28477_ (.A(\u_inv.d_reg[243] ),
    .B(\u_inv.d_reg[242] ),
    .C(_05878_),
    .X(_05879_));
 sg13g2_or3_1 _28478_ (.A(\u_inv.d_reg[245] ),
    .B(\u_inv.d_reg[244] ),
    .C(_05879_),
    .X(_05880_));
 sg13g2_nor4_1 _28479_ (.A(\u_inv.d_reg[247] ),
    .B(\u_inv.d_reg[246] ),
    .C(_05877_),
    .D(_05880_),
    .Y(_05881_));
 sg13g2_nor4_1 _28480_ (.A(\u_inv.d_reg[251] ),
    .B(\u_inv.d_reg[250] ),
    .C(\u_inv.d_reg[249] ),
    .D(\u_inv.d_reg[248] ),
    .Y(_05882_));
 sg13g2_nor2_1 _28481_ (.A(net4501),
    .B(_05881_),
    .Y(_05883_));
 sg13g2_a21o_2 _28482_ (.A2(_05882_),
    .A1(_05881_),
    .B1(net4501),
    .X(_05884_));
 sg13g2_o21ai_1 _28483_ (.B1(net4727),
    .Y(_05885_),
    .A1(\u_inv.d_reg[253] ),
    .A2(\u_inv.d_reg[252] ));
 sg13g2_nand2_1 _28484_ (.Y(_05886_),
    .A(_05884_),
    .B(_05885_));
 sg13g2_o21ai_1 _28485_ (.B1(net4727),
    .Y(_05887_),
    .A1(\u_inv.d_reg[255] ),
    .A2(\u_inv.d_reg[254] ));
 sg13g2_nand3_1 _28486_ (.B(_05885_),
    .C(_05887_),
    .A(_05884_),
    .Y(_05888_));
 sg13g2_xnor2_1 _28487_ (.Y(_05889_),
    .A(\u_inv.d_reg[256] ),
    .B(_05888_));
 sg13g2_xor2_1 _28488_ (.B(_05888_),
    .A(\u_inv.d_reg[256] ),
    .X(_05890_));
 sg13g2_nand2b_1 _28489_ (.Y(_05891_),
    .B(_05881_),
    .A_N(\u_inv.d_reg[248] ));
 sg13g2_or3_1 _28490_ (.A(\u_inv.d_reg[250] ),
    .B(\u_inv.d_reg[249] ),
    .C(_05891_),
    .X(_05892_));
 sg13g2_a21oi_1 _28491_ (.A1(\u_inv.d_reg[251] ),
    .A2(_05892_),
    .Y(_05893_),
    .B1(_05884_));
 sg13g2_a21o_2 _28492_ (.A2(\u_inv.d_reg[251] ),
    .A1(net4501),
    .B1(_05893_),
    .X(_05894_));
 sg13g2_nand2_1 _28493_ (.Y(_05895_),
    .A(net4733),
    .B(_05868_));
 sg13g2_o21ai_1 _28494_ (.B1(net4733),
    .Y(_05896_),
    .A1(_05868_),
    .A2(_05874_));
 sg13g2_o21ai_1 _28495_ (.B1(net4733),
    .Y(_05897_),
    .A1(\u_inv.d_reg[229] ),
    .A2(net4767));
 sg13g2_and2_1 _28496_ (.A(_05896_),
    .B(_05897_),
    .X(_05898_));
 sg13g2_inv_1 _28497_ (.Y(_05899_),
    .A(_05898_));
 sg13g2_a21oi_1 _28498_ (.A1(net4733),
    .A2(\u_inv.d_reg[230] ),
    .Y(_05900_),
    .B1(_05899_));
 sg13g2_xnor2_1 _28499_ (.Y(_05901_),
    .A(\u_inv.d_reg[231] ),
    .B(_05900_));
 sg13g2_and2_1 _28500_ (.A(net4731),
    .B(_05877_),
    .X(_05902_));
 sg13g2_o21ai_1 _28501_ (.B1(net4731),
    .Y(_05903_),
    .A1(_05877_),
    .A2(_05880_));
 sg13g2_inv_1 _28502_ (.Y(_05904_),
    .A(_05903_));
 sg13g2_a21oi_1 _28503_ (.A1(net4731),
    .A2(\u_inv.d_reg[246] ),
    .Y(_05905_),
    .B1(_05904_));
 sg13g2_xnor2_1 _28504_ (.Y(_05906_),
    .A(\u_inv.d_reg[247] ),
    .B(_05905_));
 sg13g2_o21ai_1 _28505_ (.B1(net4729),
    .Y(_05907_),
    .A1(_05868_),
    .A2(_05876_));
 sg13g2_o21ai_1 _28506_ (.B1(_05907_),
    .Y(_05908_),
    .A1(net4503),
    .A2(_10887_));
 sg13g2_xnor2_1 _28507_ (.Y(_05909_),
    .A(\u_inv.d_reg[233] ),
    .B(_05908_));
 sg13g2_inv_1 _28508_ (.Y(_05910_),
    .A(_05909_));
 sg13g2_xnor2_1 _28509_ (.Y(_05911_),
    .A(_10887_),
    .B(_05907_));
 sg13g2_or2_1 _28510_ (.X(_05912_),
    .B(_05911_),
    .A(_05909_));
 sg13g2_nor2b_1 _28511_ (.A(_05912_),
    .B_N(_05906_),
    .Y(_05913_));
 sg13g2_nand4_1 _28512_ (.B(_05894_),
    .C(_05901_),
    .A(net3378),
    .Y(_05914_),
    .D(_05913_));
 sg13g2_o21ai_1 _28513_ (.B1(net4738),
    .Y(_05915_),
    .A1(net4770),
    .A2(_05862_));
 sg13g2_xnor2_1 _28514_ (.Y(_05916_),
    .A(net4769),
    .B(_05915_));
 sg13g2_xor2_1 _28515_ (.B(_05915_),
    .A(\u_inv.d_reg[209] ),
    .X(_05917_));
 sg13g2_nand3b_1 _28516_ (.B(_05855_),
    .C(_05856_),
    .Y(_05918_),
    .A_N(_05852_));
 sg13g2_o21ai_1 _28517_ (.B1(net4740),
    .Y(_05919_),
    .A1(\u_inv.d_reg[200] ),
    .A2(_05918_));
 sg13g2_xnor2_1 _28518_ (.Y(_05920_),
    .A(_10896_),
    .B(_05919_));
 sg13g2_nor2_1 _28519_ (.A(_05852_),
    .B(_05860_),
    .Y(_05921_));
 sg13g2_nor2_2 _28520_ (.A(net4506),
    .B(_05921_),
    .Y(_05922_));
 sg13g2_xnor2_1 _28521_ (.Y(_05923_),
    .A(\u_inv.d_reg[204] ),
    .B(_05922_));
 sg13g2_or2_1 _28522_ (.X(_05924_),
    .B(_05850_),
    .A(_05841_));
 sg13g2_and2_1 _28523_ (.A(net4754),
    .B(_05924_),
    .X(_05925_));
 sg13g2_o21ai_1 _28524_ (.B1(net4754),
    .Y(_05926_),
    .A1(\u_inv.d_reg[180] ),
    .A2(_05924_));
 sg13g2_xnor2_1 _28525_ (.Y(_05927_),
    .A(\u_inv.d_reg[181] ),
    .B(_05926_));
 sg13g2_xor2_1 _28526_ (.B(_05925_),
    .A(\u_inv.d_reg[180] ),
    .X(_05928_));
 sg13g2_nand2_2 _28527_ (.Y(_05929_),
    .A(_05927_),
    .B(_05928_));
 sg13g2_nor4_1 _28528_ (.A(_05917_),
    .B(_05920_),
    .C(_05923_),
    .D(_05929_),
    .Y(_05930_));
 sg13g2_or2_1 _28529_ (.X(_05931_),
    .B(_05924_),
    .A(_05848_));
 sg13g2_nand2_1 _28530_ (.Y(_05932_),
    .A(net4750),
    .B(_05931_));
 sg13g2_o21ai_1 _28531_ (.B1(net4750),
    .Y(_05933_),
    .A1(\u_inv.d_reg[184] ),
    .A2(_05931_));
 sg13g2_xnor2_1 _28532_ (.Y(_05934_),
    .A(\u_inv.d_reg[185] ),
    .B(_05933_));
 sg13g2_nand4_1 _28533_ (.B(_05814_),
    .C(_05828_),
    .A(_10912_),
    .Y(_05935_),
    .D(_05831_));
 sg13g2_o21ai_1 _28534_ (.B1(net4762),
    .Y(_05936_),
    .A1(_05829_),
    .A2(_05832_));
 sg13g2_nand2_1 _28535_ (.Y(_05937_),
    .A(net4762),
    .B(_05935_));
 sg13g2_o21ai_1 _28536_ (.B1(net4758),
    .Y(_05938_),
    .A1(\u_inv.d_reg[164] ),
    .A2(_05935_));
 sg13g2_xor2_1 _28537_ (.B(_05938_),
    .A(\u_inv.d_reg[165] ),
    .X(_05939_));
 sg13g2_xor2_1 _28538_ (.B(_05937_),
    .A(\u_inv.d_reg[164] ),
    .X(_05940_));
 sg13g2_nor2_2 _28539_ (.A(_05939_),
    .B(_05940_),
    .Y(_05941_));
 sg13g2_nand2b_1 _28540_ (.Y(_05942_),
    .B(net4737),
    .A_N(_05865_));
 sg13g2_xnor2_1 _28541_ (.Y(_05943_),
    .A(_10892_),
    .B(_05942_));
 sg13g2_inv_4 _28542_ (.A(_05943_),
    .Y(_05944_));
 sg13g2_o21ai_1 _28543_ (.B1(net4750),
    .Y(_05945_),
    .A1(_05843_),
    .A2(_05931_));
 sg13g2_o21ai_1 _28544_ (.B1(net4755),
    .Y(_05946_),
    .A1(_05845_),
    .A2(_05931_));
 sg13g2_xnor2_1 _28545_ (.Y(_05947_),
    .A(net4774),
    .B(_05945_));
 sg13g2_xor2_1 _28546_ (.B(_05945_),
    .A(net4774),
    .X(_05948_));
 sg13g2_and4_1 _28547_ (.A(_05934_),
    .B(_05941_),
    .C(_05944_),
    .D(_05947_),
    .X(_05949_));
 sg13g2_a21oi_1 _28548_ (.A1(_10900_),
    .A2(_05946_),
    .Y(_05950_),
    .B1(net4508));
 sg13g2_xor2_1 _28549_ (.B(_05950_),
    .A(\u_inv.d_reg[189] ),
    .X(_05951_));
 sg13g2_xnor2_1 _28550_ (.Y(_05952_),
    .A(\u_inv.d_reg[224] ),
    .B(_05895_));
 sg13g2_nand4_1 _28551_ (.B(_05949_),
    .C(_05951_),
    .A(_05930_),
    .Y(_05953_),
    .D(_05952_));
 sg13g2_nand2_2 _28552_ (.Y(_05954_),
    .A(net3489),
    .B(_05820_));
 sg13g2_nand3_1 _28553_ (.B(_05820_),
    .C(_05823_),
    .A(net3489),
    .Y(_05955_));
 sg13g2_nand2_1 _28554_ (.Y(_05956_),
    .A(net4757),
    .B(_05955_));
 sg13g2_o21ai_1 _28555_ (.B1(net4756),
    .Y(_05957_),
    .A1(_05815_),
    .A2(_05955_));
 sg13g2_xnor2_1 _28556_ (.Y(_05958_),
    .A(net4777),
    .B(_05957_));
 sg13g2_inv_1 _28557_ (.Y(_05959_),
    .A(_05958_));
 sg13g2_or2_1 _28558_ (.X(_05960_),
    .B(_05835_),
    .A(_05829_));
 sg13g2_nand2_1 _28559_ (.Y(_05961_),
    .A(net4762),
    .B(_05960_));
 sg13g2_xnor2_1 _28560_ (.Y(_05962_),
    .A(_10910_),
    .B(_05961_));
 sg13g2_nand2_1 _28561_ (.Y(_05963_),
    .A(net4764),
    .B(_05841_));
 sg13g2_xor2_1 _28562_ (.B(_05963_),
    .A(\u_inv.d_reg[176] ),
    .X(_05964_));
 sg13g2_nand2_1 _28563_ (.Y(_05965_),
    .A(net4757),
    .B(\u_inv.d_reg[138] ));
 sg13g2_and2_1 _28564_ (.A(_05957_),
    .B(_05965_),
    .X(_05966_));
 sg13g2_xor2_1 _28565_ (.B(_05966_),
    .A(\u_inv.d_reg[139] ),
    .X(_05967_));
 sg13g2_nor4_1 _28566_ (.A(_05959_),
    .B(_05962_),
    .C(_05964_),
    .D(_05967_),
    .Y(_05968_));
 sg13g2_o21ai_1 _28567_ (.B1(net4756),
    .Y(_05969_),
    .A1(_05816_),
    .A2(_05955_));
 sg13g2_xor2_1 _28568_ (.B(_05969_),
    .A(\u_inv.d_reg[140] ),
    .X(_05970_));
 sg13g2_o21ai_1 _28569_ (.B1(net4756),
    .Y(_05971_),
    .A1(_05818_),
    .A2(_05955_));
 sg13g2_xnor2_1 _28570_ (.Y(_05972_),
    .A(_10917_),
    .B(_05971_));
 sg13g2_nand3_1 _28571_ (.B(net3489),
    .C(_05825_),
    .A(_05709_),
    .Y(_05973_));
 sg13g2_nand2_1 _28572_ (.Y(_05974_),
    .A(net4759),
    .B(_05826_));
 sg13g2_nand2_1 _28573_ (.Y(_05975_),
    .A(net4759),
    .B(_05973_));
 sg13g2_o21ai_1 _28574_ (.B1(net4759),
    .Y(_05976_),
    .A1(_05711_),
    .A2(_05973_));
 sg13g2_nand4_1 _28575_ (.B(_05713_),
    .C(net3489),
    .A(_05709_),
    .Y(_05977_),
    .D(_05825_));
 sg13g2_nand2_1 _28576_ (.Y(_05978_),
    .A(net4759),
    .B(_05977_));
 sg13g2_nor2_1 _28577_ (.A(net4508),
    .B(_05712_),
    .Y(_05979_));
 sg13g2_a21oi_1 _28578_ (.A1(net4761),
    .A2(_05977_),
    .Y(_05980_),
    .B1(_05979_));
 sg13g2_xnor2_1 _28579_ (.Y(_05981_),
    .A(_10913_),
    .B(_05980_));
 sg13g2_xor2_1 _28580_ (.B(_05978_),
    .A(\u_inv.d_reg[152] ),
    .X(_05982_));
 sg13g2_nor4_1 _28581_ (.A(_05970_),
    .B(_05972_),
    .C(_05981_),
    .D(_05982_),
    .Y(_05983_));
 sg13g2_o21ai_1 _28582_ (.B1(net4754),
    .Y(_05984_),
    .A1(_05847_),
    .A2(_05924_));
 sg13g2_xnor2_1 _28583_ (.Y(_05985_),
    .A(_10903_),
    .B(_05984_));
 sg13g2_nand2_1 _28584_ (.Y(_05986_),
    .A(net4756),
    .B(\u_inv.d_reg[140] ));
 sg13g2_and2_1 _28585_ (.A(_05969_),
    .B(_05986_),
    .X(_05987_));
 sg13g2_xor2_1 _28586_ (.B(_05987_),
    .A(\u_inv.d_reg[141] ),
    .X(_05988_));
 sg13g2_nand2_1 _28587_ (.Y(_05989_),
    .A(net4758),
    .B(_05829_));
 sg13g2_o21ai_1 _28588_ (.B1(net4758),
    .Y(_05990_),
    .A1(\u_inv.d_reg[160] ),
    .A2(_05829_));
 sg13g2_xor2_1 _28589_ (.B(_05990_),
    .A(\u_inv.d_reg[161] ),
    .X(_05991_));
 sg13g2_o21ai_1 _28590_ (.B1(net4756),
    .Y(_05992_),
    .A1(\u_inv.d_reg[136] ),
    .A2(_05955_));
 sg13g2_xnor2_1 _28591_ (.Y(_05993_),
    .A(\u_inv.d_reg[137] ),
    .B(_05992_));
 sg13g2_o21ai_1 _28592_ (.B1(net4759),
    .Y(_05994_),
    .A1(_05710_),
    .A2(_05973_));
 sg13g2_xor2_1 _28593_ (.B(_05994_),
    .A(net4776),
    .X(_05995_));
 sg13g2_xnor2_1 _28594_ (.Y(_05996_),
    .A(net4776),
    .B(_05994_));
 sg13g2_nand2_1 _28595_ (.Y(_05997_),
    .A(_05993_),
    .B(_05996_));
 sg13g2_nor4_1 _28596_ (.A(_05985_),
    .B(_05988_),
    .C(_05991_),
    .D(_05997_),
    .Y(_05998_));
 sg13g2_nand3_1 _28597_ (.B(_05983_),
    .C(_05998_),
    .A(_05968_),
    .Y(_05999_));
 sg13g2_o21ai_1 _28598_ (.B1(net4761),
    .Y(_06000_),
    .A1(_05703_),
    .A2(_05977_));
 sg13g2_xnor2_1 _28599_ (.Y(_06001_),
    .A(\u_inv.d_reg[156] ),
    .B(_06000_));
 sg13g2_o21ai_1 _28600_ (.B1(net4758),
    .Y(_06002_),
    .A1(_05829_),
    .A2(_05830_));
 sg13g2_xor2_1 _28601_ (.B(_06002_),
    .A(\u_inv.d_reg[162] ),
    .X(_06003_));
 sg13g2_xnor2_1 _28602_ (.Y(_06004_),
    .A(_10912_),
    .B(_05936_));
 sg13g2_or2_1 _28603_ (.X(_06005_),
    .B(_06004_),
    .A(_06003_));
 sg13g2_inv_1 _28604_ (.Y(_06006_),
    .A(_06005_));
 sg13g2_o21ai_1 _28605_ (.B1(net4754),
    .Y(_06007_),
    .A1(_05841_),
    .A2(_05849_));
 sg13g2_xnor2_1 _28606_ (.Y(_06008_),
    .A(\u_inv.d_reg[178] ),
    .B(_06007_));
 sg13g2_o21ai_1 _28607_ (.B1(net4760),
    .Y(_06009_),
    .A1(\u_inv.d_reg[152] ),
    .A2(_05977_));
 sg13g2_xnor2_1 _28608_ (.Y(_06010_),
    .A(\u_inv.d_reg[153] ),
    .B(_06009_));
 sg13g2_nand4_1 _28609_ (.B(_06006_),
    .C(_06008_),
    .A(_06001_),
    .Y(_06011_),
    .D(_06010_));
 sg13g2_o21ai_1 _28610_ (.B1(net4751),
    .Y(_06012_),
    .A1(_05718_),
    .A2(_05812_));
 sg13g2_nand2_1 _28611_ (.Y(_06013_),
    .A(net4751),
    .B(\u_inv.d_reg[126] ));
 sg13g2_and2_1 _28612_ (.A(_06012_),
    .B(_06013_),
    .X(_06014_));
 sg13g2_xnor2_1 _28613_ (.Y(_06015_),
    .A(\u_inv.d_reg[127] ),
    .B(_06014_));
 sg13g2_nor2_1 _28614_ (.A(net4508),
    .B(net3489),
    .Y(_06016_));
 sg13g2_xnor2_1 _28615_ (.Y(_06017_),
    .A(\u_inv.d_reg[128] ),
    .B(_06016_));
 sg13g2_nand2b_1 _28616_ (.Y(_06018_),
    .B(_06015_),
    .A_N(_06017_));
 sg13g2_nand2_1 _28617_ (.Y(_06019_),
    .A(net4751),
    .B(_05812_));
 sg13g2_xor2_1 _28618_ (.B(_06019_),
    .A(\u_inv.d_reg[120] ),
    .X(_06020_));
 sg13g2_o21ai_1 _28619_ (.B1(net4751),
    .Y(_06021_),
    .A1(\u_inv.d_reg[120] ),
    .A2(_05812_));
 sg13g2_xor2_1 _28620_ (.B(_06021_),
    .A(\u_inv.d_reg[121] ),
    .X(_06022_));
 sg13g2_inv_1 _28621_ (.Y(_06023_),
    .A(_06022_));
 sg13g2_nor2_1 _28622_ (.A(_06020_),
    .B(_06022_),
    .Y(_06024_));
 sg13g2_inv_1 _28623_ (.Y(_06025_),
    .A(_06024_));
 sg13g2_nand2_1 _28624_ (.Y(_06026_),
    .A(net4753),
    .B(_05806_));
 sg13g2_or4_1 _28625_ (.A(\u_inv.d_reg[115] ),
    .B(_05794_),
    .C(_05805_),
    .D(_05808_),
    .X(_06027_));
 sg13g2_nand2_1 _28626_ (.Y(_06028_),
    .A(net4751),
    .B(_06027_));
 sg13g2_o21ai_1 _28627_ (.B1(net4751),
    .Y(_06029_),
    .A1(\u_inv.d_reg[116] ),
    .A2(_06027_));
 sg13g2_xor2_1 _28628_ (.B(_06029_),
    .A(\u_inv.d_reg[117] ),
    .X(_06030_));
 sg13g2_xnor2_1 _28629_ (.Y(_06031_),
    .A(\u_inv.d_reg[117] ),
    .B(_06029_));
 sg13g2_xor2_1 _28630_ (.B(_06028_),
    .A(\u_inv.d_reg[116] ),
    .X(_06032_));
 sg13g2_nand2b_1 _28631_ (.Y(_06033_),
    .B(_06031_),
    .A_N(_06032_));
 sg13g2_nand4_1 _28632_ (.B(_05764_),
    .C(_05766_),
    .A(net3493),
    .Y(_06034_),
    .D(_05770_));
 sg13g2_nand2_1 _28633_ (.Y(_06035_),
    .A(net4743),
    .B(_06034_));
 sg13g2_xor2_1 _28634_ (.B(_06035_),
    .A(\u_inv.d_reg[68] ),
    .X(_06036_));
 sg13g2_nand4_1 _28635_ (.B(_05764_),
    .C(_05766_),
    .A(net3493),
    .Y(_06037_),
    .D(_05779_));
 sg13g2_nand2_1 _28636_ (.Y(_06038_),
    .A(net4745),
    .B(_06037_));
 sg13g2_xor2_1 _28637_ (.B(_06038_),
    .A(\u_inv.d_reg[80] ),
    .X(_06039_));
 sg13g2_nand4_1 _28638_ (.B(_05764_),
    .C(_05766_),
    .A(net3493),
    .Y(_06040_),
    .D(_05773_));
 sg13g2_nand2_1 _28639_ (.Y(_06041_),
    .A(net4747),
    .B(_06040_));
 sg13g2_xnor2_1 _28640_ (.Y(_06042_),
    .A(net4783),
    .B(_06041_));
 sg13g2_xor2_1 _28641_ (.B(_06041_),
    .A(net4783),
    .X(_06043_));
 sg13g2_nand2_1 _28642_ (.Y(_06044_),
    .A(net4740),
    .B(_05765_));
 sg13g2_xor2_1 _28643_ (.B(_06044_),
    .A(\u_inv.d_reg[60] ),
    .X(_06045_));
 sg13g2_o21ai_1 _28644_ (.B1(net4741),
    .Y(_06046_),
    .A1(\u_inv.d_reg[60] ),
    .A2(_05765_));
 sg13g2_xnor2_1 _28645_ (.Y(_06047_),
    .A(_10934_),
    .B(_06046_));
 sg13g2_or2_1 _28646_ (.X(_06048_),
    .B(_06047_),
    .A(_06045_));
 sg13g2_nor4_1 _28647_ (.A(_06036_),
    .B(_06039_),
    .C(_06043_),
    .D(_06048_),
    .Y(_06049_));
 sg13g2_o21ai_1 _28648_ (.B1(net4747),
    .Y(_06050_),
    .A1(_05774_),
    .A2(_06040_));
 sg13g2_o21ai_1 _28649_ (.B1(net4747),
    .Y(_06051_),
    .A1(_05775_),
    .A2(_06040_));
 sg13g2_xnor2_1 _28650_ (.Y(_06052_),
    .A(\u_inv.d_reg[75] ),
    .B(_06051_));
 sg13g2_nand2b_1 _28651_ (.Y(_06053_),
    .B(net3493),
    .A_N(\u_inv.d_reg[56] ));
 sg13g2_nand2_1 _28652_ (.Y(_06054_),
    .A(net4741),
    .B(_06053_));
 sg13g2_xnor2_1 _28653_ (.Y(_06055_),
    .A(_10936_),
    .B(_06054_));
 sg13g2_nand2_1 _28654_ (.Y(_06056_),
    .A(net4741),
    .B(_05761_));
 sg13g2_xor2_1 _28655_ (.B(_06056_),
    .A(\u_inv.d_reg[54] ),
    .X(_06057_));
 sg13g2_o21ai_1 _28656_ (.B1(net4735),
    .Y(_06058_),
    .A1(_05753_),
    .A2(_05754_));
 sg13g2_a21oi_1 _28657_ (.A1(_10943_),
    .A2(_06058_),
    .Y(_06059_),
    .B1(net4504));
 sg13g2_xnor2_1 _28658_ (.Y(_06060_),
    .A(\u_inv.d_reg[47] ),
    .B(_06059_));
 sg13g2_nand2_1 _28659_ (.Y(_06061_),
    .A(net4737),
    .B(_05756_));
 sg13g2_xor2_1 _28660_ (.B(_06061_),
    .A(\u_inv.d_reg[48] ),
    .X(_06062_));
 sg13g2_nand2_1 _28661_ (.Y(_06063_),
    .A(net4734),
    .B(_05750_));
 sg13g2_o21ai_1 _28662_ (.B1(net4735),
    .Y(_06064_),
    .A1(\u_inv.d_reg[40] ),
    .A2(_05750_));
 sg13g2_xnor2_1 _28663_ (.Y(_06065_),
    .A(\u_inv.d_reg[41] ),
    .B(_06064_));
 sg13g2_xnor2_1 _28664_ (.Y(_06066_),
    .A(\u_inv.d_reg[40] ),
    .B(_06063_));
 sg13g2_nand2_1 _28665_ (.Y(_06067_),
    .A(_06065_),
    .B(_06066_));
 sg13g2_xnor2_1 _28666_ (.Y(_06068_),
    .A(_10943_),
    .B(_06058_));
 sg13g2_or4_1 _28667_ (.A(_06060_),
    .B(_06062_),
    .C(_06067_),
    .D(_06068_),
    .X(_06069_));
 sg13g2_o21ai_1 _28668_ (.B1(net4737),
    .Y(_06070_),
    .A1(_05756_),
    .A2(_05757_));
 sg13g2_o21ai_1 _28669_ (.B1(_06070_),
    .Y(_06071_),
    .A1(net4504),
    .A2(_10940_));
 sg13g2_xnor2_1 _28670_ (.Y(_06072_),
    .A(_10939_),
    .B(_06071_));
 sg13g2_xnor2_1 _28671_ (.Y(_06073_),
    .A(\u_inv.d_reg[50] ),
    .B(_06070_));
 sg13g2_nand2_2 _28672_ (.Y(_06074_),
    .A(_06072_),
    .B(_06073_));
 sg13g2_or3_1 _28673_ (.A(\u_inv.d_reg[37] ),
    .B(_05745_),
    .C(_05748_),
    .X(_06075_));
 sg13g2_nand2_1 _28674_ (.Y(_06076_),
    .A(net4734),
    .B(_06075_));
 sg13g2_o21ai_1 _28675_ (.B1(net4734),
    .Y(_06077_),
    .A1(\u_inv.d_reg[38] ),
    .A2(_06075_));
 sg13g2_xor2_1 _28676_ (.B(_06077_),
    .A(\u_inv.d_reg[39] ),
    .X(_06078_));
 sg13g2_o21ai_1 _28677_ (.B1(net4735),
    .Y(_06079_),
    .A1(_05750_),
    .A2(_05751_));
 sg13g2_inv_1 _28678_ (.Y(_06080_),
    .A(_06079_));
 sg13g2_xor2_1 _28679_ (.B(_06079_),
    .A(net4786),
    .X(_06081_));
 sg13g2_nor2_1 _28680_ (.A(_06078_),
    .B(_06081_),
    .Y(_06082_));
 sg13g2_nor2_1 _28681_ (.A(net4505),
    .B(_05744_),
    .Y(_06083_));
 sg13g2_o21ai_1 _28682_ (.B1(net4734),
    .Y(_06084_),
    .A1(_05745_),
    .A2(_05746_));
 sg13g2_xnor2_1 _28683_ (.Y(_06085_),
    .A(_10945_),
    .B(_06084_));
 sg13g2_o21ai_1 _28684_ (.B1(_06084_),
    .Y(_06086_),
    .A1(net4505),
    .A2(_10945_));
 sg13g2_xnor2_1 _28685_ (.Y(_06087_),
    .A(\u_inv.d_reg[35] ),
    .B(_06086_));
 sg13g2_nor2_1 _28686_ (.A(_06085_),
    .B(_06087_),
    .Y(_06088_));
 sg13g2_o21ai_1 _28687_ (.B1(net4734),
    .Y(_06089_),
    .A1(_05745_),
    .A2(_05748_));
 sg13g2_xnor2_1 _28688_ (.Y(_06090_),
    .A(\u_inv.d_reg[37] ),
    .B(_06089_));
 sg13g2_o21ai_1 _28689_ (.B1(net4734),
    .Y(_06091_),
    .A1(_05745_),
    .A2(_05747_));
 sg13g2_xnor2_1 _28690_ (.Y(_06092_),
    .A(\u_inv.d_reg[36] ),
    .B(_06091_));
 sg13g2_nand4_1 _28691_ (.B(_06088_),
    .C(_06090_),
    .A(_06082_),
    .Y(_06093_),
    .D(_06092_));
 sg13g2_a21oi_1 _28692_ (.A1(net4734),
    .A2(\u_inv.d_reg[42] ),
    .Y(_06094_),
    .B1(_06080_));
 sg13g2_xor2_1 _28693_ (.B(_06094_),
    .A(\u_inv.d_reg[43] ),
    .X(_06095_));
 sg13g2_xnor2_1 _28694_ (.Y(_06096_),
    .A(\u_inv.d_reg[32] ),
    .B(_06083_));
 sg13g2_nor2_1 _28695_ (.A(net4505),
    .B(_05741_),
    .Y(_06097_));
 sg13g2_xnor2_1 _28696_ (.Y(_06098_),
    .A(\u_inv.d_reg[28] ),
    .B(_06097_));
 sg13g2_a21oi_1 _28697_ (.A1(net4736),
    .A2(\u_inv.d_reg[28] ),
    .Y(_06099_),
    .B1(_06097_));
 sg13g2_xnor2_1 _28698_ (.Y(_06100_),
    .A(\u_inv.d_reg[29] ),
    .B(_06099_));
 sg13g2_nor2b_1 _28699_ (.A(_06098_),
    .B_N(_06100_),
    .Y(_06101_));
 sg13g2_o21ai_1 _28700_ (.B1(net4733),
    .Y(_06102_),
    .A1(\u_inv.d_reg[30] ),
    .A2(_05743_));
 sg13g2_xnor2_1 _28701_ (.Y(_06103_),
    .A(_10946_),
    .B(_06102_));
 sg13g2_inv_1 _28702_ (.Y(_06104_),
    .A(_06103_));
 sg13g2_nand2_1 _28703_ (.Y(_06105_),
    .A(net4736),
    .B(_05743_));
 sg13g2_xnor2_1 _28704_ (.Y(_06106_),
    .A(_10947_),
    .B(_06105_));
 sg13g2_inv_1 _28705_ (.Y(_06107_),
    .A(_06106_));
 sg13g2_nor2_1 _28706_ (.A(net4503),
    .B(_05740_),
    .Y(_06108_));
 sg13g2_xnor2_1 _28707_ (.Y(_06109_),
    .A(\u_inv.d_reg[27] ),
    .B(_06108_));
 sg13g2_o21ai_1 _28708_ (.B1(net4729),
    .Y(_06110_),
    .A1(net4788),
    .A2(_05739_));
 sg13g2_xor2_1 _28709_ (.B(_06110_),
    .A(net4787),
    .X(_06111_));
 sg13g2_nand2_1 _28710_ (.Y(_06112_),
    .A(net4729),
    .B(_05739_));
 sg13g2_xor2_1 _28711_ (.B(_06112_),
    .A(\u_inv.d_reg[25] ),
    .X(_06113_));
 sg13g2_nand2_1 _28712_ (.Y(_06114_),
    .A(net4729),
    .B(_05738_));
 sg13g2_xnor2_1 _28713_ (.Y(_06115_),
    .A(_10949_),
    .B(_06114_));
 sg13g2_nor2_1 _28714_ (.A(_06113_),
    .B(_06115_),
    .Y(_06116_));
 sg13g2_nand2_1 _28715_ (.Y(_06117_),
    .A(net4730),
    .B(_05736_));
 sg13g2_o21ai_1 _28716_ (.B1(net4730),
    .Y(_06118_),
    .A1(net4789),
    .A2(_05736_));
 sg13g2_xor2_1 _28717_ (.B(_06118_),
    .A(\u_inv.d_reg[23] ),
    .X(_06119_));
 sg13g2_xor2_1 _28718_ (.B(_06117_),
    .A(net4789),
    .X(_06120_));
 sg13g2_or2_1 _28719_ (.X(_06121_),
    .B(_06120_),
    .A(_06119_));
 sg13g2_nand2_1 _28720_ (.Y(_06122_),
    .A(net4730),
    .B(_05734_));
 sg13g2_o21ai_1 _28721_ (.B1(net4730),
    .Y(_06123_),
    .A1(\u_inv.d_reg[20] ),
    .A2(_05734_));
 sg13g2_xnor2_1 _28722_ (.Y(_06124_),
    .A(\u_inv.d_reg[21] ),
    .B(_06123_));
 sg13g2_xor2_1 _28723_ (.B(_06122_),
    .A(\u_inv.d_reg[20] ),
    .X(_06125_));
 sg13g2_inv_1 _28724_ (.Y(_06126_),
    .A(_06125_));
 sg13g2_nand2_1 _28725_ (.Y(_06127_),
    .A(_06124_),
    .B(_06126_));
 sg13g2_nand2_1 _28726_ (.Y(_06128_),
    .A(net4727),
    .B(_05731_));
 sg13g2_xor2_1 _28727_ (.B(_06128_),
    .A(net4790),
    .X(_06129_));
 sg13g2_nor2_1 _28728_ (.A(net4501),
    .B(_05729_),
    .Y(_06130_));
 sg13g2_xnor2_1 _28729_ (.Y(_06131_),
    .A(\u_inv.d_reg[16] ),
    .B(_06130_));
 sg13g2_a21oi_1 _28730_ (.A1(_10951_),
    .A2(_05729_),
    .Y(_06132_),
    .B1(net4501));
 sg13g2_xnor2_1 _28731_ (.Y(_06133_),
    .A(net4791),
    .B(_06132_));
 sg13g2_nor2_1 _28732_ (.A(_06131_),
    .B(_06133_),
    .Y(_06134_));
 sg13g2_nand2b_1 _28733_ (.Y(_06135_),
    .B(_06134_),
    .A_N(_06129_));
 sg13g2_a21oi_1 _28734_ (.A1(_10953_),
    .A2(_05727_),
    .Y(_06136_),
    .B1(net4501));
 sg13g2_xnor2_1 _28735_ (.Y(_06137_),
    .A(_10952_),
    .B(_06136_));
 sg13g2_inv_1 _28736_ (.Y(_06138_),
    .A(_06137_));
 sg13g2_nor2_1 _28737_ (.A(net4501),
    .B(_05727_),
    .Y(_06139_));
 sg13g2_xnor2_1 _28738_ (.Y(_06140_),
    .A(\u_inv.d_reg[14] ),
    .B(_06139_));
 sg13g2_nor2_1 _28739_ (.A(net4502),
    .B(_05726_),
    .Y(_06141_));
 sg13g2_xnor2_1 _28740_ (.Y(_06142_),
    .A(\u_inv.d_reg[13] ),
    .B(_06141_));
 sg13g2_nand2_1 _28741_ (.Y(_06143_),
    .A(net4728),
    .B(_05725_));
 sg13g2_nand3_1 _28742_ (.B(net4793),
    .C(_05725_),
    .A(net4728),
    .Y(_06144_));
 sg13g2_nand2b_1 _28743_ (.Y(_06145_),
    .B(_06143_),
    .A_N(net4793));
 sg13g2_xor2_1 _28744_ (.B(_06143_),
    .A(net4793),
    .X(_06146_));
 sg13g2_nand2b_1 _28745_ (.Y(_06147_),
    .B(net4727),
    .A_N(_05723_));
 sg13g2_xnor2_1 _28746_ (.Y(_06148_),
    .A(\u_inv.d_reg[9] ),
    .B(_06147_));
 sg13g2_xnor2_1 _28747_ (.Y(_06149_),
    .A(_10955_),
    .B(_06147_));
 sg13g2_o21ai_1 _28748_ (.B1(net4728),
    .Y(_06150_),
    .A1(net4794),
    .A2(_05722_));
 sg13g2_xnor2_1 _28749_ (.Y(_06151_),
    .A(_10956_),
    .B(_06150_));
 sg13g2_xnor2_1 _28750_ (.Y(_06152_),
    .A(\u_inv.d_reg[8] ),
    .B(_06150_));
 sg13g2_and3_1 _28751_ (.X(_06153_),
    .A(net4725),
    .B(\u_inv.d_reg[3] ),
    .C(_05719_));
 sg13g2_a21oi_1 _28752_ (.A1(net4725),
    .A2(_05719_),
    .Y(_06154_),
    .B1(\u_inv.d_reg[3] ));
 sg13g2_nor2_1 _28753_ (.A(_06153_),
    .B(_06154_),
    .Y(_06155_));
 sg13g2_o21ai_1 _28754_ (.B1(net4726),
    .Y(_06156_),
    .A1(net4797),
    .A2(net4799));
 sg13g2_xor2_1 _28755_ (.B(_06156_),
    .A(net4796),
    .X(_06157_));
 sg13g2_xnor2_1 _28756_ (.Y(_06158_),
    .A(\u_inv.d_reg[2] ),
    .B(_06156_));
 sg13g2_nand3_1 _28757_ (.B(net4798),
    .C(net4800),
    .A(net4726),
    .Y(_06159_));
 sg13g2_a21o_1 _28758_ (.A2(net4800),
    .A1(net4726),
    .B1(net4798),
    .X(_06160_));
 sg13g2_nand3_1 _28759_ (.B(_06159_),
    .C(_06160_),
    .A(net4800),
    .Y(_06161_));
 sg13g2_inv_1 _28760_ (.Y(_06162_),
    .A(_06161_));
 sg13g2_nor2_1 _28761_ (.A(_06157_),
    .B(_06161_),
    .Y(_06163_));
 sg13g2_nor4_2 _28762_ (.A(_06153_),
    .B(_06154_),
    .C(_06157_),
    .Y(_06164_),
    .D(_06161_));
 sg13g2_nand2_1 _28763_ (.Y(_06165_),
    .A(net4725),
    .B(_05720_));
 sg13g2_xnor2_1 _28764_ (.Y(_06166_),
    .A(\u_inv.d_reg[4] ),
    .B(_06165_));
 sg13g2_or2_1 _28765_ (.X(_06167_),
    .B(_06166_),
    .A(_06164_));
 sg13g2_o21ai_1 _28766_ (.B1(net4725),
    .Y(_06168_),
    .A1(\u_inv.d_reg[4] ),
    .A2(_05720_));
 sg13g2_xnor2_1 _28767_ (.Y(_06169_),
    .A(\u_inv.d_reg[5] ),
    .B(_06168_));
 sg13g2_o21ai_1 _28768_ (.B1(_06169_),
    .Y(_06170_),
    .A1(_06164_),
    .A2(_06166_));
 sg13g2_o21ai_1 _28769_ (.B1(net4725),
    .Y(_06171_),
    .A1(\u_inv.d_reg[5] ),
    .A2(_05721_));
 sg13g2_xor2_1 _28770_ (.B(_06171_),
    .A(\u_inv.d_reg[6] ),
    .X(_06172_));
 sg13g2_and2_1 _28771_ (.A(_06170_),
    .B(_06172_),
    .X(_06173_));
 sg13g2_nand2_1 _28772_ (.Y(_06174_),
    .A(net4728),
    .B(_05722_));
 sg13g2_xor2_1 _28773_ (.B(_06174_),
    .A(net4794),
    .X(_06175_));
 sg13g2_and4_1 _28774_ (.A(_06149_),
    .B(_06151_),
    .C(_06173_),
    .D(_06175_),
    .X(_06176_));
 sg13g2_a21oi_1 _28775_ (.A1(_10955_),
    .A2(_05723_),
    .Y(_06177_),
    .B1(net4502));
 sg13g2_xor2_1 _28776_ (.B(_06177_),
    .A(\u_inv.d_reg[10] ),
    .X(_06178_));
 sg13g2_nor2b_1 _28777_ (.A(_06146_),
    .B_N(_06178_),
    .Y(_06179_));
 sg13g2_nand2b_2 _28778_ (.Y(_06180_),
    .B(_06179_),
    .A_N(_06176_));
 sg13g2_o21ai_1 _28779_ (.B1(net4728),
    .Y(_06181_),
    .A1(net4793),
    .A2(_05725_));
 sg13g2_xnor2_1 _28780_ (.Y(_06182_),
    .A(_10954_),
    .B(_06181_));
 sg13g2_or2_1 _28781_ (.X(_06183_),
    .B(_06182_),
    .A(_06142_));
 sg13g2_nor4_2 _28782_ (.A(_06138_),
    .B(_06140_),
    .C(_06180_),
    .Y(_06184_),
    .D(_06183_));
 sg13g2_o21ai_1 _28783_ (.B1(net4727),
    .Y(_06185_),
    .A1(net4790),
    .A2(_05731_));
 sg13g2_xor2_1 _28784_ (.B(_06185_),
    .A(\u_inv.d_reg[19] ),
    .X(_06186_));
 sg13g2_nor4_1 _28785_ (.A(_06129_),
    .B(_06131_),
    .C(_06133_),
    .D(_06186_),
    .Y(_06187_));
 sg13g2_nand2_2 _28786_ (.Y(_06188_),
    .A(_06184_),
    .B(_06187_));
 sg13g2_inv_1 _28787_ (.Y(_06189_),
    .A(_06188_));
 sg13g2_nor3_1 _28788_ (.A(_06121_),
    .B(_06127_),
    .C(_06188_),
    .Y(_06190_));
 sg13g2_nand2_1 _28789_ (.Y(_06191_),
    .A(_06116_),
    .B(_06190_));
 sg13g2_nor2_1 _28790_ (.A(_06111_),
    .B(_06191_),
    .Y(_06192_));
 sg13g2_nor3_1 _28791_ (.A(_06109_),
    .B(_06111_),
    .C(_06191_),
    .Y(_06193_));
 sg13g2_nand2b_1 _28792_ (.Y(_06194_),
    .B(_06192_),
    .A_N(_06109_));
 sg13g2_nand4_1 _28793_ (.B(_06104_),
    .C(_06107_),
    .A(_06101_),
    .Y(_06195_),
    .D(_06193_));
 sg13g2_and2_1 _28794_ (.A(_06096_),
    .B(_06195_),
    .X(_06196_));
 sg13g2_o21ai_1 _28795_ (.B1(net4734),
    .Y(_06197_),
    .A1(\u_inv.d_reg[32] ),
    .A2(_05745_));
 sg13g2_xnor2_1 _28796_ (.Y(_06198_),
    .A(\u_inv.d_reg[33] ),
    .B(_06197_));
 sg13g2_inv_2 _28797_ (.Y(_06199_),
    .A(_06198_));
 sg13g2_xor2_1 _28798_ (.B(_06076_),
    .A(\u_inv.d_reg[38] ),
    .X(_06200_));
 sg13g2_or4_1 _28799_ (.A(_06095_),
    .B(_06196_),
    .C(_06199_),
    .D(_06200_),
    .X(_06201_));
 sg13g2_o21ai_1 _28800_ (.B1(net4738),
    .Y(_06202_),
    .A1(\u_inv.d_reg[48] ),
    .A2(_05756_));
 sg13g2_xnor2_1 _28801_ (.Y(_06203_),
    .A(\u_inv.d_reg[49] ),
    .B(_06202_));
 sg13g2_inv_1 _28802_ (.Y(_06204_),
    .A(_06203_));
 sg13g2_nand2_1 _28803_ (.Y(_06205_),
    .A(net4735),
    .B(_05753_));
 sg13g2_o21ai_1 _28804_ (.B1(net4735),
    .Y(_06206_),
    .A1(\u_inv.d_reg[44] ),
    .A2(_05753_));
 sg13g2_xnor2_1 _28805_ (.Y(_06207_),
    .A(\u_inv.d_reg[45] ),
    .B(_06206_));
 sg13g2_xnor2_1 _28806_ (.Y(_06208_),
    .A(\u_inv.d_reg[44] ),
    .B(_06205_));
 sg13g2_nand2_1 _28807_ (.Y(_06209_),
    .A(_06207_),
    .B(_06208_));
 sg13g2_nand3_1 _28808_ (.B(_06207_),
    .C(_06208_),
    .A(_06203_),
    .Y(_06210_));
 sg13g2_or4_1 _28809_ (.A(_06074_),
    .B(_06093_),
    .C(_06201_),
    .D(_06210_),
    .X(_06211_));
 sg13g2_nor4_2 _28810_ (.A(_06055_),
    .B(_06057_),
    .C(_06069_),
    .Y(_06212_),
    .D(_06211_));
 sg13g2_nand2_1 _28811_ (.Y(_06213_),
    .A(net4742),
    .B(_05767_));
 sg13g2_xor2_1 _28812_ (.B(_06213_),
    .A(net4784),
    .X(_06214_));
 sg13g2_nor2_1 _28813_ (.A(net4506),
    .B(net3493),
    .Y(_06215_));
 sg13g2_xnor2_1 _28814_ (.Y(_06216_),
    .A(\u_inv.d_reg[56] ),
    .B(_06215_));
 sg13g2_o21ai_1 _28815_ (.B1(net4741),
    .Y(_06217_),
    .A1(\u_inv.d_reg[54] ),
    .A2(_05761_));
 sg13g2_xor2_1 _28816_ (.B(_06217_),
    .A(\u_inv.d_reg[55] ),
    .X(_06218_));
 sg13g2_o21ai_1 _28817_ (.B1(net4737),
    .Y(_06219_),
    .A1(_05756_),
    .A2(_05759_));
 sg13g2_xnor2_1 _28818_ (.Y(_06220_),
    .A(_10938_),
    .B(_06219_));
 sg13g2_inv_1 _28819_ (.Y(_06221_),
    .A(_06220_));
 sg13g2_o21ai_1 _28820_ (.B1(_06219_),
    .Y(_06222_),
    .A1(net4506),
    .A2(_10938_));
 sg13g2_xnor2_1 _28821_ (.Y(_06223_),
    .A(\u_inv.d_reg[53] ),
    .B(_06222_));
 sg13g2_inv_1 _28822_ (.Y(_06224_),
    .A(_06223_));
 sg13g2_nand2_1 _28823_ (.Y(_06225_),
    .A(_06221_),
    .B(_06224_));
 sg13g2_nor4_2 _28824_ (.A(_06214_),
    .B(_06216_),
    .C(_06218_),
    .Y(_06226_),
    .D(_06225_));
 sg13g2_nand4_1 _28825_ (.B(_06052_),
    .C(_06212_),
    .A(_06049_),
    .Y(_06227_),
    .D(_06226_));
 sg13g2_o21ai_1 _28826_ (.B1(net4740),
    .Y(_06228_),
    .A1(\u_inv.d_reg[62] ),
    .A2(\u_inv.d_reg[61] ));
 sg13g2_nand2_1 _28827_ (.Y(_06229_),
    .A(_06046_),
    .B(_06228_));
 sg13g2_xor2_1 _28828_ (.B(_06229_),
    .A(\u_inv.d_reg[63] ),
    .X(_06230_));
 sg13g2_o21ai_1 _28829_ (.B1(net4743),
    .Y(_06231_),
    .A1(_05767_),
    .A2(_05768_));
 sg13g2_xor2_1 _28830_ (.B(_06231_),
    .A(\u_inv.d_reg[66] ),
    .X(_06232_));
 sg13g2_inv_1 _28831_ (.Y(_06233_),
    .A(_06232_));
 sg13g2_nand4_1 _28832_ (.B(_05764_),
    .C(_05766_),
    .A(_05763_),
    .Y(_06234_),
    .D(_05790_));
 sg13g2_nand2_1 _28833_ (.Y(_06235_),
    .A(net4746),
    .B(_06234_));
 sg13g2_xnor2_1 _28834_ (.Y(_06236_),
    .A(\u_inv.d_reg[92] ),
    .B(_06235_));
 sg13g2_o21ai_1 _28835_ (.B1(net4743),
    .Y(_06237_),
    .A1(\u_inv.d_reg[64] ),
    .A2(_05767_));
 sg13g2_xor2_1 _28836_ (.B(_06237_),
    .A(\u_inv.d_reg[65] ),
    .X(_06238_));
 sg13g2_o21ai_1 _28837_ (.B1(_06046_),
    .Y(_06239_),
    .A1(net4506),
    .A2(_10934_));
 sg13g2_xor2_1 _28838_ (.B(_06239_),
    .A(\u_inv.d_reg[62] ),
    .X(_06240_));
 sg13g2_nand2b_1 _28839_ (.Y(_06241_),
    .B(_06240_),
    .A_N(_06238_));
 sg13g2_o21ai_1 _28840_ (.B1(net4743),
    .Y(_06242_),
    .A1(_05767_),
    .A2(_05769_));
 sg13g2_xnor2_1 _28841_ (.Y(_06243_),
    .A(_10933_),
    .B(_06242_));
 sg13g2_o21ai_1 _28842_ (.B1(net4740),
    .Y(_06244_),
    .A1(\u_inv.d_reg[57] ),
    .A2(_06053_));
 sg13g2_o21ai_1 _28843_ (.B1(_06244_),
    .Y(_06245_),
    .A1(net4506),
    .A2(_10935_));
 sg13g2_xnor2_1 _28844_ (.Y(_06246_),
    .A(\u_inv.d_reg[59] ),
    .B(_06245_));
 sg13g2_xor2_1 _28845_ (.B(_06244_),
    .A(net4785),
    .X(_06247_));
 sg13g2_nor4_1 _28846_ (.A(_06241_),
    .B(_06243_),
    .C(_06246_),
    .D(_06247_),
    .Y(_06248_));
 sg13g2_nand4_1 _28847_ (.B(_06233_),
    .C(_06236_),
    .A(_06230_),
    .Y(_06249_),
    .D(_06248_));
 sg13g2_o21ai_1 _28848_ (.B1(net4747),
    .Y(_06250_),
    .A1(_05771_),
    .A2(_06034_));
 sg13g2_xor2_1 _28849_ (.B(_06250_),
    .A(\u_inv.d_reg[70] ),
    .X(_06251_));
 sg13g2_o21ai_1 _28850_ (.B1(net4746),
    .Y(_06252_),
    .A1(\u_inv.d_reg[92] ),
    .A2(_06234_));
 sg13g2_xnor2_1 _28851_ (.Y(_06253_),
    .A(\u_inv.d_reg[93] ),
    .B(_06252_));
 sg13g2_nand2b_1 _28852_ (.Y(_06254_),
    .B(_06253_),
    .A_N(_06251_));
 sg13g2_nor2b_1 _28853_ (.A(net3492),
    .B_N(_05803_),
    .Y(_06255_));
 sg13g2_nand2b_2 _28854_ (.Y(_06256_),
    .B(_05803_),
    .A_N(net3492));
 sg13g2_nand2_1 _28855_ (.Y(_06257_),
    .A(net4748),
    .B(_06256_));
 sg13g2_xor2_1 _28856_ (.B(_06257_),
    .A(\u_inv.d_reg[100] ),
    .X(_06258_));
 sg13g2_nand4_1 _28857_ (.B(_05764_),
    .C(_05766_),
    .A(_05763_),
    .Y(_06259_),
    .D(_05786_));
 sg13g2_nand2_1 _28858_ (.Y(_06260_),
    .A(net4745),
    .B(_06259_));
 sg13g2_o21ai_1 _28859_ (.B1(net4746),
    .Y(_06261_),
    .A1(_05787_),
    .A2(_06259_));
 sg13g2_xnor2_1 _28860_ (.Y(_06262_),
    .A(_10928_),
    .B(_06261_));
 sg13g2_o21ai_1 _28861_ (.B1(net4747),
    .Y(_06263_),
    .A1(net4783),
    .A2(_06040_));
 sg13g2_xnor2_1 _28862_ (.Y(_06264_),
    .A(\u_inv.d_reg[73] ),
    .B(_06263_));
 sg13g2_o21ai_1 _28863_ (.B1(net4746),
    .Y(_06265_),
    .A1(_05792_),
    .A2(_06234_));
 sg13g2_xnor2_1 _28864_ (.Y(_06266_),
    .A(_10927_),
    .B(_06265_));
 sg13g2_inv_1 _28865_ (.Y(_06267_),
    .A(_06266_));
 sg13g2_o21ai_1 _28866_ (.B1(net4747),
    .Y(_06268_),
    .A1(_05772_),
    .A2(_06034_));
 sg13g2_xor2_1 _28867_ (.B(_06268_),
    .A(\u_inv.d_reg[71] ),
    .X(_06269_));
 sg13g2_xnor2_1 _28868_ (.Y(_06270_),
    .A(\u_inv.d_reg[71] ),
    .B(_06268_));
 sg13g2_o21ai_1 _28869_ (.B1(net4745),
    .Y(_06271_),
    .A1(_05780_),
    .A2(_06037_));
 sg13g2_o21ai_1 _28870_ (.B1(net4745),
    .Y(_06272_),
    .A1(_05781_),
    .A2(_06037_));
 sg13g2_xnor2_1 _28871_ (.Y(_06273_),
    .A(\u_inv.d_reg[83] ),
    .B(_06272_));
 sg13g2_nand4_1 _28872_ (.B(_06267_),
    .C(_06270_),
    .A(_06264_),
    .Y(_06274_),
    .D(_06273_));
 sg13g2_or4_1 _28873_ (.A(_06254_),
    .B(_06258_),
    .C(_06262_),
    .D(_06274_),
    .X(_06275_));
 sg13g2_o21ai_1 _28874_ (.B1(net4748),
    .Y(_06276_),
    .A1(_05799_),
    .A2(_06256_));
 sg13g2_o21ai_1 _28875_ (.B1(net4748),
    .Y(_06277_),
    .A1(_05800_),
    .A2(_06256_));
 sg13g2_xnor2_1 _28876_ (.Y(_06278_),
    .A(_10925_),
    .B(_06277_));
 sg13g2_xor2_1 _28877_ (.B(_06276_),
    .A(\u_inv.d_reg[102] ),
    .X(_06279_));
 sg13g2_nor2_1 _28878_ (.A(net4507),
    .B(_05776_),
    .Y(_06280_));
 sg13g2_a21oi_2 _28879_ (.B1(_06280_),
    .Y(_06281_),
    .A2(_06040_),
    .A1(net4747));
 sg13g2_o21ai_1 _28880_ (.B1(net4748),
    .Y(_06282_),
    .A1(net4781),
    .A2(net4782));
 sg13g2_nand2_1 _28881_ (.Y(_06283_),
    .A(_06281_),
    .B(_06282_));
 sg13g2_xnor2_1 _28882_ (.Y(_06284_),
    .A(\u_inv.d_reg[78] ),
    .B(_06283_));
 sg13g2_o21ai_1 _28883_ (.B1(_06281_),
    .Y(_06285_),
    .A1(net4507),
    .A2(_10930_));
 sg13g2_xor2_1 _28884_ (.B(_06285_),
    .A(net4781),
    .X(_06286_));
 sg13g2_o21ai_1 _28885_ (.B1(net4746),
    .Y(_06287_),
    .A1(\u_inv.d_reg[88] ),
    .A2(_06259_));
 sg13g2_xnor2_1 _28886_ (.Y(_06288_),
    .A(\u_inv.d_reg[89] ),
    .B(_06287_));
 sg13g2_xnor2_1 _28887_ (.Y(_06289_),
    .A(\u_inv.d_reg[88] ),
    .B(_06260_));
 sg13g2_and2_1 _28888_ (.A(_06288_),
    .B(_06289_),
    .X(_06290_));
 sg13g2_o21ai_1 _28889_ (.B1(net4748),
    .Y(_06291_),
    .A1(\u_inv.d_reg[100] ),
    .A2(_06256_));
 sg13g2_xnor2_1 _28890_ (.Y(_06292_),
    .A(\u_inv.d_reg[101] ),
    .B(_06291_));
 sg13g2_xor2_1 _28891_ (.B(_06291_),
    .A(\u_inv.d_reg[101] ),
    .X(_06293_));
 sg13g2_nand2_1 _28892_ (.Y(_06294_),
    .A(net4748),
    .B(\u_inv.d_reg[78] ));
 sg13g2_and3_1 _28893_ (.X(_06295_),
    .A(_06281_),
    .B(_06282_),
    .C(_06294_));
 sg13g2_xnor2_1 _28894_ (.Y(_06296_),
    .A(\u_inv.d_reg[79] ),
    .B(_06295_));
 sg13g2_xor2_1 _28895_ (.B(_06295_),
    .A(\u_inv.d_reg[79] ),
    .X(_06297_));
 sg13g2_nand4_1 _28896_ (.B(_06290_),
    .C(_06292_),
    .A(_06286_),
    .Y(_06298_),
    .D(_06296_));
 sg13g2_or4_1 _28897_ (.A(_06278_),
    .B(_06279_),
    .C(_06284_),
    .D(_06298_),
    .X(_06299_));
 sg13g2_or4_1 _28898_ (.A(_06227_),
    .B(_06249_),
    .C(_06275_),
    .D(_06299_),
    .X(_06300_));
 sg13g2_nor4_1 _28899_ (.A(_06018_),
    .B(_06025_),
    .C(_06033_),
    .D(_06300_),
    .Y(_06301_));
 sg13g2_nor2b_1 _28900_ (.A(\u_inv.d_reg[128] ),
    .B_N(net3489),
    .Y(_06302_));
 sg13g2_nor2_1 _28901_ (.A(net4509),
    .B(_06302_),
    .Y(_06303_));
 sg13g2_a21oi_1 _28902_ (.A1(_10919_),
    .A2(_06302_),
    .Y(_06304_),
    .B1(net4509));
 sg13g2_xor2_1 _28903_ (.B(_06304_),
    .A(\u_inv.d_reg[130] ),
    .X(_06305_));
 sg13g2_a21oi_2 _28904_ (.B1(net4508),
    .Y(_06306_),
    .A2(_06255_),
    .A1(_05801_));
 sg13g2_nand3_1 _28905_ (.B(_05801_),
    .C(_06255_),
    .A(_05798_),
    .Y(_06307_));
 sg13g2_nand2_1 _28906_ (.Y(_06308_),
    .A(net4750),
    .B(_06307_));
 sg13g2_o21ai_1 _28907_ (.B1(net4750),
    .Y(_06309_),
    .A1(\u_inv.d_reg[110] ),
    .A2(_06307_));
 sg13g2_xnor2_1 _28908_ (.Y(_06310_),
    .A(\u_inv.d_reg[111] ),
    .B(_06309_));
 sg13g2_xnor2_1 _28909_ (.Y(_06311_),
    .A(_10922_),
    .B(_06309_));
 sg13g2_o21ai_1 _28910_ (.B1(net4752),
    .Y(_06312_),
    .A1(_05715_),
    .A2(_05812_));
 sg13g2_o21ai_1 _28911_ (.B1(net4752),
    .Y(_06313_),
    .A1(_05716_),
    .A2(_05812_));
 sg13g2_xnor2_1 _28912_ (.Y(_06314_),
    .A(\u_inv.d_reg[123] ),
    .B(_06313_));
 sg13g2_xnor2_1 _28913_ (.Y(_06315_),
    .A(\u_inv.d_reg[122] ),
    .B(_06312_));
 sg13g2_nand2_2 _28914_ (.Y(_06316_),
    .A(_06314_),
    .B(_06315_));
 sg13g2_a21oi_1 _28915_ (.A1(net4750),
    .A2(net4780),
    .Y(_06317_),
    .B1(_06306_));
 sg13g2_xnor2_1 _28916_ (.Y(_06318_),
    .A(_10924_),
    .B(_06317_));
 sg13g2_xnor2_1 _28917_ (.Y(_06319_),
    .A(\u_inv.d_reg[105] ),
    .B(_06317_));
 sg13g2_xor2_1 _28918_ (.B(_06306_),
    .A(net4780),
    .X(_06320_));
 sg13g2_inv_1 _28919_ (.Y(_06321_),
    .A(_06320_));
 sg13g2_nand2_1 _28920_ (.Y(_06322_),
    .A(_06319_),
    .B(_06320_));
 sg13g2_nor2_1 _28921_ (.A(_05783_),
    .B(_06037_),
    .Y(_06323_));
 sg13g2_or2_1 _28922_ (.X(_06324_),
    .B(_06037_),
    .A(_05783_));
 sg13g2_nand2_1 _28923_ (.Y(_06325_),
    .A(net4745),
    .B(_06324_));
 sg13g2_o21ai_1 _28924_ (.B1(net4745),
    .Y(_06326_),
    .A1(\u_inv.d_reg[84] ),
    .A2(_06324_));
 sg13g2_xnor2_1 _28925_ (.Y(_06327_),
    .A(\u_inv.d_reg[85] ),
    .B(_06326_));
 sg13g2_xnor2_1 _28926_ (.Y(_06328_),
    .A(\u_inv.d_reg[84] ),
    .B(_06325_));
 sg13g2_nand2_2 _28927_ (.Y(_06329_),
    .A(_06327_),
    .B(_06328_));
 sg13g2_nor4_2 _28928_ (.A(_06311_),
    .B(_06316_),
    .C(_06322_),
    .Y(_06330_),
    .D(_06329_));
 sg13g2_or2_1 _28929_ (.X(_06331_),
    .B(_05812_),
    .A(_05717_));
 sg13g2_nand2_1 _28930_ (.Y(_06332_),
    .A(net4752),
    .B(_06331_));
 sg13g2_o21ai_1 _28931_ (.B1(net4751),
    .Y(_06333_),
    .A1(\u_inv.d_reg[124] ),
    .A2(_06331_));
 sg13g2_xnor2_1 _28932_ (.Y(_06334_),
    .A(\u_inv.d_reg[125] ),
    .B(_06333_));
 sg13g2_xnor2_1 _28933_ (.Y(_06335_),
    .A(\u_inv.d_reg[124] ),
    .B(_06332_));
 sg13g2_nand2_1 _28934_ (.Y(_06336_),
    .A(_06334_),
    .B(_06335_));
 sg13g2_xnor2_1 _28935_ (.Y(_06337_),
    .A(\u_inv.d_reg[129] ),
    .B(_06303_));
 sg13g2_nand2_1 _28936_ (.Y(_06338_),
    .A(net4756),
    .B(_05954_));
 sg13g2_xor2_1 _28937_ (.B(_06338_),
    .A(\u_inv.d_reg[132] ),
    .X(_06339_));
 sg13g2_a21oi_1 _28938_ (.A1(_05819_),
    .A2(_06302_),
    .Y(_06340_),
    .B1(net4509));
 sg13g2_xor2_1 _28939_ (.B(_06340_),
    .A(\u_inv.d_reg[131] ),
    .X(_06341_));
 sg13g2_nand2b_1 _28940_ (.Y(_06342_),
    .B(_06341_),
    .A_N(_06339_));
 sg13g2_xnor2_1 _28941_ (.Y(_06343_),
    .A(\u_inv.d_reg[110] ),
    .B(_06308_));
 sg13g2_nand2_1 _28942_ (.Y(_06344_),
    .A(net4748),
    .B(net3492));
 sg13g2_o21ai_1 _28943_ (.B1(net4748),
    .Y(_06345_),
    .A1(\u_inv.d_reg[96] ),
    .A2(net3492));
 sg13g2_xnor2_1 _28944_ (.Y(_06346_),
    .A(\u_inv.d_reg[97] ),
    .B(_06345_));
 sg13g2_inv_1 _28945_ (.Y(_06347_),
    .A(_06346_));
 sg13g2_o21ai_1 _28946_ (.B1(net4749),
    .Y(_06348_),
    .A1(net3492),
    .A2(_05802_));
 sg13g2_xnor2_1 _28947_ (.Y(_06349_),
    .A(_10926_),
    .B(_06348_));
 sg13g2_inv_1 _28948_ (.Y(_06350_),
    .A(_06349_));
 sg13g2_xor2_1 _28949_ (.B(_06344_),
    .A(\u_inv.d_reg[96] ),
    .X(_06351_));
 sg13g2_inv_2 _28950_ (.Y(_06352_),
    .A(_06351_));
 sg13g2_nor3_1 _28951_ (.A(_06347_),
    .B(_06349_),
    .C(_06351_),
    .Y(_06353_));
 sg13g2_and2_1 _28952_ (.A(_06343_),
    .B(_06353_),
    .X(_06354_));
 sg13g2_nor2_1 _28953_ (.A(net4508),
    .B(_05796_),
    .Y(_06355_));
 sg13g2_or2_1 _28954_ (.X(_06356_),
    .B(_06355_),
    .A(_06306_));
 sg13g2_xor2_1 _28955_ (.B(_06356_),
    .A(\u_inv.d_reg[108] ),
    .X(_06357_));
 sg13g2_o21ai_1 _28956_ (.B1(net4753),
    .Y(_06358_),
    .A1(_05809_),
    .A2(_06027_));
 sg13g2_xor2_1 _28957_ (.B(_06358_),
    .A(\u_inv.d_reg[118] ),
    .X(_06359_));
 sg13g2_nor2b_1 _28958_ (.A(_06359_),
    .B_N(_06357_),
    .Y(_06360_));
 sg13g2_xnor2_1 _28959_ (.Y(_06361_),
    .A(\u_inv.d_reg[82] ),
    .B(_06271_));
 sg13g2_o21ai_1 _28960_ (.B1(net4743),
    .Y(_06362_),
    .A1(\u_inv.d_reg[68] ),
    .A2(_06034_));
 sg13g2_xnor2_1 _28961_ (.Y(_06363_),
    .A(_10932_),
    .B(_06362_));
 sg13g2_o21ai_1 _28962_ (.B1(net4746),
    .Y(_06364_),
    .A1(_05791_),
    .A2(_06234_));
 sg13g2_xnor2_1 _28963_ (.Y(_06365_),
    .A(\u_inv.d_reg[94] ),
    .B(_06364_));
 sg13g2_nand3b_1 _28964_ (.B(_06365_),
    .C(_06361_),
    .Y(_06366_),
    .A_N(_06363_));
 sg13g2_xor2_1 _28965_ (.B(_06050_),
    .A(\u_inv.d_reg[74] ),
    .X(_06367_));
 sg13g2_inv_1 _28966_ (.Y(_06368_),
    .A(_06367_));
 sg13g2_a21oi_1 _28967_ (.A1(_05784_),
    .A2(_06323_),
    .Y(_06369_),
    .B1(net4507));
 sg13g2_xor2_1 _28968_ (.B(_06369_),
    .A(\u_inv.d_reg[87] ),
    .X(_06370_));
 sg13g2_xnor2_1 _28969_ (.Y(_06371_),
    .A(net4782),
    .B(_06281_));
 sg13g2_o21ai_1 _28970_ (.B1(net4745),
    .Y(_06372_),
    .A1(\u_inv.d_reg[80] ),
    .A2(_06037_));
 sg13g2_xnor2_1 _28971_ (.Y(_06373_),
    .A(\u_inv.d_reg[81] ),
    .B(_06372_));
 sg13g2_nand4_1 _28972_ (.B(_06370_),
    .C(_06371_),
    .A(_06368_),
    .Y(_06374_),
    .D(_06373_));
 sg13g2_xnor2_1 _28973_ (.Y(_06375_),
    .A(\u_inv.d_reg[126] ),
    .B(_06012_));
 sg13g2_o21ai_1 _28974_ (.B1(net4745),
    .Y(_06376_),
    .A1(_05782_),
    .A2(_06324_));
 sg13g2_xnor2_1 _28975_ (.Y(_06377_),
    .A(\u_inv.d_reg[86] ),
    .B(_06376_));
 sg13g2_nand2_1 _28976_ (.Y(_06378_),
    .A(_06375_),
    .B(_06377_));
 sg13g2_nor3_1 _28977_ (.A(_06366_),
    .B(_06374_),
    .C(_06378_),
    .Y(_06379_));
 sg13g2_a21oi_1 _28978_ (.A1(_10926_),
    .A2(_06348_),
    .Y(_06380_),
    .B1(net4508));
 sg13g2_xor2_1 _28979_ (.B(_06380_),
    .A(\u_inv.d_reg[99] ),
    .X(_06381_));
 sg13g2_a21oi_1 _28980_ (.A1(net4750),
    .A2(_05797_),
    .Y(_06382_),
    .B1(_06306_));
 sg13g2_xnor2_1 _28981_ (.Y(_06383_),
    .A(\u_inv.d_reg[109] ),
    .B(_06382_));
 sg13g2_o21ai_1 _28982_ (.B1(net4751),
    .Y(_06384_),
    .A1(_05810_),
    .A2(_06027_));
 sg13g2_xnor2_1 _28983_ (.Y(_06385_),
    .A(\u_inv.d_reg[119] ),
    .B(_06384_));
 sg13g2_xor2_1 _28984_ (.B(_06384_),
    .A(\u_inv.d_reg[119] ),
    .X(_06386_));
 sg13g2_a21oi_1 _28985_ (.A1(_10928_),
    .A2(_06261_),
    .Y(_06387_),
    .B1(net4507));
 sg13g2_xor2_1 _28986_ (.B(_06387_),
    .A(\u_inv.d_reg[91] ),
    .X(_06388_));
 sg13g2_nand4_1 _28987_ (.B(_06383_),
    .C(_06385_),
    .A(_06381_),
    .Y(_06389_),
    .D(_06388_));
 sg13g2_o21ai_1 _28988_ (.B1(net4753),
    .Y(_06390_),
    .A1(\u_inv.d_reg[112] ),
    .A2(_05806_));
 sg13g2_xor2_1 _28989_ (.B(_06390_),
    .A(\u_inv.d_reg[113] ),
    .X(_06391_));
 sg13g2_xor2_1 _28990_ (.B(_06026_),
    .A(\u_inv.d_reg[112] ),
    .X(_06392_));
 sg13g2_nor2_1 _28991_ (.A(_06391_),
    .B(_06392_),
    .Y(_06393_));
 sg13g2_o21ai_1 _28992_ (.B1(net4753),
    .Y(_06394_),
    .A1(_05806_),
    .A2(_05807_));
 sg13g2_o21ai_1 _28993_ (.B1(net4753),
    .Y(_06395_),
    .A1(_05806_),
    .A2(_05808_));
 sg13g2_xor2_1 _28994_ (.B(_06395_),
    .A(\u_inv.d_reg[115] ),
    .X(_06396_));
 sg13g2_inv_1 _28995_ (.Y(_06397_),
    .A(_06396_));
 sg13g2_xor2_1 _28996_ (.B(_06394_),
    .A(\u_inv.d_reg[114] ),
    .X(_06398_));
 sg13g2_nor2_1 _28997_ (.A(_06396_),
    .B(_06398_),
    .Y(_06399_));
 sg13g2_nand2_2 _28998_ (.Y(_06400_),
    .A(_06393_),
    .B(_06399_));
 sg13g2_o21ai_1 _28999_ (.B1(net4749),
    .Y(_06401_),
    .A1(\u_inv.d_reg[105] ),
    .A2(\u_inv.d_reg[104] ));
 sg13g2_nor2b_1 _29000_ (.A(_06306_),
    .B_N(_06401_),
    .Y(_06402_));
 sg13g2_a21oi_1 _29001_ (.A1(net4750),
    .A2(_05795_),
    .Y(_06403_),
    .B1(_06306_));
 sg13g2_xor2_1 _29002_ (.B(_06403_),
    .A(\u_inv.d_reg[107] ),
    .X(_06404_));
 sg13g2_xor2_1 _29003_ (.B(_06402_),
    .A(\u_inv.d_reg[106] ),
    .X(_06405_));
 sg13g2_nor4_1 _29004_ (.A(_06389_),
    .B(_06400_),
    .C(_06404_),
    .D(_06405_),
    .Y(_06406_));
 sg13g2_nand4_1 _29005_ (.B(_06360_),
    .C(_06379_),
    .A(_06354_),
    .Y(_06407_),
    .D(_06406_));
 sg13g2_nor4_1 _29006_ (.A(_06336_),
    .B(_06337_),
    .C(_06342_),
    .D(_06407_),
    .Y(_06408_));
 sg13g2_nand4_1 _29007_ (.B(_06305_),
    .C(_06330_),
    .A(_06301_),
    .Y(_06409_),
    .D(_06408_));
 sg13g2_o21ai_1 _29008_ (.B1(net4756),
    .Y(_06410_),
    .A1(_05822_),
    .A2(_05954_));
 sg13g2_xnor2_1 _29009_ (.Y(_06411_),
    .A(_10918_),
    .B(_06410_));
 sg13g2_xnor2_1 _29010_ (.Y(_06412_),
    .A(_10916_),
    .B(_05976_));
 sg13g2_xor2_1 _29011_ (.B(_05956_),
    .A(\u_inv.d_reg[136] ),
    .X(_06413_));
 sg13g2_xor2_1 _29012_ (.B(_05989_),
    .A(\u_inv.d_reg[160] ),
    .X(_06414_));
 sg13g2_nor4_1 _29013_ (.A(_06411_),
    .B(_06412_),
    .C(_06413_),
    .D(_06414_),
    .Y(_06415_));
 sg13g2_o21ai_1 _29014_ (.B1(net4757),
    .Y(_06416_),
    .A1(\u_inv.d_reg[132] ),
    .A2(_05954_));
 sg13g2_xnor2_1 _29015_ (.Y(_06417_),
    .A(\u_inv.d_reg[133] ),
    .B(_06416_));
 sg13g2_xor2_1 _29016_ (.B(_06416_),
    .A(\u_inv.d_reg[133] ),
    .X(_06418_));
 sg13g2_xor2_1 _29017_ (.B(_05975_),
    .A(\u_inv.d_reg[148] ),
    .X(_06419_));
 sg13g2_o21ai_1 _29018_ (.B1(net4756),
    .Y(_06420_),
    .A1(_05821_),
    .A2(_05954_));
 sg13g2_xor2_1 _29019_ (.B(_06420_),
    .A(\u_inv.d_reg[134] ),
    .X(_06421_));
 sg13g2_o21ai_1 _29020_ (.B1(net4759),
    .Y(_06422_),
    .A1(_05707_),
    .A2(_05826_));
 sg13g2_o21ai_1 _29021_ (.B1(net4759),
    .Y(_06423_),
    .A1(_05708_),
    .A2(_05826_));
 sg13g2_xor2_1 _29022_ (.B(_06423_),
    .A(\u_inv.d_reg[147] ),
    .X(_06424_));
 sg13g2_nor4_1 _29023_ (.A(_06418_),
    .B(_06419_),
    .C(_06421_),
    .D(_06424_),
    .Y(_06425_));
 sg13g2_nand2_1 _29024_ (.Y(_06426_),
    .A(_06415_),
    .B(_06425_));
 sg13g2_nor4_2 _29025_ (.A(_05999_),
    .B(_06011_),
    .C(_06409_),
    .Y(_06427_),
    .D(_06426_));
 sg13g2_nand2_1 _29026_ (.Y(_06428_),
    .A(net4740),
    .B(_05918_));
 sg13g2_xor2_1 _29027_ (.B(_06428_),
    .A(\u_inv.d_reg[200] ),
    .X(_06429_));
 sg13g2_o21ai_1 _29028_ (.B1(net4742),
    .Y(_06430_),
    .A1(_05852_),
    .A2(_05853_));
 sg13g2_xnor2_1 _29029_ (.Y(_06431_),
    .A(_10898_),
    .B(_06430_));
 sg13g2_nand2_1 _29030_ (.Y(_06432_),
    .A(net4738),
    .B(_05862_));
 sg13g2_xor2_1 _29031_ (.B(_06432_),
    .A(net4770),
    .X(_06433_));
 sg13g2_xnor2_1 _29032_ (.Y(_06434_),
    .A(\u_inv.d_reg[208] ),
    .B(_06432_));
 sg13g2_xor2_1 _29033_ (.B(_05932_),
    .A(\u_inv.d_reg[184] ),
    .X(_06435_));
 sg13g2_nor4_1 _29034_ (.A(_06429_),
    .B(_06431_),
    .C(_06433_),
    .D(_06435_),
    .Y(_06436_));
 sg13g2_nand2_1 _29035_ (.Y(_06437_),
    .A(net4742),
    .B(_05852_));
 sg13g2_o21ai_1 _29036_ (.B1(net4742),
    .Y(_06438_),
    .A1(_05852_),
    .A2(_05854_));
 sg13g2_xnor2_1 _29037_ (.Y(_06439_),
    .A(\u_inv.d_reg[195] ),
    .B(_06438_));
 sg13g2_inv_1 _29038_ (.Y(_06440_),
    .A(_06439_));
 sg13g2_or2_1 _29039_ (.X(_06441_),
    .B(_05837_),
    .A(_05829_));
 sg13g2_nand2_1 _29040_ (.Y(_06442_),
    .A(net4762),
    .B(_06441_));
 sg13g2_o21ai_1 _29041_ (.B1(net4763),
    .Y(_06443_),
    .A1(\u_inv.d_reg[172] ),
    .A2(_06441_));
 sg13g2_xnor2_1 _29042_ (.Y(_06444_),
    .A(_10906_),
    .B(_06443_));
 sg13g2_xnor2_1 _29043_ (.Y(_06445_),
    .A(_10907_),
    .B(_06442_));
 sg13g2_or2_1 _29044_ (.X(_06446_),
    .B(_06445_),
    .A(_06444_));
 sg13g2_o21ai_1 _29045_ (.B1(net4742),
    .Y(_06447_),
    .A1(\u_inv.d_reg[192] ),
    .A2(_05852_));
 sg13g2_xor2_1 _29046_ (.B(_06447_),
    .A(\u_inv.d_reg[193] ),
    .X(_06448_));
 sg13g2_o21ai_1 _29047_ (.B1(net4760),
    .Y(_06449_),
    .A1(_05701_),
    .A2(_05977_));
 sg13g2_xor2_1 _29048_ (.B(_06449_),
    .A(\u_inv.d_reg[154] ),
    .X(_06450_));
 sg13g2_o21ai_1 _29049_ (.B1(net4760),
    .Y(_06451_),
    .A1(_05702_),
    .A2(_05977_));
 sg13g2_xnor2_1 _29050_ (.Y(_06452_),
    .A(_10915_),
    .B(_06451_));
 sg13g2_or2_1 _29051_ (.X(_06453_),
    .B(_06452_),
    .A(_06450_));
 sg13g2_nor4_1 _29052_ (.A(_06440_),
    .B(_06446_),
    .C(_06448_),
    .D(_06453_),
    .Y(_06454_));
 sg13g2_o21ai_1 _29053_ (.B1(_06438_),
    .Y(_06455_),
    .A1(net4506),
    .A2(_10897_));
 sg13g2_o21ai_1 _29054_ (.B1(net4742),
    .Y(_06456_),
    .A1(net4772),
    .A2(net4773));
 sg13g2_nor2b_1 _29055_ (.A(_06455_),
    .B_N(_06456_),
    .Y(_06457_));
 sg13g2_nand2_1 _29056_ (.Y(_06458_),
    .A(net4742),
    .B(net4771));
 sg13g2_and2_1 _29057_ (.A(_06457_),
    .B(_06458_),
    .X(_06459_));
 sg13g2_xor2_1 _29058_ (.B(_06459_),
    .A(\u_inv.d_reg[199] ),
    .X(_06460_));
 sg13g2_xnor2_1 _29059_ (.Y(_06461_),
    .A(\u_inv.d_reg[188] ),
    .B(_05946_));
 sg13g2_nand2b_1 _29060_ (.Y(_06462_),
    .B(_06461_),
    .A_N(_06460_));
 sg13g2_xor2_1 _29061_ (.B(_06457_),
    .A(net4771),
    .X(_06463_));
 sg13g2_o21ai_1 _29062_ (.B1(net4755),
    .Y(_06464_),
    .A1(_05842_),
    .A2(_05931_));
 sg13g2_xor2_1 _29063_ (.B(_06464_),
    .A(\u_inv.d_reg[186] ),
    .X(_06465_));
 sg13g2_xor2_1 _29064_ (.B(_06422_),
    .A(\u_inv.d_reg[146] ),
    .X(_06466_));
 sg13g2_xor2_1 _29065_ (.B(_05974_),
    .A(\u_inv.d_reg[144] ),
    .X(_06467_));
 sg13g2_o21ai_1 _29066_ (.B1(net4760),
    .Y(_06468_),
    .A1(\u_inv.d_reg[144] ),
    .A2(_05826_));
 sg13g2_xor2_1 _29067_ (.B(_06468_),
    .A(\u_inv.d_reg[145] ),
    .X(_06469_));
 sg13g2_or3_1 _29068_ (.A(_06466_),
    .B(_06467_),
    .C(_06469_),
    .X(_06470_));
 sg13g2_o21ai_1 _29069_ (.B1(net4762),
    .Y(_06471_),
    .A1(\u_inv.d_reg[168] ),
    .A2(_05960_));
 sg13g2_xnor2_1 _29070_ (.Y(_06472_),
    .A(_10909_),
    .B(_06471_));
 sg13g2_o21ai_1 _29071_ (.B1(net4759),
    .Y(_06473_),
    .A1(\u_inv.d_reg[148] ),
    .A2(_05973_));
 sg13g2_xor2_1 _29072_ (.B(_06473_),
    .A(\u_inv.d_reg[149] ),
    .X(_06474_));
 sg13g2_o21ai_1 _29073_ (.B1(net4762),
    .Y(_06475_),
    .A1(_05836_),
    .A2(_05960_));
 sg13g2_xor2_1 _29074_ (.B(_06475_),
    .A(\u_inv.d_reg[170] ),
    .X(_06476_));
 sg13g2_nor4_1 _29075_ (.A(_06470_),
    .B(_06472_),
    .C(_06474_),
    .D(_06476_),
    .Y(_06477_));
 sg13g2_o21ai_1 _29076_ (.B1(net4764),
    .Y(_06478_),
    .A1(\u_inv.d_reg[176] ),
    .A2(_05841_));
 sg13g2_xor2_1 _29077_ (.B(_06478_),
    .A(\u_inv.d_reg[177] ),
    .X(_06479_));
 sg13g2_o21ai_1 _29078_ (.B1(net4761),
    .Y(_06480_),
    .A1(_05706_),
    .A2(_05977_));
 sg13g2_xor2_1 _29079_ (.B(_06480_),
    .A(\u_inv.d_reg[158] ),
    .X(_06481_));
 sg13g2_xor2_1 _29080_ (.B(_06437_),
    .A(\u_inv.d_reg[192] ),
    .X(_06482_));
 sg13g2_o21ai_1 _29081_ (.B1(net4762),
    .Y(_06483_),
    .A1(_05839_),
    .A2(_06441_));
 sg13g2_xor2_1 _29082_ (.B(_06483_),
    .A(\u_inv.d_reg[175] ),
    .X(_06484_));
 sg13g2_nor4_1 _29083_ (.A(_06479_),
    .B(_06481_),
    .C(_06482_),
    .D(_06484_),
    .Y(_06485_));
 sg13g2_o21ai_1 _29084_ (.B1(net4754),
    .Y(_06486_),
    .A1(_05846_),
    .A2(_05931_));
 sg13g2_xnor2_1 _29085_ (.Y(_06487_),
    .A(\u_inv.d_reg[191] ),
    .B(_06486_));
 sg13g2_o21ai_1 _29086_ (.B1(net4763),
    .Y(_06488_),
    .A1(_05838_),
    .A2(_06441_));
 sg13g2_xor2_1 _29087_ (.B(_06488_),
    .A(\u_inv.d_reg[174] ),
    .X(_06489_));
 sg13g2_o21ai_1 _29088_ (.B1(net4761),
    .Y(_06490_),
    .A1(_05704_),
    .A2(_05977_));
 sg13g2_xnor2_1 _29089_ (.Y(_06491_),
    .A(_10914_),
    .B(_06490_));
 sg13g2_nand2_1 _29090_ (.Y(_06492_),
    .A(net4762),
    .B(\u_inv.d_reg[170] ));
 sg13g2_and2_1 _29091_ (.A(_06475_),
    .B(_06492_),
    .X(_06493_));
 sg13g2_xnor2_1 _29092_ (.Y(_06494_),
    .A(_10908_),
    .B(_06493_));
 sg13g2_nor3_1 _29093_ (.A(_06489_),
    .B(_06491_),
    .C(_06494_),
    .Y(_06495_));
 sg13g2_nand4_1 _29094_ (.B(_06485_),
    .C(_06487_),
    .A(_06477_),
    .Y(_06496_),
    .D(_06495_));
 sg13g2_nor4_1 _29095_ (.A(_06462_),
    .B(_06463_),
    .C(_06465_),
    .D(_06496_),
    .Y(_06497_));
 sg13g2_nand4_1 _29096_ (.B(_06436_),
    .C(_06454_),
    .A(_06427_),
    .Y(_06498_),
    .D(_06497_));
 sg13g2_o21ai_1 _29097_ (.B1(_05907_),
    .Y(_06499_),
    .A1(net4503),
    .A2(_05869_));
 sg13g2_o21ai_1 _29098_ (.B1(net4729),
    .Y(_06500_),
    .A1(\u_inv.d_reg[237] ),
    .A2(\u_inv.d_reg[236] ));
 sg13g2_nor2b_1 _29099_ (.A(_06499_),
    .B_N(_06500_),
    .Y(_06501_));
 sg13g2_o21ai_1 _29100_ (.B1(_06501_),
    .Y(_06502_),
    .A1(net4503),
    .A2(_10886_));
 sg13g2_xnor2_1 _29101_ (.Y(_06503_),
    .A(\u_inv.d_reg[239] ),
    .B(_06502_));
 sg13g2_a21o_1 _29102_ (.A2(_05867_),
    .A1(_05865_),
    .B1(net4504),
    .X(_06504_));
 sg13g2_o21ai_1 _29103_ (.B1(_06504_),
    .Y(_06505_),
    .A1(net4504),
    .A2(_10889_));
 sg13g2_xnor2_1 _29104_ (.Y(_06506_),
    .A(_10888_),
    .B(_06505_));
 sg13g2_o21ai_1 _29105_ (.B1(net4738),
    .Y(_06507_),
    .A1(_05862_),
    .A2(_05863_));
 sg13g2_inv_1 _29106_ (.Y(_06508_),
    .A(_06507_));
 sg13g2_nor3_1 _29107_ (.A(net4769),
    .B(net4770),
    .C(_05862_),
    .Y(_06509_));
 sg13g2_a21oi_1 _29108_ (.A1(_10895_),
    .A2(_06509_),
    .Y(_06510_),
    .B1(_10894_));
 sg13g2_nand2_1 _29109_ (.Y(_06511_),
    .A(net4504),
    .B(\u_inv.d_reg[211] ));
 sg13g2_o21ai_1 _29110_ (.B1(_06511_),
    .Y(_06512_),
    .A1(_06507_),
    .A2(_06510_));
 sg13g2_nand2_1 _29111_ (.Y(_06513_),
    .A(_06506_),
    .B(_06512_));
 sg13g2_nand3_1 _29112_ (.B(_10892_),
    .C(_05865_),
    .A(_10891_),
    .Y(_06514_));
 sg13g2_o21ai_1 _29113_ (.B1(net4737),
    .Y(_06515_),
    .A1(\u_inv.d_reg[218] ),
    .A2(_06514_));
 sg13g2_nand2_1 _29114_ (.Y(_06516_),
    .A(net4737),
    .B(_05866_));
 sg13g2_and2_1 _29115_ (.A(_05942_),
    .B(_06516_),
    .X(_06517_));
 sg13g2_xor2_1 _29116_ (.B(_06515_),
    .A(\u_inv.d_reg[219] ),
    .X(_06518_));
 sg13g2_inv_1 _29117_ (.Y(_06519_),
    .A(_06518_));
 sg13g2_nand2_1 _29118_ (.Y(_06520_),
    .A(net4737),
    .B(_06514_));
 sg13g2_xor2_1 _29119_ (.B(_06520_),
    .A(\u_inv.d_reg[218] ),
    .X(_06521_));
 sg13g2_or2_1 _29120_ (.X(_06522_),
    .B(_06521_),
    .A(_06518_));
 sg13g2_or3_1 _29121_ (.A(\u_inv.d_reg[201] ),
    .B(\u_inv.d_reg[200] ),
    .C(_05918_),
    .X(_06523_));
 sg13g2_o21ai_1 _29122_ (.B1(\u_inv.d_reg[203] ),
    .Y(_06524_),
    .A1(\u_inv.d_reg[202] ),
    .A2(_06523_));
 sg13g2_a22oi_1 _29123_ (.Y(_06525_),
    .B1(_05922_),
    .B2(_06524_),
    .A2(\u_inv.d_reg[203] ),
    .A1(net4506));
 sg13g2_or4_1 _29124_ (.A(_06503_),
    .B(_06513_),
    .C(_06522_),
    .D(_06525_),
    .X(_06526_));
 sg13g2_o21ai_1 _29125_ (.B1(net4733),
    .Y(_06527_),
    .A1(_05868_),
    .A2(_05872_));
 sg13g2_xnor2_1 _29126_ (.Y(_06528_),
    .A(net4768),
    .B(_06527_));
 sg13g2_o21ai_1 _29127_ (.B1(_06517_),
    .Y(_06529_),
    .A1(net4504),
    .A2(_10890_));
 sg13g2_xor2_1 _29128_ (.B(_06529_),
    .A(\u_inv.d_reg[221] ),
    .X(_06530_));
 sg13g2_xnor2_1 _29129_ (.Y(_06531_),
    .A(\u_inv.d_reg[221] ),
    .B(_06529_));
 sg13g2_xnor2_1 _29130_ (.Y(_06532_),
    .A(\u_inv.d_reg[212] ),
    .B(_06507_));
 sg13g2_a21oi_1 _29131_ (.A1(net4738),
    .A2(\u_inv.d_reg[212] ),
    .Y(_06533_),
    .B1(_06508_));
 sg13g2_xnor2_1 _29132_ (.Y(_06534_),
    .A(\u_inv.d_reg[213] ),
    .B(_06533_));
 sg13g2_and2_1 _29133_ (.A(_06532_),
    .B(_06534_),
    .X(_06535_));
 sg13g2_o21ai_1 _29134_ (.B1(_06533_),
    .Y(_06536_),
    .A1(net4504),
    .A2(_10893_));
 sg13g2_xor2_1 _29135_ (.B(_06536_),
    .A(\u_inv.d_reg[214] ),
    .X(_06537_));
 sg13g2_and3_1 _29136_ (.X(_06538_),
    .A(_06530_),
    .B(_06535_),
    .C(_06537_));
 sg13g2_nand2_1 _29137_ (.Y(_06539_),
    .A(net4740),
    .B(_06523_));
 sg13g2_xor2_1 _29138_ (.B(_06539_),
    .A(\u_inv.d_reg[202] ),
    .X(_06540_));
 sg13g2_inv_1 _29139_ (.Y(_06541_),
    .A(_06540_));
 sg13g2_o21ai_1 _29140_ (.B1(net4755),
    .Y(_06542_),
    .A1(\u_inv.d_reg[189] ),
    .A2(\u_inv.d_reg[188] ));
 sg13g2_nand2_1 _29141_ (.Y(_06543_),
    .A(_05946_),
    .B(_06542_));
 sg13g2_xor2_1 _29142_ (.B(_06543_),
    .A(\u_inv.d_reg[190] ),
    .X(_06544_));
 sg13g2_nor2_1 _29143_ (.A(net4505),
    .B(_06509_),
    .Y(_06545_));
 sg13g2_xnor2_1 _29144_ (.Y(_06546_),
    .A(_10895_),
    .B(_06545_));
 sg13g2_a21o_1 _29145_ (.A2(\u_inv.d_reg[196] ),
    .A1(net4742),
    .B1(_06455_),
    .X(_06547_));
 sg13g2_xnor2_1 _29146_ (.Y(_06548_),
    .A(net4772),
    .B(_06547_));
 sg13g2_xnor2_1 _29147_ (.Y(_06549_),
    .A(net4773),
    .B(_06455_));
 sg13g2_nor2_2 _29148_ (.A(_06548_),
    .B(_06549_),
    .Y(_06550_));
 sg13g2_nand4_1 _29149_ (.B(_06544_),
    .C(_06546_),
    .A(_06541_),
    .Y(_06551_),
    .D(_06550_));
 sg13g2_xnor2_1 _29150_ (.Y(_06552_),
    .A(\u_inv.d_reg[220] ),
    .B(_06517_));
 sg13g2_nor3_1 _29151_ (.A(\u_inv.d_reg[178] ),
    .B(_05841_),
    .C(_05849_),
    .Y(_06553_));
 sg13g2_nand2b_1 _29152_ (.Y(_06554_),
    .B(\u_inv.d_reg[179] ),
    .A_N(_06553_));
 sg13g2_a22oi_1 _29153_ (.Y(_06555_),
    .B1(_05925_),
    .B2(_06554_),
    .A2(\u_inv.d_reg[179] ),
    .A1(net4509));
 sg13g2_o21ai_1 _29154_ (.B1(_05984_),
    .Y(_06556_),
    .A1(net4508),
    .A2(_10903_));
 sg13g2_xnor2_1 _29155_ (.Y(_06557_),
    .A(\u_inv.d_reg[183] ),
    .B(_06556_));
 sg13g2_o21ai_1 _29156_ (.B1(_05971_),
    .Y(_06558_),
    .A1(net4509),
    .A2(_10917_));
 sg13g2_xnor2_1 _29157_ (.Y(_06559_),
    .A(\u_inv.d_reg[143] ),
    .B(_06558_));
 sg13g2_o21ai_1 _29158_ (.B1(net4758),
    .Y(_06560_),
    .A1(_05833_),
    .A2(_05935_));
 sg13g2_xnor2_1 _29159_ (.Y(_06561_),
    .A(_10911_),
    .B(_06560_));
 sg13g2_nor4_2 _29160_ (.A(_06555_),
    .B(_06557_),
    .C(_06559_),
    .Y(_06562_),
    .D(_06561_));
 sg13g2_a21oi_1 _29161_ (.A1(_10892_),
    .A2(_05865_),
    .Y(_06563_),
    .B1(net4504));
 sg13g2_xnor2_1 _29162_ (.Y(_06564_),
    .A(_10891_),
    .B(_06563_));
 sg13g2_a21oi_1 _29163_ (.A1(_05857_),
    .A2(_05921_),
    .Y(_06565_),
    .B1(net4506));
 sg13g2_xor2_1 _29164_ (.B(_06565_),
    .A(\u_inv.d_reg[206] ),
    .X(_06566_));
 sg13g2_nand4_1 _29165_ (.B(_06562_),
    .C(_06564_),
    .A(_06552_),
    .Y(_06567_),
    .D(_06566_));
 sg13g2_o21ai_1 _29166_ (.B1(net4733),
    .Y(_06568_),
    .A1(\u_inv.d_reg[224] ),
    .A2(_05868_));
 sg13g2_xnor2_1 _29167_ (.Y(_06569_),
    .A(\u_inv.d_reg[225] ),
    .B(_06568_));
 sg13g2_xnor2_1 _29168_ (.Y(_06570_),
    .A(_10889_),
    .B(_06504_));
 sg13g2_a21oi_1 _29169_ (.A1(net4740),
    .A2(_05858_),
    .Y(_06571_),
    .B1(_05922_));
 sg13g2_xor2_1 _29170_ (.B(_06571_),
    .A(\u_inv.d_reg[207] ),
    .X(_06572_));
 sg13g2_a21o_1 _29171_ (.A2(\u_inv.d_reg[204] ),
    .A1(net4740),
    .B1(_05922_),
    .X(_06573_));
 sg13g2_xnor2_1 _29172_ (.Y(_06574_),
    .A(\u_inv.d_reg[205] ),
    .B(_06573_));
 sg13g2_a21oi_1 _29173_ (.A1(_10911_),
    .A2(_06560_),
    .Y(_06575_),
    .B1(net4508));
 sg13g2_xnor2_1 _29174_ (.Y(_06576_),
    .A(\u_inv.d_reg[167] ),
    .B(_06575_));
 sg13g2_nor4_1 _29175_ (.A(_06570_),
    .B(_06572_),
    .C(_06574_),
    .D(_06576_),
    .Y(_06577_));
 sg13g2_nand2_1 _29176_ (.Y(_06578_),
    .A(_06569_),
    .B(_06577_));
 sg13g2_nor3_1 _29177_ (.A(_06551_),
    .B(_06567_),
    .C(_06578_),
    .Y(_06579_));
 sg13g2_nand3_1 _29178_ (.B(_06538_),
    .C(_06579_),
    .A(_06528_),
    .Y(_06580_));
 sg13g2_nor4_2 _29179_ (.A(_05953_),
    .B(_06498_),
    .C(_06526_),
    .Y(_06581_),
    .D(_06580_));
 sg13g2_o21ai_1 _29180_ (.B1(net4737),
    .Y(_06582_),
    .A1(\u_inv.d_reg[214] ),
    .A2(_06536_));
 sg13g2_xor2_1 _29181_ (.B(_06582_),
    .A(\u_inv.d_reg[215] ),
    .X(_06583_));
 sg13g2_xnor2_1 _29182_ (.Y(_06584_),
    .A(\u_inv.d_reg[246] ),
    .B(_05903_));
 sg13g2_inv_2 _29183_ (.Y(_06585_),
    .A(_06584_));
 sg13g2_o21ai_1 _29184_ (.B1(net4731),
    .Y(_06586_),
    .A1(_05877_),
    .A2(_05878_));
 sg13g2_xor2_1 _29185_ (.B(_06586_),
    .A(\u_inv.d_reg[242] ),
    .X(_06587_));
 sg13g2_or3_1 _29186_ (.A(net4768),
    .B(_05868_),
    .C(_05872_),
    .X(_06588_));
 sg13g2_a21oi_1 _29187_ (.A1(\u_inv.d_reg[227] ),
    .A2(_06588_),
    .Y(_06589_),
    .B1(_05896_));
 sg13g2_a21oi_2 _29188_ (.B1(_06589_),
    .Y(_06590_),
    .A2(\u_inv.d_reg[227] ),
    .A1(net4505));
 sg13g2_xnor2_1 _29189_ (.Y(_06591_),
    .A(\u_inv.d_reg[236] ),
    .B(_06499_));
 sg13g2_xor2_1 _29190_ (.B(_05898_),
    .A(\u_inv.d_reg[230] ),
    .X(_06592_));
 sg13g2_or4_1 _29191_ (.A(\u_inv.d_reg[233] ),
    .B(\u_inv.d_reg[232] ),
    .C(_05868_),
    .D(_05876_),
    .X(_06593_));
 sg13g2_nand2_1 _29192_ (.Y(_06594_),
    .A(net4729),
    .B(_06593_));
 sg13g2_xor2_1 _29193_ (.B(_06594_),
    .A(\u_inv.d_reg[234] ),
    .X(_06595_));
 sg13g2_or4_1 _29194_ (.A(_06590_),
    .B(_06591_),
    .C(_06592_),
    .D(_06595_),
    .X(_06596_));
 sg13g2_nor4_1 _29195_ (.A(_06583_),
    .B(_06585_),
    .C(_06587_),
    .D(_06596_),
    .Y(_06597_));
 sg13g2_a21o_2 _29196_ (.A2(_05879_),
    .A1(net4731),
    .B1(_05902_),
    .X(_06598_));
 sg13g2_a21oi_1 _29197_ (.A1(net4731),
    .A2(\u_inv.d_reg[244] ),
    .Y(_06599_),
    .B1(_06598_));
 sg13g2_xnor2_1 _29198_ (.Y(_06600_),
    .A(\u_inv.d_reg[245] ),
    .B(_06599_));
 sg13g2_xnor2_1 _29199_ (.Y(_06601_),
    .A(\u_inv.d_reg[244] ),
    .B(_06598_));
 sg13g2_nand2b_1 _29200_ (.Y(_06602_),
    .B(_06600_),
    .A_N(_06601_));
 sg13g2_a21oi_1 _29201_ (.A1(net4729),
    .A2(\u_inv.d_reg[236] ),
    .Y(_06603_),
    .B1(_06499_));
 sg13g2_xor2_1 _29202_ (.B(_06603_),
    .A(\u_inv.d_reg[237] ),
    .X(_06604_));
 sg13g2_xnor2_1 _29203_ (.Y(_06605_),
    .A(_10886_),
    .B(_06501_));
 sg13g2_o21ai_1 _29204_ (.B1(\u_inv.d_reg[235] ),
    .Y(_06606_),
    .A1(\u_inv.d_reg[234] ),
    .A2(_06593_));
 sg13g2_a22oi_1 _29205_ (.Y(_06607_),
    .B1(_06499_),
    .B2(_06606_),
    .A2(\u_inv.d_reg[235] ),
    .A1(net4503));
 sg13g2_inv_1 _29206_ (.Y(_06608_),
    .A(_06607_));
 sg13g2_nor4_1 _29207_ (.A(_06602_),
    .B(_06604_),
    .C(_06605_),
    .D(_06607_),
    .Y(_06609_));
 sg13g2_nor3_1 _29208_ (.A(\u_inv.d_reg[242] ),
    .B(_05877_),
    .C(_05878_),
    .Y(_06610_));
 sg13g2_nand2b_1 _29209_ (.Y(_06611_),
    .B(\u_inv.d_reg[243] ),
    .A_N(_06610_));
 sg13g2_a22oi_1 _29210_ (.Y(_06612_),
    .B1(_06598_),
    .B2(_06611_),
    .A2(\u_inv.d_reg[243] ),
    .A1(net4503));
 sg13g2_nand2_1 _29211_ (.Y(_06613_),
    .A(net4733),
    .B(net4767));
 sg13g2_and2_1 _29212_ (.A(_05896_),
    .B(_06613_),
    .X(_06614_));
 sg13g2_xnor2_1 _29213_ (.Y(_06615_),
    .A(net4766),
    .B(_06614_));
 sg13g2_xor2_1 _29214_ (.B(_06614_),
    .A(net4766),
    .X(_06616_));
 sg13g2_xor2_1 _29215_ (.B(_05896_),
    .A(net4767),
    .X(_06617_));
 sg13g2_nor2_2 _29216_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sg13g2_inv_1 _29217_ (.Y(_06619_),
    .A(_06618_));
 sg13g2_xor2_1 _29218_ (.B(_05902_),
    .A(\u_inv.d_reg[240] ),
    .X(_06620_));
 sg13g2_o21ai_1 _29219_ (.B1(net4731),
    .Y(_06621_),
    .A1(\u_inv.d_reg[240] ),
    .A2(_05877_));
 sg13g2_xnor2_1 _29220_ (.Y(_06622_),
    .A(\u_inv.d_reg[241] ),
    .B(_06621_));
 sg13g2_nand2_1 _29221_ (.Y(_06623_),
    .A(_06620_),
    .B(_06622_));
 sg13g2_xnor2_1 _29222_ (.Y(_06624_),
    .A(_10884_),
    .B(_05884_));
 sg13g2_nor4_1 _29223_ (.A(_06612_),
    .B(_06619_),
    .C(_06623_),
    .D(_06624_),
    .Y(_06625_));
 sg13g2_nand4_1 _29224_ (.B(_06597_),
    .C(_06609_),
    .A(_06581_),
    .Y(_06626_),
    .D(_06625_));
 sg13g2_o21ai_1 _29225_ (.B1(net4727),
    .Y(_06627_),
    .A1(\u_inv.d_reg[254] ),
    .A2(_05886_));
 sg13g2_xor2_1 _29226_ (.B(_06627_),
    .A(\u_inv.d_reg[255] ),
    .X(_06628_));
 sg13g2_o21ai_1 _29227_ (.B1(net4727),
    .Y(_06629_),
    .A1(\u_inv.d_reg[249] ),
    .A2(_05891_));
 sg13g2_xnor2_1 _29228_ (.Y(_06630_),
    .A(\u_inv.d_reg[250] ),
    .B(_06629_));
 sg13g2_nand2_1 _29229_ (.Y(_06631_),
    .A(net4727),
    .B(_05891_));
 sg13g2_xor2_1 _29230_ (.B(_06631_),
    .A(\u_inv.d_reg[249] ),
    .X(_06632_));
 sg13g2_xnor2_1 _29231_ (.Y(_06633_),
    .A(\u_inv.d_reg[248] ),
    .B(_05883_));
 sg13g2_nor2_1 _29232_ (.A(_06632_),
    .B(_06633_),
    .Y(_06634_));
 sg13g2_xor2_1 _29233_ (.B(_05886_),
    .A(\u_inv.d_reg[254] ),
    .X(_06635_));
 sg13g2_o21ai_1 _29234_ (.B1(_05884_),
    .Y(_06636_),
    .A1(net4501),
    .A2(_10884_));
 sg13g2_xnor2_1 _29235_ (.Y(_06637_),
    .A(\u_inv.d_reg[253] ),
    .B(_06636_));
 sg13g2_inv_1 _29236_ (.Y(_06638_),
    .A(_06637_));
 sg13g2_nand4_1 _29237_ (.B(_06634_),
    .C(_06635_),
    .A(_06630_),
    .Y(_06639_),
    .D(_06638_));
 sg13g2_nor4_2 _29238_ (.A(_05914_),
    .B(_06626_),
    .C(_06628_),
    .Y(_06640_),
    .D(_06639_));
 sg13g2_inv_1 _29239_ (.Y(_06641_),
    .A(net3332));
 sg13g2_nor2_1 _29240_ (.A(net3353),
    .B(net3338),
    .Y(_06642_));
 sg13g2_nand2b_2 _29241_ (.Y(_06643_),
    .B(net3379),
    .A_N(net3334));
 sg13g2_xnor2_1 _29242_ (.Y(_06644_),
    .A(net4800),
    .B(net3310));
 sg13g2_nor2_1 _29243_ (.A(net1427),
    .B(net4174),
    .Y(_06645_));
 sg13g2_a21oi_1 _29244_ (.A1(net4174),
    .A2(_06644_),
    .Y(_01048_),
    .B1(_06645_));
 sg13g2_a21oi_1 _29245_ (.A1(_06159_),
    .A2(_06160_),
    .Y(_06646_),
    .B1(net3310));
 sg13g2_o21ai_1 _29246_ (.B1(_06161_),
    .Y(_06647_),
    .A1(net4798),
    .A2(net4800));
 sg13g2_nor2_1 _29247_ (.A(net3345),
    .B(_06647_),
    .Y(_06648_));
 sg13g2_a21oi_1 _29248_ (.A1(net3331),
    .A2(_06647_),
    .Y(_06649_),
    .B1(_06648_));
 sg13g2_nor3_1 _29249_ (.A(net4145),
    .B(_06646_),
    .C(_06649_),
    .Y(_06650_));
 sg13g2_a21o_1 _29250_ (.A2(net4145),
    .A1(net1548),
    .B1(_06650_),
    .X(_01049_));
 sg13g2_a22oi_1 _29251_ (.Y(_06651_),
    .B1(_06162_),
    .B2(net3332),
    .A2(_06158_),
    .A1(net3376));
 sg13g2_a21oi_1 _29252_ (.A1(_06163_),
    .A2(net3332),
    .Y(_06652_),
    .B1(_06651_));
 sg13g2_o21ai_1 _29253_ (.B1(_06158_),
    .Y(_06653_),
    .A1(net4798),
    .A2(net4800));
 sg13g2_a21oi_1 _29254_ (.A1(_05719_),
    .A2(_06653_),
    .Y(_06654_),
    .B1(net3376));
 sg13g2_nor3_1 _29255_ (.A(net4145),
    .B(_06652_),
    .C(_06654_),
    .Y(_06655_));
 sg13g2_a21oi_1 _29256_ (.A1(_10985_),
    .A2(net4146),
    .Y(_01050_),
    .B1(_06655_));
 sg13g2_a21oi_1 _29257_ (.A1(_06163_),
    .A2(net3332),
    .Y(_06656_),
    .B1(_06155_));
 sg13g2_a21oi_1 _29258_ (.A1(_06164_),
    .A2(net3332),
    .Y(_06657_),
    .B1(net3345));
 sg13g2_nand2b_1 _29259_ (.Y(_06658_),
    .B(_06657_),
    .A_N(_06656_));
 sg13g2_nand2_1 _29260_ (.Y(_06659_),
    .A(_05719_),
    .B(_06155_));
 sg13g2_nand2_1 _29261_ (.Y(_06660_),
    .A(_05720_),
    .B(_06659_));
 sg13g2_a21oi_1 _29262_ (.A1(net3345),
    .A2(_06660_),
    .Y(_06661_),
    .B1(net4145));
 sg13g2_a22oi_1 _29263_ (.Y(_01051_),
    .B1(_06658_),
    .B2(_06661_),
    .A2(net4145),
    .A1(_10986_));
 sg13g2_nor2_1 _29264_ (.A(_06164_),
    .B(net3331),
    .Y(_06662_));
 sg13g2_a21oi_1 _29265_ (.A1(_06166_),
    .A2(_06662_),
    .Y(_06663_),
    .B1(net3345));
 sg13g2_o21ai_1 _29266_ (.B1(_06663_),
    .Y(_06664_),
    .A1(_06166_),
    .A2(_06662_));
 sg13g2_a21oi_1 _29267_ (.A1(_05720_),
    .A2(_06166_),
    .Y(_06665_),
    .B1(net3376));
 sg13g2_a21oi_1 _29268_ (.A1(_05721_),
    .A2(_06665_),
    .Y(_06666_),
    .B1(net4145));
 sg13g2_a22oi_1 _29269_ (.Y(_01052_),
    .B1(_06664_),
    .B2(_06666_),
    .A2(net4145),
    .A1(_10987_));
 sg13g2_a21oi_1 _29270_ (.A1(_06167_),
    .A2(net3332),
    .Y(_06667_),
    .B1(_06665_));
 sg13g2_xnor2_1 _29271_ (.Y(_06668_),
    .A(_06169_),
    .B(_06667_));
 sg13g2_mux2_1 _29272_ (.A0(net2070),
    .A1(_06668_),
    .S(net4174),
    .X(_01053_));
 sg13g2_nor2_1 _29273_ (.A(net1426),
    .B(net4174),
    .Y(_06669_));
 sg13g2_nand2_1 _29274_ (.Y(_06670_),
    .A(_06170_),
    .B(net3332));
 sg13g2_a21oi_1 _29275_ (.A1(_05720_),
    .A2(_06166_),
    .Y(_06671_),
    .B1(_06169_));
 sg13g2_o21ai_1 _29276_ (.B1(_06670_),
    .Y(_06672_),
    .A1(net3376),
    .A2(_06671_));
 sg13g2_xor2_1 _29277_ (.B(_06672_),
    .A(net1451),
    .X(_06673_));
 sg13g2_a21oi_1 _29278_ (.A1(net4175),
    .A2(_06673_),
    .Y(_01054_),
    .B1(_06669_));
 sg13g2_or2_1 _29279_ (.X(_06674_),
    .B(_06671_),
    .A(_06172_));
 sg13g2_nor2_1 _29280_ (.A(net3376),
    .B(_06674_),
    .Y(_06675_));
 sg13g2_a21oi_1 _29281_ (.A1(_06173_),
    .A2(net3332),
    .Y(_06676_),
    .B1(_06675_));
 sg13g2_xnor2_1 _29282_ (.Y(_06677_),
    .A(_06175_),
    .B(_06676_));
 sg13g2_nand2_1 _29283_ (.Y(_06678_),
    .A(net1117),
    .B(net4146));
 sg13g2_o21ai_1 _29284_ (.B1(_06678_),
    .Y(_01055_),
    .A1(net4145),
    .A2(_06677_));
 sg13g2_nor2_1 _29285_ (.A(net1547),
    .B(net4174),
    .Y(_06679_));
 sg13g2_nor2_1 _29286_ (.A(_06175_),
    .B(_06674_),
    .Y(_06680_));
 sg13g2_nand2_1 _29287_ (.Y(_06681_),
    .A(net3345),
    .B(_06680_));
 sg13g2_nand3_1 _29288_ (.B(_06175_),
    .C(net3333),
    .A(_06173_),
    .Y(_06682_));
 sg13g2_nand2_1 _29289_ (.Y(_06683_),
    .A(_06681_),
    .B(_06682_));
 sg13g2_xnor2_1 _29290_ (.Y(_06684_),
    .A(_06152_),
    .B(_06683_));
 sg13g2_a21oi_1 _29291_ (.A1(net4175),
    .A2(_06684_),
    .Y(_01056_),
    .B1(_06679_));
 sg13g2_nor2_1 _29292_ (.A(net1206),
    .B(net4174),
    .Y(_06685_));
 sg13g2_nor4_1 _29293_ (.A(_06151_),
    .B(_06172_),
    .C(_06175_),
    .D(_06671_),
    .Y(_06686_));
 sg13g2_nand2_1 _29294_ (.Y(_06687_),
    .A(_06152_),
    .B(_06680_));
 sg13g2_a22oi_1 _29295_ (.Y(_06688_),
    .B1(_06682_),
    .B2(_06687_),
    .A2(_06152_),
    .A1(net3376));
 sg13g2_xnor2_1 _29296_ (.Y(_06689_),
    .A(_06148_),
    .B(_06688_));
 sg13g2_a21oi_1 _29297_ (.A1(net4174),
    .A2(_06689_),
    .Y(_01057_),
    .B1(_06685_));
 sg13g2_nor2_1 _29298_ (.A(net1677),
    .B(net4176),
    .Y(_06690_));
 sg13g2_nor2_1 _29299_ (.A(_06149_),
    .B(_06687_),
    .Y(_06691_));
 sg13g2_a21o_1 _29300_ (.A2(_06176_),
    .A1(net3376),
    .B1(net3318),
    .X(_06692_));
 sg13g2_a21oi_1 _29301_ (.A1(net3345),
    .A2(_06691_),
    .Y(_06693_),
    .B1(_06692_));
 sg13g2_xnor2_1 _29302_ (.Y(_06694_),
    .A(_06178_),
    .B(_06693_));
 sg13g2_a21oi_1 _29303_ (.A1(net4176),
    .A2(_06694_),
    .Y(_01058_),
    .B1(_06690_));
 sg13g2_nor2_1 _29304_ (.A(net1518),
    .B(net4174),
    .Y(_06695_));
 sg13g2_nor2_1 _29305_ (.A(_06178_),
    .B(_06691_),
    .Y(_06696_));
 sg13g2_nor2_1 _29306_ (.A(net3377),
    .B(_06696_),
    .Y(_06697_));
 sg13g2_nor2_1 _29307_ (.A(net3345),
    .B(_06178_),
    .Y(_06698_));
 sg13g2_nor3_1 _29308_ (.A(_06692_),
    .B(_06697_),
    .C(_06698_),
    .Y(_06699_));
 sg13g2_xor2_1 _29309_ (.B(_06699_),
    .A(_06146_),
    .X(_06700_));
 sg13g2_a21oi_1 _29310_ (.A1(net4175),
    .A2(_06700_),
    .Y(_01059_),
    .B1(_06695_));
 sg13g2_nor2_1 _29311_ (.A(net2089),
    .B(net4176),
    .Y(_06701_));
 sg13g2_a221oi_1 _29312_ (.B2(_06686_),
    .C1(_06178_),
    .B1(_06148_),
    .A1(_06144_),
    .Y(_06702_),
    .A2(_06145_));
 sg13g2_nand2_1 _29313_ (.Y(_06703_),
    .A(_06146_),
    .B(_06696_));
 sg13g2_nand2b_1 _29314_ (.Y(_06704_),
    .B(net3333),
    .A_N(_06180_));
 sg13g2_o21ai_1 _29315_ (.B1(_06704_),
    .Y(_06705_),
    .A1(net3377),
    .A2(_06703_));
 sg13g2_xor2_1 _29316_ (.B(_06705_),
    .A(_06182_),
    .X(_06706_));
 sg13g2_a21oi_1 _29317_ (.A1(net4176),
    .A2(_06706_),
    .Y(_01060_),
    .B1(_06701_));
 sg13g2_nor2_1 _29318_ (.A(net1646),
    .B(net4176),
    .Y(_06707_));
 sg13g2_and2_1 _29319_ (.A(_06182_),
    .B(_06702_),
    .X(_06708_));
 sg13g2_nand2_1 _29320_ (.Y(_06709_),
    .A(_06182_),
    .B(_06702_));
 sg13g2_a22oi_1 _29321_ (.Y(_06710_),
    .B1(_06704_),
    .B2(_06709_),
    .A2(_06182_),
    .A1(net3377));
 sg13g2_xor2_1 _29322_ (.B(_06710_),
    .A(_06142_),
    .X(_06711_));
 sg13g2_a21oi_1 _29323_ (.A1(net4176),
    .A2(_06711_),
    .Y(_01061_),
    .B1(_06707_));
 sg13g2_nor2_1 _29324_ (.A(net1734),
    .B(net4177),
    .Y(_06712_));
 sg13g2_nand3_1 _29325_ (.B(_06142_),
    .C(_06708_),
    .A(net3345),
    .Y(_06713_));
 sg13g2_or4_1 _29326_ (.A(_06142_),
    .B(_06180_),
    .C(_06182_),
    .D(net3331),
    .X(_06714_));
 sg13g2_nand2_1 _29327_ (.Y(_06715_),
    .A(_06713_),
    .B(_06714_));
 sg13g2_xor2_1 _29328_ (.B(_06715_),
    .A(_06140_),
    .X(_06716_));
 sg13g2_a21oi_1 _29329_ (.A1(net4176),
    .A2(_06716_),
    .Y(_01062_),
    .B1(_06712_));
 sg13g2_nor2_1 _29330_ (.A(net1560),
    .B(net4177),
    .Y(_06717_));
 sg13g2_and4_1 _29331_ (.A(_06140_),
    .B(_06142_),
    .C(_06182_),
    .D(_06702_),
    .X(_06718_));
 sg13g2_nand3_1 _29332_ (.B(_06142_),
    .C(_06708_),
    .A(_06140_),
    .Y(_06719_));
 sg13g2_a22oi_1 _29333_ (.Y(_06720_),
    .B1(_06714_),
    .B2(_06719_),
    .A2(_06140_),
    .A1(net3377));
 sg13g2_xnor2_1 _29334_ (.Y(_06721_),
    .A(_06137_),
    .B(_06720_));
 sg13g2_a21oi_1 _29335_ (.A1(net4176),
    .A2(_06721_),
    .Y(_01063_),
    .B1(_06717_));
 sg13g2_nor2_1 _29336_ (.A(net1453),
    .B(net4177),
    .Y(_06722_));
 sg13g2_nor2_1 _29337_ (.A(_06137_),
    .B(_06719_),
    .Y(_06723_));
 sg13g2_nand2_1 _29338_ (.Y(_06724_),
    .A(net3346),
    .B(_06723_));
 sg13g2_nand2_1 _29339_ (.Y(_06725_),
    .A(_06184_),
    .B(net3333));
 sg13g2_nand2_1 _29340_ (.Y(_06726_),
    .A(_06724_),
    .B(_06725_));
 sg13g2_xor2_1 _29341_ (.B(_06726_),
    .A(_06131_),
    .X(_06727_));
 sg13g2_a21oi_1 _29342_ (.A1(net4177),
    .A2(_06727_),
    .Y(_01064_),
    .B1(_06722_));
 sg13g2_o21ai_1 _29343_ (.B1(_06133_),
    .Y(_06728_),
    .A1(_06131_),
    .A2(_06725_));
 sg13g2_nand3_1 _29344_ (.B(_06184_),
    .C(net3333),
    .A(_06134_),
    .Y(_06729_));
 sg13g2_nand2_1 _29345_ (.Y(_06730_),
    .A(_06728_),
    .B(_06729_));
 sg13g2_and4_1 _29346_ (.A(_06131_),
    .B(_06133_),
    .C(_06138_),
    .D(_06718_),
    .X(_06731_));
 sg13g2_nor2_1 _29347_ (.A(net3377),
    .B(_06731_),
    .Y(_06732_));
 sg13g2_a21o_1 _29348_ (.A2(_06723_),
    .A1(_06131_),
    .B1(_06133_),
    .X(_06733_));
 sg13g2_a221oi_1 _29349_ (.B2(_06733_),
    .C1(net4146),
    .B1(_06732_),
    .A1(net3376),
    .Y(_06734_),
    .A2(_06730_));
 sg13g2_a21o_1 _29350_ (.A2(net4146),
    .A1(net2063),
    .B1(_06734_),
    .X(_01065_));
 sg13g2_nor2_1 _29351_ (.A(net1647),
    .B(net4177),
    .Y(_06735_));
 sg13g2_a21oi_1 _29352_ (.A1(net3380),
    .A2(_06729_),
    .Y(_06736_),
    .B1(_06732_));
 sg13g2_xor2_1 _29353_ (.B(_06736_),
    .A(_06129_),
    .X(_06737_));
 sg13g2_a21oi_1 _29354_ (.A1(net4177),
    .A2(_06737_),
    .Y(_01066_),
    .B1(_06735_));
 sg13g2_nor2_1 _29355_ (.A(net1668),
    .B(net4180),
    .Y(_06738_));
 sg13g2_nand3_1 _29356_ (.B(_06129_),
    .C(_06731_),
    .A(net3351),
    .Y(_06739_));
 sg13g2_o21ai_1 _29357_ (.B1(_06739_),
    .Y(_06740_),
    .A1(_06135_),
    .A2(_06725_));
 sg13g2_xor2_1 _29358_ (.B(_06740_),
    .A(_06186_),
    .X(_06741_));
 sg13g2_a21oi_1 _29359_ (.A1(net4177),
    .A2(_06741_),
    .Y(_01067_),
    .B1(_06738_));
 sg13g2_nor2_1 _29360_ (.A(net1342),
    .B(net4182),
    .Y(_06742_));
 sg13g2_nand3_1 _29361_ (.B(_06186_),
    .C(_06731_),
    .A(_06129_),
    .Y(_06743_));
 sg13g2_a21oi_1 _29362_ (.A1(_06189_),
    .A2(net3334),
    .Y(_06744_),
    .B1(net3348));
 sg13g2_a21oi_1 _29363_ (.A1(net3348),
    .A2(_06743_),
    .Y(_06745_),
    .B1(_06744_));
 sg13g2_xnor2_1 _29364_ (.Y(_06746_),
    .A(_06126_),
    .B(_06745_));
 sg13g2_a21oi_1 _29365_ (.A1(net4182),
    .A2(_06746_),
    .Y(_01068_),
    .B1(_06742_));
 sg13g2_nor2b_1 _29366_ (.A(_06124_),
    .B_N(_06744_),
    .Y(_06747_));
 sg13g2_nand2b_2 _29367_ (.Y(_06748_),
    .B(_06125_),
    .A_N(_06124_));
 sg13g2_nand4_1 _29368_ (.B(_06126_),
    .C(_06189_),
    .A(_06124_),
    .Y(_06749_),
    .D(net3334));
 sg13g2_a21oi_1 _29369_ (.A1(_06748_),
    .A2(_06749_),
    .Y(_06750_),
    .B1(net3349));
 sg13g2_o21ai_1 _29370_ (.B1(net3349),
    .Y(_06751_),
    .A1(_06743_),
    .A2(_06748_));
 sg13g2_nand2_1 _29371_ (.Y(_06752_),
    .A(_06124_),
    .B(_06743_));
 sg13g2_nand2_1 _29372_ (.Y(_06753_),
    .A(_06127_),
    .B(_06752_));
 sg13g2_o21ai_1 _29373_ (.B1(net4182),
    .Y(_06754_),
    .A1(_06751_),
    .A2(_06753_));
 sg13g2_nor3_1 _29374_ (.A(_06747_),
    .B(_06750_),
    .C(_06754_),
    .Y(_06755_));
 sg13g2_a21o_1 _29375_ (.A2(net4148),
    .A1(net1701),
    .B1(_06755_),
    .X(_01069_));
 sg13g2_nor2_1 _29376_ (.A(net1552),
    .B(net4182),
    .Y(_06756_));
 sg13g2_nand2_1 _29377_ (.Y(_06757_),
    .A(net3379),
    .B(_06749_));
 sg13g2_and2_1 _29378_ (.A(_06751_),
    .B(_06757_),
    .X(_06758_));
 sg13g2_xor2_1 _29379_ (.B(_06758_),
    .A(_06120_),
    .X(_06759_));
 sg13g2_a21oi_1 _29380_ (.A1(net4182),
    .A2(_06759_),
    .Y(_01070_),
    .B1(_06756_));
 sg13g2_nor2_1 _29381_ (.A(net1321),
    .B(net4182),
    .Y(_06760_));
 sg13g2_xnor2_1 _29382_ (.Y(_06761_),
    .A(net3349),
    .B(_06120_));
 sg13g2_nand2_1 _29383_ (.Y(_06762_),
    .A(_06758_),
    .B(_06761_));
 sg13g2_xnor2_1 _29384_ (.Y(_06763_),
    .A(_06119_),
    .B(_06762_));
 sg13g2_a21oi_1 _29385_ (.A1(net4182),
    .A2(_06763_),
    .Y(_01071_),
    .B1(_06760_));
 sg13g2_nor2_1 _29386_ (.A(net2174),
    .B(net4183),
    .Y(_06764_));
 sg13g2_nand2_1 _29387_ (.Y(_06765_),
    .A(_06119_),
    .B(_06120_));
 sg13g2_nor3_1 _29388_ (.A(_06743_),
    .B(_06748_),
    .C(_06765_),
    .Y(_06766_));
 sg13g2_nor2_1 _29389_ (.A(_06121_),
    .B(_06749_),
    .Y(_06767_));
 sg13g2_a21oi_1 _29390_ (.A1(net3349),
    .A2(_06766_),
    .Y(_06768_),
    .B1(_06767_));
 sg13g2_xnor2_1 _29391_ (.Y(_06769_),
    .A(_06115_),
    .B(_06768_));
 sg13g2_a21oi_1 _29392_ (.A1(net4182),
    .A2(_06769_),
    .Y(_01072_),
    .B1(_06764_));
 sg13g2_o21ai_1 _29393_ (.B1(_06113_),
    .Y(_06770_),
    .A1(_06121_),
    .A2(_06749_));
 sg13g2_nand2_1 _29394_ (.Y(_06771_),
    .A(_06113_),
    .B(_06115_));
 sg13g2_nand2b_1 _29395_ (.Y(_06772_),
    .B(net3334),
    .A_N(_06191_));
 sg13g2_nand3_1 _29396_ (.B(_06771_),
    .C(_06772_),
    .A(_06770_),
    .Y(_06773_));
 sg13g2_nor4_2 _29397_ (.A(_06743_),
    .B(_06748_),
    .C(_06765_),
    .Y(_06774_),
    .D(_06771_));
 sg13g2_nor2_1 _29398_ (.A(net3379),
    .B(_06774_),
    .Y(_06775_));
 sg13g2_a21o_1 _29399_ (.A2(_06766_),
    .A1(_06115_),
    .B1(_06113_),
    .X(_06776_));
 sg13g2_a221oi_1 _29400_ (.B2(_06776_),
    .C1(net4149),
    .B1(_06775_),
    .A1(net3379),
    .Y(_06777_),
    .A2(_06773_));
 sg13g2_a21o_1 _29401_ (.A2(net4149),
    .A1(net2416),
    .B1(_06777_),
    .X(_01073_));
 sg13g2_nor2_1 _29402_ (.A(net1883),
    .B(net4185),
    .Y(_06778_));
 sg13g2_a21oi_1 _29403_ (.A1(net3379),
    .A2(_06772_),
    .Y(_06779_),
    .B1(_06775_));
 sg13g2_xor2_1 _29404_ (.B(_06779_),
    .A(_06111_),
    .X(_06780_));
 sg13g2_a21oi_1 _29405_ (.A1(net4185),
    .A2(_06780_),
    .Y(_01074_),
    .B1(_06778_));
 sg13g2_a21oi_1 _29406_ (.A1(_06192_),
    .A2(net3334),
    .Y(_06781_),
    .B1(_06109_));
 sg13g2_nor2_1 _29407_ (.A(net3350),
    .B(_06781_),
    .Y(_06782_));
 sg13g2_nand3_1 _29408_ (.B(_06192_),
    .C(net3334),
    .A(_06109_),
    .Y(_06783_));
 sg13g2_nand3_1 _29409_ (.B(_06111_),
    .C(_06774_),
    .A(_06109_),
    .Y(_06784_));
 sg13g2_a21o_1 _29410_ (.A2(_06774_),
    .A1(_06111_),
    .B1(_06109_),
    .X(_06785_));
 sg13g2_and2_1 _29411_ (.A(_06784_),
    .B(_06785_),
    .X(_06786_));
 sg13g2_a221oi_1 _29412_ (.B2(net3350),
    .C1(net4149),
    .B1(_06786_),
    .A1(_06782_),
    .Y(_06787_),
    .A2(_06783_));
 sg13g2_a21o_1 _29413_ (.A2(net4149),
    .A1(net2371),
    .B1(_06787_),
    .X(_01075_));
 sg13g2_nor2_1 _29414_ (.A(net2229),
    .B(net4185),
    .Y(_06788_));
 sg13g2_nor2_1 _29415_ (.A(_06194_),
    .B(net3331),
    .Y(_06789_));
 sg13g2_nand2_1 _29416_ (.Y(_06790_),
    .A(_06193_),
    .B(net3335));
 sg13g2_o21ai_1 _29417_ (.B1(_06790_),
    .Y(_06791_),
    .A1(net3379),
    .A2(_06784_));
 sg13g2_xor2_1 _29418_ (.B(_06791_),
    .A(_06098_),
    .X(_06792_));
 sg13g2_a21oi_1 _29419_ (.A1(net4184),
    .A2(_06792_),
    .Y(_01076_),
    .B1(_06788_));
 sg13g2_nor2_1 _29420_ (.A(net2050),
    .B(net4185),
    .Y(_06793_));
 sg13g2_nand4_1 _29421_ (.B(_06109_),
    .C(_06111_),
    .A(_06098_),
    .Y(_06794_),
    .D(_06774_));
 sg13g2_a22oi_1 _29422_ (.Y(_06795_),
    .B1(_06790_),
    .B2(_06794_),
    .A2(_06098_),
    .A1(net3380));
 sg13g2_xnor2_1 _29423_ (.Y(_06796_),
    .A(_06100_),
    .B(_06795_));
 sg13g2_a21oi_1 _29424_ (.A1(net4184),
    .A2(_06796_),
    .Y(_01077_),
    .B1(_06793_));
 sg13g2_nor2_1 _29425_ (.A(net2043),
    .B(net4184),
    .Y(_06797_));
 sg13g2_nor2_1 _29426_ (.A(_06100_),
    .B(_06794_),
    .Y(_06798_));
 sg13g2_a22oi_1 _29427_ (.Y(_06799_),
    .B1(_06798_),
    .B2(net3350),
    .A2(_06789_),
    .A1(_06101_));
 sg13g2_xnor2_1 _29428_ (.Y(_06800_),
    .A(_06106_),
    .B(_06799_));
 sg13g2_a21oi_1 _29429_ (.A1(net4184),
    .A2(_06800_),
    .Y(_01078_),
    .B1(_06797_));
 sg13g2_nor2_1 _29430_ (.A(net2095),
    .B(net4184),
    .Y(_06801_));
 sg13g2_a22oi_1 _29431_ (.Y(_06802_),
    .B1(_06798_),
    .B2(_06106_),
    .A2(_06789_),
    .A1(_06101_));
 sg13g2_a21oi_1 _29432_ (.A1(net3380),
    .A2(_06106_),
    .Y(_06803_),
    .B1(_06802_));
 sg13g2_xnor2_1 _29433_ (.Y(_06804_),
    .A(_06104_),
    .B(_06803_));
 sg13g2_a21oi_1 _29434_ (.A1(net4184),
    .A2(_06804_),
    .Y(_01079_),
    .B1(_06801_));
 sg13g2_nor2_1 _29435_ (.A(net1184),
    .B(net4188),
    .Y(_06805_));
 sg13g2_nor4_1 _29436_ (.A(_06100_),
    .B(_06104_),
    .C(_06107_),
    .D(_06794_),
    .Y(_06806_));
 sg13g2_nor2_1 _29437_ (.A(net3382),
    .B(_06806_),
    .Y(_06807_));
 sg13g2_a21oi_1 _29438_ (.A1(_06195_),
    .A2(net3338),
    .Y(_06808_),
    .B1(_06807_));
 sg13g2_xnor2_1 _29439_ (.Y(_06809_),
    .A(_06096_),
    .B(_06808_));
 sg13g2_a21oi_1 _29440_ (.A1(net4189),
    .A2(_06809_),
    .Y(_01080_),
    .B1(_06805_));
 sg13g2_nor2_1 _29441_ (.A(net1390),
    .B(net4186),
    .Y(_06810_));
 sg13g2_or2_1 _29442_ (.X(_06811_),
    .B(_06806_),
    .A(_06096_));
 sg13g2_a21oi_1 _29443_ (.A1(net3353),
    .A2(_06811_),
    .Y(_06812_),
    .B1(net3338));
 sg13g2_and2_1 _29444_ (.A(_06199_),
    .B(_06811_),
    .X(_06813_));
 sg13g2_xnor2_1 _29445_ (.Y(_06814_),
    .A(_06199_),
    .B(_06812_));
 sg13g2_a21oi_1 _29446_ (.A1(net4186),
    .A2(_06814_),
    .Y(_01081_),
    .B1(_06810_));
 sg13g2_nor2_1 _29447_ (.A(net1493),
    .B(net4189),
    .Y(_06815_));
 sg13g2_o21ai_1 _29448_ (.B1(net3311),
    .Y(_06816_),
    .A1(net3382),
    .A2(_06813_));
 sg13g2_xnor2_1 _29449_ (.Y(_06817_),
    .A(_06085_),
    .B(_06816_));
 sg13g2_a21oi_1 _29450_ (.A1(net4188),
    .A2(_06817_),
    .Y(_01082_),
    .B1(_06815_));
 sg13g2_nand2_1 _29451_ (.Y(_06818_),
    .A(net1074),
    .B(net4152));
 sg13g2_and3_1 _29452_ (.X(_06819_),
    .A(_06085_),
    .B(_06087_),
    .C(_06199_));
 sg13g2_o21ai_1 _29453_ (.B1(_06819_),
    .Y(_06820_),
    .A1(_06096_),
    .A2(_06806_));
 sg13g2_nand2_1 _29454_ (.Y(_06821_),
    .A(net3352),
    .B(_06820_));
 sg13g2_a21oi_1 _29455_ (.A1(_06085_),
    .A2(_06813_),
    .Y(_06822_),
    .B1(_06087_));
 sg13g2_a21oi_1 _29456_ (.A1(net3382),
    .A2(_06087_),
    .Y(_06823_),
    .B1(net4151));
 sg13g2_o21ai_1 _29457_ (.B1(_06823_),
    .Y(_06824_),
    .A1(_06821_),
    .A2(_06822_));
 sg13g2_o21ai_1 _29458_ (.B1(_06818_),
    .Y(_01083_),
    .A1(net3338),
    .A2(_06824_));
 sg13g2_nor2_1 _29459_ (.A(net1595),
    .B(net4188),
    .Y(_06825_));
 sg13g2_nand2_1 _29460_ (.Y(_06826_),
    .A(net3311),
    .B(_06821_));
 sg13g2_xor2_1 _29461_ (.B(_06826_),
    .A(_06092_),
    .X(_06827_));
 sg13g2_a21oi_1 _29462_ (.A1(net4189),
    .A2(_06827_),
    .Y(_01084_),
    .B1(_06825_));
 sg13g2_nand2_1 _29463_ (.Y(_06828_),
    .A(net1072),
    .B(net4152));
 sg13g2_or2_1 _29464_ (.X(_06829_),
    .B(_06092_),
    .A(_06090_));
 sg13g2_nor2_1 _29465_ (.A(_06820_),
    .B(_06829_),
    .Y(_06830_));
 sg13g2_nor2_1 _29466_ (.A(net3382),
    .B(_06830_),
    .Y(_06831_));
 sg13g2_o21ai_1 _29467_ (.B1(_06090_),
    .Y(_06832_),
    .A1(_06092_),
    .A2(_06820_));
 sg13g2_o21ai_1 _29468_ (.B1(net4188),
    .Y(_06833_),
    .A1(net3352),
    .A2(_06090_));
 sg13g2_a21o_1 _29469_ (.A2(_06832_),
    .A1(_06831_),
    .B1(_06833_),
    .X(_06834_));
 sg13g2_o21ai_1 _29470_ (.B1(_06828_),
    .Y(_01085_),
    .A1(net3338),
    .A2(_06834_));
 sg13g2_nor2_1 _29471_ (.A(net1610),
    .B(net4188),
    .Y(_06835_));
 sg13g2_nor2_1 _29472_ (.A(net3320),
    .B(_06831_),
    .Y(_06836_));
 sg13g2_xor2_1 _29473_ (.B(_06836_),
    .A(_06200_),
    .X(_06837_));
 sg13g2_a21oi_1 _29474_ (.A1(net4188),
    .A2(_06837_),
    .Y(_01086_),
    .B1(_06835_));
 sg13g2_nor2_1 _29475_ (.A(net2246),
    .B(net4188),
    .Y(_06838_));
 sg13g2_xnor2_1 _29476_ (.Y(_06839_),
    .A(net3352),
    .B(_06200_));
 sg13g2_nand2_1 _29477_ (.Y(_06840_),
    .A(_06836_),
    .B(_06839_));
 sg13g2_xnor2_1 _29478_ (.Y(_06841_),
    .A(_06078_),
    .B(_06840_));
 sg13g2_a21oi_1 _29479_ (.A1(net4188),
    .A2(_06841_),
    .Y(_01087_),
    .B1(_06838_));
 sg13g2_nand2_1 _29480_ (.Y(_06842_),
    .A(_06078_),
    .B(_06200_));
 sg13g2_nand3_1 _29481_ (.B(_06200_),
    .C(_06830_),
    .A(_06078_),
    .Y(_06843_));
 sg13g2_a21oi_1 _29482_ (.A1(net3352),
    .A2(_06843_),
    .Y(_06844_),
    .B1(net3320));
 sg13g2_xnor2_1 _29483_ (.Y(_06845_),
    .A(_06066_),
    .B(_06844_));
 sg13g2_nand2_1 _29484_ (.Y(_06846_),
    .A(net1223),
    .B(net4151));
 sg13g2_o21ai_1 _29485_ (.B1(_06846_),
    .Y(_01088_),
    .A1(net4152),
    .A2(_06845_));
 sg13g2_nor2_1 _29486_ (.A(_06065_),
    .B(net3311),
    .Y(_06847_));
 sg13g2_or2_1 _29487_ (.X(_06848_),
    .B(_06066_),
    .A(_06065_));
 sg13g2_or4_1 _29488_ (.A(_06820_),
    .B(_06829_),
    .C(_06842_),
    .D(_06848_),
    .X(_06849_));
 sg13g2_o21ai_1 _29489_ (.B1(_06065_),
    .Y(_06850_),
    .A1(_06066_),
    .A2(_06843_));
 sg13g2_and3_1 _29490_ (.X(_06851_),
    .A(net3352),
    .B(_06849_),
    .C(_06850_));
 sg13g2_o21ai_1 _29491_ (.B1(net4200),
    .Y(_06852_),
    .A1(net3352),
    .A2(_06848_));
 sg13g2_nor4_1 _29492_ (.A(net3338),
    .B(_06847_),
    .C(_06851_),
    .D(_06852_),
    .Y(_06853_));
 sg13g2_a21o_1 _29493_ (.A2(net4151),
    .A1(net2214),
    .B1(_06853_),
    .X(_01089_));
 sg13g2_a21o_1 _29494_ (.A2(_06849_),
    .A1(net3352),
    .B1(net3320),
    .X(_06854_));
 sg13g2_xnor2_1 _29495_ (.Y(_06855_),
    .A(_06081_),
    .B(_06854_));
 sg13g2_nand2_1 _29496_ (.Y(_06856_),
    .A(net1078),
    .B(net4152));
 sg13g2_o21ai_1 _29497_ (.B1(_06856_),
    .Y(_01090_),
    .A1(net4152),
    .A2(_06855_));
 sg13g2_nand2_1 _29498_ (.Y(_06857_),
    .A(net1077),
    .B(net4152));
 sg13g2_nor2b_1 _29499_ (.A(_06849_),
    .B_N(_06081_),
    .Y(_06858_));
 sg13g2_nand2_2 _29500_ (.Y(_06859_),
    .A(_06081_),
    .B(_06095_));
 sg13g2_nor2_1 _29501_ (.A(_06849_),
    .B(_06859_),
    .Y(_06860_));
 sg13g2_nor2_1 _29502_ (.A(net3382),
    .B(_06860_),
    .Y(_06861_));
 sg13g2_o21ai_1 _29503_ (.B1(_06861_),
    .Y(_06862_),
    .A1(_06095_),
    .A2(_06858_));
 sg13g2_a21oi_1 _29504_ (.A1(net3382),
    .A2(_06095_),
    .Y(_06863_),
    .B1(net4151));
 sg13g2_nand2_1 _29505_ (.Y(_06864_),
    .A(_06862_),
    .B(_06863_));
 sg13g2_o21ai_1 _29506_ (.B1(_06857_),
    .Y(_01091_),
    .A1(net3338),
    .A2(_06864_));
 sg13g2_nor2_1 _29507_ (.A(net1255),
    .B(net4192),
    .Y(_06865_));
 sg13g2_nor2_1 _29508_ (.A(net3320),
    .B(_06861_),
    .Y(_06866_));
 sg13g2_xnor2_1 _29509_ (.Y(_06867_),
    .A(_06208_),
    .B(_06866_));
 sg13g2_a21oi_1 _29510_ (.A1(net4192),
    .A2(_06867_),
    .Y(_01092_),
    .B1(_06865_));
 sg13g2_nor2_1 _29511_ (.A(_06207_),
    .B(_06208_),
    .Y(_06868_));
 sg13g2_inv_2 _29512_ (.Y(_06869_),
    .A(_06868_));
 sg13g2_a21oi_1 _29513_ (.A1(_06860_),
    .A2(_06868_),
    .Y(_06870_),
    .B1(net3382));
 sg13g2_o21ai_1 _29514_ (.B1(_06207_),
    .Y(_06871_),
    .A1(_06849_),
    .A2(_06859_));
 sg13g2_and3_1 _29515_ (.X(_06872_),
    .A(_06209_),
    .B(_06870_),
    .C(_06871_));
 sg13g2_o21ai_1 _29516_ (.B1(net4191),
    .Y(_06873_),
    .A1(net3353),
    .A2(_06869_));
 sg13g2_nor3_1 _29517_ (.A(net3338),
    .B(_06872_),
    .C(_06873_),
    .Y(_06874_));
 sg13g2_o21ai_1 _29518_ (.B1(_06874_),
    .Y(_06875_),
    .A1(_06207_),
    .A2(net3311));
 sg13g2_o21ai_1 _29519_ (.B1(_06875_),
    .Y(_01093_),
    .A1(_10996_),
    .A2(net4191));
 sg13g2_nor2_1 _29520_ (.A(net3320),
    .B(_06870_),
    .Y(_06876_));
 sg13g2_xor2_1 _29521_ (.B(_06876_),
    .A(_06068_),
    .X(_06877_));
 sg13g2_nand2_1 _29522_ (.Y(_06878_),
    .A(net1502),
    .B(net4153));
 sg13g2_o21ai_1 _29523_ (.B1(_06878_),
    .Y(_01094_),
    .A1(net4153),
    .A2(_06877_));
 sg13g2_nor2_1 _29524_ (.A(net1778),
    .B(net4192),
    .Y(_06879_));
 sg13g2_xnor2_1 _29525_ (.Y(_06880_),
    .A(net3353),
    .B(_06068_));
 sg13g2_nand2_1 _29526_ (.Y(_06881_),
    .A(_06876_),
    .B(_06880_));
 sg13g2_xnor2_1 _29527_ (.Y(_06882_),
    .A(_06060_),
    .B(_06881_));
 sg13g2_a21oi_1 _29528_ (.A1(net4192),
    .A2(_06882_),
    .Y(_01095_),
    .B1(_06879_));
 sg13g2_nand2_1 _29529_ (.Y(_06883_),
    .A(_06060_),
    .B(_06068_));
 sg13g2_nor4_2 _29530_ (.A(_06849_),
    .B(_06859_),
    .C(_06869_),
    .Y(_06884_),
    .D(_06883_));
 sg13g2_or4_1 _29531_ (.A(_06849_),
    .B(_06859_),
    .C(_06869_),
    .D(_06883_),
    .X(_06885_));
 sg13g2_a21oi_1 _29532_ (.A1(net3353),
    .A2(_06885_),
    .Y(_06886_),
    .B1(net3320));
 sg13g2_xor2_1 _29533_ (.B(_06886_),
    .A(_06062_),
    .X(_06887_));
 sg13g2_nand2_1 _29534_ (.Y(_06888_),
    .A(net1141),
    .B(net4153));
 sg13g2_o21ai_1 _29535_ (.B1(_06888_),
    .Y(_01096_),
    .A1(net4153),
    .A2(_06887_));
 sg13g2_nand2_1 _29536_ (.Y(_06889_),
    .A(_06062_),
    .B(_06884_));
 sg13g2_nand3_1 _29537_ (.B(_06204_),
    .C(_06884_),
    .A(_06062_),
    .Y(_06890_));
 sg13g2_nand2_1 _29538_ (.Y(_06891_),
    .A(net3357),
    .B(_06890_));
 sg13g2_a21oi_1 _29539_ (.A1(_06203_),
    .A2(_06889_),
    .Y(_06892_),
    .B1(_06891_));
 sg13g2_o21ai_1 _29540_ (.B1(net4196),
    .Y(_06893_),
    .A1(net3357),
    .A2(_06203_));
 sg13g2_nor3_1 _29541_ (.A(net3336),
    .B(_06892_),
    .C(_06893_),
    .Y(_06894_));
 sg13g2_a21o_1 _29542_ (.A2(net4154),
    .A1(net2233),
    .B1(_06894_),
    .X(_01097_));
 sg13g2_nor2_1 _29543_ (.A(net2253),
    .B(net4196),
    .Y(_06895_));
 sg13g2_nand2_1 _29544_ (.Y(_06896_),
    .A(net3312),
    .B(_06891_));
 sg13g2_xor2_1 _29545_ (.B(_06896_),
    .A(_06073_),
    .X(_06897_));
 sg13g2_a21oi_1 _29546_ (.A1(net4196),
    .A2(_06897_),
    .Y(_01098_),
    .B1(_06895_));
 sg13g2_nand2_1 _29547_ (.Y(_06898_),
    .A(_06062_),
    .B(_06204_));
 sg13g2_or3_1 _29548_ (.A(_06072_),
    .B(_06073_),
    .C(_06898_),
    .X(_06899_));
 sg13g2_or2_1 _29549_ (.X(_06900_),
    .B(_06899_),
    .A(_06885_));
 sg13g2_nand3_1 _29550_ (.B(_06074_),
    .C(_06900_),
    .A(net3357),
    .Y(_06901_));
 sg13g2_a21oi_1 _29551_ (.A1(_06072_),
    .A2(_06890_),
    .Y(_06902_),
    .B1(_06901_));
 sg13g2_o21ai_1 _29552_ (.B1(net4196),
    .Y(_06903_),
    .A1(net3357),
    .A2(_06072_));
 sg13g2_nor3_1 _29553_ (.A(net3336),
    .B(_06902_),
    .C(_06903_),
    .Y(_06904_));
 sg13g2_a21o_1 _29554_ (.A2(net4157),
    .A1(net2357),
    .B1(_06904_),
    .X(_01099_));
 sg13g2_a21oi_1 _29555_ (.A1(net3358),
    .A2(_06900_),
    .Y(_06905_),
    .B1(net3322));
 sg13g2_xnor2_1 _29556_ (.Y(_06906_),
    .A(_06221_),
    .B(_06905_));
 sg13g2_nand2_1 _29557_ (.Y(_06907_),
    .A(net1256),
    .B(net4155));
 sg13g2_o21ai_1 _29558_ (.B1(_06907_),
    .Y(_01100_),
    .A1(net4155),
    .A2(_06906_));
 sg13g2_nand2_2 _29559_ (.Y(_06908_),
    .A(_06220_),
    .B(_06223_));
 sg13g2_nor2_1 _29560_ (.A(_06900_),
    .B(_06908_),
    .Y(_06909_));
 sg13g2_or2_1 _29561_ (.X(_06910_),
    .B(_06909_),
    .A(net3381));
 sg13g2_o21ai_1 _29562_ (.B1(_06224_),
    .Y(_06911_),
    .A1(_06221_),
    .A2(_06900_));
 sg13g2_nor2b_1 _29563_ (.A(_06910_),
    .B_N(_06911_),
    .Y(_06912_));
 sg13g2_o21ai_1 _29564_ (.B1(net4199),
    .Y(_06913_),
    .A1(net3358),
    .A2(_06908_));
 sg13g2_nor3_1 _29565_ (.A(net3336),
    .B(_06912_),
    .C(_06913_),
    .Y(_06914_));
 sg13g2_o21ai_1 _29566_ (.B1(_06914_),
    .Y(_06915_),
    .A1(_06224_),
    .A2(net3311));
 sg13g2_o21ai_1 _29567_ (.B1(_06915_),
    .Y(_01101_),
    .A1(_10997_),
    .A2(net4196));
 sg13g2_nand2_1 _29568_ (.Y(_06916_),
    .A(net3311),
    .B(_06910_));
 sg13g2_xnor2_1 _29569_ (.Y(_06917_),
    .A(_06057_),
    .B(_06916_));
 sg13g2_nand2_1 _29570_ (.Y(_06918_),
    .A(net1094),
    .B(net4156));
 sg13g2_o21ai_1 _29571_ (.B1(_06918_),
    .Y(_01102_),
    .A1(net4155),
    .A2(_06917_));
 sg13g2_nor2_1 _29572_ (.A(net1994),
    .B(net4199),
    .Y(_06919_));
 sg13g2_xnor2_1 _29573_ (.Y(_06920_),
    .A(net3381),
    .B(_06057_));
 sg13g2_nor2_1 _29574_ (.A(_06916_),
    .B(_06920_),
    .Y(_06921_));
 sg13g2_xor2_1 _29575_ (.B(_06921_),
    .A(_06218_),
    .X(_06922_));
 sg13g2_a21oi_1 _29576_ (.A1(net4199),
    .A2(_06922_),
    .Y(_01103_),
    .B1(_06919_));
 sg13g2_nand2_1 _29577_ (.Y(_06923_),
    .A(_06057_),
    .B(_06218_));
 sg13g2_nor4_2 _29578_ (.A(_06885_),
    .B(_06899_),
    .C(_06908_),
    .Y(_06924_),
    .D(_06923_));
 sg13g2_nand3_1 _29579_ (.B(_06218_),
    .C(_06909_),
    .A(_06057_),
    .Y(_06925_));
 sg13g2_a21oi_1 _29580_ (.A1(net3358),
    .A2(_06925_),
    .Y(_06926_),
    .B1(net3321));
 sg13g2_xor2_1 _29581_ (.B(_06926_),
    .A(_06216_),
    .X(_06927_));
 sg13g2_nand2_1 _29582_ (.Y(_06928_),
    .A(net1080),
    .B(net4155));
 sg13g2_o21ai_1 _29583_ (.B1(_06928_),
    .Y(_01104_),
    .A1(net4156),
    .A2(_06927_));
 sg13g2_nand2_1 _29584_ (.Y(_06929_),
    .A(net1508),
    .B(net4155));
 sg13g2_a21oi_1 _29585_ (.A1(_06216_),
    .A2(_06924_),
    .Y(_06930_),
    .B1(_06055_));
 sg13g2_and3_1 _29586_ (.X(_06931_),
    .A(_06055_),
    .B(_06216_),
    .C(_06924_));
 sg13g2_nor2_1 _29587_ (.A(net3384),
    .B(_06931_),
    .Y(_06932_));
 sg13g2_nand2b_1 _29588_ (.Y(_06933_),
    .B(_06932_),
    .A_N(_06930_));
 sg13g2_a21oi_1 _29589_ (.A1(net3381),
    .A2(_06055_),
    .Y(_06934_),
    .B1(net4155));
 sg13g2_nand2_1 _29590_ (.Y(_06935_),
    .A(_06933_),
    .B(_06934_));
 sg13g2_o21ai_1 _29591_ (.B1(_06929_),
    .Y(_01105_),
    .A1(net3336),
    .A2(_06935_));
 sg13g2_nor2_1 _29592_ (.A(net2190),
    .B(net4197),
    .Y(_06936_));
 sg13g2_nor2_1 _29593_ (.A(net3321),
    .B(_06932_),
    .Y(_06937_));
 sg13g2_xor2_1 _29594_ (.B(_06937_),
    .A(_06247_),
    .X(_06938_));
 sg13g2_a21oi_1 _29595_ (.A1(net4197),
    .A2(_06938_),
    .Y(_01106_),
    .B1(_06936_));
 sg13g2_nand2_1 _29596_ (.Y(_06939_),
    .A(net1299),
    .B(net4155));
 sg13g2_nand4_1 _29597_ (.B(_06216_),
    .C(_06246_),
    .A(_06055_),
    .Y(_06940_),
    .D(_06247_));
 sg13g2_inv_1 _29598_ (.Y(_06941_),
    .A(_06940_));
 sg13g2_nor2_1 _29599_ (.A(_06925_),
    .B(_06940_),
    .Y(_06942_));
 sg13g2_or2_1 _29600_ (.X(_06943_),
    .B(_06942_),
    .A(net3384));
 sg13g2_a21oi_1 _29601_ (.A1(_06247_),
    .A2(_06931_),
    .Y(_06944_),
    .B1(_06246_));
 sg13g2_a21oi_1 _29602_ (.A1(net3384),
    .A2(_06246_),
    .Y(_06945_),
    .B1(net4158));
 sg13g2_o21ai_1 _29603_ (.B1(_06945_),
    .Y(_06946_),
    .A1(_06943_),
    .A2(_06944_));
 sg13g2_o21ai_1 _29604_ (.B1(_06939_),
    .Y(_01107_),
    .A1(net3337),
    .A2(_06946_));
 sg13g2_nor2_1 _29605_ (.A(net1794),
    .B(net4197),
    .Y(_06947_));
 sg13g2_nand2_1 _29606_ (.Y(_06948_),
    .A(net3313),
    .B(_06943_));
 sg13g2_xnor2_1 _29607_ (.Y(_06949_),
    .A(_06045_),
    .B(_06948_));
 sg13g2_a21oi_1 _29608_ (.A1(net4198),
    .A2(_06949_),
    .Y(_01108_),
    .B1(_06947_));
 sg13g2_nand2_1 _29609_ (.Y(_06950_),
    .A(net1377),
    .B(net4155));
 sg13g2_nand2_1 _29610_ (.Y(_06951_),
    .A(_06045_),
    .B(_06047_));
 sg13g2_nand3_1 _29611_ (.B(_06047_),
    .C(_06942_),
    .A(_06045_),
    .Y(_06952_));
 sg13g2_nand2_1 _29612_ (.Y(_06953_),
    .A(net3364),
    .B(_06952_));
 sg13g2_a21oi_1 _29613_ (.A1(_06045_),
    .A2(_06942_),
    .Y(_06954_),
    .B1(_06047_));
 sg13g2_a21oi_1 _29614_ (.A1(net3384),
    .A2(_06047_),
    .Y(_06955_),
    .B1(net4158));
 sg13g2_o21ai_1 _29615_ (.B1(_06955_),
    .Y(_06956_),
    .A1(_06953_),
    .A2(_06954_));
 sg13g2_o21ai_1 _29616_ (.B1(_06950_),
    .Y(_01109_),
    .A1(net3337),
    .A2(_06956_));
 sg13g2_nand2_1 _29617_ (.Y(_06957_),
    .A(net3313),
    .B(_06953_));
 sg13g2_xor2_1 _29618_ (.B(_06957_),
    .A(_06240_),
    .X(_06958_));
 sg13g2_nand2_1 _29619_ (.Y(_06959_),
    .A(net1095),
    .B(net4158));
 sg13g2_o21ai_1 _29620_ (.B1(_06959_),
    .Y(_01110_),
    .A1(net4158),
    .A2(_06958_));
 sg13g2_nor2_1 _29621_ (.A(net1700),
    .B(net4198),
    .Y(_06960_));
 sg13g2_xnor2_1 _29622_ (.Y(_06961_),
    .A(net3364),
    .B(_06240_));
 sg13g2_nor2_1 _29623_ (.A(_06957_),
    .B(_06961_),
    .Y(_06962_));
 sg13g2_xnor2_1 _29624_ (.Y(_06963_),
    .A(_06230_),
    .B(_06962_));
 sg13g2_a21oi_1 _29625_ (.A1(net4197),
    .A2(_06963_),
    .Y(_01111_),
    .B1(_06960_));
 sg13g2_nor2_1 _29626_ (.A(net1393),
    .B(net4197),
    .Y(_06964_));
 sg13g2_nor3_1 _29627_ (.A(_06230_),
    .B(_06240_),
    .C(_06951_),
    .Y(_06965_));
 sg13g2_nand3_1 _29628_ (.B(_06941_),
    .C(_06965_),
    .A(_06924_),
    .Y(_06966_));
 sg13g2_nor2_1 _29629_ (.A(net3384),
    .B(_06966_),
    .Y(_06967_));
 sg13g2_nor2_1 _29630_ (.A(net3340),
    .B(_06967_),
    .Y(_06968_));
 sg13g2_xnor2_1 _29631_ (.Y(_06969_),
    .A(_06214_),
    .B(_06968_));
 sg13g2_a21oi_1 _29632_ (.A1(net4197),
    .A2(_06969_),
    .Y(_01112_),
    .B1(_06964_));
 sg13g2_nand2_1 _29633_ (.Y(_06970_),
    .A(net1236),
    .B(net4158));
 sg13g2_nor2b_1 _29634_ (.A(_06966_),
    .B_N(_06214_),
    .Y(_06971_));
 sg13g2_a21oi_1 _29635_ (.A1(_06238_),
    .A2(_06971_),
    .Y(_06972_),
    .B1(net3384));
 sg13g2_o21ai_1 _29636_ (.B1(_06972_),
    .Y(_06973_),
    .A1(_06238_),
    .A2(_06971_));
 sg13g2_a21oi_1 _29637_ (.A1(net3384),
    .A2(_06238_),
    .Y(_06974_),
    .B1(net4158));
 sg13g2_nand2_1 _29638_ (.Y(_06975_),
    .A(_06973_),
    .B(_06974_));
 sg13g2_o21ai_1 _29639_ (.B1(_06970_),
    .Y(_01113_),
    .A1(net3340),
    .A2(_06975_));
 sg13g2_nor2_1 _29640_ (.A(net1653),
    .B(net4205),
    .Y(_06976_));
 sg13g2_nor2_1 _29641_ (.A(net3324),
    .B(_06972_),
    .Y(_06977_));
 sg13g2_xnor2_1 _29642_ (.Y(_06978_),
    .A(_06233_),
    .B(_06977_));
 sg13g2_a21oi_1 _29643_ (.A1(net4205),
    .A2(_06978_),
    .Y(_01114_),
    .B1(_06976_));
 sg13g2_nor2_1 _29644_ (.A(net1693),
    .B(net4198),
    .Y(_06979_));
 sg13g2_nand4_1 _29645_ (.B(_06232_),
    .C(_06238_),
    .A(_06214_),
    .Y(_06980_),
    .D(_06967_));
 sg13g2_nor2b_1 _29646_ (.A(net3340),
    .B_N(_06980_),
    .Y(_06981_));
 sg13g2_xnor2_1 _29647_ (.Y(_06982_),
    .A(_06243_),
    .B(_06981_));
 sg13g2_a21oi_1 _29648_ (.A1(net4198),
    .A2(_06982_),
    .Y(_01115_),
    .B1(_06979_));
 sg13g2_nor2_1 _29649_ (.A(net1578),
    .B(net4205),
    .Y(_06983_));
 sg13g2_nand4_1 _29650_ (.B(_06232_),
    .C(_06238_),
    .A(_06214_),
    .Y(_06984_),
    .D(_06243_));
 sg13g2_nor2_1 _29651_ (.A(_06966_),
    .B(_06984_),
    .Y(_06985_));
 sg13g2_a21oi_1 _29652_ (.A1(net3359),
    .A2(_06985_),
    .Y(_06986_),
    .B1(net3341));
 sg13g2_xnor2_1 _29653_ (.Y(_06987_),
    .A(_06036_),
    .B(_06986_));
 sg13g2_a21oi_1 _29654_ (.A1(net4205),
    .A2(_06987_),
    .Y(_01116_),
    .B1(_06983_));
 sg13g2_nand3_1 _29655_ (.B(_06363_),
    .C(_06985_),
    .A(_06036_),
    .Y(_06988_));
 sg13g2_a21o_1 _29656_ (.A2(_06985_),
    .A1(_06036_),
    .B1(_06363_),
    .X(_06989_));
 sg13g2_nand2_1 _29657_ (.Y(_06990_),
    .A(_06988_),
    .B(_06989_));
 sg13g2_a21oi_1 _29658_ (.A1(net3359),
    .A2(_06990_),
    .Y(_06991_),
    .B1(net4159));
 sg13g2_o21ai_1 _29659_ (.B1(_06991_),
    .Y(_06992_),
    .A1(_06363_),
    .A2(net3313));
 sg13g2_o21ai_1 _29660_ (.B1(_06992_),
    .Y(_06993_),
    .A1(net2668),
    .A2(net4205));
 sg13g2_inv_1 _29661_ (.Y(_01117_),
    .A(_06993_));
 sg13g2_nor2_1 _29662_ (.A(net1185),
    .B(net4204),
    .Y(_06994_));
 sg13g2_a21oi_1 _29663_ (.A1(net3359),
    .A2(_06988_),
    .Y(_06995_),
    .B1(net3324));
 sg13g2_xor2_1 _29664_ (.B(_06995_),
    .A(_06251_),
    .X(_06996_));
 sg13g2_a21oi_1 _29665_ (.A1(net4204),
    .A2(_06996_),
    .Y(_01118_),
    .B1(_06994_));
 sg13g2_nor2_1 _29666_ (.A(net1432),
    .B(net4204),
    .Y(_06997_));
 sg13g2_xnor2_1 _29667_ (.Y(_06998_),
    .A(net3359),
    .B(_06251_));
 sg13g2_nand2_1 _29668_ (.Y(_06999_),
    .A(_06995_),
    .B(_06998_));
 sg13g2_xnor2_1 _29669_ (.Y(_07000_),
    .A(_06269_),
    .B(_06999_));
 sg13g2_a21oi_1 _29670_ (.A1(net4204),
    .A2(_07000_),
    .Y(_01119_),
    .B1(_06997_));
 sg13g2_nor2_1 _29671_ (.A(net1713),
    .B(net4203),
    .Y(_07001_));
 sg13g2_nand4_1 _29672_ (.B(_06251_),
    .C(_06269_),
    .A(_06036_),
    .Y(_07002_),
    .D(_06363_));
 sg13g2_or2_1 _29673_ (.X(_07003_),
    .B(_07002_),
    .A(_06984_));
 sg13g2_nor2_1 _29674_ (.A(_06966_),
    .B(_07003_),
    .Y(_07004_));
 sg13g2_a21oi_1 _29675_ (.A1(net3360),
    .A2(_07004_),
    .Y(_07005_),
    .B1(net3340));
 sg13g2_xnor2_1 _29676_ (.Y(_07006_),
    .A(_06043_),
    .B(_07005_));
 sg13g2_a21oi_1 _29677_ (.A1(net4203),
    .A2(_07006_),
    .Y(_01120_),
    .B1(_07001_));
 sg13g2_nor2_1 _29678_ (.A(net1641),
    .B(net4204),
    .Y(_07007_));
 sg13g2_nand2_1 _29679_ (.Y(_07008_),
    .A(_06043_),
    .B(_07004_));
 sg13g2_or2_1 _29680_ (.X(_07009_),
    .B(_07008_),
    .A(_06264_));
 sg13g2_xnor2_1 _29681_ (.Y(_07010_),
    .A(_06264_),
    .B(_07008_));
 sg13g2_a22oi_1 _29682_ (.Y(_07011_),
    .B1(_07010_),
    .B2(net3360),
    .A2(net3324),
    .A1(_06264_));
 sg13g2_a21oi_1 _29683_ (.A1(net4203),
    .A2(_07011_),
    .Y(_01121_),
    .B1(_07007_));
 sg13g2_nor2_1 _29684_ (.A(net3385),
    .B(_07009_),
    .Y(_07012_));
 sg13g2_nor3_1 _29685_ (.A(_06367_),
    .B(net3340),
    .C(_07012_),
    .Y(_07013_));
 sg13g2_nor3_1 _29686_ (.A(net3385),
    .B(_06368_),
    .C(_07009_),
    .Y(_07014_));
 sg13g2_nor2_1 _29687_ (.A(_07013_),
    .B(_07014_),
    .Y(_07015_));
 sg13g2_nand2_1 _29688_ (.Y(_07016_),
    .A(net1101),
    .B(net4159));
 sg13g2_o21ai_1 _29689_ (.B1(_07016_),
    .Y(_01122_),
    .A1(net4159),
    .A2(_07015_));
 sg13g2_nor2_1 _29690_ (.A(net1623),
    .B(net4208),
    .Y(_07017_));
 sg13g2_nor2_1 _29691_ (.A(net3340),
    .B(_07014_),
    .Y(_07018_));
 sg13g2_nor2_1 _29692_ (.A(_06042_),
    .B(_06264_),
    .Y(_07019_));
 sg13g2_nand2_1 _29693_ (.Y(_07020_),
    .A(_06367_),
    .B(_07019_));
 sg13g2_nor3_1 _29694_ (.A(_06966_),
    .B(_07003_),
    .C(_07020_),
    .Y(_07021_));
 sg13g2_xor2_1 _29695_ (.B(_07018_),
    .A(_06052_),
    .X(_07022_));
 sg13g2_a21oi_1 _29696_ (.A1(net4208),
    .A2(_07022_),
    .Y(_01123_),
    .B1(_07017_));
 sg13g2_nor2_1 _29697_ (.A(net1760),
    .B(net4208),
    .Y(_07023_));
 sg13g2_nor4_1 _29698_ (.A(net3385),
    .B(_06052_),
    .C(_06368_),
    .D(_07009_),
    .Y(_07024_));
 sg13g2_nor2_1 _29699_ (.A(net3340),
    .B(_07024_),
    .Y(_07025_));
 sg13g2_xor2_1 _29700_ (.B(_07025_),
    .A(_06371_),
    .X(_07026_));
 sg13g2_a21oi_1 _29701_ (.A1(net4208),
    .A2(_07026_),
    .Y(_01124_),
    .B1(_07023_));
 sg13g2_nor2_1 _29702_ (.A(net1665),
    .B(net4202),
    .Y(_07027_));
 sg13g2_nor2_1 _29703_ (.A(_06052_),
    .B(_06371_),
    .Y(_07028_));
 sg13g2_nand2_1 _29704_ (.Y(_07029_),
    .A(_06367_),
    .B(_07028_));
 sg13g2_nand2_1 _29705_ (.Y(_07030_),
    .A(_07021_),
    .B(_07028_));
 sg13g2_nand2b_1 _29706_ (.Y(_07031_),
    .B(_07019_),
    .A_N(_06286_));
 sg13g2_nor2_1 _29707_ (.A(_06286_),
    .B(_07030_),
    .Y(_07032_));
 sg13g2_xnor2_1 _29708_ (.Y(_07033_),
    .A(_06286_),
    .B(_07030_));
 sg13g2_a22oi_1 _29709_ (.Y(_07034_),
    .B1(_07033_),
    .B2(net3361),
    .A2(net3324),
    .A1(_06286_));
 sg13g2_a21oi_1 _29710_ (.A1(net4202),
    .A2(_07034_),
    .Y(_01125_),
    .B1(_07027_));
 sg13g2_nor2_1 _29711_ (.A(net2029),
    .B(net4209),
    .Y(_07035_));
 sg13g2_o21ai_1 _29712_ (.B1(net3313),
    .Y(_07036_),
    .A1(net3386),
    .A2(_07032_));
 sg13g2_xnor2_1 _29713_ (.Y(_07037_),
    .A(_06284_),
    .B(_07036_));
 sg13g2_a21oi_1 _29714_ (.A1(net4209),
    .A2(_07037_),
    .Y(_01126_),
    .B1(_07035_));
 sg13g2_nor2_1 _29715_ (.A(net1821),
    .B(net4209),
    .Y(_07038_));
 sg13g2_xnor2_1 _29716_ (.Y(_07039_),
    .A(net3387),
    .B(_06284_));
 sg13g2_nor2_1 _29717_ (.A(_07036_),
    .B(_07039_),
    .Y(_07040_));
 sg13g2_xnor2_1 _29718_ (.Y(_07041_),
    .A(_06296_),
    .B(_07040_));
 sg13g2_a21oi_1 _29719_ (.A1(net4210),
    .A2(_07041_),
    .Y(_01127_),
    .B1(_07038_));
 sg13g2_and3_2 _29720_ (.X(_07042_),
    .A(_06284_),
    .B(_06297_),
    .C(_07032_));
 sg13g2_a21oi_1 _29721_ (.A1(net3360),
    .A2(_07042_),
    .Y(_07043_),
    .B1(net3340));
 sg13g2_nand2_1 _29722_ (.Y(_07044_),
    .A(_06039_),
    .B(_07042_));
 sg13g2_xnor2_1 _29723_ (.Y(_07045_),
    .A(_06039_),
    .B(_07043_));
 sg13g2_nand2_1 _29724_ (.Y(_07046_),
    .A(net1134),
    .B(net4159));
 sg13g2_o21ai_1 _29725_ (.B1(_07046_),
    .Y(_01128_),
    .A1(net4159),
    .A2(_07045_));
 sg13g2_nor2b_2 _29726_ (.A(_06373_),
    .B_N(_06039_),
    .Y(_07047_));
 sg13g2_nand2_2 _29727_ (.Y(_07048_),
    .A(_07042_),
    .B(_07047_));
 sg13g2_xnor2_1 _29728_ (.Y(_07049_),
    .A(_06373_),
    .B(_07044_));
 sg13g2_a221oi_1 _29729_ (.B2(net3360),
    .C1(net4160),
    .B1(_07049_),
    .A1(_06373_),
    .Y(_07050_),
    .A2(net3324));
 sg13g2_a21oi_1 _29730_ (.A1(_10998_),
    .A2(net4159),
    .Y(_01129_),
    .B1(_07050_));
 sg13g2_nor2_1 _29731_ (.A(net1667),
    .B(net4207),
    .Y(_07051_));
 sg13g2_a21oi_1 _29732_ (.A1(net3361),
    .A2(_07048_),
    .Y(_07052_),
    .B1(net3323));
 sg13g2_xnor2_1 _29733_ (.Y(_07053_),
    .A(_06361_),
    .B(_07052_));
 sg13g2_a21oi_1 _29734_ (.A1(net4206),
    .A2(_07053_),
    .Y(_01130_),
    .B1(_07051_));
 sg13g2_or2_1 _29735_ (.X(_07054_),
    .B(_06361_),
    .A(_06273_));
 sg13g2_o21ai_1 _29736_ (.B1(_06273_),
    .Y(_07055_),
    .A1(_06361_),
    .A2(_07048_));
 sg13g2_o21ai_1 _29737_ (.B1(_07055_),
    .Y(_07056_),
    .A1(_07048_),
    .A2(_07054_));
 sg13g2_a221oi_1 _29738_ (.B2(net3361),
    .C1(net4161),
    .B1(_07056_),
    .A1(_06273_),
    .Y(_07057_),
    .A2(net3323));
 sg13g2_a21oi_1 _29739_ (.A1(_10999_),
    .A2(net4160),
    .Y(_01131_),
    .B1(_07057_));
 sg13g2_nor2_1 _29740_ (.A(net1580),
    .B(net4206),
    .Y(_07058_));
 sg13g2_o21ai_1 _29741_ (.B1(net3361),
    .Y(_07059_),
    .A1(_07048_),
    .A2(_07054_));
 sg13g2_nand2_1 _29742_ (.Y(_07060_),
    .A(net3317),
    .B(_07059_));
 sg13g2_xor2_1 _29743_ (.B(_07060_),
    .A(_06328_),
    .X(_07061_));
 sg13g2_a21oi_1 _29744_ (.A1(net4206),
    .A2(_07061_),
    .Y(_01132_),
    .B1(_07058_));
 sg13g2_or3_1 _29745_ (.A(_06327_),
    .B(_06328_),
    .C(_07054_),
    .X(_07062_));
 sg13g2_or2_1 _29746_ (.X(_07063_),
    .B(_07062_),
    .A(_07048_));
 sg13g2_nand2_1 _29747_ (.Y(_07064_),
    .A(_06329_),
    .B(_07063_));
 sg13g2_a221oi_1 _29748_ (.B2(net3361),
    .C1(net4161),
    .B1(_07064_),
    .A1(_06327_),
    .Y(_07065_),
    .A2(_07060_));
 sg13g2_a21oi_1 _29749_ (.A1(_11000_),
    .A2(net4159),
    .Y(_01133_),
    .B1(_07065_));
 sg13g2_nor2_1 _29750_ (.A(net1434),
    .B(net4206),
    .Y(_07066_));
 sg13g2_a21o_1 _29751_ (.A2(_07063_),
    .A1(net3361),
    .B1(net3323),
    .X(_07067_));
 sg13g2_xor2_1 _29752_ (.B(_07067_),
    .A(_06377_),
    .X(_07068_));
 sg13g2_a21oi_1 _29753_ (.A1(net4206),
    .A2(_07068_),
    .Y(_01134_),
    .B1(_07066_));
 sg13g2_nor2_1 _29754_ (.A(net1526),
    .B(net4207),
    .Y(_07069_));
 sg13g2_xnor2_1 _29755_ (.Y(_07070_),
    .A(net3361),
    .B(_06377_));
 sg13g2_nor2_1 _29756_ (.A(_07067_),
    .B(_07070_),
    .Y(_07071_));
 sg13g2_xnor2_1 _29757_ (.Y(_07072_),
    .A(_06370_),
    .B(_07071_));
 sg13g2_a21oi_1 _29758_ (.A1(net4206),
    .A2(_07072_),
    .Y(_01135_),
    .B1(_07069_));
 sg13g2_nor2_1 _29759_ (.A(net1724),
    .B(net4209),
    .Y(_07073_));
 sg13g2_or2_1 _29760_ (.X(_07074_),
    .B(_06377_),
    .A(_06370_));
 sg13g2_nor2_1 _29761_ (.A(_07063_),
    .B(_07074_),
    .Y(_07075_));
 sg13g2_o21ai_1 _29762_ (.B1(net3317),
    .Y(_07076_),
    .A1(net3386),
    .A2(_07075_));
 sg13g2_xor2_1 _29763_ (.B(_07076_),
    .A(_06289_),
    .X(_07077_));
 sg13g2_a21oi_1 _29764_ (.A1(net4209),
    .A2(_07077_),
    .Y(_01136_),
    .B1(_07073_));
 sg13g2_nor2_1 _29765_ (.A(_06288_),
    .B(_06289_),
    .Y(_07078_));
 sg13g2_and2_1 _29766_ (.A(_07075_),
    .B(_07078_),
    .X(_07079_));
 sg13g2_o21ai_1 _29767_ (.B1(net3363),
    .Y(_07080_),
    .A1(_06290_),
    .A2(_07079_));
 sg13g2_a21oi_1 _29768_ (.A1(_06288_),
    .A2(_07076_),
    .Y(_07081_),
    .B1(net4161));
 sg13g2_a22oi_1 _29769_ (.Y(_01137_),
    .B1(_07080_),
    .B2(_07081_),
    .A2(net4161),
    .A1(_11001_));
 sg13g2_nor2_1 _29770_ (.A(net1523),
    .B(net4210),
    .Y(_07082_));
 sg13g2_a21oi_1 _29771_ (.A1(net3363),
    .A2(_07079_),
    .Y(_07083_),
    .B1(net3341));
 sg13g2_xnor2_1 _29772_ (.Y(_07084_),
    .A(_06262_),
    .B(_07083_));
 sg13g2_a21oi_1 _29773_ (.A1(net4209),
    .A2(_07084_),
    .Y(_01138_),
    .B1(_07082_));
 sg13g2_nor2_1 _29774_ (.A(net1177),
    .B(net4210),
    .Y(_07085_));
 sg13g2_nand2_1 _29775_ (.Y(_07086_),
    .A(_06262_),
    .B(_07079_));
 sg13g2_o21ai_1 _29776_ (.B1(net3330),
    .Y(_07087_),
    .A1(net3386),
    .A2(_07086_));
 sg13g2_xnor2_1 _29777_ (.Y(_07088_),
    .A(_06388_),
    .B(_07087_));
 sg13g2_a21oi_1 _29778_ (.A1(net4210),
    .A2(_07088_),
    .Y(_01139_),
    .B1(_07085_));
 sg13g2_nor2_1 _29779_ (.A(net1510),
    .B(net4207),
    .Y(_07089_));
 sg13g2_nor2_1 _29780_ (.A(_06388_),
    .B(_07086_),
    .Y(_07090_));
 sg13g2_o21ai_1 _29781_ (.B1(net3317),
    .Y(_07091_),
    .A1(net3386),
    .A2(_07090_));
 sg13g2_xor2_1 _29782_ (.B(_07091_),
    .A(_06236_),
    .X(_07092_));
 sg13g2_a21oi_1 _29783_ (.A1(net4206),
    .A2(_07092_),
    .Y(_01140_),
    .B1(_07089_));
 sg13g2_nor3_1 _29784_ (.A(_06236_),
    .B(_06388_),
    .C(_07086_),
    .Y(_07093_));
 sg13g2_nor2_1 _29785_ (.A(_06236_),
    .B(_06253_),
    .Y(_07094_));
 sg13g2_xor2_1 _29786_ (.B(_07093_),
    .A(_06253_),
    .X(_07095_));
 sg13g2_a221oi_1 _29787_ (.B2(net3361),
    .C1(net4161),
    .B1(_07095_),
    .A1(_06253_),
    .Y(_07096_),
    .A2(net3323));
 sg13g2_a21oi_1 _29788_ (.A1(_11002_),
    .A2(net4161),
    .Y(_01141_),
    .B1(_07096_));
 sg13g2_nor2_1 _29789_ (.A(net1538),
    .B(net4209),
    .Y(_07097_));
 sg13g2_a21oi_1 _29790_ (.A1(_07090_),
    .A2(_07094_),
    .Y(_07098_),
    .B1(net3386));
 sg13g2_nor2_1 _29791_ (.A(net3323),
    .B(_07098_),
    .Y(_07099_));
 sg13g2_xnor2_1 _29792_ (.Y(_07100_),
    .A(_06365_),
    .B(_07099_));
 sg13g2_a21oi_1 _29793_ (.A1(net4209),
    .A2(_07100_),
    .Y(_01142_),
    .B1(_07097_));
 sg13g2_nor2_1 _29794_ (.A(net1551),
    .B(net4207),
    .Y(_07101_));
 sg13g2_xnor2_1 _29795_ (.Y(_07102_),
    .A(net3386),
    .B(_06365_));
 sg13g2_nand2_1 _29796_ (.Y(_07103_),
    .A(_07099_),
    .B(_07102_));
 sg13g2_xnor2_1 _29797_ (.Y(_07104_),
    .A(_06266_),
    .B(_07103_));
 sg13g2_a21oi_1 _29798_ (.A1(net4206),
    .A2(_07104_),
    .Y(_01143_),
    .B1(_07101_));
 sg13g2_nor2_1 _29799_ (.A(net1636),
    .B(net4212),
    .Y(_07105_));
 sg13g2_nand3_1 _29800_ (.B(_07078_),
    .C(_07094_),
    .A(_07047_),
    .Y(_07106_));
 sg13g2_nand3b_1 _29801_ (.B(_06266_),
    .C(_06262_),
    .Y(_07107_),
    .A_N(_06365_));
 sg13g2_or2_1 _29802_ (.X(_07108_),
    .B(_07107_),
    .A(_06388_));
 sg13g2_nor4_2 _29803_ (.A(_07062_),
    .B(_07074_),
    .C(_07106_),
    .Y(_07109_),
    .D(_07108_));
 sg13g2_nand2_2 _29804_ (.Y(_07110_),
    .A(_07042_),
    .B(_07109_));
 sg13g2_a21oi_1 _29805_ (.A1(net3362),
    .A2(_07110_),
    .Y(_07111_),
    .B1(net3323));
 sg13g2_xnor2_1 _29806_ (.Y(_07112_),
    .A(_06352_),
    .B(_07111_));
 sg13g2_a21oi_1 _29807_ (.A1(net4213),
    .A2(_07112_),
    .Y(_01144_),
    .B1(_07105_));
 sg13g2_nor3_1 _29808_ (.A(net3387),
    .B(_06352_),
    .C(_07110_),
    .Y(_07113_));
 sg13g2_or3_1 _29809_ (.A(_06347_),
    .B(net3341),
    .C(_07113_),
    .X(_07114_));
 sg13g2_nor3_1 _29810_ (.A(_06346_),
    .B(_06352_),
    .C(_07110_),
    .Y(_07115_));
 sg13g2_a21oi_1 _29811_ (.A1(net3362),
    .A2(_07115_),
    .Y(_07116_),
    .B1(net4162));
 sg13g2_a22oi_1 _29812_ (.Y(_01145_),
    .B1(_07114_),
    .B2(_07116_),
    .A2(net4162),
    .A1(_11003_));
 sg13g2_nor2_1 _29813_ (.A(net1757),
    .B(net4213),
    .Y(_07117_));
 sg13g2_o21ai_1 _29814_ (.B1(net3313),
    .Y(_07118_),
    .A1(net3387),
    .A2(_07115_));
 sg13g2_xnor2_1 _29815_ (.Y(_07119_),
    .A(_06349_),
    .B(_07118_));
 sg13g2_a21oi_1 _29816_ (.A1(net4213),
    .A2(_07119_),
    .Y(_01146_),
    .B1(_07117_));
 sg13g2_nor2_1 _29817_ (.A(net1735),
    .B(net4213),
    .Y(_07120_));
 sg13g2_nand2_1 _29818_ (.Y(_07121_),
    .A(net3387),
    .B(_06353_));
 sg13g2_o21ai_1 _29819_ (.B1(_07121_),
    .Y(_07122_),
    .A1(_06350_),
    .A2(_07118_));
 sg13g2_and2_1 _29820_ (.A(net3313),
    .B(_07122_),
    .X(_07123_));
 sg13g2_xnor2_1 _29821_ (.Y(_07124_),
    .A(_06381_),
    .B(_07123_));
 sg13g2_a21oi_1 _29822_ (.A1(net4211),
    .A2(_07124_),
    .Y(_01147_),
    .B1(_07120_));
 sg13g2_nor2_1 _29823_ (.A(net1605),
    .B(net4211),
    .Y(_07125_));
 sg13g2_nor2_1 _29824_ (.A(_06350_),
    .B(_06381_),
    .Y(_07126_));
 sg13g2_and2_1 _29825_ (.A(_07115_),
    .B(_07126_),
    .X(_07127_));
 sg13g2_a21oi_1 _29826_ (.A1(net3362),
    .A2(_07127_),
    .Y(_07128_),
    .B1(net3341));
 sg13g2_xnor2_1 _29827_ (.Y(_07129_),
    .A(_06258_),
    .B(_07128_));
 sg13g2_a21oi_1 _29828_ (.A1(net4211),
    .A2(_07129_),
    .Y(_01148_),
    .B1(_07125_));
 sg13g2_nor2_1 _29829_ (.A(net1692),
    .B(net4211),
    .Y(_07130_));
 sg13g2_nand2_1 _29830_ (.Y(_07131_),
    .A(_06258_),
    .B(_07127_));
 sg13g2_xnor2_1 _29831_ (.Y(_07132_),
    .A(_06292_),
    .B(_07131_));
 sg13g2_a22oi_1 _29832_ (.Y(_07133_),
    .B1(_07132_),
    .B2(net3362),
    .A2(net3323),
    .A1(_06292_));
 sg13g2_a21oi_1 _29833_ (.A1(net4211),
    .A2(_07133_),
    .Y(_01149_),
    .B1(_07130_));
 sg13g2_o21ai_1 _29834_ (.B1(net3362),
    .Y(_07134_),
    .A1(_06292_),
    .A2(_07131_));
 sg13g2_and2_1 _29835_ (.A(net3313),
    .B(_07134_),
    .X(_07135_));
 sg13g2_xor2_1 _29836_ (.B(_07135_),
    .A(_06279_),
    .X(_07136_));
 sg13g2_nand2_1 _29837_ (.Y(_07137_),
    .A(net1135),
    .B(net4161));
 sg13g2_o21ai_1 _29838_ (.B1(_07137_),
    .Y(_01150_),
    .A1(net4161),
    .A2(_07136_));
 sg13g2_nor2_1 _29839_ (.A(net1921),
    .B(net4211),
    .Y(_07138_));
 sg13g2_xnor2_1 _29840_ (.Y(_07139_),
    .A(net3362),
    .B(_06279_));
 sg13g2_nand2_1 _29841_ (.Y(_07140_),
    .A(_07135_),
    .B(_07139_));
 sg13g2_xnor2_1 _29842_ (.Y(_07141_),
    .A(_06278_),
    .B(_07140_));
 sg13g2_a21oi_1 _29843_ (.A1(net4211),
    .A2(_07141_),
    .Y(_01151_),
    .B1(_07138_));
 sg13g2_nor2_1 _29844_ (.A(net1574),
    .B(net4212),
    .Y(_07142_));
 sg13g2_and4_1 _29845_ (.A(_06278_),
    .B(_06279_),
    .C(_06347_),
    .D(_06351_),
    .X(_07143_));
 sg13g2_nand4_1 _29846_ (.B(_06293_),
    .C(_07126_),
    .A(_06258_),
    .Y(_07144_),
    .D(_07143_));
 sg13g2_nor2_1 _29847_ (.A(_07110_),
    .B(_07144_),
    .Y(_07145_));
 sg13g2_o21ai_1 _29848_ (.B1(net3313),
    .Y(_07146_),
    .A1(net3387),
    .A2(_07145_));
 sg13g2_xnor2_1 _29849_ (.Y(_07147_),
    .A(_06321_),
    .B(_07146_));
 sg13g2_a21oi_1 _29850_ (.A1(net4212),
    .A2(_07147_),
    .Y(_01152_),
    .B1(_07142_));
 sg13g2_nor2_1 _29851_ (.A(net1944),
    .B(net4214),
    .Y(_07148_));
 sg13g2_nor4_1 _29852_ (.A(_06319_),
    .B(_06320_),
    .C(_07110_),
    .D(_07144_),
    .Y(_07149_));
 sg13g2_nand2_1 _29853_ (.Y(_07150_),
    .A(net3362),
    .B(_07149_));
 sg13g2_o21ai_1 _29854_ (.B1(_07150_),
    .Y(_07151_),
    .A1(net3386),
    .A2(_06322_));
 sg13g2_a21oi_1 _29855_ (.A1(_06319_),
    .A2(_07146_),
    .Y(_07152_),
    .B1(_07151_));
 sg13g2_a21oi_1 _29856_ (.A1(net4212),
    .A2(_07152_),
    .Y(_01153_),
    .B1(_07148_));
 sg13g2_nand2_1 _29857_ (.Y(_07153_),
    .A(net3330),
    .B(_07150_));
 sg13g2_nor2_1 _29858_ (.A(_06405_),
    .B(net3344),
    .Y(_07154_));
 sg13g2_a221oi_1 _29859_ (.B2(_07150_),
    .C1(net4162),
    .B1(_07154_),
    .A1(_06405_),
    .Y(_07155_),
    .A2(_07153_));
 sg13g2_a21oi_1 _29860_ (.A1(_11004_),
    .A2(net4162),
    .Y(_01154_),
    .B1(_07155_));
 sg13g2_o21ai_1 _29861_ (.B1(_07153_),
    .Y(_07156_),
    .A1(_06405_),
    .A2(net3341));
 sg13g2_xor2_1 _29862_ (.B(_07156_),
    .A(_06404_),
    .X(_07157_));
 sg13g2_mux2_1 _29863_ (.A0(net2481),
    .A1(_07157_),
    .S(net4213),
    .X(_01155_));
 sg13g2_nor2_1 _29864_ (.A(net1964),
    .B(net4214),
    .Y(_07158_));
 sg13g2_nand3_1 _29865_ (.B(_06405_),
    .C(_07149_),
    .A(_06404_),
    .Y(_07159_));
 sg13g2_a21oi_1 _29866_ (.A1(net3362),
    .A2(_07159_),
    .Y(_07160_),
    .B1(net3323));
 sg13g2_xnor2_1 _29867_ (.Y(_07161_),
    .A(_06357_),
    .B(_07160_));
 sg13g2_a21oi_1 _29868_ (.A1(net4212),
    .A2(_07161_),
    .Y(_01156_),
    .B1(_07158_));
 sg13g2_or2_1 _29869_ (.X(_07162_),
    .B(_06383_),
    .A(_06357_));
 sg13g2_o21ai_1 _29870_ (.B1(_06383_),
    .Y(_07163_),
    .A1(_06357_),
    .A2(_07159_));
 sg13g2_o21ai_1 _29871_ (.B1(_07163_),
    .Y(_07164_),
    .A1(_07159_),
    .A2(_07162_));
 sg13g2_a221oi_1 _29872_ (.B2(net3365),
    .C1(net4162),
    .B1(_07164_),
    .A1(_06383_),
    .Y(_07165_),
    .A2(net3325));
 sg13g2_a21oi_1 _29873_ (.A1(_11005_),
    .A2(net4165),
    .Y(_01157_),
    .B1(_07165_));
 sg13g2_nor2_1 _29874_ (.A(net1581),
    .B(net4214),
    .Y(_07166_));
 sg13g2_o21ai_1 _29875_ (.B1(net3365),
    .Y(_07167_),
    .A1(_07159_),
    .A2(_07162_));
 sg13g2_and2_1 _29876_ (.A(net3316),
    .B(_07167_),
    .X(_07168_));
 sg13g2_xnor2_1 _29877_ (.Y(_07169_),
    .A(_06343_),
    .B(_07168_));
 sg13g2_a21oi_1 _29878_ (.A1(net4214),
    .A2(_07169_),
    .Y(_01158_),
    .B1(_07166_));
 sg13g2_nor2_1 _29879_ (.A(net1511),
    .B(net4214),
    .Y(_07170_));
 sg13g2_xnor2_1 _29880_ (.Y(_07171_),
    .A(net3386),
    .B(_06343_));
 sg13g2_nand2_1 _29881_ (.Y(_07172_),
    .A(_07168_),
    .B(_07171_));
 sg13g2_xnor2_1 _29882_ (.Y(_07173_),
    .A(_06311_),
    .B(_07172_));
 sg13g2_a21oi_1 _29883_ (.A1(net4214),
    .A2(_07173_),
    .Y(_01159_),
    .B1(_07170_));
 sg13g2_nor2_1 _29884_ (.A(net1437),
    .B(net4218),
    .Y(_07174_));
 sg13g2_or2_1 _29885_ (.X(_07175_),
    .B(_06343_),
    .A(_06310_));
 sg13g2_nand4_1 _29886_ (.B(_06321_),
    .C(_06404_),
    .A(_06318_),
    .Y(_07176_),
    .D(_06405_));
 sg13g2_or4_1 _29887_ (.A(_07144_),
    .B(_07162_),
    .C(_07175_),
    .D(_07176_),
    .X(_07177_));
 sg13g2_nor2_1 _29888_ (.A(_07110_),
    .B(_07177_),
    .Y(_07178_));
 sg13g2_o21ai_1 _29889_ (.B1(net3316),
    .Y(_07179_),
    .A1(net3391),
    .A2(_07178_));
 sg13g2_xnor2_1 _29890_ (.Y(_07180_),
    .A(_06392_),
    .B(_07179_));
 sg13g2_a21oi_1 _29891_ (.A1(net4218),
    .A2(_07180_),
    .Y(_01160_),
    .B1(_07174_));
 sg13g2_nand2b_1 _29892_ (.Y(_07181_),
    .B(_07179_),
    .A_N(_06391_));
 sg13g2_nand2_1 _29893_ (.Y(_07182_),
    .A(_06391_),
    .B(_06392_));
 sg13g2_nor3_1 _29894_ (.A(_07110_),
    .B(_07177_),
    .C(_07182_),
    .Y(_07183_));
 sg13g2_o21ai_1 _29895_ (.B1(net3366),
    .Y(_07184_),
    .A1(_06393_),
    .A2(_07183_));
 sg13g2_nand3_1 _29896_ (.B(_07181_),
    .C(_07184_),
    .A(net4217),
    .Y(_07185_));
 sg13g2_o21ai_1 _29897_ (.B1(_07185_),
    .Y(_07186_),
    .A1(net2898),
    .A2(net4217));
 sg13g2_inv_1 _29898_ (.Y(_01161_),
    .A(_07186_));
 sg13g2_o21ai_1 _29899_ (.B1(net3316),
    .Y(_07187_),
    .A1(net3391),
    .A2(_07183_));
 sg13g2_xnor2_1 _29900_ (.Y(_07188_),
    .A(_06398_),
    .B(_07187_));
 sg13g2_nand2_1 _29901_ (.Y(_07189_),
    .A(net1082),
    .B(net4164));
 sg13g2_o21ai_1 _29902_ (.B1(_07189_),
    .Y(_01162_),
    .A1(net4164),
    .A2(_07188_));
 sg13g2_and3_1 _29903_ (.X(_07190_),
    .A(_06396_),
    .B(_06398_),
    .C(_07183_));
 sg13g2_o21ai_1 _29904_ (.B1(net3366),
    .Y(_07191_),
    .A1(_06399_),
    .A2(_07190_));
 sg13g2_a21oi_1 _29905_ (.A1(_06397_),
    .A2(_07187_),
    .Y(_07192_),
    .B1(net4163));
 sg13g2_a22oi_1 _29906_ (.Y(_01163_),
    .B1(_07191_),
    .B2(_07192_),
    .A2(net4163),
    .A1(_11006_));
 sg13g2_nor2_1 _29907_ (.A(net1591),
    .B(net4226),
    .Y(_07193_));
 sg13g2_o21ai_1 _29908_ (.B1(net3316),
    .Y(_07194_),
    .A1(net3391),
    .A2(_07190_));
 sg13g2_xnor2_1 _29909_ (.Y(_07195_),
    .A(_06032_),
    .B(_07194_));
 sg13g2_a21oi_1 _29910_ (.A1(net4230),
    .A2(_07195_),
    .Y(_01164_),
    .B1(_07193_));
 sg13g2_nand4_1 _29911_ (.B(_06032_),
    .C(_06396_),
    .A(_06030_),
    .Y(_07196_),
    .D(_06398_));
 sg13g2_or4_1 _29912_ (.A(_07110_),
    .B(_07177_),
    .C(_07182_),
    .D(_07196_),
    .X(_07197_));
 sg13g2_nand2_1 _29913_ (.Y(_07198_),
    .A(_06033_),
    .B(_07197_));
 sg13g2_a221oi_1 _29914_ (.B2(net3366),
    .C1(net4163),
    .B1(_07198_),
    .A1(_06031_),
    .Y(_07199_),
    .A2(_07194_));
 sg13g2_a21oi_1 _29915_ (.A1(_11007_),
    .A2(net4170),
    .Y(_01165_),
    .B1(_07199_));
 sg13g2_a21o_1 _29916_ (.A2(_07197_),
    .A1(net3366),
    .B1(net3325),
    .X(_07200_));
 sg13g2_xnor2_1 _29917_ (.Y(_07201_),
    .A(_06359_),
    .B(_07200_));
 sg13g2_nand2_1 _29918_ (.Y(_07202_),
    .A(net1120),
    .B(net4163));
 sg13g2_o21ai_1 _29919_ (.B1(_07202_),
    .Y(_01166_),
    .A1(net4163),
    .A2(_07201_));
 sg13g2_nor2_1 _29920_ (.A(net2300),
    .B(net4217),
    .Y(_07203_));
 sg13g2_xnor2_1 _29921_ (.Y(_07204_),
    .A(net3391),
    .B(_06359_));
 sg13g2_nor2_1 _29922_ (.A(_07200_),
    .B(_07204_),
    .Y(_07205_));
 sg13g2_xnor2_1 _29923_ (.Y(_07206_),
    .A(_06385_),
    .B(_07205_));
 sg13g2_a21oi_1 _29924_ (.A1(net4217),
    .A2(_07206_),
    .Y(_01167_),
    .B1(_07203_));
 sg13g2_nor2_1 _29925_ (.A(net1914),
    .B(net4231),
    .Y(_07207_));
 sg13g2_nand2_1 _29926_ (.Y(_07208_),
    .A(_06359_),
    .B(_06386_));
 sg13g2_o21ai_1 _29927_ (.B1(net3366),
    .Y(_07209_),
    .A1(_07197_),
    .A2(_07208_));
 sg13g2_nand2_1 _29928_ (.Y(_07210_),
    .A(net3316),
    .B(_07209_));
 sg13g2_xnor2_1 _29929_ (.Y(_07211_),
    .A(_06020_),
    .B(_07210_));
 sg13g2_a21oi_1 _29930_ (.A1(net4231),
    .A2(_07211_),
    .Y(_01168_),
    .B1(_07207_));
 sg13g2_nand4_1 _29931_ (.B(_06022_),
    .C(_06359_),
    .A(_06020_),
    .Y(_07212_),
    .D(_06386_));
 sg13g2_nor2_2 _29932_ (.A(_07197_),
    .B(_07212_),
    .Y(_07213_));
 sg13g2_o21ai_1 _29933_ (.B1(net3366),
    .Y(_07214_),
    .A1(_06024_),
    .A2(_07213_));
 sg13g2_a21oi_1 _29934_ (.A1(_06023_),
    .A2(_07210_),
    .Y(_07215_),
    .B1(net4163));
 sg13g2_a22oi_1 _29935_ (.Y(_01169_),
    .B1(_07214_),
    .B2(_07215_),
    .A2(net4164),
    .A1(_11008_));
 sg13g2_nor2_1 _29936_ (.A(net2087),
    .B(net4230),
    .Y(_07216_));
 sg13g2_o21ai_1 _29937_ (.B1(net3315),
    .Y(_07217_),
    .A1(net3392),
    .A2(_07213_));
 sg13g2_xor2_1 _29938_ (.B(_07217_),
    .A(_06315_),
    .X(_07218_));
 sg13g2_a21oi_1 _29939_ (.A1(net4230),
    .A2(_07218_),
    .Y(_01170_),
    .B1(_07216_));
 sg13g2_or4_1 _29940_ (.A(_06314_),
    .B(_06315_),
    .C(_07197_),
    .D(_07212_),
    .X(_07219_));
 sg13g2_nand2_1 _29941_ (.Y(_07220_),
    .A(_06316_),
    .B(_07219_));
 sg13g2_a221oi_1 _29942_ (.B2(net3367),
    .C1(net4163),
    .B1(_07220_),
    .A1(_06314_),
    .Y(_07221_),
    .A2(_07217_));
 sg13g2_a21oi_1 _29943_ (.A1(_11009_),
    .A2(net4164),
    .Y(_01171_),
    .B1(_07221_));
 sg13g2_nor2_1 _29944_ (.A(net1743),
    .B(net4229),
    .Y(_07222_));
 sg13g2_a21o_1 _29945_ (.A2(_07219_),
    .A1(net3367),
    .B1(net3328),
    .X(_07223_));
 sg13g2_xor2_1 _29946_ (.B(_07223_),
    .A(_06335_),
    .X(_07224_));
 sg13g2_a21oi_1 _29947_ (.A1(net4231),
    .A2(_07224_),
    .Y(_01172_),
    .B1(_07222_));
 sg13g2_nor4_2 _29948_ (.A(_06314_),
    .B(_06315_),
    .C(_06334_),
    .Y(_07225_),
    .D(_06335_));
 sg13g2_nand2_1 _29949_ (.Y(_07226_),
    .A(_07213_),
    .B(_07225_));
 sg13g2_nand2_1 _29950_ (.Y(_07227_),
    .A(_06336_),
    .B(_07226_));
 sg13g2_a221oi_1 _29951_ (.B2(net3367),
    .C1(net4163),
    .B1(_07227_),
    .A1(_06334_),
    .Y(_07228_),
    .A2(_07223_));
 sg13g2_a21oi_1 _29952_ (.A1(_11010_),
    .A2(net4171),
    .Y(_01173_),
    .B1(_07228_));
 sg13g2_nand3_1 _29953_ (.B(_07213_),
    .C(_07225_),
    .A(net3367),
    .Y(_07229_));
 sg13g2_nand2_1 _29954_ (.Y(_07230_),
    .A(net3330),
    .B(_07229_));
 sg13g2_xnor2_1 _29955_ (.Y(_07231_),
    .A(_06375_),
    .B(_07230_));
 sg13g2_nand2_1 _29956_ (.Y(_07232_),
    .A(net1111),
    .B(net4170));
 sg13g2_o21ai_1 _29957_ (.B1(_07232_),
    .Y(_01174_),
    .A1(net4171),
    .A2(_07231_));
 sg13g2_nor2_1 _29958_ (.A(net1703),
    .B(net4227),
    .Y(_07233_));
 sg13g2_a22oi_1 _29959_ (.Y(_07234_),
    .B1(net3330),
    .B2(_07229_),
    .A2(_06375_),
    .A1(net3367));
 sg13g2_xnor2_1 _29960_ (.Y(_07235_),
    .A(_06015_),
    .B(_07234_));
 sg13g2_a21oi_1 _29961_ (.A1(net4227),
    .A2(_07235_),
    .Y(_01175_),
    .B1(_07233_));
 sg13g2_nand3b_1 _29962_ (.B(_06284_),
    .C(_06297_),
    .Y(_07236_),
    .A_N(_06375_));
 sg13g2_nor4_1 _29963_ (.A(_07182_),
    .B(_07196_),
    .C(_07212_),
    .D(_07236_),
    .Y(_07237_));
 sg13g2_nor4_2 _29964_ (.A(_06015_),
    .B(_07003_),
    .C(_07029_),
    .Y(_07238_),
    .D(_07031_));
 sg13g2_nand4_1 _29965_ (.B(_07225_),
    .C(_07237_),
    .A(_07109_),
    .Y(_07239_),
    .D(_07238_));
 sg13g2_nor3_2 _29966_ (.A(_06966_),
    .B(_07177_),
    .C(_07239_),
    .Y(_07240_));
 sg13g2_or3_1 _29967_ (.A(_06966_),
    .B(_07177_),
    .C(_07239_),
    .X(_07241_));
 sg13g2_a21oi_1 _29968_ (.A1(net3370),
    .A2(_07240_),
    .Y(_07242_),
    .B1(net3343));
 sg13g2_xnor2_1 _29969_ (.Y(_07243_),
    .A(_06017_),
    .B(_07242_));
 sg13g2_nand2_1 _29970_ (.Y(_07244_),
    .A(net1334),
    .B(net4170));
 sg13g2_o21ai_1 _29971_ (.B1(_07244_),
    .Y(_01176_),
    .A1(net4169),
    .A2(_07243_));
 sg13g2_nor2_1 _29972_ (.A(net1672),
    .B(net4226),
    .Y(_07245_));
 sg13g2_nor2_1 _29973_ (.A(_06337_),
    .B(net3314),
    .Y(_07246_));
 sg13g2_nand3_1 _29974_ (.B(_06337_),
    .C(_07240_),
    .A(_06017_),
    .Y(_07247_));
 sg13g2_a21o_1 _29975_ (.A2(_07240_),
    .A1(_06017_),
    .B1(_06337_),
    .X(_07248_));
 sg13g2_a21oi_1 _29976_ (.A1(_07247_),
    .A2(_07248_),
    .Y(_07249_),
    .B1(net3389));
 sg13g2_nor2_1 _29977_ (.A(_07246_),
    .B(_07249_),
    .Y(_07250_));
 sg13g2_a21oi_1 _29978_ (.A1(net4219),
    .A2(_07250_),
    .Y(_01177_),
    .B1(_07245_));
 sg13g2_nor2_1 _29979_ (.A(net1664),
    .B(net4223),
    .Y(_07251_));
 sg13g2_a21oi_1 _29980_ (.A1(net3370),
    .A2(_07247_),
    .Y(_07252_),
    .B1(net3326));
 sg13g2_xnor2_1 _29981_ (.Y(_07253_),
    .A(_06305_),
    .B(_07252_));
 sg13g2_a21oi_1 _29982_ (.A1(net4223),
    .A2(_07253_),
    .Y(_01178_),
    .B1(_07251_));
 sg13g2_or2_1 _29983_ (.X(_07254_),
    .B(_07247_),
    .A(_06305_));
 sg13g2_nor2_1 _29984_ (.A(_06341_),
    .B(_07254_),
    .Y(_07255_));
 sg13g2_xnor2_1 _29985_ (.Y(_07256_),
    .A(_06341_),
    .B(_07254_));
 sg13g2_a221oi_1 _29986_ (.B2(net3369),
    .C1(net4168),
    .B1(_07256_),
    .A1(_06341_),
    .Y(_07257_),
    .A2(net3326));
 sg13g2_a21oi_1 _29987_ (.A1(_11011_),
    .A2(net4168),
    .Y(_01179_),
    .B1(_07257_));
 sg13g2_nor2_1 _29988_ (.A(net1166),
    .B(net4221),
    .Y(_07258_));
 sg13g2_a21oi_1 _29989_ (.A1(net3369),
    .A2(_07255_),
    .Y(_07259_),
    .B1(net3342));
 sg13g2_xnor2_1 _29990_ (.Y(_07260_),
    .A(_06339_),
    .B(_07259_));
 sg13g2_a21oi_1 _29991_ (.A1(net4220),
    .A2(_07260_),
    .Y(_01180_),
    .B1(_07258_));
 sg13g2_nand2_1 _29992_ (.Y(_07261_),
    .A(_06339_),
    .B(_07255_));
 sg13g2_nor2_1 _29993_ (.A(_06417_),
    .B(_07261_),
    .Y(_07262_));
 sg13g2_xnor2_1 _29994_ (.Y(_07263_),
    .A(_06417_),
    .B(_07261_));
 sg13g2_a221oi_1 _29995_ (.B2(net3368),
    .C1(net4168),
    .B1(_07263_),
    .A1(_06417_),
    .Y(_07264_),
    .A2(net3326));
 sg13g2_a21oi_1 _29996_ (.A1(_11012_),
    .A2(net4166),
    .Y(_01181_),
    .B1(_07264_));
 sg13g2_nor2_1 _29997_ (.A(net1176),
    .B(net4222),
    .Y(_07265_));
 sg13g2_o21ai_1 _29998_ (.B1(net3314),
    .Y(_07266_),
    .A1(net3390),
    .A2(_07262_));
 sg13g2_xnor2_1 _29999_ (.Y(_07267_),
    .A(_06421_),
    .B(_07266_));
 sg13g2_a21oi_1 _30000_ (.A1(net4222),
    .A2(_07267_),
    .Y(_01182_),
    .B1(_07265_));
 sg13g2_nor2_1 _30001_ (.A(net1611),
    .B(net4220),
    .Y(_07268_));
 sg13g2_xnor2_1 _30002_ (.Y(_07269_),
    .A(net3390),
    .B(_06421_));
 sg13g2_nor2_1 _30003_ (.A(_07266_),
    .B(_07269_),
    .Y(_07270_));
 sg13g2_xor2_1 _30004_ (.B(_07270_),
    .A(_06411_),
    .X(_07271_));
 sg13g2_a21oi_1 _30005_ (.A1(net4220),
    .A2(_07271_),
    .Y(_01183_),
    .B1(_07268_));
 sg13g2_and4_1 _30006_ (.A(_06339_),
    .B(_06411_),
    .C(_06418_),
    .D(_06421_),
    .X(_07272_));
 sg13g2_and2_1 _30007_ (.A(_07255_),
    .B(_07272_),
    .X(_07273_));
 sg13g2_a21oi_1 _30008_ (.A1(net3369),
    .A2(_07273_),
    .Y(_07274_),
    .B1(net3342));
 sg13g2_nand2_1 _30009_ (.Y(_07275_),
    .A(_06413_),
    .B(_07273_));
 sg13g2_xnor2_1 _30010_ (.Y(_07276_),
    .A(_06413_),
    .B(_07274_));
 sg13g2_nand2_1 _30011_ (.Y(_07277_),
    .A(net1363),
    .B(net4168));
 sg13g2_o21ai_1 _30012_ (.B1(_07277_),
    .Y(_01184_),
    .A1(net4168),
    .A2(_07276_));
 sg13g2_or2_1 _30013_ (.X(_07278_),
    .B(_07275_),
    .A(_05993_));
 sg13g2_xnor2_1 _30014_ (.Y(_07279_),
    .A(_05993_),
    .B(_07275_));
 sg13g2_a221oi_1 _30015_ (.B2(net3369),
    .C1(net4168),
    .B1(_07279_),
    .A1(_05993_),
    .Y(_07280_),
    .A2(net3326));
 sg13g2_a21oi_1 _30016_ (.A1(_11013_),
    .A2(net4168),
    .Y(_01185_),
    .B1(_07280_));
 sg13g2_nor2_1 _30017_ (.A(net1458),
    .B(net4224),
    .Y(_07281_));
 sg13g2_a21oi_1 _30018_ (.A1(net3369),
    .A2(_07278_),
    .Y(_07282_),
    .B1(net3326));
 sg13g2_xnor2_1 _30019_ (.Y(_07283_),
    .A(_05958_),
    .B(_07282_));
 sg13g2_a21oi_1 _30020_ (.A1(net4223),
    .A2(_07283_),
    .Y(_01186_),
    .B1(_07281_));
 sg13g2_nor2_1 _30021_ (.A(net1576),
    .B(net4224),
    .Y(_07284_));
 sg13g2_nor3_1 _30022_ (.A(net3390),
    .B(_05958_),
    .C(_07278_),
    .Y(_07285_));
 sg13g2_nor2_1 _30023_ (.A(net3342),
    .B(_07285_),
    .Y(_07286_));
 sg13g2_xnor2_1 _30024_ (.Y(_07287_),
    .A(_05967_),
    .B(_07286_));
 sg13g2_a21oi_1 _30025_ (.A1(net4223),
    .A2(_07287_),
    .Y(_01187_),
    .B1(_07284_));
 sg13g2_nor2_1 _30026_ (.A(net1263),
    .B(net4220),
    .Y(_07288_));
 sg13g2_nand2_1 _30027_ (.Y(_07289_),
    .A(_05959_),
    .B(_05967_));
 sg13g2_nor2_1 _30028_ (.A(_07278_),
    .B(_07289_),
    .Y(_07290_));
 sg13g2_a21oi_1 _30029_ (.A1(net3368),
    .A2(_07290_),
    .Y(_07291_),
    .B1(net3342));
 sg13g2_xnor2_1 _30030_ (.Y(_07292_),
    .A(_05970_),
    .B(_07291_));
 sg13g2_a21oi_1 _30031_ (.A1(net4221),
    .A2(_07292_),
    .Y(_01188_),
    .B1(_07288_));
 sg13g2_nand2_1 _30032_ (.Y(_07293_),
    .A(_05970_),
    .B(_05988_));
 sg13g2_nand3_1 _30033_ (.B(_05988_),
    .C(_07290_),
    .A(_05970_),
    .Y(_07294_));
 sg13g2_a21o_1 _30034_ (.A2(_07290_),
    .A1(_05970_),
    .B1(_05988_),
    .X(_07295_));
 sg13g2_nand2_1 _30035_ (.Y(_07296_),
    .A(_07294_),
    .B(_07295_));
 sg13g2_o21ai_1 _30036_ (.B1(net4225),
    .Y(_07297_),
    .A1(_05988_),
    .A2(net3314));
 sg13g2_a21oi_1 _30037_ (.A1(net3368),
    .A2(_07296_),
    .Y(_07298_),
    .B1(_07297_));
 sg13g2_a21oi_1 _30038_ (.A1(_11014_),
    .A2(net4166),
    .Y(_01189_),
    .B1(_07298_));
 sg13g2_nor2_1 _30039_ (.A(net1553),
    .B(net4220),
    .Y(_07299_));
 sg13g2_a21oi_1 _30040_ (.A1(net3368),
    .A2(_07294_),
    .Y(_07300_),
    .B1(net3326));
 sg13g2_xor2_1 _30041_ (.B(_07300_),
    .A(_05972_),
    .X(_07301_));
 sg13g2_a21oi_1 _30042_ (.A1(net4222),
    .A2(_07301_),
    .Y(_01190_),
    .B1(_07299_));
 sg13g2_nor2_1 _30043_ (.A(net1918),
    .B(net4219),
    .Y(_07302_));
 sg13g2_xnor2_1 _30044_ (.Y(_07303_),
    .A(net3368),
    .B(_05972_));
 sg13g2_nand2_1 _30045_ (.Y(_07304_),
    .A(_07300_),
    .B(_07303_));
 sg13g2_xnor2_1 _30046_ (.Y(_07305_),
    .A(_06559_),
    .B(_07304_));
 sg13g2_a21oi_1 _30047_ (.A1(net4219),
    .A2(_07305_),
    .Y(_01191_),
    .B1(_07302_));
 sg13g2_nor2_1 _30048_ (.A(net1566),
    .B(net4222),
    .Y(_07306_));
 sg13g2_nand4_1 _30049_ (.B(_06017_),
    .C(_06337_),
    .A(_05972_),
    .Y(_07307_),
    .D(_06413_));
 sg13g2_or3_1 _30050_ (.A(_07289_),
    .B(_07293_),
    .C(_07307_),
    .X(_07308_));
 sg13g2_nor3_1 _30051_ (.A(_05993_),
    .B(_06305_),
    .C(_06341_),
    .Y(_07309_));
 sg13g2_nand3_1 _30052_ (.B(_07272_),
    .C(_07309_),
    .A(_06559_),
    .Y(_07310_));
 sg13g2_or3_1 _30053_ (.A(_07241_),
    .B(_07308_),
    .C(_07310_),
    .X(_07311_));
 sg13g2_a21oi_1 _30054_ (.A1(net3368),
    .A2(_07311_),
    .Y(_07312_),
    .B1(net3326));
 sg13g2_nand2_1 _30055_ (.Y(_07313_),
    .A(_06467_),
    .B(_07312_));
 sg13g2_xor2_1 _30056_ (.B(_07312_),
    .A(_06467_),
    .X(_07314_));
 sg13g2_a21oi_1 _30057_ (.A1(net4222),
    .A2(_07314_),
    .Y(_01192_),
    .B1(_07306_));
 sg13g2_nor2_1 _30058_ (.A(_06469_),
    .B(net3342),
    .Y(_07315_));
 sg13g2_nand2_1 _30059_ (.Y(_07316_),
    .A(_06467_),
    .B(_06469_));
 sg13g2_nor3_1 _30060_ (.A(net3390),
    .B(_07311_),
    .C(_07316_),
    .Y(_07317_));
 sg13g2_or3_1 _30061_ (.A(net3390),
    .B(_07311_),
    .C(_07316_),
    .X(_07318_));
 sg13g2_a21oi_1 _30062_ (.A1(_07313_),
    .A2(_07315_),
    .Y(_07319_),
    .B1(net4166));
 sg13g2_a22oi_1 _30063_ (.Y(_01193_),
    .B1(_07318_),
    .B2(_07319_),
    .A2(net4166),
    .A1(_11015_));
 sg13g2_nor2_1 _30064_ (.A(net1352),
    .B(net4220),
    .Y(_07320_));
 sg13g2_nor2_1 _30065_ (.A(net3343),
    .B(_07317_),
    .Y(_07321_));
 sg13g2_xnor2_1 _30066_ (.Y(_07322_),
    .A(_06466_),
    .B(_07321_));
 sg13g2_a21oi_1 _30067_ (.A1(net4220),
    .A2(_07322_),
    .Y(_01194_),
    .B1(_07320_));
 sg13g2_nand2_1 _30068_ (.Y(_07323_),
    .A(_06424_),
    .B(_06466_));
 sg13g2_nor2_1 _30069_ (.A(_07316_),
    .B(_07323_),
    .Y(_07324_));
 sg13g2_nor2b_1 _30070_ (.A(_07311_),
    .B_N(_07324_),
    .Y(_07325_));
 sg13g2_o21ai_1 _30071_ (.B1(net3314),
    .Y(_07326_),
    .A1(net3390),
    .A2(_06466_));
 sg13g2_a21oi_1 _30072_ (.A1(_06470_),
    .A2(_07318_),
    .Y(_07327_),
    .B1(_07326_));
 sg13g2_xor2_1 _30073_ (.B(_07327_),
    .A(_06424_),
    .X(_07328_));
 sg13g2_nand2_1 _30074_ (.Y(_07329_),
    .A(net1224),
    .B(net4167));
 sg13g2_o21ai_1 _30075_ (.B1(_07329_),
    .Y(_01195_),
    .A1(net4166),
    .A2(_07328_));
 sg13g2_nor2_1 _30076_ (.A(net1431),
    .B(net4220),
    .Y(_07330_));
 sg13g2_a21oi_1 _30077_ (.A1(net3368),
    .A2(_07325_),
    .Y(_07331_),
    .B1(net3342));
 sg13g2_xnor2_1 _30078_ (.Y(_07332_),
    .A(_06419_),
    .B(_07331_));
 sg13g2_a21oi_1 _30079_ (.A1(net4221),
    .A2(_07332_),
    .Y(_01196_),
    .B1(_07330_));
 sg13g2_nand3_1 _30080_ (.B(_06474_),
    .C(_07325_),
    .A(_06419_),
    .Y(_07333_));
 sg13g2_a21o_1 _30081_ (.A2(_07325_),
    .A1(_06419_),
    .B1(_06474_),
    .X(_07334_));
 sg13g2_nand2_1 _30082_ (.Y(_07335_),
    .A(_07333_),
    .B(_07334_));
 sg13g2_a21oi_1 _30083_ (.A1(net3369),
    .A2(_07335_),
    .Y(_07336_),
    .B1(net4166));
 sg13g2_o21ai_1 _30084_ (.B1(_07336_),
    .Y(_07337_),
    .A1(_06474_),
    .A2(net3314));
 sg13g2_o21ai_1 _30085_ (.B1(_07337_),
    .Y(_07338_),
    .A1(net2556),
    .A2(net4219));
 sg13g2_inv_1 _30086_ (.Y(_01197_),
    .A(_07338_));
 sg13g2_nor2_1 _30087_ (.A(net1187),
    .B(net4219),
    .Y(_07339_));
 sg13g2_a21oi_1 _30088_ (.A1(net3369),
    .A2(_07333_),
    .Y(_07340_),
    .B1(net3326));
 sg13g2_xnor2_1 _30089_ (.Y(_07341_),
    .A(_05996_),
    .B(_07340_));
 sg13g2_a21oi_1 _30090_ (.A1(net4219),
    .A2(_07341_),
    .Y(_01198_),
    .B1(_07339_));
 sg13g2_nor2_1 _30091_ (.A(net1506),
    .B(net4219),
    .Y(_07342_));
 sg13g2_xnor2_1 _30092_ (.Y(_07343_),
    .A(net3368),
    .B(_05995_));
 sg13g2_nand2_1 _30093_ (.Y(_07344_),
    .A(_07340_),
    .B(_07343_));
 sg13g2_xnor2_1 _30094_ (.Y(_07345_),
    .A(_06412_),
    .B(_07344_));
 sg13g2_a21oi_1 _30095_ (.A1(net4219),
    .A2(_07345_),
    .Y(_01199_),
    .B1(_07342_));
 sg13g2_nor2_1 _30096_ (.A(net1484),
    .B(net4223),
    .Y(_07346_));
 sg13g2_nand4_1 _30097_ (.B(_06412_),
    .C(_06419_),
    .A(_05995_),
    .Y(_07347_),
    .D(_06474_));
 sg13g2_nor4_1 _30098_ (.A(_07311_),
    .B(_07316_),
    .C(_07323_),
    .D(_07347_),
    .Y(_07348_));
 sg13g2_a21oi_1 _30099_ (.A1(net3369),
    .A2(_07348_),
    .Y(_07349_),
    .B1(net3342));
 sg13g2_xnor2_1 _30100_ (.Y(_07350_),
    .A(_05982_),
    .B(_07349_));
 sg13g2_a21oi_1 _30101_ (.A1(net4223),
    .A2(_07350_),
    .Y(_01200_),
    .B1(_07346_));
 sg13g2_nand2_1 _30102_ (.Y(_07351_),
    .A(_05982_),
    .B(_07348_));
 sg13g2_o21ai_1 _30103_ (.B1(_06010_),
    .Y(_07352_),
    .A1(net3390),
    .A2(_07351_));
 sg13g2_or2_1 _30104_ (.X(_07353_),
    .B(_07352_),
    .A(net3342));
 sg13g2_nor2_1 _30105_ (.A(_06010_),
    .B(_07351_),
    .Y(_07354_));
 sg13g2_a21oi_1 _30106_ (.A1(net3370),
    .A2(_07354_),
    .Y(_07355_),
    .B1(net4167));
 sg13g2_a22oi_1 _30107_ (.Y(_01201_),
    .B1(_07353_),
    .B2(_07355_),
    .A2(net4167),
    .A1(_11016_));
 sg13g2_nor2_1 _30108_ (.A(net1613),
    .B(net4223),
    .Y(_07356_));
 sg13g2_o21ai_1 _30109_ (.B1(net3314),
    .Y(_07357_),
    .A1(net3389),
    .A2(_07354_));
 sg13g2_xnor2_1 _30110_ (.Y(_07358_),
    .A(_06450_),
    .B(_07357_));
 sg13g2_a21oi_1 _30111_ (.A1(net4225),
    .A2(_07358_),
    .Y(_01202_),
    .B1(_07356_));
 sg13g2_nand2b_1 _30112_ (.Y(_07359_),
    .B(_07357_),
    .A_N(_06452_));
 sg13g2_nand2_1 _30113_ (.Y(_07360_),
    .A(_06450_),
    .B(_06452_));
 sg13g2_nand3_1 _30114_ (.B(_06452_),
    .C(_07354_),
    .A(_06450_),
    .Y(_07361_));
 sg13g2_a21oi_1 _30115_ (.A1(_06453_),
    .A2(_07361_),
    .Y(_07362_),
    .B1(net3389));
 sg13g2_nor2_1 _30116_ (.A(net4166),
    .B(_07362_),
    .Y(_07363_));
 sg13g2_a22oi_1 _30117_ (.Y(_01203_),
    .B1(_07359_),
    .B2(_07363_),
    .A2(net4166),
    .A1(_11017_));
 sg13g2_nor2_1 _30118_ (.A(net1759),
    .B(net4229),
    .Y(_07364_));
 sg13g2_a21oi_1 _30119_ (.A1(net3371),
    .A2(_07361_),
    .Y(_07365_),
    .B1(net3327));
 sg13g2_xnor2_1 _30120_ (.Y(_07366_),
    .A(_06001_),
    .B(_07365_));
 sg13g2_a21oi_1 _30121_ (.A1(net4223),
    .A2(_07366_),
    .Y(_01204_),
    .B1(_07364_));
 sg13g2_nor2_1 _30122_ (.A(_06001_),
    .B(_07361_),
    .Y(_07367_));
 sg13g2_xnor2_1 _30123_ (.Y(_07368_),
    .A(_06491_),
    .B(_07367_));
 sg13g2_a21oi_1 _30124_ (.A1(net3370),
    .A2(_07368_),
    .Y(_07369_),
    .B1(net4167));
 sg13g2_o21ai_1 _30125_ (.B1(_07369_),
    .Y(_07370_),
    .A1(_06491_),
    .A2(net3314));
 sg13g2_o21ai_1 _30126_ (.B1(_07370_),
    .Y(_07371_),
    .A1(net2808),
    .A2(net4226));
 sg13g2_inv_1 _30127_ (.Y(_01205_),
    .A(_07371_));
 sg13g2_a21oi_1 _30128_ (.A1(_06491_),
    .A2(_07367_),
    .Y(_07372_),
    .B1(net3391));
 sg13g2_nor2_1 _30129_ (.A(net3327),
    .B(_07372_),
    .Y(_07373_));
 sg13g2_xor2_1 _30130_ (.B(_07373_),
    .A(_06481_),
    .X(_07374_));
 sg13g2_nor2_1 _30131_ (.A(net1457),
    .B(net4227),
    .Y(_07375_));
 sg13g2_a21oi_1 _30132_ (.A1(net4226),
    .A2(_07374_),
    .Y(_01206_),
    .B1(_07375_));
 sg13g2_nor2_1 _30133_ (.A(net1409),
    .B(net4229),
    .Y(_07376_));
 sg13g2_xnor2_1 _30134_ (.Y(_07377_),
    .A(net3370),
    .B(_06481_));
 sg13g2_nand2_1 _30135_ (.Y(_07378_),
    .A(_07373_),
    .B(_07377_));
 sg13g2_xnor2_1 _30136_ (.Y(_07379_),
    .A(_05981_),
    .B(_07378_));
 sg13g2_a21oi_1 _30137_ (.A1(net4229),
    .A2(_07379_),
    .Y(_01207_),
    .B1(_07376_));
 sg13g2_nor2_1 _30138_ (.A(net1373),
    .B(net4229),
    .Y(_07380_));
 sg13g2_nor2b_1 _30139_ (.A(_06010_),
    .B_N(_06481_),
    .Y(_07381_));
 sg13g2_nand2_1 _30140_ (.Y(_07382_),
    .A(_05981_),
    .B(_05982_));
 sg13g2_nor4_1 _30141_ (.A(_06001_),
    .B(_07347_),
    .C(_07360_),
    .D(_07382_),
    .Y(_07383_));
 sg13g2_nand4_1 _30142_ (.B(_07324_),
    .C(_07381_),
    .A(_06491_),
    .Y(_07384_),
    .D(_07383_));
 sg13g2_nor4_2 _30143_ (.A(_07241_),
    .B(_07308_),
    .C(_07310_),
    .Y(_07385_),
    .D(_07384_));
 sg13g2_a21oi_1 _30144_ (.A1(net3370),
    .A2(_07385_),
    .Y(_07386_),
    .B1(net3343));
 sg13g2_xnor2_1 _30145_ (.Y(_07387_),
    .A(_06414_),
    .B(_07386_));
 sg13g2_a21oi_1 _30146_ (.A1(net4229),
    .A2(_07387_),
    .Y(_01208_),
    .B1(_07380_));
 sg13g2_and2_1 _30147_ (.A(_05991_),
    .B(_06414_),
    .X(_07388_));
 sg13g2_and2_1 _30148_ (.A(_07385_),
    .B(_07388_),
    .X(_07389_));
 sg13g2_a21oi_1 _30149_ (.A1(_06414_),
    .A2(_07385_),
    .Y(_07390_),
    .B1(_05991_));
 sg13g2_or2_1 _30150_ (.X(_07391_),
    .B(_07390_),
    .A(_07389_));
 sg13g2_a21oi_1 _30151_ (.A1(net3370),
    .A2(_07391_),
    .Y(_07392_),
    .B1(net4169));
 sg13g2_o21ai_1 _30152_ (.B1(_07392_),
    .Y(_07393_),
    .A1(_05991_),
    .A2(net3315));
 sg13g2_o21ai_1 _30153_ (.B1(_07393_),
    .Y(_07394_),
    .A1(net2506),
    .A2(net4229));
 sg13g2_inv_1 _30154_ (.Y(_01209_),
    .A(_07394_));
 sg13g2_nor2_1 _30155_ (.A(net1448),
    .B(net4227),
    .Y(_07395_));
 sg13g2_o21ai_1 _30156_ (.B1(net3315),
    .Y(_07396_),
    .A1(net3389),
    .A2(_07389_));
 sg13g2_xnor2_1 _30157_ (.Y(_07397_),
    .A(_06003_),
    .B(_07396_));
 sg13g2_a21oi_1 _30158_ (.A1(net4226),
    .A2(_07397_),
    .Y(_01210_),
    .B1(_07395_));
 sg13g2_nand2b_1 _30159_ (.Y(_07398_),
    .B(_07396_),
    .A_N(_06004_));
 sg13g2_nand4_1 _30160_ (.B(_06004_),
    .C(_07385_),
    .A(_06003_),
    .Y(_07399_),
    .D(_07388_));
 sg13g2_nand2_1 _30161_ (.Y(_07400_),
    .A(_06005_),
    .B(_07399_));
 sg13g2_a21oi_1 _30162_ (.A1(net3370),
    .A2(_07400_),
    .Y(_07401_),
    .B1(net4169));
 sg13g2_a22oi_1 _30163_ (.Y(_01211_),
    .B1(_07398_),
    .B2(_07401_),
    .A2(net4169),
    .A1(_11018_));
 sg13g2_nor2_1 _30164_ (.A(net1309),
    .B(net4226),
    .Y(_07402_));
 sg13g2_a21oi_1 _30165_ (.A1(net3371),
    .A2(_07399_),
    .Y(_07403_),
    .B1(net3327));
 sg13g2_xor2_1 _30166_ (.B(_07403_),
    .A(_05940_),
    .X(_07404_));
 sg13g2_a21oi_1 _30167_ (.A1(net4226),
    .A2(_07404_),
    .Y(_01212_),
    .B1(_07402_));
 sg13g2_nand2_1 _30168_ (.Y(_07405_),
    .A(_05939_),
    .B(_05940_));
 sg13g2_nor2_1 _30169_ (.A(_07399_),
    .B(_07405_),
    .Y(_07406_));
 sg13g2_or2_1 _30170_ (.X(_07407_),
    .B(_07406_),
    .A(_05941_));
 sg13g2_a21oi_1 _30171_ (.A1(net3371),
    .A2(_07407_),
    .Y(_07408_),
    .B1(net4169));
 sg13g2_o21ai_1 _30172_ (.B1(_07408_),
    .Y(_07409_),
    .A1(_05939_),
    .A2(_07403_));
 sg13g2_o21ai_1 _30173_ (.B1(_07409_),
    .Y(_07410_),
    .A1(net2609),
    .A2(net4226));
 sg13g2_inv_1 _30174_ (.Y(_01213_),
    .A(_07410_));
 sg13g2_o21ai_1 _30175_ (.B1(net3371),
    .Y(_07411_),
    .A1(_07399_),
    .A2(_07405_));
 sg13g2_nand2_1 _30176_ (.Y(_07412_),
    .A(net3314),
    .B(_07411_));
 sg13g2_xnor2_1 _30177_ (.Y(_07413_),
    .A(_06561_),
    .B(_07412_));
 sg13g2_nand2_1 _30178_ (.Y(_07414_),
    .A(net1096),
    .B(net4170));
 sg13g2_o21ai_1 _30179_ (.B1(_07414_),
    .Y(_01214_),
    .A1(net4170),
    .A2(_07413_));
 sg13g2_nor2_1 _30180_ (.A(net1445),
    .B(net4228),
    .Y(_07415_));
 sg13g2_xnor2_1 _30181_ (.Y(_07416_),
    .A(net3389),
    .B(_06561_));
 sg13g2_nor2_1 _30182_ (.A(_07412_),
    .B(_07416_),
    .Y(_07417_));
 sg13g2_xor2_1 _30183_ (.B(_07417_),
    .A(_06576_),
    .X(_07418_));
 sg13g2_a21oi_1 _30184_ (.A1(net4228),
    .A2(_07418_),
    .Y(_01215_),
    .B1(_07415_));
 sg13g2_nor2_1 _30185_ (.A(net1240),
    .B(net4228),
    .Y(_07419_));
 sg13g2_nand4_1 _30186_ (.B(_06004_),
    .C(_06561_),
    .A(_06003_),
    .Y(_07420_),
    .D(_07388_));
 sg13g2_nor2_1 _30187_ (.A(_07405_),
    .B(_07420_),
    .Y(_07421_));
 sg13g2_and2_1 _30188_ (.A(_06576_),
    .B(_07421_),
    .X(_07422_));
 sg13g2_a21oi_1 _30189_ (.A1(_07385_),
    .A2(_07422_),
    .Y(_07423_),
    .B1(net3389));
 sg13g2_nor2_1 _30190_ (.A(net3327),
    .B(_07423_),
    .Y(_07424_));
 sg13g2_xor2_1 _30191_ (.B(_07424_),
    .A(_05962_),
    .X(_07425_));
 sg13g2_a21oi_1 _30192_ (.A1(net4228),
    .A2(_07425_),
    .Y(_01216_),
    .B1(_07419_));
 sg13g2_and3_2 _30193_ (.X(_07426_),
    .A(_05962_),
    .B(_07385_),
    .C(_07422_));
 sg13g2_a21o_1 _30194_ (.A2(_07426_),
    .A1(net3372),
    .B1(_06472_),
    .X(_07427_));
 sg13g2_and3_1 _30195_ (.X(_07428_),
    .A(net3372),
    .B(_06472_),
    .C(_07426_));
 sg13g2_nor2_1 _30196_ (.A(net4169),
    .B(_07428_),
    .Y(_07429_));
 sg13g2_o21ai_1 _30197_ (.B1(_07429_),
    .Y(_07430_),
    .A1(net3343),
    .A2(_07427_));
 sg13g2_o21ai_1 _30198_ (.B1(_07430_),
    .Y(_07431_),
    .A1(net2330),
    .A2(net4230));
 sg13g2_inv_1 _30199_ (.Y(_01217_),
    .A(_07431_));
 sg13g2_nor2_1 _30200_ (.A(net3343),
    .B(_07428_),
    .Y(_07432_));
 sg13g2_xnor2_1 _30201_ (.Y(_07433_),
    .A(_06476_),
    .B(_07432_));
 sg13g2_nand2_1 _30202_ (.Y(_07434_),
    .A(net1093),
    .B(net4169));
 sg13g2_o21ai_1 _30203_ (.B1(_07434_),
    .Y(_01218_),
    .A1(net4169),
    .A2(_07433_));
 sg13g2_a21oi_1 _30204_ (.A1(_06476_),
    .A2(_07428_),
    .Y(_07435_),
    .B1(_06494_));
 sg13g2_and4_1 _30205_ (.A(_06472_),
    .B(_06476_),
    .C(_06494_),
    .D(_07426_),
    .X(_07436_));
 sg13g2_a221oi_1 _30206_ (.B2(net3372),
    .C1(net4172),
    .B1(_07436_),
    .A1(net3330),
    .Y(_07437_),
    .A2(_07435_));
 sg13g2_a21oi_1 _30207_ (.A1(_11019_),
    .A2(net4172),
    .Y(_01219_),
    .B1(_07437_));
 sg13g2_o21ai_1 _30208_ (.B1(net3315),
    .Y(_07438_),
    .A1(net3389),
    .A2(_07436_));
 sg13g2_xnor2_1 _30209_ (.Y(_07439_),
    .A(_06445_),
    .B(_07438_));
 sg13g2_nand2_1 _30210_ (.Y(_07440_),
    .A(net1085),
    .B(net4170));
 sg13g2_o21ai_1 _30211_ (.B1(_07440_),
    .Y(_01220_),
    .A1(net4170),
    .A2(_07439_));
 sg13g2_nand2b_1 _30212_ (.Y(_07441_),
    .B(_07438_),
    .A_N(_06444_));
 sg13g2_and4_1 _30213_ (.A(_06444_),
    .B(_06445_),
    .C(_06476_),
    .D(_06494_),
    .X(_07442_));
 sg13g2_nand3_1 _30214_ (.B(_07426_),
    .C(_07442_),
    .A(_06472_),
    .Y(_07443_));
 sg13g2_a21oi_1 _30215_ (.A1(_06446_),
    .A2(_07443_),
    .Y(_07444_),
    .B1(net3389));
 sg13g2_nor2_1 _30216_ (.A(net4172),
    .B(_07444_),
    .Y(_07445_));
 sg13g2_a22oi_1 _30217_ (.Y(_01221_),
    .B1(_07441_),
    .B2(_07445_),
    .A2(net4172),
    .A1(_11020_));
 sg13g2_nor2_1 _30218_ (.A(net1308),
    .B(net4230),
    .Y(_07446_));
 sg13g2_a21oi_1 _30219_ (.A1(net3372),
    .A2(_07443_),
    .Y(_07447_),
    .B1(net3327));
 sg13g2_xor2_1 _30220_ (.B(_07447_),
    .A(_06489_),
    .X(_07448_));
 sg13g2_a21oi_1 _30221_ (.A1(net4230),
    .A2(_07448_),
    .Y(_01222_),
    .B1(_07446_));
 sg13g2_nor2_1 _30222_ (.A(net1411),
    .B(net4230),
    .Y(_07449_));
 sg13g2_xnor2_1 _30223_ (.Y(_07450_),
    .A(net3372),
    .B(_06489_));
 sg13g2_nand2_1 _30224_ (.Y(_07451_),
    .A(_07447_),
    .B(_07450_));
 sg13g2_xnor2_1 _30225_ (.Y(_07452_),
    .A(_06484_),
    .B(_07451_));
 sg13g2_a21oi_1 _30226_ (.A1(net4230),
    .A2(_07452_),
    .Y(_01223_),
    .B1(_07449_));
 sg13g2_and4_1 _30227_ (.A(_05962_),
    .B(_06472_),
    .C(_06484_),
    .D(_06489_),
    .X(_07453_));
 sg13g2_and4_1 _30228_ (.A(_07385_),
    .B(_07422_),
    .C(_07442_),
    .D(_07453_),
    .X(_07454_));
 sg13g2_mux2_1 _30229_ (.A0(net3344),
    .A1(_07454_),
    .S(net3367),
    .X(_07455_));
 sg13g2_xnor2_1 _30230_ (.Y(_07456_),
    .A(_05964_),
    .B(_07455_));
 sg13g2_mux2_1 _30231_ (.A0(net2080),
    .A1(_07456_),
    .S(net4217),
    .X(_01224_));
 sg13g2_and2_1 _30232_ (.A(_05964_),
    .B(_07454_),
    .X(_07457_));
 sg13g2_nand2_1 _30233_ (.Y(_07458_),
    .A(_06479_),
    .B(_07457_));
 sg13g2_xnor2_1 _30234_ (.Y(_07459_),
    .A(_06479_),
    .B(_07457_));
 sg13g2_a21oi_1 _30235_ (.A1(net3373),
    .A2(_07459_),
    .Y(_07460_),
    .B1(net4165));
 sg13g2_o21ai_1 _30236_ (.B1(_07460_),
    .Y(_07461_),
    .A1(_06479_),
    .A2(net3315));
 sg13g2_o21ai_1 _30237_ (.B1(_07461_),
    .Y(_07462_),
    .A1(net2491),
    .A2(net4216));
 sg13g2_inv_1 _30238_ (.Y(_01225_),
    .A(_07462_));
 sg13g2_nor2_1 _30239_ (.A(net1543),
    .B(net4216),
    .Y(_07463_));
 sg13g2_a21oi_1 _30240_ (.A1(net3373),
    .A2(_07458_),
    .Y(_07464_),
    .B1(net3325));
 sg13g2_xnor2_1 _30241_ (.Y(_07465_),
    .A(_06008_),
    .B(_07464_));
 sg13g2_a21oi_1 _30242_ (.A1(net4217),
    .A2(_07465_),
    .Y(_01226_),
    .B1(_07463_));
 sg13g2_nor2_1 _30243_ (.A(_06008_),
    .B(_07458_),
    .Y(_07466_));
 sg13g2_a21oi_1 _30244_ (.A1(net3367),
    .A2(_07466_),
    .Y(_07467_),
    .B1(_06555_));
 sg13g2_and2_1 _30245_ (.A(_06555_),
    .B(_07466_),
    .X(_07468_));
 sg13g2_a221oi_1 _30246_ (.B2(net3367),
    .C1(net4165),
    .B1(_07468_),
    .A1(net3330),
    .Y(_07469_),
    .A2(_07467_));
 sg13g2_a21oi_1 _30247_ (.A1(_11021_),
    .A2(net4164),
    .Y(_01227_),
    .B1(_07469_));
 sg13g2_nor2_1 _30248_ (.A(net1410),
    .B(net4216),
    .Y(_07470_));
 sg13g2_a21oi_1 _30249_ (.A1(_06555_),
    .A2(_07466_),
    .Y(_07471_),
    .B1(net3391));
 sg13g2_nor2_1 _30250_ (.A(net3325),
    .B(_07471_),
    .Y(_07472_));
 sg13g2_xnor2_1 _30251_ (.Y(_07473_),
    .A(_05928_),
    .B(_07472_));
 sg13g2_a21oi_1 _30252_ (.A1(net4216),
    .A2(_07473_),
    .Y(_01228_),
    .B1(_07470_));
 sg13g2_o21ai_1 _30253_ (.B1(_05927_),
    .Y(_07474_),
    .A1(net3325),
    .A2(_07471_));
 sg13g2_nor2_1 _30254_ (.A(_05927_),
    .B(_06008_),
    .Y(_07475_));
 sg13g2_nand3b_1 _30255_ (.B(_06555_),
    .C(_07475_),
    .Y(_07476_),
    .A_N(_05928_));
 sg13g2_or2_1 _30256_ (.X(_07477_),
    .B(_07476_),
    .A(_07458_));
 sg13g2_a21oi_1 _30257_ (.A1(_05929_),
    .A2(_07477_),
    .Y(_07478_),
    .B1(net3391));
 sg13g2_nor2_1 _30258_ (.A(net4164),
    .B(_07478_),
    .Y(_07479_));
 sg13g2_a22oi_1 _30259_ (.Y(_01229_),
    .B1(_07474_),
    .B2(_07479_),
    .A2(net4164),
    .A1(_11022_));
 sg13g2_a21oi_1 _30260_ (.A1(net3366),
    .A2(_07477_),
    .Y(_07480_),
    .B1(net3328));
 sg13g2_xor2_1 _30261_ (.B(_07480_),
    .A(_05985_),
    .X(_07481_));
 sg13g2_nor2_1 _30262_ (.A(net1416),
    .B(net4216),
    .Y(_07482_));
 sg13g2_a21oi_1 _30263_ (.A1(net4216),
    .A2(_07481_),
    .Y(_01230_),
    .B1(_07482_));
 sg13g2_nor2_1 _30264_ (.A(net1400),
    .B(net4216),
    .Y(_07483_));
 sg13g2_xnor2_1 _30265_ (.Y(_07484_),
    .A(net3366),
    .B(_05985_));
 sg13g2_nand2_1 _30266_ (.Y(_07485_),
    .A(_07480_),
    .B(_07484_));
 sg13g2_xnor2_1 _30267_ (.Y(_07486_),
    .A(_06557_),
    .B(_07485_));
 sg13g2_a21oi_1 _30268_ (.A1(net4216),
    .A2(_07486_),
    .Y(_01231_),
    .B1(_07483_));
 sg13g2_nor2_1 _30269_ (.A(net1338),
    .B(net4218),
    .Y(_07487_));
 sg13g2_nand2_1 _30270_ (.Y(_07488_),
    .A(_05985_),
    .B(_06557_));
 sg13g2_nor2_1 _30271_ (.A(_07477_),
    .B(_07488_),
    .Y(_07489_));
 sg13g2_a21oi_1 _30272_ (.A1(net3365),
    .A2(_07489_),
    .Y(_07490_),
    .B1(net3344));
 sg13g2_xnor2_1 _30273_ (.Y(_07491_),
    .A(_06435_),
    .B(_07490_));
 sg13g2_a21oi_1 _30274_ (.A1(net4218),
    .A2(_07491_),
    .Y(_01232_),
    .B1(_07487_));
 sg13g2_nor2_1 _30275_ (.A(net1293),
    .B(net4214),
    .Y(_07492_));
 sg13g2_nand2_1 _30276_ (.Y(_07493_),
    .A(_06435_),
    .B(_07489_));
 sg13g2_nor2_2 _30277_ (.A(_05934_),
    .B(_07493_),
    .Y(_07494_));
 sg13g2_xnor2_1 _30278_ (.Y(_07495_),
    .A(_05934_),
    .B(_07493_));
 sg13g2_a22oi_1 _30279_ (.Y(_07496_),
    .B1(_07495_),
    .B2(net3365),
    .A2(net3325),
    .A1(_05934_));
 sg13g2_a21oi_1 _30280_ (.A1(net4215),
    .A2(_07496_),
    .Y(_01233_),
    .B1(_07492_));
 sg13g2_nor2_1 _30281_ (.A(net1535),
    .B(net4213),
    .Y(_07497_));
 sg13g2_o21ai_1 _30282_ (.B1(net3316),
    .Y(_07498_),
    .A1(net3387),
    .A2(_07494_));
 sg13g2_xnor2_1 _30283_ (.Y(_07499_),
    .A(_06465_),
    .B(_07498_));
 sg13g2_a21oi_1 _30284_ (.A1(net4212),
    .A2(_07499_),
    .Y(_01234_),
    .B1(_07497_));
 sg13g2_and2_1 _30285_ (.A(_05948_),
    .B(_06465_),
    .X(_07500_));
 sg13g2_nand2_1 _30286_ (.Y(_07501_),
    .A(_07494_),
    .B(_07500_));
 sg13g2_a21oi_1 _30287_ (.A1(_06465_),
    .A2(_07494_),
    .Y(_07502_),
    .B1(_05948_));
 sg13g2_a21o_1 _30288_ (.A2(_07500_),
    .A1(_07494_),
    .B1(_07502_),
    .X(_07503_));
 sg13g2_a221oi_1 _30289_ (.B2(net3365),
    .C1(net4162),
    .B1(_07503_),
    .A1(_05947_),
    .Y(_07504_),
    .A2(net3325));
 sg13g2_a21oi_1 _30290_ (.A1(_11023_),
    .A2(net4165),
    .Y(_01235_),
    .B1(_07504_));
 sg13g2_nor2_1 _30291_ (.A(net1467),
    .B(net4212),
    .Y(_07505_));
 sg13g2_a21oi_1 _30292_ (.A1(net3363),
    .A2(_07501_),
    .Y(_07506_),
    .B1(net3329));
 sg13g2_xnor2_1 _30293_ (.Y(_07507_),
    .A(_06461_),
    .B(_07506_));
 sg13g2_a21oi_1 _30294_ (.A1(net4212),
    .A2(_07507_),
    .Y(_01236_),
    .B1(_07505_));
 sg13g2_nor2_1 _30295_ (.A(_06461_),
    .B(_07501_),
    .Y(_07508_));
 sg13g2_nor2_1 _30296_ (.A(_05951_),
    .B(_06461_),
    .Y(_07509_));
 sg13g2_xor2_1 _30297_ (.B(_07508_),
    .A(_05951_),
    .X(_07510_));
 sg13g2_a221oi_1 _30298_ (.B2(net3365),
    .C1(net4162),
    .B1(_07510_),
    .A1(_05951_),
    .Y(_07511_),
    .A2(net3325));
 sg13g2_a21oi_1 _30299_ (.A1(_11024_),
    .A2(net4162),
    .Y(_01237_),
    .B1(_07511_));
 sg13g2_nor2_1 _30300_ (.A(net1290),
    .B(net4218),
    .Y(_07512_));
 sg13g2_nand4_1 _30301_ (.B(_07494_),
    .C(_07500_),
    .A(net3365),
    .Y(_07513_),
    .D(_07509_));
 sg13g2_nand2_1 _30302_ (.Y(_07514_),
    .A(net3331),
    .B(_07513_));
 sg13g2_xnor2_1 _30303_ (.Y(_07515_),
    .A(_06544_),
    .B(_07514_));
 sg13g2_a21oi_1 _30304_ (.A1(net4218),
    .A2(_07515_),
    .Y(_01238_),
    .B1(_07512_));
 sg13g2_nor2_1 _30305_ (.A(net1656),
    .B(net4218),
    .Y(_07516_));
 sg13g2_a22oi_1 _30306_ (.Y(_07517_),
    .B1(net3331),
    .B2(_07513_),
    .A2(_06544_),
    .A1(net3365));
 sg13g2_xnor2_1 _30307_ (.Y(_07518_),
    .A(_06487_),
    .B(_07517_));
 sg13g2_a21oi_1 _30308_ (.A1(net4218),
    .A2(_07518_),
    .Y(_01239_),
    .B1(_07516_));
 sg13g2_nand3_1 _30309_ (.B(_06435_),
    .C(_06479_),
    .A(_05964_),
    .Y(_07519_));
 sg13g2_nor2_1 _30310_ (.A(_06544_),
    .B(_07476_),
    .Y(_07520_));
 sg13g2_nand2b_1 _30311_ (.Y(_07521_),
    .B(_07500_),
    .A_N(_07488_));
 sg13g2_nor4_1 _30312_ (.A(_05934_),
    .B(_06487_),
    .C(_07519_),
    .D(_07521_),
    .Y(_07522_));
 sg13g2_and4_1 _30313_ (.A(_07454_),
    .B(_07509_),
    .C(_07520_),
    .D(_07522_),
    .X(_07523_));
 sg13g2_a21oi_1 _30314_ (.A1(net3360),
    .A2(_07523_),
    .Y(_07524_),
    .B1(_06482_));
 sg13g2_and3_1 _30315_ (.X(_07525_),
    .A(net3359),
    .B(_06482_),
    .C(_07523_));
 sg13g2_nand2_1 _30316_ (.Y(_07526_),
    .A(_06482_),
    .B(_07523_));
 sg13g2_nor2_1 _30317_ (.A(net3384),
    .B(_07526_),
    .Y(_07527_));
 sg13g2_nand2b_1 _30318_ (.Y(_07528_),
    .B(net4202),
    .A_N(_07525_));
 sg13g2_a21oi_1 _30319_ (.A1(net3330),
    .A2(_07524_),
    .Y(_07529_),
    .B1(_07528_));
 sg13g2_a21oi_1 _30320_ (.A1(_11025_),
    .A2(net4158),
    .Y(_01240_),
    .B1(_07529_));
 sg13g2_nor2_1 _30321_ (.A(_06448_),
    .B(_07525_),
    .Y(_07530_));
 sg13g2_a22oi_1 _30322_ (.Y(_07531_),
    .B1(_07530_),
    .B2(net3330),
    .A2(_07527_),
    .A1(_06448_));
 sg13g2_nand2_1 _30323_ (.Y(_07532_),
    .A(net1084),
    .B(net4158));
 sg13g2_o21ai_1 _30324_ (.B1(_07532_),
    .Y(_01241_),
    .A1(net4160),
    .A2(_07531_));
 sg13g2_nor2_1 _30325_ (.A(net1468),
    .B(net4205),
    .Y(_07533_));
 sg13g2_a21oi_1 _30326_ (.A1(_06448_),
    .A2(_07525_),
    .Y(_07534_),
    .B1(net3341));
 sg13g2_xnor2_1 _30327_ (.Y(_07535_),
    .A(_06431_),
    .B(_07534_));
 sg13g2_a21oi_1 _30328_ (.A1(net4205),
    .A2(_07535_),
    .Y(_01242_),
    .B1(_07533_));
 sg13g2_nand2_1 _30329_ (.Y(_07536_),
    .A(net1145),
    .B(net4159));
 sg13g2_nand2_1 _30330_ (.Y(_07537_),
    .A(_06431_),
    .B(_06448_));
 sg13g2_nor2b_1 _30331_ (.A(_07537_),
    .B_N(_06482_),
    .Y(_07538_));
 sg13g2_o21ai_1 _30332_ (.B1(_06439_),
    .Y(_07539_),
    .A1(_07526_),
    .A2(_07537_));
 sg13g2_nor3_1 _30333_ (.A(_06439_),
    .B(_07526_),
    .C(_07537_),
    .Y(_07540_));
 sg13g2_nor2_1 _30334_ (.A(net3385),
    .B(_07540_),
    .Y(_07541_));
 sg13g2_o21ai_1 _30335_ (.B1(net4203),
    .Y(_07542_),
    .A1(net3359),
    .A2(_06439_));
 sg13g2_a21o_1 _30336_ (.A2(_07541_),
    .A1(_07539_),
    .B1(_07542_),
    .X(_07543_));
 sg13g2_o21ai_1 _30337_ (.B1(_07536_),
    .Y(_01243_),
    .A1(net3341),
    .A2(_07543_));
 sg13g2_nor2_1 _30338_ (.A(net1497),
    .B(net4202),
    .Y(_07544_));
 sg13g2_nor2_1 _30339_ (.A(net3324),
    .B(_07541_),
    .Y(_07545_));
 sg13g2_xor2_1 _30340_ (.B(_07545_),
    .A(_06549_),
    .X(_07546_));
 sg13g2_a21oi_1 _30341_ (.A1(net4202),
    .A2(_07546_),
    .Y(_01244_),
    .B1(_07544_));
 sg13g2_nand3_1 _30342_ (.B(_06549_),
    .C(_07540_),
    .A(_06548_),
    .Y(_07547_));
 sg13g2_nand2b_1 _30343_ (.Y(_07548_),
    .B(_07547_),
    .A_N(_06550_));
 sg13g2_a21oi_1 _30344_ (.A1(net3359),
    .A2(_07548_),
    .Y(_07549_),
    .B1(net4160));
 sg13g2_o21ai_1 _30345_ (.B1(_07549_),
    .Y(_07550_),
    .A1(_06548_),
    .A2(_07545_));
 sg13g2_o21ai_1 _30346_ (.B1(_07550_),
    .Y(_07551_),
    .A1(net2577),
    .A2(net4202));
 sg13g2_inv_1 _30347_ (.Y(_01245_),
    .A(_07551_));
 sg13g2_nor2_1 _30348_ (.A(net1349),
    .B(net4202),
    .Y(_07552_));
 sg13g2_a21o_1 _30349_ (.A2(_07547_),
    .A1(net3359),
    .B1(net3324),
    .X(_07553_));
 sg13g2_xnor2_1 _30350_ (.Y(_07554_),
    .A(_06463_),
    .B(_07553_));
 sg13g2_a21oi_1 _30351_ (.A1(net4202),
    .A2(_07554_),
    .Y(_01246_),
    .B1(_07552_));
 sg13g2_nor2_1 _30352_ (.A(net1654),
    .B(net4208),
    .Y(_07555_));
 sg13g2_xnor2_1 _30353_ (.Y(_07556_),
    .A(net3385),
    .B(_06463_));
 sg13g2_nor2_1 _30354_ (.A(_07553_),
    .B(_07556_),
    .Y(_07557_));
 sg13g2_xor2_1 _30355_ (.B(_07557_),
    .A(_06460_),
    .X(_07558_));
 sg13g2_a21oi_1 _30356_ (.A1(net4208),
    .A2(_07558_),
    .Y(_01247_),
    .B1(_07555_));
 sg13g2_nor2_1 _30357_ (.A(net1374),
    .B(net4197),
    .Y(_07559_));
 sg13g2_and4_1 _30358_ (.A(_06440_),
    .B(_06460_),
    .C(_06463_),
    .D(_07538_),
    .X(_07560_));
 sg13g2_and4_1 _30359_ (.A(_06548_),
    .B(_06549_),
    .C(_07523_),
    .D(_07560_),
    .X(_07561_));
 sg13g2_a21oi_1 _30360_ (.A1(net3358),
    .A2(_07561_),
    .Y(_07562_),
    .B1(net3336));
 sg13g2_xnor2_1 _30361_ (.Y(_07563_),
    .A(_06429_),
    .B(_07562_));
 sg13g2_a21oi_1 _30362_ (.A1(net4197),
    .A2(_07563_),
    .Y(_01248_),
    .B1(_07559_));
 sg13g2_nand2_1 _30363_ (.Y(_07564_),
    .A(_05920_),
    .B(_06429_));
 sg13g2_nand3_1 _30364_ (.B(_06429_),
    .C(_07561_),
    .A(_05920_),
    .Y(_07565_));
 sg13g2_nor2_1 _30365_ (.A(net3381),
    .B(_07565_),
    .Y(_07566_));
 sg13g2_a21o_1 _30366_ (.A2(_07561_),
    .A1(_06429_),
    .B1(_05920_),
    .X(_07567_));
 sg13g2_a21o_1 _30367_ (.A2(_07567_),
    .A1(_07565_),
    .B1(net3381),
    .X(_07568_));
 sg13g2_o21ai_1 _30368_ (.B1(_07568_),
    .Y(_07569_),
    .A1(_05920_),
    .A2(net3311));
 sg13g2_mux2_1 _30369_ (.A0(net2001),
    .A1(_07569_),
    .S(net4200),
    .X(_01249_));
 sg13g2_nor3_1 _30370_ (.A(_06540_),
    .B(net3337),
    .C(_07566_),
    .Y(_07570_));
 sg13g2_nor3_1 _30371_ (.A(net3383),
    .B(_06541_),
    .C(_07565_),
    .Y(_07571_));
 sg13g2_nor2_1 _30372_ (.A(_07570_),
    .B(_07571_),
    .Y(_07572_));
 sg13g2_nand2_1 _30373_ (.Y(_07573_),
    .A(net1081),
    .B(net4156));
 sg13g2_o21ai_1 _30374_ (.B1(_07573_),
    .Y(_01250_),
    .A1(net4156),
    .A2(_07572_));
 sg13g2_or3_1 _30375_ (.A(_06525_),
    .B(net3337),
    .C(_07571_),
    .X(_07574_));
 sg13g2_nand2_1 _30376_ (.Y(_07575_),
    .A(_06525_),
    .B(_06540_));
 sg13g2_nor2_1 _30377_ (.A(_07565_),
    .B(_07575_),
    .Y(_07576_));
 sg13g2_a21oi_1 _30378_ (.A1(net3358),
    .A2(_07576_),
    .Y(_07577_),
    .B1(net4156));
 sg13g2_a22oi_1 _30379_ (.Y(_01251_),
    .B1(_07574_),
    .B2(_07577_),
    .A2(net4156),
    .A1(_11026_));
 sg13g2_nor2_1 _30380_ (.A(net1368),
    .B(net4196),
    .Y(_07578_));
 sg13g2_a21oi_1 _30381_ (.A1(net3358),
    .A2(_07576_),
    .Y(_07579_),
    .B1(net3337));
 sg13g2_xnor2_1 _30382_ (.Y(_07580_),
    .A(_05923_),
    .B(_07579_));
 sg13g2_a21oi_1 _30383_ (.A1(net4195),
    .A2(_07580_),
    .Y(_01252_),
    .B1(_07578_));
 sg13g2_and2_1 _30384_ (.A(_05923_),
    .B(_07576_),
    .X(_07581_));
 sg13g2_nand2_1 _30385_ (.Y(_07582_),
    .A(_06574_),
    .B(_07581_));
 sg13g2_xnor2_1 _30386_ (.Y(_07583_),
    .A(_06574_),
    .B(_07581_));
 sg13g2_o21ai_1 _30387_ (.B1(net4195),
    .Y(_07584_),
    .A1(_06574_),
    .A2(net3312));
 sg13g2_a21oi_1 _30388_ (.A1(net3357),
    .A2(_07583_),
    .Y(_07585_),
    .B1(_07584_));
 sg13g2_a21oi_1 _30389_ (.A1(_11027_),
    .A2(net4154),
    .Y(_01253_),
    .B1(_07585_));
 sg13g2_nor2_1 _30390_ (.A(net1586),
    .B(net4195),
    .Y(_07586_));
 sg13g2_a21oi_1 _30391_ (.A1(net3356),
    .A2(_07582_),
    .Y(_07587_),
    .B1(net3321));
 sg13g2_xnor2_1 _30392_ (.Y(_07588_),
    .A(_06566_),
    .B(_07587_));
 sg13g2_a21oi_1 _30393_ (.A1(net4195),
    .A2(_07588_),
    .Y(_01254_),
    .B1(_07586_));
 sg13g2_nor2_1 _30394_ (.A(net1507),
    .B(net4194),
    .Y(_07589_));
 sg13g2_xnor2_1 _30395_ (.Y(_07590_),
    .A(net3381),
    .B(_06566_));
 sg13g2_nand2_1 _30396_ (.Y(_07591_),
    .A(_07587_),
    .B(_07590_));
 sg13g2_xnor2_1 _30397_ (.Y(_07592_),
    .A(_06572_),
    .B(_07591_));
 sg13g2_a21oi_1 _30398_ (.A1(net4194),
    .A2(_07592_),
    .Y(_01255_),
    .B1(_07589_));
 sg13g2_nor2_1 _30399_ (.A(net1455),
    .B(net4193),
    .Y(_07593_));
 sg13g2_nand3_1 _30400_ (.B(_06572_),
    .C(_06574_),
    .A(_05923_),
    .Y(_07594_));
 sg13g2_nor4_2 _30401_ (.A(_06566_),
    .B(_07564_),
    .C(_07575_),
    .Y(_07595_),
    .D(_07594_));
 sg13g2_nand2_1 _30402_ (.Y(_07596_),
    .A(_07561_),
    .B(_07595_));
 sg13g2_a21oi_1 _30403_ (.A1(net3354),
    .A2(_07596_),
    .Y(_07597_),
    .B1(net3322));
 sg13g2_xnor2_1 _30404_ (.Y(_07598_),
    .A(_06434_),
    .B(_07597_));
 sg13g2_a21oi_1 _30405_ (.A1(net4193),
    .A2(_07598_),
    .Y(_01256_),
    .B1(_07593_));
 sg13g2_nor2_1 _30406_ (.A(net1689),
    .B(net4193),
    .Y(_07599_));
 sg13g2_nand3_1 _30407_ (.B(_07561_),
    .C(_07595_),
    .A(_06433_),
    .Y(_07600_));
 sg13g2_nand2b_2 _30408_ (.Y(_07601_),
    .B(_05917_),
    .A_N(_07600_));
 sg13g2_xnor2_1 _30409_ (.Y(_07602_),
    .A(_05916_),
    .B(_07600_));
 sg13g2_a22oi_1 _30410_ (.Y(_07603_),
    .B1(_07602_),
    .B2(net3356),
    .A2(net3321),
    .A1(_05916_));
 sg13g2_a21oi_1 _30411_ (.A1(net4194),
    .A2(_07603_),
    .Y(_01257_),
    .B1(_07599_));
 sg13g2_a21oi_1 _30412_ (.A1(net3356),
    .A2(_07601_),
    .Y(_07604_),
    .B1(net3321));
 sg13g2_xnor2_1 _30413_ (.Y(_07605_),
    .A(_06546_),
    .B(_07604_));
 sg13g2_nand2_1 _30414_ (.Y(_07606_),
    .A(net1092),
    .B(net4154));
 sg13g2_o21ai_1 _30415_ (.B1(_07606_),
    .Y(_01258_),
    .A1(net4154),
    .A2(_07605_));
 sg13g2_nor3_1 _30416_ (.A(_06512_),
    .B(_06546_),
    .C(_07601_),
    .Y(_07607_));
 sg13g2_o21ai_1 _30417_ (.B1(_06512_),
    .Y(_07608_),
    .A1(_06546_),
    .A2(_07601_));
 sg13g2_nand2b_1 _30418_ (.Y(_07609_),
    .B(_07608_),
    .A_N(_07607_));
 sg13g2_a221oi_1 _30419_ (.B2(net3356),
    .C1(net4154),
    .B1(_07609_),
    .A1(_06512_),
    .Y(_07610_),
    .A2(net3321));
 sg13g2_a21oi_1 _30420_ (.A1(_11028_),
    .A2(net4154),
    .Y(_01259_),
    .B1(_07610_));
 sg13g2_nor2_1 _30421_ (.A(net1335),
    .B(net4194),
    .Y(_07611_));
 sg13g2_o21ai_1 _30422_ (.B1(net3311),
    .Y(_07612_),
    .A1(net3381),
    .A2(_07607_));
 sg13g2_xor2_1 _30423_ (.B(_07612_),
    .A(_06532_),
    .X(_07613_));
 sg13g2_a21oi_1 _30424_ (.A1(net4193),
    .A2(_07613_),
    .Y(_01260_),
    .B1(_07611_));
 sg13g2_or4_1 _30425_ (.A(_06512_),
    .B(_06532_),
    .C(_06534_),
    .D(_06546_),
    .X(_07614_));
 sg13g2_nor2_1 _30426_ (.A(_07601_),
    .B(_07614_),
    .Y(_07615_));
 sg13g2_or2_1 _30427_ (.X(_07616_),
    .B(_07615_),
    .A(_06535_));
 sg13g2_a221oi_1 _30428_ (.B2(net3354),
    .C1(net4154),
    .B1(_07616_),
    .A1(_06534_),
    .Y(_07617_),
    .A2(_07612_));
 sg13g2_a21oi_1 _30429_ (.A1(_11029_),
    .A2(net4154),
    .Y(_01261_),
    .B1(_07617_));
 sg13g2_nor2_1 _30430_ (.A(net1577),
    .B(net4193),
    .Y(_07618_));
 sg13g2_a21oi_1 _30431_ (.A1(net3355),
    .A2(_07615_),
    .Y(_07619_),
    .B1(net3336));
 sg13g2_xor2_1 _30432_ (.B(_07619_),
    .A(_06537_),
    .X(_07620_));
 sg13g2_a21oi_1 _30433_ (.A1(net4193),
    .A2(_07620_),
    .Y(_01262_),
    .B1(_07618_));
 sg13g2_nor2_1 _30434_ (.A(net1575),
    .B(net4193),
    .Y(_07621_));
 sg13g2_a21oi_1 _30435_ (.A1(net3355),
    .A2(_06537_),
    .Y(_07622_),
    .B1(_07619_));
 sg13g2_xor2_1 _30436_ (.B(_07622_),
    .A(_06583_),
    .X(_07623_));
 sg13g2_a21oi_1 _30437_ (.A1(net4193),
    .A2(_07623_),
    .Y(_01263_),
    .B1(_07621_));
 sg13g2_nor2_1 _30438_ (.A(net1739),
    .B(net4190),
    .Y(_07624_));
 sg13g2_nor4_1 _30439_ (.A(_05916_),
    .B(_06434_),
    .C(_06537_),
    .D(_07614_),
    .Y(_07625_));
 sg13g2_nand2_1 _30440_ (.Y(_07626_),
    .A(_06583_),
    .B(_07625_));
 sg13g2_nor2_1 _30441_ (.A(_07596_),
    .B(_07626_),
    .Y(_07627_));
 sg13g2_a21oi_1 _30442_ (.A1(net3354),
    .A2(_07627_),
    .Y(_07628_),
    .B1(net3336));
 sg13g2_xnor2_1 _30443_ (.Y(_07629_),
    .A(_05943_),
    .B(_07628_));
 sg13g2_a21oi_1 _30444_ (.A1(net4190),
    .A2(_07629_),
    .Y(_01264_),
    .B1(_07624_));
 sg13g2_nor2_1 _30445_ (.A(net1392),
    .B(net4190),
    .Y(_07630_));
 sg13g2_nand2_1 _30446_ (.Y(_07631_),
    .A(_05943_),
    .B(_07627_));
 sg13g2_xnor2_1 _30447_ (.Y(_07632_),
    .A(_06564_),
    .B(_07631_));
 sg13g2_a22oi_1 _30448_ (.Y(_07633_),
    .B1(_07632_),
    .B2(net3354),
    .A2(net3320),
    .A1(_06564_));
 sg13g2_a21oi_1 _30449_ (.A1(net4190),
    .A2(_07633_),
    .Y(_01265_),
    .B1(_07630_));
 sg13g2_nor2_1 _30450_ (.A(net1322),
    .B(net4191),
    .Y(_07634_));
 sg13g2_o21ai_1 _30451_ (.B1(net3354),
    .Y(_07635_),
    .A1(_06564_),
    .A2(_07631_));
 sg13g2_nand2_1 _30452_ (.Y(_07636_),
    .A(net3312),
    .B(_07635_));
 sg13g2_xnor2_1 _30453_ (.Y(_07637_),
    .A(_06521_),
    .B(_07636_));
 sg13g2_a21oi_1 _30454_ (.A1(net4190),
    .A2(_07637_),
    .Y(_01266_),
    .B1(_07634_));
 sg13g2_nor2_1 _30455_ (.A(net1816),
    .B(net4190),
    .Y(_07638_));
 sg13g2_nor2_1 _30456_ (.A(_05944_),
    .B(_06564_),
    .Y(_07639_));
 sg13g2_nand4_1 _30457_ (.B(_06521_),
    .C(_07595_),
    .A(_06518_),
    .Y(_07640_),
    .D(_07639_));
 sg13g2_nor2_1 _30458_ (.A(_07626_),
    .B(_07640_),
    .Y(_07641_));
 sg13g2_and2_1 _30459_ (.A(_07561_),
    .B(_07641_),
    .X(_07642_));
 sg13g2_inv_1 _30460_ (.Y(_07643_),
    .A(_07642_));
 sg13g2_nand2_1 _30461_ (.Y(_07644_),
    .A(_06522_),
    .B(_07643_));
 sg13g2_a22oi_1 _30462_ (.Y(_07645_),
    .B1(_07644_),
    .B2(net3354),
    .A2(_07636_),
    .A1(_06519_));
 sg13g2_a21oi_1 _30463_ (.A1(net4191),
    .A2(_07645_),
    .Y(_01267_),
    .B1(_07638_));
 sg13g2_nor2_1 _30464_ (.A(net1598),
    .B(net4190),
    .Y(_07646_));
 sg13g2_a21oi_1 _30465_ (.A1(net3354),
    .A2(_07642_),
    .Y(_07647_),
    .B1(net3336));
 sg13g2_xor2_1 _30466_ (.B(_07647_),
    .A(_06552_),
    .X(_07648_));
 sg13g2_a21oi_1 _30467_ (.A1(net4190),
    .A2(_07648_),
    .Y(_01268_),
    .B1(_07646_));
 sg13g2_nor2_1 _30468_ (.A(_06552_),
    .B(_07643_),
    .Y(_07649_));
 sg13g2_xnor2_1 _30469_ (.Y(_07650_),
    .A(_06531_),
    .B(_07649_));
 sg13g2_a221oi_1 _30470_ (.B2(net3355),
    .C1(net4157),
    .B1(_07650_),
    .A1(_06530_),
    .Y(_07651_),
    .A2(net3320));
 sg13g2_a21oi_1 _30471_ (.A1(_11030_),
    .A2(net4153),
    .Y(_01269_),
    .B1(_07651_));
 sg13g2_a21oi_1 _30472_ (.A1(_06531_),
    .A2(_07649_),
    .Y(_07652_),
    .B1(net3381));
 sg13g2_nor2_1 _30473_ (.A(net3321),
    .B(_07652_),
    .Y(_07653_));
 sg13g2_xor2_1 _30474_ (.B(_07653_),
    .A(_06570_),
    .X(_07654_));
 sg13g2_nand2_1 _30475_ (.Y(_07655_),
    .A(net1083),
    .B(net4153));
 sg13g2_o21ai_1 _30476_ (.B1(_07655_),
    .Y(_01270_),
    .A1(net4157),
    .A2(_07654_));
 sg13g2_nor2_1 _30477_ (.A(net1935),
    .B(net4191),
    .Y(_07656_));
 sg13g2_xnor2_1 _30478_ (.Y(_07657_),
    .A(net3354),
    .B(_06570_));
 sg13g2_nand2_1 _30479_ (.Y(_07658_),
    .A(_07653_),
    .B(_07657_));
 sg13g2_xor2_1 _30480_ (.B(_07658_),
    .A(_06506_),
    .X(_07659_));
 sg13g2_a21oi_1 _30481_ (.A1(net4191),
    .A2(_07659_),
    .Y(_01271_),
    .B1(_07656_));
 sg13g2_nand2b_1 _30482_ (.Y(_07660_),
    .B(_06570_),
    .A_N(_06552_));
 sg13g2_nor3_2 _30483_ (.A(_06506_),
    .B(_06530_),
    .C(_07660_),
    .Y(_07661_));
 sg13g2_nand2_2 _30484_ (.Y(_07662_),
    .A(_07642_),
    .B(_07661_));
 sg13g2_a21oi_1 _30485_ (.A1(net3352),
    .A2(_07662_),
    .Y(_07663_),
    .B1(net3319));
 sg13g2_xnor2_1 _30486_ (.Y(_07664_),
    .A(_05952_),
    .B(_07663_));
 sg13g2_nand2_1 _30487_ (.Y(_07665_),
    .A(net1073),
    .B(net4151));
 sg13g2_o21ai_1 _30488_ (.B1(_07665_),
    .Y(_01272_),
    .A1(net4151),
    .A2(_07664_));
 sg13g2_nor2_2 _30489_ (.A(_05952_),
    .B(_06569_),
    .Y(_07666_));
 sg13g2_nand3_1 _30490_ (.B(_07661_),
    .C(_07666_),
    .A(_07642_),
    .Y(_07667_));
 sg13g2_o21ai_1 _30491_ (.B1(_06569_),
    .Y(_07668_),
    .A1(_05952_),
    .A2(_07662_));
 sg13g2_a21o_1 _30492_ (.A2(_07668_),
    .A1(_07667_),
    .B1(net3382),
    .X(_07669_));
 sg13g2_a21oi_1 _30493_ (.A1(_06569_),
    .A2(net3319),
    .Y(_07670_),
    .B1(net4151));
 sg13g2_a22oi_1 _30494_ (.Y(_01273_),
    .B1(_07669_),
    .B2(_07670_),
    .A2(net4151),
    .A1(_11031_));
 sg13g2_nor2_1 _30495_ (.A(net1532),
    .B(net4187),
    .Y(_07671_));
 sg13g2_a21oi_1 _30496_ (.A1(net3350),
    .A2(_07667_),
    .Y(_07672_),
    .B1(net3319));
 sg13g2_xnor2_1 _30497_ (.Y(_07673_),
    .A(_06528_),
    .B(_07672_));
 sg13g2_a21oi_1 _30498_ (.A1(net4187),
    .A2(_07673_),
    .Y(_01274_),
    .B1(_07671_));
 sg13g2_nor2_1 _30499_ (.A(_06528_),
    .B(_07667_),
    .Y(_07674_));
 sg13g2_nand2b_1 _30500_ (.Y(_07675_),
    .B(_06590_),
    .A_N(_06528_));
 sg13g2_xnor2_1 _30501_ (.Y(_07676_),
    .A(_06590_),
    .B(_07674_));
 sg13g2_o21ai_1 _30502_ (.B1(net4187),
    .Y(_07677_),
    .A1(_06590_),
    .A2(net3312));
 sg13g2_a21oi_1 _30503_ (.A1(net3350),
    .A2(_07676_),
    .Y(_07678_),
    .B1(_07677_));
 sg13g2_a21oi_1 _30504_ (.A1(_11032_),
    .A2(net4149),
    .Y(_01275_),
    .B1(_07678_));
 sg13g2_nor2_1 _30505_ (.A(net1643),
    .B(net4187),
    .Y(_07679_));
 sg13g2_o21ai_1 _30506_ (.B1(net3350),
    .Y(_07680_),
    .A1(_07667_),
    .A2(_07675_));
 sg13g2_nand2_1 _30507_ (.Y(_07681_),
    .A(net3310),
    .B(_07680_));
 sg13g2_xnor2_1 _30508_ (.Y(_07682_),
    .A(_06617_),
    .B(_07681_));
 sg13g2_a21oi_1 _30509_ (.A1(net4187),
    .A2(_07682_),
    .Y(_01276_),
    .B1(_07679_));
 sg13g2_nand2_1 _30510_ (.Y(_07683_),
    .A(_06616_),
    .B(_06617_));
 sg13g2_nor3_1 _30511_ (.A(_07667_),
    .B(_07675_),
    .C(_07683_),
    .Y(_07684_));
 sg13g2_or2_1 _30512_ (.X(_07685_),
    .B(_07684_),
    .A(_06618_));
 sg13g2_a221oi_1 _30513_ (.B2(net3351),
    .C1(net4149),
    .B1(_07685_),
    .A1(_06615_),
    .Y(_07686_),
    .A2(_07681_));
 sg13g2_a21oi_1 _30514_ (.A1(_11033_),
    .A2(net4150),
    .Y(_01277_),
    .B1(_07686_));
 sg13g2_a21o_1 _30515_ (.A2(_07684_),
    .A1(net3351),
    .B1(net3335),
    .X(_07687_));
 sg13g2_xor2_1 _30516_ (.B(_07687_),
    .A(_06592_),
    .X(_07688_));
 sg13g2_nand2_1 _30517_ (.Y(_07689_),
    .A(net1071),
    .B(net4149));
 sg13g2_o21ai_1 _30518_ (.B1(_07689_),
    .Y(_01278_),
    .A1(net4150),
    .A2(_07688_));
 sg13g2_nor2_1 _30519_ (.A(net1454),
    .B(net4184),
    .Y(_07690_));
 sg13g2_o21ai_1 _30520_ (.B1(_07687_),
    .Y(_07691_),
    .A1(net3380),
    .A2(_06592_));
 sg13g2_xor2_1 _30521_ (.B(_07691_),
    .A(_05901_),
    .X(_07692_));
 sg13g2_a21oi_1 _30522_ (.A1(net4184),
    .A2(_07692_),
    .Y(_01279_),
    .B1(_07690_));
 sg13g2_nor2_1 _30523_ (.A(net2007),
    .B(net4183),
    .Y(_07693_));
 sg13g2_nand2_1 _30524_ (.Y(_07694_),
    .A(_06592_),
    .B(_07666_));
 sg13g2_or4_1 _30525_ (.A(_05901_),
    .B(_07675_),
    .C(_07683_),
    .D(_07694_),
    .X(_07695_));
 sg13g2_nor2_1 _30526_ (.A(_07662_),
    .B(_07695_),
    .Y(_07696_));
 sg13g2_a21oi_1 _30527_ (.A1(net3348),
    .A2(_07696_),
    .Y(_07697_),
    .B1(net3334));
 sg13g2_xnor2_1 _30528_ (.Y(_07698_),
    .A(_05911_),
    .B(_07697_));
 sg13g2_a21oi_1 _30529_ (.A1(net4181),
    .A2(_07698_),
    .Y(_01280_),
    .B1(_07693_));
 sg13g2_and2_1 _30530_ (.A(_05909_),
    .B(_05911_),
    .X(_07699_));
 sg13g2_and2_1 _30531_ (.A(_07696_),
    .B(_07699_),
    .X(_07700_));
 sg13g2_o21ai_1 _30532_ (.B1(_05912_),
    .Y(_07701_),
    .A1(_05909_),
    .A2(_07696_));
 sg13g2_o21ai_1 _30533_ (.B1(net3348),
    .Y(_07702_),
    .A1(_07700_),
    .A2(_07701_));
 sg13g2_a21oi_1 _30534_ (.A1(_05910_),
    .A2(net3319),
    .Y(_07703_),
    .B1(net4148));
 sg13g2_a22oi_1 _30535_ (.Y(_01281_),
    .B1(_07702_),
    .B2(_07703_),
    .A2(net4148),
    .A1(_11034_));
 sg13g2_a21oi_1 _30536_ (.A1(net3348),
    .A2(_07700_),
    .Y(_07704_),
    .B1(net3334));
 sg13g2_xnor2_1 _30537_ (.Y(_07705_),
    .A(_06595_),
    .B(_07704_));
 sg13g2_nand2_1 _30538_ (.Y(_07706_),
    .A(net1676),
    .B(net4148));
 sg13g2_o21ai_1 _30539_ (.B1(_07706_),
    .Y(_01282_),
    .A1(net4148),
    .A2(_07705_));
 sg13g2_nand2_1 _30540_ (.Y(_07707_),
    .A(_06595_),
    .B(_06607_));
 sg13g2_inv_1 _30541_ (.Y(_07708_),
    .A(_07707_));
 sg13g2_and2_1 _30542_ (.A(_07700_),
    .B(_07708_),
    .X(_07709_));
 sg13g2_a21oi_1 _30543_ (.A1(_06595_),
    .A2(_07700_),
    .Y(_07710_),
    .B1(_06607_));
 sg13g2_o21ai_1 _30544_ (.B1(net3348),
    .Y(_07711_),
    .A1(_07709_),
    .A2(_07710_));
 sg13g2_a21oi_1 _30545_ (.A1(_06608_),
    .A2(net3318),
    .Y(_07712_),
    .B1(net4148));
 sg13g2_a22oi_1 _30546_ (.Y(_01283_),
    .B1(_07711_),
    .B2(_07712_),
    .A2(net4148),
    .A1(_11035_));
 sg13g2_nor2_1 _30547_ (.A(net2036),
    .B(net4181),
    .Y(_07713_));
 sg13g2_o21ai_1 _30548_ (.B1(net3312),
    .Y(_07714_),
    .A1(net3379),
    .A2(_07709_));
 sg13g2_xnor2_1 _30549_ (.Y(_07715_),
    .A(_06591_),
    .B(_07714_));
 sg13g2_a21oi_1 _30550_ (.A1(net4181),
    .A2(_07715_),
    .Y(_01284_),
    .B1(_07713_));
 sg13g2_and2_1 _30551_ (.A(_06591_),
    .B(_06604_),
    .X(_07716_));
 sg13g2_nand2_1 _30552_ (.Y(_07717_),
    .A(_07708_),
    .B(_07716_));
 sg13g2_a21oi_1 _30553_ (.A1(_06591_),
    .A2(_07709_),
    .Y(_07718_),
    .B1(_06604_));
 sg13g2_a21o_1 _30554_ (.A2(_07716_),
    .A1(_07709_),
    .B1(_07718_),
    .X(_07719_));
 sg13g2_o21ai_1 _30555_ (.B1(net4181),
    .Y(_07720_),
    .A1(_06604_),
    .A2(net3312));
 sg13g2_a21oi_1 _30556_ (.A1(net3348),
    .A2(_07719_),
    .Y(_07721_),
    .B1(_07720_));
 sg13g2_a21oi_1 _30557_ (.A1(_11036_),
    .A2(net4148),
    .Y(_01285_),
    .B1(_07721_));
 sg13g2_nor2_1 _30558_ (.A(net2069),
    .B(net4181),
    .Y(_07722_));
 sg13g2_a21oi_1 _30559_ (.A1(_07709_),
    .A2(_07716_),
    .Y(_07723_),
    .B1(net3379));
 sg13g2_nor2_1 _30560_ (.A(net3318),
    .B(_07723_),
    .Y(_07724_));
 sg13g2_xor2_1 _30561_ (.B(_07724_),
    .A(_06605_),
    .X(_07725_));
 sg13g2_a21oi_1 _30562_ (.A1(net4181),
    .A2(_07725_),
    .Y(_01286_),
    .B1(_07722_));
 sg13g2_nor2_1 _30563_ (.A(net2055),
    .B(net4181),
    .Y(_07726_));
 sg13g2_xnor2_1 _30564_ (.Y(_07727_),
    .A(net3348),
    .B(_06605_));
 sg13g2_nand2_1 _30565_ (.Y(_07728_),
    .A(_07724_),
    .B(_07727_));
 sg13g2_xnor2_1 _30566_ (.Y(_07729_),
    .A(_06503_),
    .B(_07728_));
 sg13g2_a21oi_1 _30567_ (.A1(net4181),
    .A2(_07729_),
    .Y(_01287_),
    .B1(_07726_));
 sg13g2_nor2_1 _30568_ (.A(net2032),
    .B(net4179),
    .Y(_07730_));
 sg13g2_nand3_1 _30569_ (.B(_06605_),
    .C(_07699_),
    .A(_06503_),
    .Y(_07731_));
 sg13g2_nor4_2 _30570_ (.A(_07662_),
    .B(_07695_),
    .C(_07717_),
    .Y(_07732_),
    .D(_07731_));
 sg13g2_a21oi_1 _30571_ (.A1(net3347),
    .A2(_07732_),
    .Y(_07733_),
    .B1(net3335));
 sg13g2_xor2_1 _30572_ (.B(_07733_),
    .A(_06620_),
    .X(_07734_));
 sg13g2_a21oi_1 _30573_ (.A1(net4179),
    .A2(_07734_),
    .Y(_01288_),
    .B1(_07730_));
 sg13g2_nor2_1 _30574_ (.A(_06620_),
    .B(_06622_),
    .Y(_07735_));
 sg13g2_nand2_2 _30575_ (.Y(_07736_),
    .A(_07732_),
    .B(_07735_));
 sg13g2_nand2b_1 _30576_ (.Y(_07737_),
    .B(_06622_),
    .A_N(_07732_));
 sg13g2_nand3_1 _30577_ (.B(_07736_),
    .C(_07737_),
    .A(_06623_),
    .Y(_07738_));
 sg13g2_a221oi_1 _30578_ (.B2(net3347),
    .C1(net4150),
    .B1(_07738_),
    .A1(_06622_),
    .Y(_07739_),
    .A2(net3318));
 sg13g2_a21oi_1 _30579_ (.A1(_11037_),
    .A2(net4147),
    .Y(_01289_),
    .B1(_07739_));
 sg13g2_a21oi_1 _30580_ (.A1(net3347),
    .A2(_07736_),
    .Y(_07740_),
    .B1(net3319));
 sg13g2_xor2_1 _30581_ (.B(_07740_),
    .A(_06587_),
    .X(_07741_));
 sg13g2_nand2_1 _30582_ (.Y(_07742_),
    .A(net1583),
    .B(net4147));
 sg13g2_o21ai_1 _30583_ (.B1(_07742_),
    .Y(_01290_),
    .A1(net4147),
    .A2(_07741_));
 sg13g2_nand3_1 _30584_ (.B(_07732_),
    .C(_07735_),
    .A(_06587_),
    .Y(_07743_));
 sg13g2_nand2_1 _30585_ (.Y(_07744_),
    .A(_06587_),
    .B(_06612_));
 sg13g2_xor2_1 _30586_ (.B(_07743_),
    .A(_06612_),
    .X(_07745_));
 sg13g2_o21ai_1 _30587_ (.B1(net4179),
    .Y(_07746_),
    .A1(_06612_),
    .A2(net3310));
 sg13g2_a21oi_1 _30588_ (.A1(net3347),
    .A2(_07745_),
    .Y(_07747_),
    .B1(_07746_));
 sg13g2_a21oi_1 _30589_ (.A1(_11038_),
    .A2(net4147),
    .Y(_01291_),
    .B1(_07747_));
 sg13g2_o21ai_1 _30590_ (.B1(net3347),
    .Y(_07748_),
    .A1(_07736_),
    .A2(_07744_));
 sg13g2_nand2_1 _30591_ (.Y(_07749_),
    .A(net3310),
    .B(_07748_));
 sg13g2_xnor2_1 _30592_ (.Y(_07750_),
    .A(_06601_),
    .B(_07749_));
 sg13g2_nand2_1 _30593_ (.Y(_07751_),
    .A(net1375),
    .B(net4147));
 sg13g2_o21ai_1 _30594_ (.B1(_07751_),
    .Y(_01292_),
    .A1(net4150),
    .A2(_07750_));
 sg13g2_nor2_1 _30595_ (.A(net2345),
    .B(net4179),
    .Y(_07752_));
 sg13g2_nand2b_1 _30596_ (.Y(_07753_),
    .B(_06601_),
    .A_N(_06600_));
 sg13g2_or3_1 _30597_ (.A(_07736_),
    .B(_07744_),
    .C(_07753_),
    .X(_07754_));
 sg13g2_nand2_1 _30598_ (.Y(_07755_),
    .A(_06602_),
    .B(_07754_));
 sg13g2_a22oi_1 _30599_ (.Y(_07756_),
    .B1(_07755_),
    .B2(net3347),
    .A2(_07749_),
    .A1(_06600_));
 sg13g2_a21oi_1 _30600_ (.A1(net4179),
    .A2(_07756_),
    .Y(_01293_),
    .B1(_07752_));
 sg13g2_a21oi_1 _30601_ (.A1(net3347),
    .A2(_07754_),
    .Y(_07757_),
    .B1(net3318));
 sg13g2_xnor2_1 _30602_ (.Y(_07758_),
    .A(_06584_),
    .B(_07757_));
 sg13g2_nor2_1 _30603_ (.A(net2106),
    .B(net4179),
    .Y(_07759_));
 sg13g2_a21oi_1 _30604_ (.A1(net4179),
    .A2(_07758_),
    .Y(_01294_),
    .B1(_07759_));
 sg13g2_nor2_1 _30605_ (.A(net2137),
    .B(net4178),
    .Y(_07760_));
 sg13g2_xnor2_1 _30606_ (.Y(_07761_),
    .A(net3347),
    .B(_06585_));
 sg13g2_nand2_1 _30607_ (.Y(_07762_),
    .A(_07757_),
    .B(_07761_));
 sg13g2_xor2_1 _30608_ (.B(_07762_),
    .A(_05906_),
    .X(_07763_));
 sg13g2_a21oi_1 _30609_ (.A1(net4179),
    .A2(_07763_),
    .Y(_01295_),
    .B1(_07760_));
 sg13g2_nand2_1 _30610_ (.Y(_07764_),
    .A(_06585_),
    .B(_07735_));
 sg13g2_nor4_1 _30611_ (.A(_05906_),
    .B(_07744_),
    .C(_07753_),
    .D(_07764_),
    .Y(_07765_));
 sg13g2_and2_1 _30612_ (.A(_07732_),
    .B(_07765_),
    .X(_07766_));
 sg13g2_o21ai_1 _30613_ (.B1(net3310),
    .Y(_07767_),
    .A1(net3378),
    .A2(_07766_));
 sg13g2_xnor2_1 _30614_ (.Y(_07768_),
    .A(_06633_),
    .B(_07767_));
 sg13g2_nand2_1 _30615_ (.Y(_07769_),
    .A(net1609),
    .B(net4144));
 sg13g2_o21ai_1 _30616_ (.B1(_07769_),
    .Y(_01296_),
    .A1(net4144),
    .A2(_07768_));
 sg13g2_nand2b_1 _30617_ (.Y(_07770_),
    .B(_07767_),
    .A_N(_06632_));
 sg13g2_and3_2 _30618_ (.X(_07771_),
    .A(_06632_),
    .B(_06633_),
    .C(_07766_));
 sg13g2_o21ai_1 _30619_ (.B1(net3346),
    .Y(_07772_),
    .A1(_06634_),
    .A2(_07771_));
 sg13g2_nand3_1 _30620_ (.B(_07770_),
    .C(_07772_),
    .A(net4178),
    .Y(_07773_));
 sg13g2_o21ai_1 _30621_ (.B1(_07773_),
    .Y(_07774_),
    .A1(net3170),
    .A2(net4178));
 sg13g2_inv_1 _30622_ (.Y(_01297_),
    .A(_07774_));
 sg13g2_o21ai_1 _30623_ (.B1(net3310),
    .Y(_07775_),
    .A1(net3378),
    .A2(_07771_));
 sg13g2_xor2_1 _30624_ (.B(_07775_),
    .A(_06630_),
    .X(_07776_));
 sg13g2_nand2_1 _30625_ (.Y(_07777_),
    .A(net1936),
    .B(net4144));
 sg13g2_o21ai_1 _30626_ (.B1(_07777_),
    .Y(_01298_),
    .A1(net4144),
    .A2(_07776_));
 sg13g2_nand2b_1 _30627_ (.Y(_07778_),
    .B(_07771_),
    .A_N(_06630_));
 sg13g2_nor2_1 _30628_ (.A(_05894_),
    .B(_06630_),
    .Y(_07779_));
 sg13g2_and2_1 _30629_ (.A(_07771_),
    .B(_07779_),
    .X(_07780_));
 sg13g2_a21o_1 _30630_ (.A2(_07778_),
    .A1(_05894_),
    .B1(_07780_),
    .X(_07781_));
 sg13g2_a221oi_1 _30631_ (.B2(net3346),
    .C1(net4144),
    .B1(_07781_),
    .A1(_05894_),
    .Y(_07782_),
    .A2(net3318));
 sg13g2_a21oi_1 _30632_ (.A1(_11039_),
    .A2(net4144),
    .Y(_01299_),
    .B1(_07782_));
 sg13g2_nor2_1 _30633_ (.A(net2249),
    .B(net4178),
    .Y(_07783_));
 sg13g2_o21ai_1 _30634_ (.B1(net3310),
    .Y(_07784_),
    .A1(net3378),
    .A2(_07780_));
 sg13g2_xnor2_1 _30635_ (.Y(_07785_),
    .A(_06624_),
    .B(_07784_));
 sg13g2_a21oi_1 _30636_ (.A1(net4178),
    .A2(_07785_),
    .Y(_01300_),
    .B1(_07783_));
 sg13g2_and2_1 _30637_ (.A(_06624_),
    .B(_07780_),
    .X(_07786_));
 sg13g2_nand4_1 _30638_ (.B(_06624_),
    .C(_06637_),
    .A(net3346),
    .Y(_07787_),
    .D(_07780_));
 sg13g2_nand3_1 _30639_ (.B(_06637_),
    .C(_07780_),
    .A(_06624_),
    .Y(_07788_));
 sg13g2_o21ai_1 _30640_ (.B1(_07788_),
    .Y(_07789_),
    .A1(_06637_),
    .A2(_07786_));
 sg13g2_a221oi_1 _30641_ (.B2(net3346),
    .C1(net4147),
    .B1(_07789_),
    .A1(_06638_),
    .Y(_07790_),
    .A2(net3318));
 sg13g2_a21oi_1 _30642_ (.A1(_11040_),
    .A2(net4144),
    .Y(_01301_),
    .B1(_07790_));
 sg13g2_nor2_1 _30643_ (.A(net2284),
    .B(net4178),
    .Y(_07791_));
 sg13g2_a21oi_1 _30644_ (.A1(net3346),
    .A2(_07788_),
    .Y(_07792_),
    .B1(net3318));
 sg13g2_xnor2_1 _30645_ (.Y(_07793_),
    .A(_06635_),
    .B(_07792_));
 sg13g2_a21oi_1 _30646_ (.A1(net4178),
    .A2(_07793_),
    .Y(_01302_),
    .B1(_07791_));
 sg13g2_nand2_1 _30647_ (.Y(_07794_),
    .A(net2116),
    .B(net4144));
 sg13g2_nor2_1 _30648_ (.A(_06635_),
    .B(_07787_),
    .Y(_07795_));
 sg13g2_nor3_1 _30649_ (.A(_06628_),
    .B(_06635_),
    .C(_07787_),
    .Y(_07796_));
 sg13g2_nor2_1 _30650_ (.A(_06628_),
    .B(net3335),
    .Y(_07797_));
 sg13g2_o21ai_1 _30651_ (.B1(net4178),
    .Y(_07798_),
    .A1(_07795_),
    .A2(_07797_));
 sg13g2_o21ai_1 _30652_ (.B1(_07794_),
    .Y(_01303_),
    .A1(_07796_),
    .A2(_07798_));
 sg13g2_nand2_1 _30653_ (.Y(_07799_),
    .A(net1297),
    .B(net3742));
 sg13g2_xnor2_1 _30654_ (.Y(_07800_),
    .A(_12676_),
    .B(_12677_));
 sg13g2_nand2_1 _30655_ (.Y(_07801_),
    .A(net4639),
    .B(_07800_));
 sg13g2_o21ai_1 _30656_ (.B1(_07801_),
    .Y(_07802_),
    .A1(\u_inv.f_next[1] ),
    .A2(net4639));
 sg13g2_xnor2_1 _30657_ (.Y(_07803_),
    .A(_07799_),
    .B(_07802_));
 sg13g2_a21oi_1 _30658_ (.A1(net4379),
    .A2(_07803_),
    .Y(_07804_),
    .B1(net3915));
 sg13g2_o21ai_1 _30659_ (.B1(_07804_),
    .Y(_07805_),
    .A1(net4601),
    .A2(net3233));
 sg13g2_o21ai_1 _30660_ (.B1(_07805_),
    .Y(_01304_),
    .A1(net4528),
    .A2(net4000));
 sg13g2_xnor2_1 _30661_ (.Y(_07806_),
    .A(_11132_),
    .B(_12678_));
 sg13g2_nor2_1 _30662_ (.A(net2399),
    .B(net4639),
    .Y(_07807_));
 sg13g2_a21oi_1 _30663_ (.A1(net4639),
    .A2(_07806_),
    .Y(_07808_),
    .B1(_07807_));
 sg13g2_nand2b_1 _30664_ (.Y(_07809_),
    .B(_11132_),
    .A_N(_11136_));
 sg13g2_nand3b_1 _30665_ (.B(net3689),
    .C(_07809_),
    .Y(_07810_),
    .A_N(_11137_));
 sg13g2_a221oi_1 _30666_ (.B2(_07808_),
    .C1(net3917),
    .B1(net3711),
    .A1(net1529),
    .Y(_07811_),
    .A2(net4436));
 sg13g2_a22oi_1 _30667_ (.Y(_01305_),
    .B1(_07810_),
    .B2(_07811_),
    .A2(net3917),
    .A1(_10576_));
 sg13g2_xnor2_1 _30668_ (.Y(_07812_),
    .A(_11127_),
    .B(_12679_));
 sg13g2_nor2_1 _30669_ (.A(net4527),
    .B(_07812_),
    .Y(_07813_));
 sg13g2_a21oi_1 _30670_ (.A1(net2186),
    .A2(net4527),
    .Y(_07814_),
    .B1(_07813_));
 sg13g2_or3_1 _30671_ (.A(_11127_),
    .B(_11128_),
    .C(_11137_),
    .X(_07815_));
 sg13g2_and2_1 _30672_ (.A(_11138_),
    .B(_07815_),
    .X(_07816_));
 sg13g2_a21oi_1 _30673_ (.A1(_10957_),
    .A2(net4436),
    .Y(_07817_),
    .B1(net3918));
 sg13g2_o21ai_1 _30674_ (.B1(_07817_),
    .Y(_07818_),
    .A1(net3679),
    .A2(_07816_));
 sg13g2_a21oi_1 _30675_ (.A1(net3711),
    .A2(_07814_),
    .Y(_07819_),
    .B1(_07818_));
 sg13g2_a21o_1 _30676_ (.A2(net3918),
    .A1(net2399),
    .B1(_07819_),
    .X(_01306_));
 sg13g2_xor2_1 _30677_ (.B(_12680_),
    .A(_11124_),
    .X(_07820_));
 sg13g2_nand2_1 _30678_ (.Y(_07821_),
    .A(net4640),
    .B(_07820_));
 sg13g2_a21oi_1 _30679_ (.A1(net2933),
    .A2(net4527),
    .Y(_07822_),
    .B1(net3701));
 sg13g2_nand3_1 _30680_ (.B(_11125_),
    .C(_11138_),
    .A(_11124_),
    .Y(_07823_));
 sg13g2_nand2b_1 _30681_ (.Y(_07824_),
    .B(_07823_),
    .A_N(_11139_));
 sg13g2_o21ai_1 _30682_ (.B1(net4002),
    .Y(_07825_),
    .A1(net4602),
    .A2(net1267));
 sg13g2_a221oi_1 _30683_ (.B2(net3689),
    .C1(_07825_),
    .B1(_07824_),
    .A1(_07821_),
    .Y(_07826_),
    .A2(_07822_));
 sg13g2_a21o_1 _30684_ (.A2(net3918),
    .A1(net2186),
    .B1(_07826_),
    .X(_01307_));
 sg13g2_o21ai_1 _30685_ (.B1(net4640),
    .Y(_07827_),
    .A1(_11122_),
    .A2(_12681_));
 sg13g2_a21oi_1 _30686_ (.A1(_11122_),
    .A2(_12681_),
    .Y(_07828_),
    .B1(_07827_));
 sg13g2_a21oi_1 _30687_ (.A1(net2122),
    .A2(net4527),
    .Y(_07829_),
    .B1(_07828_));
 sg13g2_or3_1 _30688_ (.A(_11122_),
    .B(_11123_),
    .C(_11139_),
    .X(_07830_));
 sg13g2_nand2_1 _30689_ (.Y(_07831_),
    .A(_11140_),
    .B(_07830_));
 sg13g2_nor2_1 _30690_ (.A(net4602),
    .B(net1214),
    .Y(_07832_));
 sg13g2_a221oi_1 _30691_ (.B2(net3689),
    .C1(_07832_),
    .B1(_07831_),
    .A1(net3711),
    .Y(_07833_),
    .A2(_07829_));
 sg13g2_mux2_1 _30692_ (.A0(net2933),
    .A1(_07833_),
    .S(net4002),
    .X(_01308_));
 sg13g2_xor2_1 _30693_ (.B(_12682_),
    .A(_11119_),
    .X(_07834_));
 sg13g2_nor2_1 _30694_ (.A(_10572_),
    .B(net4640),
    .Y(_07835_));
 sg13g2_a21oi_1 _30695_ (.A1(net4640),
    .A2(_07834_),
    .Y(_07836_),
    .B1(_07835_));
 sg13g2_nand3_1 _30696_ (.B(_11120_),
    .C(_11140_),
    .A(_11119_),
    .Y(_07837_));
 sg13g2_nand2b_1 _30697_ (.Y(_07838_),
    .B(_07837_),
    .A_N(_11141_));
 sg13g2_o21ai_1 _30698_ (.B1(net4002),
    .Y(_07839_),
    .A1(net4602),
    .A2(net1300));
 sg13g2_a221oi_1 _30699_ (.B2(net3689),
    .C1(_07839_),
    .B1(_07838_),
    .A1(net3711),
    .Y(_07840_),
    .A2(_07836_));
 sg13g2_a21o_1 _30700_ (.A2(net3918),
    .A1(net2122),
    .B1(_07840_),
    .X(_01309_));
 sg13g2_xor2_1 _30701_ (.B(_12683_),
    .A(_11117_),
    .X(_07841_));
 sg13g2_mux2_1 _30702_ (.A0(net2705),
    .A1(_07841_),
    .S(net4640),
    .X(_07842_));
 sg13g2_or3_1 _30703_ (.A(_11117_),
    .B(_11118_),
    .C(_11141_),
    .X(_07843_));
 sg13g2_nand2_1 _30704_ (.Y(_07844_),
    .A(_11142_),
    .B(_07843_));
 sg13g2_o21ai_1 _30705_ (.B1(net4002),
    .Y(_07845_),
    .A1(net4602),
    .A2(net3257));
 sg13g2_a21oi_1 _30706_ (.A1(net3689),
    .A2(_07844_),
    .Y(_07846_),
    .B1(_07845_));
 sg13g2_o21ai_1 _30707_ (.B1(_07846_),
    .Y(_07847_),
    .A1(net3701),
    .A2(_07842_));
 sg13g2_o21ai_1 _30708_ (.B1(_07847_),
    .Y(_01310_),
    .A1(_10572_),
    .A2(net4002));
 sg13g2_nor2_1 _30709_ (.A(net2705),
    .B(net4002),
    .Y(_07848_));
 sg13g2_xnor2_1 _30710_ (.Y(_07849_),
    .A(_11114_),
    .B(_12684_));
 sg13g2_o21ai_1 _30711_ (.B1(net3711),
    .Y(_07850_),
    .A1(\u_inv.f_next[8] ),
    .A2(net4641));
 sg13g2_a21oi_1 _30712_ (.A1(net4641),
    .A2(_07849_),
    .Y(_07851_),
    .B1(_07850_));
 sg13g2_nand3_1 _30713_ (.B(_11115_),
    .C(_11142_),
    .A(_11114_),
    .Y(_07852_));
 sg13g2_and2_1 _30714_ (.A(_11143_),
    .B(_07852_),
    .X(_07853_));
 sg13g2_a221oi_1 _30715_ (.B2(_07853_),
    .C1(_07851_),
    .B1(net3690),
    .A1(net4512),
    .Y(_07854_),
    .A2(net1670));
 sg13g2_a21oi_1 _30716_ (.A1(net4003),
    .A2(_07854_),
    .Y(_01311_),
    .B1(_07848_));
 sg13g2_xnor2_1 _30717_ (.Y(_07855_),
    .A(_11112_),
    .B(_12685_));
 sg13g2_nand2_1 _30718_ (.Y(_07856_),
    .A(net4641),
    .B(_07855_));
 sg13g2_a21oi_1 _30719_ (.A1(net2394),
    .A2(net4527),
    .Y(_07857_),
    .B1(net3701));
 sg13g2_o21ai_1 _30720_ (.B1(net4002),
    .Y(_07858_),
    .A1(net4608),
    .A2(net2059));
 sg13g2_nand3_1 _30721_ (.B(_11143_),
    .C(_11144_),
    .A(_11112_),
    .Y(_07859_));
 sg13g2_nand2b_1 _30722_ (.Y(_07860_),
    .B(_07859_),
    .A_N(_11145_));
 sg13g2_a221oi_1 _30723_ (.B2(net3690),
    .C1(_07858_),
    .B1(_07860_),
    .A1(_07856_),
    .Y(_07861_),
    .A2(_07857_));
 sg13g2_a21o_1 _30724_ (.A2(net3919),
    .A1(net3025),
    .B1(_07861_),
    .X(_01312_));
 sg13g2_nand2_1 _30725_ (.Y(_07862_),
    .A(net2394),
    .B(net3918));
 sg13g2_o21ai_1 _30726_ (.B1(_11109_),
    .Y(_07863_),
    .A1(_11111_),
    .A2(_12686_));
 sg13g2_a21oi_1 _30727_ (.A1(_12687_),
    .A2(_07863_),
    .Y(_07864_),
    .B1(net4527));
 sg13g2_a21oi_1 _30728_ (.A1(_10571_),
    .A2(net4527),
    .Y(_07865_),
    .B1(_07864_));
 sg13g2_nor3_1 _30729_ (.A(_11109_),
    .B(_11110_),
    .C(_11145_),
    .Y(_07866_));
 sg13g2_o21ai_1 _30730_ (.B1(net4379),
    .Y(_07867_),
    .A1(_11147_),
    .A2(_07866_));
 sg13g2_a22oi_1 _30731_ (.Y(_07868_),
    .B1(_07867_),
    .B2(net3701),
    .A2(_07865_),
    .A1(net3828));
 sg13g2_o21ai_1 _30732_ (.B1(net4003),
    .Y(_07869_),
    .A1(net4608),
    .A2(net1815));
 sg13g2_o21ai_1 _30733_ (.B1(_07862_),
    .Y(_01313_),
    .A1(_07868_),
    .A2(_07869_));
 sg13g2_a21oi_1 _30734_ (.A1(_10570_),
    .A2(net4527),
    .Y(_07870_),
    .B1(net3743));
 sg13g2_xnor2_1 _30735_ (.Y(_07871_),
    .A(_12688_),
    .B(_12690_));
 sg13g2_o21ai_1 _30736_ (.B1(_07870_),
    .Y(_07872_),
    .A1(net4528),
    .A2(_07871_));
 sg13g2_xor2_1 _30737_ (.B(_12690_),
    .A(_11148_),
    .X(_07873_));
 sg13g2_a21oi_1 _30738_ (.A1(net3743),
    .A2(_07873_),
    .Y(_07874_),
    .B1(net4436));
 sg13g2_a21oi_1 _30739_ (.A1(_07872_),
    .A2(_07874_),
    .Y(_07875_),
    .B1(net3918));
 sg13g2_o21ai_1 _30740_ (.B1(_07875_),
    .Y(_07876_),
    .A1(net4602),
    .A2(net1999));
 sg13g2_o21ai_1 _30741_ (.B1(_07876_),
    .Y(_01314_),
    .A1(_10571_),
    .A2(net4003));
 sg13g2_xnor2_1 _30742_ (.Y(_07877_),
    .A(_11153_),
    .B(_12692_));
 sg13g2_o21ai_1 _30743_ (.B1(net3711),
    .Y(_07878_),
    .A1(_10569_),
    .A2(net4640));
 sg13g2_a21oi_1 _30744_ (.A1(net4640),
    .A2(_07877_),
    .Y(_07879_),
    .B1(_07878_));
 sg13g2_nand2_1 _30745_ (.Y(_07880_),
    .A(_11151_),
    .B(_11153_));
 sg13g2_a21oi_1 _30746_ (.A1(_11155_),
    .A2(_07880_),
    .Y(_07881_),
    .B1(net3679));
 sg13g2_o21ai_1 _30747_ (.B1(net4003),
    .Y(_07882_),
    .A1(net4602),
    .A2(net1963));
 sg13g2_nor3_1 _30748_ (.A(_07879_),
    .B(_07881_),
    .C(_07882_),
    .Y(_07883_));
 sg13g2_a21o_1 _30749_ (.A2(net3918),
    .A1(net3044),
    .B1(_07883_),
    .X(_01315_));
 sg13g2_nand2_1 _30750_ (.Y(_07884_),
    .A(net2528),
    .B(net3918));
 sg13g2_nand2_1 _30751_ (.Y(_07885_),
    .A(\u_inv.f_next[13] ),
    .B(net3828));
 sg13g2_o21ai_1 _30752_ (.B1(_11152_),
    .Y(_07886_),
    .A1(_11154_),
    .A2(_12692_));
 sg13g2_xor2_1 _30753_ (.B(_07886_),
    .A(_11106_),
    .X(_07887_));
 sg13g2_a22oi_1 _30754_ (.Y(_07888_),
    .B1(_07887_),
    .B2(net4640),
    .A2(_07885_),
    .A1(net3723));
 sg13g2_o21ai_1 _30755_ (.B1(_11155_),
    .Y(_07889_),
    .A1(_10569_),
    .A2(\u_inv.f_reg[12] ));
 sg13g2_o21ai_1 _30756_ (.B1(net3743),
    .Y(_07890_),
    .A1(_11106_),
    .A2(_07889_));
 sg13g2_a21oi_1 _30757_ (.A1(_11106_),
    .A2(_07889_),
    .Y(_07891_),
    .B1(_07890_));
 sg13g2_nor3_1 _30758_ (.A(net4436),
    .B(_07888_),
    .C(_07891_),
    .Y(_07892_));
 sg13g2_o21ai_1 _30759_ (.B1(net4002),
    .Y(_07893_),
    .A1(net4604),
    .A2(net1862));
 sg13g2_o21ai_1 _30760_ (.B1(_07884_),
    .Y(_01316_),
    .A1(_07892_),
    .A2(_07893_));
 sg13g2_nor2_1 _30761_ (.A(_10568_),
    .B(net4008),
    .Y(_07894_));
 sg13g2_xnor2_1 _30762_ (.Y(_07895_),
    .A(_11102_),
    .B(_12694_));
 sg13g2_a21oi_1 _30763_ (.A1(net3297),
    .A2(net4536),
    .Y(_07896_),
    .B1(net3701));
 sg13g2_o21ai_1 _30764_ (.B1(_07896_),
    .Y(_07897_),
    .A1(net4536),
    .A2(_07895_));
 sg13g2_o21ai_1 _30765_ (.B1(net4008),
    .Y(_07898_),
    .A1(net4606),
    .A2(net1875));
 sg13g2_and2_1 _30766_ (.A(_11156_),
    .B(_11162_),
    .X(_07899_));
 sg13g2_xnor2_1 _30767_ (.Y(_07900_),
    .A(_11102_),
    .B(_07899_));
 sg13g2_a21oi_1 _30768_ (.A1(net3689),
    .A2(_07900_),
    .Y(_07901_),
    .B1(_07898_));
 sg13g2_a21o_1 _30769_ (.A2(_07901_),
    .A1(_07897_),
    .B1(_07894_),
    .X(_01317_));
 sg13g2_nand2_1 _30770_ (.Y(_07902_),
    .A(net3064),
    .B(net3832));
 sg13g2_a21oi_1 _30771_ (.A1(_11102_),
    .A2(_12694_),
    .Y(_07903_),
    .B1(_11101_));
 sg13g2_xnor2_1 _30772_ (.Y(_07904_),
    .A(_11100_),
    .B(_07903_));
 sg13g2_a22oi_1 _30773_ (.Y(_07905_),
    .B1(_07904_),
    .B2(net4650),
    .A2(_07902_),
    .A1(net3729));
 sg13g2_o21ai_1 _30774_ (.B1(_11159_),
    .Y(_07906_),
    .A1(_11102_),
    .A2(_07899_));
 sg13g2_xnor2_1 _30775_ (.Y(_07907_),
    .A(_11100_),
    .B(_07906_));
 sg13g2_o21ai_1 _30776_ (.B1(net4378),
    .Y(_07908_),
    .A1(net3832),
    .A2(_07907_));
 sg13g2_a21oi_1 _30777_ (.A1(net4511),
    .A2(_10958_),
    .Y(_07909_),
    .B1(net3927));
 sg13g2_o21ai_1 _30778_ (.B1(_07909_),
    .Y(_07910_),
    .A1(_07905_),
    .A2(_07908_));
 sg13g2_o21ai_1 _30779_ (.B1(_07910_),
    .Y(_01318_),
    .A1(_10567_),
    .A2(net4008));
 sg13g2_a21oi_1 _30780_ (.A1(_11168_),
    .A2(_12699_),
    .Y(_07911_),
    .B1(net4536));
 sg13g2_o21ai_1 _30781_ (.B1(_07911_),
    .Y(_07912_),
    .A1(_11168_),
    .A2(_12699_));
 sg13g2_a21oi_1 _30782_ (.A1(\u_inv.f_next[16] ),
    .A2(net4536),
    .Y(_07913_),
    .B1(net3701));
 sg13g2_xnor2_1 _30783_ (.Y(_07914_),
    .A(_11166_),
    .B(_11168_));
 sg13g2_o21ai_1 _30784_ (.B1(net4008),
    .Y(_07915_),
    .A1(net4606),
    .A2(net1785));
 sg13g2_a221oi_1 _30785_ (.B2(net3689),
    .C1(_07915_),
    .B1(_07914_),
    .A1(_07912_),
    .Y(_07916_),
    .A2(_07913_));
 sg13g2_a21o_1 _30786_ (.A2(net3927),
    .A1(net3064),
    .B1(_07916_),
    .X(_01319_));
 sg13g2_nand2_1 _30787_ (.Y(_07917_),
    .A(net1744),
    .B(net3832));
 sg13g2_a21oi_1 _30788_ (.A1(_11168_),
    .A2(_12699_),
    .Y(_07918_),
    .B1(_11167_));
 sg13g2_xor2_1 _30789_ (.B(_07918_),
    .A(_11094_),
    .X(_07919_));
 sg13g2_a22oi_1 _30790_ (.Y(_07920_),
    .B1(_07919_),
    .B2(net4650),
    .A2(_07917_),
    .A1(net3724));
 sg13g2_a21oi_1 _30791_ (.A1(_11170_),
    .A2(_11176_),
    .Y(_07921_),
    .B1(_11094_));
 sg13g2_nand3_1 _30792_ (.B(_11170_),
    .C(_11176_),
    .A(_11094_),
    .Y(_07922_));
 sg13g2_nand2_1 _30793_ (.Y(_07923_),
    .A(net3752),
    .B(_07922_));
 sg13g2_o21ai_1 _30794_ (.B1(net4378),
    .Y(_07924_),
    .A1(_07921_),
    .A2(_07923_));
 sg13g2_a21oi_1 _30795_ (.A1(net4511),
    .A2(_10959_),
    .Y(_07925_),
    .B1(net3927));
 sg13g2_o21ai_1 _30796_ (.B1(_07925_),
    .Y(_07926_),
    .A1(_07920_),
    .A2(_07924_));
 sg13g2_o21ai_1 _30797_ (.B1(_07926_),
    .Y(_01320_),
    .A1(_10565_),
    .A2(net4008));
 sg13g2_nand2_1 _30798_ (.Y(_07927_),
    .A(net1744),
    .B(net3927));
 sg13g2_nor3_1 _30799_ (.A(_11093_),
    .B(_11175_),
    .C(_07921_),
    .Y(_07928_));
 sg13g2_o21ai_1 _30800_ (.B1(_11093_),
    .Y(_07929_),
    .A1(_11175_),
    .A2(_07921_));
 sg13g2_nor2b_1 _30801_ (.A(_07928_),
    .B_N(_07929_),
    .Y(_07930_));
 sg13g2_o21ai_1 _30802_ (.B1(net4009),
    .Y(_07931_),
    .A1(net4606),
    .A2(\u_inv.input_reg[17] ));
 sg13g2_or2_1 _30803_ (.X(_07932_),
    .B(_12704_),
    .A(_12701_));
 sg13g2_nand2_1 _30804_ (.Y(_07933_),
    .A(_11092_),
    .B(_07932_));
 sg13g2_xnor2_1 _30805_ (.Y(_07934_),
    .A(_11092_),
    .B(_07932_));
 sg13g2_a21oi_1 _30806_ (.A1(\u_inv.f_next[18] ),
    .A2(net4536),
    .Y(_07935_),
    .B1(net3702));
 sg13g2_o21ai_1 _30807_ (.B1(_07935_),
    .Y(_07936_),
    .A1(net4536),
    .A2(_07934_));
 sg13g2_o21ai_1 _30808_ (.B1(_07936_),
    .Y(_07937_),
    .A1(net3680),
    .A2(_07930_));
 sg13g2_o21ai_1 _30809_ (.B1(_07927_),
    .Y(_01321_),
    .A1(_07931_),
    .A2(_07937_));
 sg13g2_and2_1 _30810_ (.A(_11091_),
    .B(_07933_),
    .X(_07938_));
 sg13g2_xnor2_1 _30811_ (.Y(_07939_),
    .A(_11098_),
    .B(_07938_));
 sg13g2_o21ai_1 _30812_ (.B1(net3712),
    .Y(_07940_),
    .A1(net2812),
    .A2(net4650));
 sg13g2_a21oi_1 _30813_ (.A1(net4651),
    .A2(_07939_),
    .Y(_07941_),
    .B1(_07940_));
 sg13g2_and2_1 _30814_ (.A(_11174_),
    .B(_07929_),
    .X(_07942_));
 sg13g2_o21ai_1 _30815_ (.B1(net3691),
    .Y(_07943_),
    .A1(_11097_),
    .A2(_07942_));
 sg13g2_a21oi_1 _30816_ (.A1(_11097_),
    .A2(_07942_),
    .Y(_07944_),
    .B1(_07943_));
 sg13g2_nor2b_1 _30817_ (.A(net4604),
    .B_N(net1619),
    .Y(_07945_));
 sg13g2_nor4_1 _30818_ (.A(net3927),
    .B(_07941_),
    .C(_07944_),
    .D(_07945_),
    .Y(_07946_));
 sg13g2_a21oi_1 _30819_ (.A1(_10563_),
    .A2(net3927),
    .Y(_01322_),
    .B1(_07946_));
 sg13g2_and2_1 _30820_ (.A(_11183_),
    .B(_12707_),
    .X(_07947_));
 sg13g2_o21ai_1 _30821_ (.B1(net4650),
    .Y(_07948_),
    .A1(_11183_),
    .A2(_12707_));
 sg13g2_a21oi_1 _30822_ (.A1(net2622),
    .A2(net4536),
    .Y(_07949_),
    .B1(net3701));
 sg13g2_o21ai_1 _30823_ (.B1(_07949_),
    .Y(_07950_),
    .A1(_07947_),
    .A2(_07948_));
 sg13g2_nand3_1 _30824_ (.B(_11180_),
    .C(_11182_),
    .A(_11172_),
    .Y(_07951_));
 sg13g2_nand2b_1 _30825_ (.Y(_07952_),
    .B(_07951_),
    .A_N(_11184_));
 sg13g2_o21ai_1 _30826_ (.B1(net4009),
    .Y(_07953_),
    .A1(net4604),
    .A2(net1855));
 sg13g2_a21oi_1 _30827_ (.A1(net3691),
    .A2(_07952_),
    .Y(_07954_),
    .B1(_07953_));
 sg13g2_nand2_1 _30828_ (.Y(_07955_),
    .A(_07950_),
    .B(_07954_));
 sg13g2_o21ai_1 _30829_ (.B1(_07955_),
    .Y(_01323_),
    .A1(_10562_),
    .A2(net4008));
 sg13g2_nand2_1 _30830_ (.Y(_07956_),
    .A(net2622),
    .B(net3927));
 sg13g2_a21oi_1 _30831_ (.A1(_10560_),
    .A2(net4538),
    .Y(_07957_),
    .B1(net3753));
 sg13g2_o21ai_1 _30832_ (.B1(_11181_),
    .Y(_07958_),
    .A1(_11183_),
    .A2(_12707_));
 sg13g2_o21ai_1 _30833_ (.B1(net4650),
    .Y(_07959_),
    .A1(_11187_),
    .A2(_07958_));
 sg13g2_a21o_1 _30834_ (.A2(_07958_),
    .A1(_11187_),
    .B1(_07959_),
    .X(_07960_));
 sg13g2_nor2_1 _30835_ (.A(_11184_),
    .B(_11196_),
    .Y(_07961_));
 sg13g2_o21ai_1 _30836_ (.B1(_11187_),
    .Y(_07962_),
    .A1(_11184_),
    .A2(_11196_));
 sg13g2_xnor2_1 _30837_ (.Y(_07963_),
    .A(_11187_),
    .B(_07961_));
 sg13g2_a221oi_1 _30838_ (.B2(net3753),
    .C1(net4438),
    .B1(_07963_),
    .A1(_07957_),
    .Y(_07964_),
    .A2(_07960_));
 sg13g2_o21ai_1 _30839_ (.B1(net4008),
    .Y(_07965_),
    .A1(net4604),
    .A2(net2065));
 sg13g2_o21ai_1 _30840_ (.B1(_07956_),
    .Y(_01324_),
    .A1(_07964_),
    .A2(_07965_));
 sg13g2_nand2_1 _30841_ (.Y(_07966_),
    .A(_11195_),
    .B(_07962_));
 sg13g2_a21oi_1 _30842_ (.A1(_11195_),
    .A2(_07962_),
    .Y(_07967_),
    .B1(_11186_));
 sg13g2_xnor2_1 _30843_ (.Y(_07968_),
    .A(_11186_),
    .B(_07966_));
 sg13g2_nor2_1 _30844_ (.A(net3679),
    .B(_07968_),
    .Y(_07969_));
 sg13g2_nor3_1 _30845_ (.A(_11183_),
    .B(_11187_),
    .C(_12707_),
    .Y(_07970_));
 sg13g2_o21ai_1 _30846_ (.B1(_11186_),
    .Y(_07971_),
    .A1(_12713_),
    .A2(_07970_));
 sg13g2_or3_1 _30847_ (.A(_11186_),
    .B(_12713_),
    .C(_07970_),
    .X(_07972_));
 sg13g2_and2_1 _30848_ (.A(_07971_),
    .B(_07972_),
    .X(_07973_));
 sg13g2_o21ai_1 _30849_ (.B1(net3712),
    .Y(_07974_),
    .A1(_10559_),
    .A2(net4650));
 sg13g2_a21oi_1 _30850_ (.A1(net4650),
    .A2(_07973_),
    .Y(_07975_),
    .B1(_07974_));
 sg13g2_nor3_1 _30851_ (.A(net3927),
    .B(_07969_),
    .C(_07975_),
    .Y(_07976_));
 sg13g2_o21ai_1 _30852_ (.B1(_07976_),
    .Y(_07977_),
    .A1(net4606),
    .A2(net1962));
 sg13g2_o21ai_1 _30853_ (.B1(_07977_),
    .Y(_01325_),
    .A1(_10560_),
    .A2(net4009));
 sg13g2_nand2_1 _30854_ (.Y(_07978_),
    .A(net2961),
    .B(net3832));
 sg13g2_nand2_1 _30855_ (.Y(_07979_),
    .A(_11185_),
    .B(_07971_));
 sg13g2_xnor2_1 _30856_ (.Y(_07980_),
    .A(_11188_),
    .B(_07979_));
 sg13g2_a22oi_1 _30857_ (.Y(_07981_),
    .B1(_07980_),
    .B2(net4650),
    .A2(_07978_),
    .A1(net3724));
 sg13g2_nor2_1 _30858_ (.A(_11194_),
    .B(_07967_),
    .Y(_07982_));
 sg13g2_xnor2_1 _30859_ (.Y(_07983_),
    .A(_11189_),
    .B(_07982_));
 sg13g2_a21oi_1 _30860_ (.A1(net3753),
    .A2(_07983_),
    .Y(_07984_),
    .B1(_07981_));
 sg13g2_o21ai_1 _30861_ (.B1(net4011),
    .Y(_07985_),
    .A1(net4606),
    .A2(net1937));
 sg13g2_a21o_1 _30862_ (.A2(_07984_),
    .A1(net4378),
    .B1(_07985_),
    .X(_07986_));
 sg13g2_o21ai_1 _30863_ (.B1(_07986_),
    .Y(_01326_),
    .A1(_10559_),
    .A2(net4009));
 sg13g2_nand2_1 _30864_ (.Y(_07987_),
    .A(_11202_),
    .B(_12715_));
 sg13g2_xnor2_1 _30865_ (.Y(_07988_),
    .A(_11201_),
    .B(_12715_));
 sg13g2_o21ai_1 _30866_ (.B1(net3712),
    .Y(_07989_),
    .A1(_10557_),
    .A2(net4652));
 sg13g2_a21oi_1 _30867_ (.A1(net4652),
    .A2(_07988_),
    .Y(_07990_),
    .B1(_07989_));
 sg13g2_xnor2_1 _30868_ (.Y(_07991_),
    .A(_11200_),
    .B(_11202_));
 sg13g2_o21ai_1 _30869_ (.B1(net4011),
    .Y(_07992_),
    .A1(net4605),
    .A2(net1912));
 sg13g2_a21oi_1 _30870_ (.A1(net3691),
    .A2(_07991_),
    .Y(_07993_),
    .B1(_07992_));
 sg13g2_nand2b_1 _30871_ (.Y(_07994_),
    .B(_07993_),
    .A_N(_07990_));
 sg13g2_o21ai_1 _30872_ (.B1(_07994_),
    .Y(_01327_),
    .A1(_10558_),
    .A2(net4008));
 sg13g2_nand2_1 _30873_ (.Y(_07995_),
    .A(net1754),
    .B(net3929));
 sg13g2_a21oi_1 _30874_ (.A1(_10556_),
    .A2(net4539),
    .Y(_07996_),
    .B1(net3754));
 sg13g2_o21ai_1 _30875_ (.B1(_07987_),
    .Y(_07997_),
    .A1(_10557_),
    .A2(_10865_));
 sg13g2_a21oi_1 _30876_ (.A1(_11204_),
    .A2(_07997_),
    .Y(_07998_),
    .B1(net4538));
 sg13g2_o21ai_1 _30877_ (.B1(_07998_),
    .Y(_07999_),
    .A1(_11204_),
    .A2(_07997_));
 sg13g2_o21ai_1 _30878_ (.B1(_11216_),
    .Y(_08000_),
    .A1(_11200_),
    .A2(_11202_));
 sg13g2_xnor2_1 _30879_ (.Y(_08001_),
    .A(_11203_),
    .B(_08000_));
 sg13g2_a221oi_1 _30880_ (.B2(net3754),
    .C1(net4438),
    .B1(_08001_),
    .A1(_07996_),
    .Y(_08002_),
    .A2(_07999_));
 sg13g2_o21ai_1 _30881_ (.B1(net4011),
    .Y(_08003_),
    .A1(net4605),
    .A2(\u_inv.input_reg[24] ));
 sg13g2_o21ai_1 _30882_ (.B1(_07995_),
    .Y(_01328_),
    .A1(_08002_),
    .A2(_08003_));
 sg13g2_o21ai_1 _30883_ (.B1(_12723_),
    .Y(_08004_),
    .A1(_11204_),
    .A2(_07987_));
 sg13g2_o21ai_1 _30884_ (.B1(net4652),
    .Y(_08005_),
    .A1(_11207_),
    .A2(_08004_));
 sg13g2_a21o_1 _30885_ (.A2(_08004_),
    .A1(_11207_),
    .B1(_08005_),
    .X(_08006_));
 sg13g2_a21oi_1 _30886_ (.A1(\u_inv.f_next[26] ),
    .A2(net4538),
    .Y(_08007_),
    .B1(net3702));
 sg13g2_a21oi_1 _30887_ (.A1(_11204_),
    .A2(_08000_),
    .Y(_08008_),
    .B1(_11220_));
 sg13g2_xnor2_1 _30888_ (.Y(_08009_),
    .A(_11207_),
    .B(_08008_));
 sg13g2_a221oi_1 _30889_ (.B2(net3691),
    .C1(net3929),
    .B1(_08009_),
    .A1(_08006_),
    .Y(_08010_),
    .A2(_08007_));
 sg13g2_o21ai_1 _30890_ (.B1(_08010_),
    .Y(_08011_),
    .A1(net4605),
    .A2(net1737));
 sg13g2_o21ai_1 _30891_ (.B1(_08011_),
    .Y(_01329_),
    .A1(_10556_),
    .A2(net4011));
 sg13g2_a21oi_1 _30892_ (.A1(_11207_),
    .A2(_08004_),
    .Y(_08012_),
    .B1(_11205_));
 sg13g2_xor2_1 _30893_ (.B(_08012_),
    .A(_11208_),
    .X(_08013_));
 sg13g2_nand2_1 _30894_ (.Y(_08014_),
    .A(net3133),
    .B(net3833));
 sg13g2_a22oi_1 _30895_ (.Y(_08015_),
    .B1(_08014_),
    .B2(net3724),
    .A2(_08013_),
    .A1(net4652));
 sg13g2_o21ai_1 _30896_ (.B1(_11217_),
    .Y(_08016_),
    .A1(_11207_),
    .A2(_08008_));
 sg13g2_xor2_1 _30897_ (.B(_08016_),
    .A(_11208_),
    .X(_08017_));
 sg13g2_o21ai_1 _30898_ (.B1(net4378),
    .Y(_08018_),
    .A1(net3833),
    .A2(_08017_));
 sg13g2_a21oi_1 _30899_ (.A1(net4512),
    .A2(_10960_),
    .Y(_08019_),
    .B1(net3930));
 sg13g2_o21ai_1 _30900_ (.B1(_08019_),
    .Y(_08020_),
    .A1(_08015_),
    .A2(_08018_));
 sg13g2_o21ai_1 _30901_ (.B1(_08020_),
    .Y(_01330_),
    .A1(_10555_),
    .A2(net4011));
 sg13g2_a21oi_2 _30902_ (.B1(_12725_),
    .Y(_08021_),
    .A2(_08004_),
    .A1(_12719_));
 sg13g2_xnor2_1 _30903_ (.Y(_08022_),
    .A(_11088_),
    .B(_08021_));
 sg13g2_o21ai_1 _30904_ (.B1(net3712),
    .Y(_08023_),
    .A1(_10553_),
    .A2(net4652));
 sg13g2_a21oi_1 _30905_ (.A1(net4652),
    .A2(_08022_),
    .Y(_08024_),
    .B1(_08023_));
 sg13g2_or2_1 _30906_ (.X(_08025_),
    .B(_11223_),
    .A(_11211_));
 sg13g2_xnor2_1 _30907_ (.Y(_08026_),
    .A(_11088_),
    .B(_08025_));
 sg13g2_o21ai_1 _30908_ (.B1(net4012),
    .Y(_08027_),
    .A1(net4605),
    .A2(net1837));
 sg13g2_nor2_1 _30909_ (.A(_08024_),
    .B(_08027_),
    .Y(_08028_));
 sg13g2_o21ai_1 _30910_ (.B1(_08028_),
    .Y(_08029_),
    .A1(net3679),
    .A2(_08026_));
 sg13g2_o21ai_1 _30911_ (.B1(_08029_),
    .Y(_01331_),
    .A1(_10554_),
    .A2(net4011));
 sg13g2_o21ai_1 _30912_ (.B1(_11087_),
    .Y(_08030_),
    .A1(_11089_),
    .A2(_08021_));
 sg13g2_xnor2_1 _30913_ (.Y(_08031_),
    .A(_11086_),
    .B(_08030_));
 sg13g2_o21ai_1 _30914_ (.B1(net3712),
    .Y(_08032_),
    .A1(_10552_),
    .A2(net4653));
 sg13g2_a21oi_1 _30915_ (.A1(net4653),
    .A2(_08031_),
    .Y(_08033_),
    .B1(_08032_));
 sg13g2_a21oi_1 _30916_ (.A1(_11089_),
    .A2(_08025_),
    .Y(_08034_),
    .B1(_11215_));
 sg13g2_xnor2_1 _30917_ (.Y(_08035_),
    .A(_11086_),
    .B(_08034_));
 sg13g2_o21ai_1 _30918_ (.B1(net4011),
    .Y(_08036_),
    .A1(net4605),
    .A2(net1784));
 sg13g2_nor2_1 _30919_ (.A(_08033_),
    .B(_08036_),
    .Y(_08037_));
 sg13g2_o21ai_1 _30920_ (.B1(_08037_),
    .Y(_08038_),
    .A1(net3680),
    .A2(_08035_));
 sg13g2_o21ai_1 _30921_ (.B1(_08038_),
    .Y(_01332_),
    .A1(_10553_),
    .A2(net4011));
 sg13g2_or2_1 _30922_ (.X(_08039_),
    .B(_08021_),
    .A(_12717_));
 sg13g2_a21oi_1 _30923_ (.A1(_12729_),
    .A2(_08039_),
    .Y(_08040_),
    .B1(_11083_));
 sg13g2_nand3_1 _30924_ (.B(_12729_),
    .C(_08039_),
    .A(_11083_),
    .Y(_08041_));
 sg13g2_nand3b_1 _30925_ (.B(_08041_),
    .C(net4653),
    .Y(_08042_),
    .A_N(_08040_));
 sg13g2_a21oi_1 _30926_ (.A1(\u_inv.f_next[30] ),
    .A2(net4538),
    .Y(_08043_),
    .B1(net3702));
 sg13g2_o21ai_1 _30927_ (.B1(_11214_),
    .Y(_08044_),
    .A1(_11085_),
    .A2(_08034_));
 sg13g2_xnor2_1 _30928_ (.Y(_08045_),
    .A(_11083_),
    .B(_08044_));
 sg13g2_o21ai_1 _30929_ (.B1(net4012),
    .Y(_08046_),
    .A1(net4605),
    .A2(net1747));
 sg13g2_a221oi_1 _30930_ (.B2(net3691),
    .C1(_08046_),
    .B1(_08045_),
    .A1(_08042_),
    .Y(_08047_),
    .A2(_08043_));
 sg13g2_a21o_1 _30931_ (.A2(net3930),
    .A1(net3119),
    .B1(_08047_),
    .X(_01333_));
 sg13g2_nand2_1 _30932_ (.Y(_08048_),
    .A(net2712),
    .B(net3833));
 sg13g2_a21oi_1 _30933_ (.A1(\u_inv.f_next[30] ),
    .A2(\u_inv.f_reg[30] ),
    .Y(_08049_),
    .B1(_08040_));
 sg13g2_xnor2_1 _30934_ (.Y(_08050_),
    .A(_11080_),
    .B(_08049_));
 sg13g2_a22oi_1 _30935_ (.Y(_08051_),
    .B1(_08050_),
    .B2(net4653),
    .A2(_08048_),
    .A1(net3724));
 sg13g2_a21oi_1 _30936_ (.A1(_11083_),
    .A2(_08044_),
    .Y(_08052_),
    .B1(_11226_));
 sg13g2_xnor2_1 _30937_ (.Y(_08053_),
    .A(_11079_),
    .B(_08052_));
 sg13g2_o21ai_1 _30938_ (.B1(net4382),
    .Y(_08054_),
    .A1(net3833),
    .A2(_08053_));
 sg13g2_a21oi_1 _30939_ (.A1(net4512),
    .A2(_10961_),
    .Y(_08055_),
    .B1(net3930));
 sg13g2_o21ai_1 _30940_ (.B1(_08055_),
    .Y(_08056_),
    .A1(_08051_),
    .A2(_08054_));
 sg13g2_o21ai_1 _30941_ (.B1(_08056_),
    .Y(_01334_),
    .A1(_10551_),
    .A2(net4012));
 sg13g2_nand2b_1 _30942_ (.Y(_08057_),
    .B(_11236_),
    .A_N(_12733_));
 sg13g2_xnor2_1 _30943_ (.Y(_08058_),
    .A(_11235_),
    .B(_12733_));
 sg13g2_o21ai_1 _30944_ (.B1(net3712),
    .Y(_08059_),
    .A1(net2280),
    .A2(net4652));
 sg13g2_a21oi_1 _30945_ (.A1(net4652),
    .A2(_08058_),
    .Y(_08060_),
    .B1(_08059_));
 sg13g2_nand2_1 _30946_ (.Y(_08061_),
    .A(_11230_),
    .B(_11235_));
 sg13g2_o21ai_1 _30947_ (.B1(net3691),
    .Y(_08062_),
    .A1(_11230_),
    .A2(_11235_));
 sg13g2_nor2b_1 _30948_ (.A(_08062_),
    .B_N(_08061_),
    .Y(_08063_));
 sg13g2_nor2b_1 _30949_ (.A(net4610),
    .B_N(net1663),
    .Y(_08064_));
 sg13g2_nor4_1 _30950_ (.A(net3930),
    .B(_08060_),
    .C(_08063_),
    .D(_08064_),
    .Y(_08065_));
 sg13g2_a21oi_1 _30951_ (.A1(_10550_),
    .A2(net3930),
    .Y(_01335_),
    .B1(_08065_));
 sg13g2_a21oi_1 _30952_ (.A1(_11257_),
    .A2(_08061_),
    .Y(_08066_),
    .B1(_11239_));
 sg13g2_nand3_1 _30953_ (.B(_11257_),
    .C(_08061_),
    .A(_11239_),
    .Y(_08067_));
 sg13g2_nand2_1 _30954_ (.Y(_08068_),
    .A(net3691),
    .B(_08067_));
 sg13g2_and2_1 _30955_ (.A(_11234_),
    .B(_08057_),
    .X(_08069_));
 sg13g2_xnor2_1 _30956_ (.Y(_08070_),
    .A(_11240_),
    .B(_08069_));
 sg13g2_o21ai_1 _30957_ (.B1(net3713),
    .Y(_08071_),
    .A1(\u_inv.f_next[33] ),
    .A2(net4662));
 sg13g2_a21oi_1 _30958_ (.A1(net4662),
    .A2(_08070_),
    .Y(_08072_),
    .B1(_08071_));
 sg13g2_nand2_1 _30959_ (.Y(_08073_),
    .A(net4512),
    .B(net1694));
 sg13g2_o21ai_1 _30960_ (.B1(_08073_),
    .Y(_08074_),
    .A1(_08066_),
    .A2(_08068_));
 sg13g2_nor3_1 _30961_ (.A(net3936),
    .B(_08072_),
    .C(_08074_),
    .Y(_08075_));
 sg13g2_a21oi_1 _30962_ (.A1(_10549_),
    .A2(net3936),
    .Y(_01336_),
    .B1(_08075_));
 sg13g2_nor2_1 _30963_ (.A(_11256_),
    .B(_08066_),
    .Y(_08076_));
 sg13g2_nor2_1 _30964_ (.A(_11232_),
    .B(_08076_),
    .Y(_08077_));
 sg13g2_a21oi_1 _30965_ (.A1(_11232_),
    .A2(_08076_),
    .Y(_08078_),
    .B1(net3680));
 sg13g2_nor2b_1 _30966_ (.A(_08077_),
    .B_N(_08078_),
    .Y(_08079_));
 sg13g2_o21ai_1 _30967_ (.B1(_11238_),
    .Y(_08080_),
    .A1(_11237_),
    .A2(_08069_));
 sg13g2_nand2_1 _30968_ (.Y(_08081_),
    .A(_11232_),
    .B(_08080_));
 sg13g2_xnor2_1 _30969_ (.Y(_08082_),
    .A(_11232_),
    .B(_08080_));
 sg13g2_a21oi_1 _30970_ (.A1(net4662),
    .A2(_08082_),
    .Y(_08083_),
    .B1(net3702));
 sg13g2_o21ai_1 _30971_ (.B1(_08083_),
    .Y(_08084_),
    .A1(net2896),
    .A2(net4662));
 sg13g2_nor2b_1 _30972_ (.A(net4610),
    .B_N(net1717),
    .Y(_08085_));
 sg13g2_nor3_1 _30973_ (.A(net3936),
    .B(_08079_),
    .C(_08085_),
    .Y(_08086_));
 sg13g2_a22oi_1 _30974_ (.Y(_01337_),
    .B1(_08084_),
    .B2(_08086_),
    .A2(net3936),
    .A1(_10548_));
 sg13g2_nand2_1 _30975_ (.Y(_08087_),
    .A(net2801),
    .B(net3840));
 sg13g2_o21ai_1 _30976_ (.B1(_08081_),
    .Y(_08088_),
    .A1(_10547_),
    .A2(_10856_));
 sg13g2_xnor2_1 _30977_ (.Y(_08089_),
    .A(_11231_),
    .B(_08088_));
 sg13g2_a22oi_1 _30978_ (.Y(_08090_),
    .B1(_08089_),
    .B2(net4662),
    .A2(_08087_),
    .A1(net3725));
 sg13g2_nor2_1 _30979_ (.A(_11255_),
    .B(_08077_),
    .Y(_08091_));
 sg13g2_xnor2_1 _30980_ (.Y(_08092_),
    .A(_11231_),
    .B(_08091_));
 sg13g2_o21ai_1 _30981_ (.B1(net4380),
    .Y(_08093_),
    .A1(net3840),
    .A2(_08092_));
 sg13g2_a21oi_1 _30982_ (.A1(net4512),
    .A2(_10962_),
    .Y(_08094_),
    .B1(net3936));
 sg13g2_o21ai_1 _30983_ (.B1(_08094_),
    .Y(_08095_),
    .A1(_08090_),
    .A2(_08093_));
 sg13g2_o21ai_1 _30984_ (.B1(_08095_),
    .Y(_01338_),
    .A1(_10547_),
    .A2(net4015));
 sg13g2_a21oi_1 _30985_ (.A1(_12659_),
    .A2(_08080_),
    .Y(_08096_),
    .B1(_12661_));
 sg13g2_nand2b_1 _30986_ (.Y(_08097_),
    .B(_08096_),
    .A_N(_11243_));
 sg13g2_nand2b_1 _30987_ (.Y(_08098_),
    .B(_11243_),
    .A_N(_08096_));
 sg13g2_nand3_1 _30988_ (.B(_08097_),
    .C(_08098_),
    .A(net4663),
    .Y(_08099_));
 sg13g2_a21oi_1 _30989_ (.A1(net2077),
    .A2(net4546),
    .Y(_08100_),
    .B1(net3702));
 sg13g2_a21oi_1 _30990_ (.A1(_11230_),
    .A2(_11241_),
    .Y(_08101_),
    .B1(_11261_));
 sg13g2_or2_1 _30991_ (.X(_08102_),
    .B(_08101_),
    .A(_11243_));
 sg13g2_xnor2_1 _30992_ (.Y(_08103_),
    .A(_11243_),
    .B(_08101_));
 sg13g2_o21ai_1 _30993_ (.B1(net4015),
    .Y(_08104_),
    .A1(net4610),
    .A2(net1795));
 sg13g2_a221oi_1 _30994_ (.B2(net3692),
    .C1(_08104_),
    .B1(_08103_),
    .A1(_08099_),
    .Y(_08105_),
    .A2(_08100_));
 sg13g2_a21o_1 _30995_ (.A2(net3936),
    .A1(net2801),
    .B1(_08105_),
    .X(_01339_));
 sg13g2_nand2_1 _30996_ (.Y(_08106_),
    .A(net2077),
    .B(net3936));
 sg13g2_nand2_1 _30997_ (.Y(_08107_),
    .A(\u_inv.f_next[37] ),
    .B(net3840));
 sg13g2_o21ai_1 _30998_ (.B1(_08098_),
    .Y(_08108_),
    .A1(_10545_),
    .A2(_10854_));
 sg13g2_xnor2_1 _30999_ (.Y(_08109_),
    .A(_11242_),
    .B(_08108_));
 sg13g2_a22oi_1 _31000_ (.Y(_08110_),
    .B1(_08109_),
    .B2(net4663),
    .A2(_08107_),
    .A1(net3725));
 sg13g2_and3_1 _31001_ (.X(_08111_),
    .A(_11242_),
    .B(_11262_),
    .C(_08102_));
 sg13g2_a21oi_1 _31002_ (.A1(_11262_),
    .A2(_08102_),
    .Y(_08112_),
    .B1(_11242_));
 sg13g2_o21ai_1 _31003_ (.B1(net4380),
    .Y(_08113_),
    .A1(_08111_),
    .A2(_08112_));
 sg13g2_a21oi_1 _31004_ (.A1(net3702),
    .A2(_08113_),
    .Y(_08114_),
    .B1(_08110_));
 sg13g2_o21ai_1 _31005_ (.B1(net4015),
    .Y(_08115_),
    .A1(net4610),
    .A2(net1940));
 sg13g2_o21ai_1 _31006_ (.B1(_08106_),
    .Y(_01340_),
    .A1(_08114_),
    .A2(_08115_));
 sg13g2_o21ai_1 _31007_ (.B1(_12664_),
    .Y(_08116_),
    .A1(_12657_),
    .A2(_08096_));
 sg13g2_xnor2_1 _31008_ (.Y(_08117_),
    .A(_11250_),
    .B(_08116_));
 sg13g2_o21ai_1 _31009_ (.B1(net3714),
    .Y(_08118_),
    .A1(_10543_),
    .A2(net4662));
 sg13g2_a21oi_1 _31010_ (.A1(net4662),
    .A2(_08117_),
    .Y(_08119_),
    .B1(_08118_));
 sg13g2_o21ai_1 _31011_ (.B1(_11250_),
    .Y(_08120_),
    .A1(_11263_),
    .A2(_08112_));
 sg13g2_or3_1 _31012_ (.A(_11250_),
    .B(_11263_),
    .C(_08112_),
    .X(_08121_));
 sg13g2_and2_1 _31013_ (.A(_08120_),
    .B(_08121_),
    .X(_08122_));
 sg13g2_o21ai_1 _31014_ (.B1(net4015),
    .Y(_08123_),
    .A1(net4610),
    .A2(net1802));
 sg13g2_nor2_1 _31015_ (.A(_08119_),
    .B(_08123_),
    .Y(_08124_));
 sg13g2_o21ai_1 _31016_ (.B1(_08124_),
    .Y(_08125_),
    .A1(net3680),
    .A2(_08122_));
 sg13g2_o21ai_1 _31017_ (.B1(_08125_),
    .Y(_01341_),
    .A1(_10544_),
    .A2(net4015));
 sg13g2_nand2_1 _31018_ (.Y(_08126_),
    .A(net2513),
    .B(net3838));
 sg13g2_a21oi_1 _31019_ (.A1(_11249_),
    .A2(_08116_),
    .Y(_08127_),
    .B1(_11248_));
 sg13g2_xnor2_1 _31020_ (.Y(_08128_),
    .A(_11247_),
    .B(_08127_));
 sg13g2_a22oi_1 _31021_ (.Y(_08129_),
    .B1(_08128_),
    .B2(net4662),
    .A2(_08126_),
    .A1(net3725));
 sg13g2_o21ai_1 _31022_ (.B1(_08120_),
    .Y(_08130_),
    .A1(_10543_),
    .A2(\u_inv.f_reg[38] ));
 sg13g2_xnor2_1 _31023_ (.Y(_08131_),
    .A(_11247_),
    .B(_08130_));
 sg13g2_o21ai_1 _31024_ (.B1(net4380),
    .Y(_08132_),
    .A1(net3838),
    .A2(_08131_));
 sg13g2_a21oi_1 _31025_ (.A1(net4514),
    .A2(_10963_),
    .Y(_08133_),
    .B1(net3936));
 sg13g2_o21ai_1 _31026_ (.B1(_08133_),
    .Y(_08134_),
    .A1(_08129_),
    .A2(_08132_));
 sg13g2_o21ai_1 _31027_ (.B1(_08134_),
    .Y(_01342_),
    .A1(_10543_),
    .A2(net4015));
 sg13g2_nor2b_1 _31028_ (.A(_11277_),
    .B_N(_12736_),
    .Y(_08135_));
 sg13g2_xor2_1 _31029_ (.B(_12736_),
    .A(_11277_),
    .X(_08136_));
 sg13g2_nor2_1 _31030_ (.A(net2156),
    .B(net4663),
    .Y(_08137_));
 sg13g2_a21oi_1 _31031_ (.A1(net4669),
    .A2(_08136_),
    .Y(_08138_),
    .B1(_08137_));
 sg13g2_and2_1 _31032_ (.A(_11270_),
    .B(_11277_),
    .X(_08139_));
 sg13g2_nor2_1 _31033_ (.A(net3681),
    .B(_08139_),
    .Y(_08140_));
 sg13g2_o21ai_1 _31034_ (.B1(_08140_),
    .Y(_08141_),
    .A1(_11270_),
    .A2(_11277_));
 sg13g2_a221oi_1 _31035_ (.B2(_08138_),
    .C1(net3937),
    .B1(net3714),
    .A1(net4514),
    .Y(_08142_),
    .A2(net1993));
 sg13g2_a22oi_1 _31036_ (.Y(_01343_),
    .B1(_08141_),
    .B2(_08142_),
    .A2(net3937),
    .A1(_10542_));
 sg13g2_nand2_1 _31037_ (.Y(_08143_),
    .A(net2156),
    .B(net3937));
 sg13g2_nand2_1 _31038_ (.Y(_08144_),
    .A(net1905),
    .B(net3838));
 sg13g2_a21oi_1 _31039_ (.A1(\u_inv.f_next[40] ),
    .A2(\u_inv.f_reg[40] ),
    .Y(_08145_),
    .B1(_08135_));
 sg13g2_xnor2_1 _31040_ (.Y(_08146_),
    .A(_11278_),
    .B(_08145_));
 sg13g2_a22oi_1 _31041_ (.Y(_08147_),
    .B1(_08146_),
    .B2(net4663),
    .A2(_08144_),
    .A1(net3725));
 sg13g2_or2_1 _31042_ (.X(_08148_),
    .B(_08139_),
    .A(_11293_));
 sg13g2_and2_1 _31043_ (.A(_11278_),
    .B(_08148_),
    .X(_08149_));
 sg13g2_o21ai_1 _31044_ (.B1(net3762),
    .Y(_08150_),
    .A1(_11278_),
    .A2(_08148_));
 sg13g2_o21ai_1 _31045_ (.B1(net4380),
    .Y(_08151_),
    .A1(_08149_),
    .A2(_08150_));
 sg13g2_nor2_1 _31046_ (.A(net4611),
    .B(net1767),
    .Y(_08152_));
 sg13g2_o21ai_1 _31047_ (.B1(net4015),
    .Y(_08153_),
    .A1(_08147_),
    .A2(_08151_));
 sg13g2_o21ai_1 _31048_ (.B1(_08143_),
    .Y(_01344_),
    .A1(_08152_),
    .A2(_08153_));
 sg13g2_nand2_1 _31049_ (.Y(_08154_),
    .A(net1905),
    .B(net3937));
 sg13g2_nor3_1 _31050_ (.A(_11273_),
    .B(_11292_),
    .C(_08149_),
    .Y(_08155_));
 sg13g2_o21ai_1 _31051_ (.B1(_11273_),
    .Y(_08156_),
    .A1(_11292_),
    .A2(_08149_));
 sg13g2_nor2_1 _31052_ (.A(net3838),
    .B(_08155_),
    .Y(_08157_));
 sg13g2_a21oi_2 _31053_ (.B1(_12641_),
    .Y(_08158_),
    .A2(_08135_),
    .A1(_11279_));
 sg13g2_xnor2_1 _31054_ (.Y(_08159_),
    .A(_11273_),
    .B(_08158_));
 sg13g2_nor2_1 _31055_ (.A(\u_inv.f_next[42] ),
    .B(net4663),
    .Y(_08160_));
 sg13g2_a21oi_1 _31056_ (.A1(net4663),
    .A2(_08159_),
    .Y(_08161_),
    .B1(_08160_));
 sg13g2_a221oi_1 _31057_ (.B2(net3838),
    .C1(net4440),
    .B1(_08161_),
    .A1(_08156_),
    .Y(_08162_),
    .A2(_08157_));
 sg13g2_o21ai_1 _31058_ (.B1(net4016),
    .Y(_08163_),
    .A1(net4610),
    .A2(net1902));
 sg13g2_o21ai_1 _31059_ (.B1(_08154_),
    .Y(_01345_),
    .A1(_08162_),
    .A2(_08163_));
 sg13g2_nand2_1 _31060_ (.Y(_08164_),
    .A(net2306),
    .B(net3937));
 sg13g2_nand2_1 _31061_ (.Y(_08165_),
    .A(_11296_),
    .B(_08156_));
 sg13g2_xnor2_1 _31062_ (.Y(_08166_),
    .A(_11275_),
    .B(_08165_));
 sg13g2_o21ai_1 _31063_ (.B1(_11272_),
    .Y(_08167_),
    .A1(_11273_),
    .A2(_08158_));
 sg13g2_a21oi_1 _31064_ (.A1(_11276_),
    .A2(_08167_),
    .Y(_08168_),
    .B1(net4546));
 sg13g2_o21ai_1 _31065_ (.B1(_08168_),
    .Y(_08169_),
    .A1(_11276_),
    .A2(_08167_));
 sg13g2_o21ai_1 _31066_ (.B1(_08169_),
    .Y(_08170_),
    .A1(\u_inv.f_next[43] ),
    .A2(net4663));
 sg13g2_o21ai_1 _31067_ (.B1(net4380),
    .Y(_08171_),
    .A1(net3762),
    .A2(_08170_));
 sg13g2_a21oi_1 _31068_ (.A1(net3764),
    .A2(_08166_),
    .Y(_08172_),
    .B1(_08171_));
 sg13g2_o21ai_1 _31069_ (.B1(net4016),
    .Y(_08173_),
    .A1(net4610),
    .A2(net1860));
 sg13g2_o21ai_1 _31070_ (.B1(_08164_),
    .Y(_01346_),
    .A1(_08172_),
    .A2(_08173_));
 sg13g2_o21ai_1 _31071_ (.B1(_12649_),
    .Y(_08174_),
    .A1(_12645_),
    .A2(_08158_));
 sg13g2_nor2b_1 _31072_ (.A(_11282_),
    .B_N(_08174_),
    .Y(_08175_));
 sg13g2_xnor2_1 _31073_ (.Y(_08176_),
    .A(_11282_),
    .B(_08174_));
 sg13g2_o21ai_1 _31074_ (.B1(net3714),
    .Y(_08177_),
    .A1(_10537_),
    .A2(net4667));
 sg13g2_a21oi_1 _31075_ (.A1(net4667),
    .A2(_08176_),
    .Y(_08178_),
    .B1(_08177_));
 sg13g2_o21ai_1 _31076_ (.B1(_11299_),
    .Y(_08179_),
    .A1(_11271_),
    .A2(_11280_));
 sg13g2_xor2_1 _31077_ (.B(_08179_),
    .A(_11282_),
    .X(_08180_));
 sg13g2_o21ai_1 _31078_ (.B1(net4018),
    .Y(_08181_),
    .A1(net4611),
    .A2(net1863));
 sg13g2_nor2_1 _31079_ (.A(_08178_),
    .B(_08181_),
    .Y(_08182_));
 sg13g2_o21ai_1 _31080_ (.B1(_08182_),
    .Y(_08183_),
    .A1(net3681),
    .A2(_08180_));
 sg13g2_o21ai_1 _31081_ (.B1(_08183_),
    .Y(_01347_),
    .A1(_10538_),
    .A2(net4015));
 sg13g2_a21oi_1 _31082_ (.A1(\u_inv.f_next[44] ),
    .A2(\u_inv.f_reg[44] ),
    .Y(_08184_),
    .B1(_08175_));
 sg13g2_xnor2_1 _31083_ (.Y(_08185_),
    .A(_11281_),
    .B(_08184_));
 sg13g2_o21ai_1 _31084_ (.B1(net3714),
    .Y(_08186_),
    .A1(net2593),
    .A2(net4667));
 sg13g2_a21o_1 _31085_ (.A2(_08185_),
    .A1(net4667),
    .B1(_08186_),
    .X(_08187_));
 sg13g2_a21oi_1 _31086_ (.A1(_11282_),
    .A2(_08179_),
    .Y(_08188_),
    .B1(_11300_));
 sg13g2_inv_1 _31087_ (.Y(_08189_),
    .A(_08188_));
 sg13g2_nand2_1 _31088_ (.Y(_08190_),
    .A(_11281_),
    .B(_08189_));
 sg13g2_xnor2_1 _31089_ (.Y(_08191_),
    .A(_11281_),
    .B(_08188_));
 sg13g2_a221oi_1 _31090_ (.B2(_08191_),
    .C1(net3941),
    .B1(net3694),
    .A1(net4514),
    .Y(_08192_),
    .A2(net2015));
 sg13g2_a22oi_1 _31091_ (.Y(_01348_),
    .B1(_08187_),
    .B2(_08192_),
    .A2(net3941),
    .A1(_10537_));
 sg13g2_a21oi_1 _31092_ (.A1(_12643_),
    .A2(_08174_),
    .Y(_08193_),
    .B1(_12653_));
 sg13g2_a21oi_1 _31093_ (.A1(_11288_),
    .A2(_08193_),
    .Y(_08194_),
    .B1(net4546));
 sg13g2_o21ai_1 _31094_ (.B1(_08194_),
    .Y(_08195_),
    .A1(_11288_),
    .A2(_08193_));
 sg13g2_a21oi_1 _31095_ (.A1(net2831),
    .A2(net4547),
    .Y(_08196_),
    .B1(net3703));
 sg13g2_nand2_1 _31096_ (.Y(_08197_),
    .A(_11301_),
    .B(_08190_));
 sg13g2_xnor2_1 _31097_ (.Y(_08198_),
    .A(_11288_),
    .B(_08197_));
 sg13g2_o21ai_1 _31098_ (.B1(net4018),
    .Y(_08199_),
    .A1(net4610),
    .A2(net1978));
 sg13g2_a221oi_1 _31099_ (.B2(net3694),
    .C1(_08199_),
    .B1(_08198_),
    .A1(_08195_),
    .Y(_08200_),
    .A2(_08196_));
 sg13g2_a21o_1 _31100_ (.A2(net3941),
    .A1(net2593),
    .B1(_08200_),
    .X(_01349_));
 sg13g2_nand2_1 _31101_ (.Y(_08201_),
    .A(net3135),
    .B(net3840));
 sg13g2_o21ai_1 _31102_ (.B1(_11286_),
    .Y(_08202_),
    .A1(_11288_),
    .A2(_08193_));
 sg13g2_xnor2_1 _31103_ (.Y(_08203_),
    .A(_11284_),
    .B(_08202_));
 sg13g2_a22oi_1 _31104_ (.Y(_08204_),
    .B1(_08203_),
    .B2(net4667),
    .A2(_08201_),
    .A1(net3726));
 sg13g2_a21oi_1 _31105_ (.A1(_11288_),
    .A2(_08197_),
    .Y(_08205_),
    .B1(_11304_));
 sg13g2_xnor2_1 _31106_ (.Y(_08206_),
    .A(_11284_),
    .B(_08205_));
 sg13g2_o21ai_1 _31107_ (.B1(net4380),
    .Y(_08207_),
    .A1(net3840),
    .A2(_08206_));
 sg13g2_a21oi_1 _31108_ (.A1(net4514),
    .A2(_10964_),
    .Y(_08208_),
    .B1(net3941));
 sg13g2_o21ai_1 _31109_ (.B1(_08208_),
    .Y(_08209_),
    .A1(_08204_),
    .A2(_08207_));
 sg13g2_o21ai_1 _31110_ (.B1(_08209_),
    .Y(_01350_),
    .A1(_10535_),
    .A2(net4018));
 sg13g2_or2_1 _31111_ (.X(_08210_),
    .B(_12738_),
    .A(_11323_));
 sg13g2_a21oi_1 _31112_ (.A1(_11323_),
    .A2(_12738_),
    .Y(_08211_),
    .B1(net4546));
 sg13g2_nand2_1 _31113_ (.Y(_08212_),
    .A(_08210_),
    .B(_08211_));
 sg13g2_a21oi_1 _31114_ (.A1(net2485),
    .A2(net4546),
    .Y(_08213_),
    .B1(net3703));
 sg13g2_xnor2_1 _31115_ (.Y(_08214_),
    .A(_11308_),
    .B(_11323_));
 sg13g2_o21ai_1 _31116_ (.B1(net4018),
    .Y(_08215_),
    .A1(net4611),
    .A2(net1803));
 sg13g2_a221oi_1 _31117_ (.B2(net3694),
    .C1(_08215_),
    .B1(_08214_),
    .A1(_08212_),
    .Y(_08216_),
    .A2(_08213_));
 sg13g2_a21o_1 _31118_ (.A2(net3941),
    .A1(net3135),
    .B1(_08216_),
    .X(_01351_));
 sg13g2_nand2_1 _31119_ (.Y(_08217_),
    .A(net3015),
    .B(net3839));
 sg13g2_o21ai_1 _31120_ (.B1(_08210_),
    .Y(_08218_),
    .A1(_10533_),
    .A2(_10842_));
 sg13g2_xor2_1 _31121_ (.B(_08218_),
    .A(_11333_),
    .X(_08219_));
 sg13g2_a22oi_1 _31122_ (.Y(_08220_),
    .B1(_08219_),
    .B2(net4667),
    .A2(_08217_),
    .A1(net3725));
 sg13g2_a21o_1 _31123_ (.A2(_11323_),
    .A1(_11308_),
    .B1(_11342_),
    .X(_08221_));
 sg13g2_and2_1 _31124_ (.A(_11333_),
    .B(_08221_),
    .X(_08222_));
 sg13g2_o21ai_1 _31125_ (.B1(net3764),
    .Y(_08223_),
    .A1(_11333_),
    .A2(_08221_));
 sg13g2_o21ai_1 _31126_ (.B1(net4380),
    .Y(_08224_),
    .A1(_08222_),
    .A2(_08223_));
 sg13g2_a21oi_1 _31127_ (.A1(net4514),
    .A2(_10965_),
    .Y(_08225_),
    .B1(net3947));
 sg13g2_o21ai_1 _31128_ (.B1(_08225_),
    .Y(_08226_),
    .A1(_08220_),
    .A2(_08224_));
 sg13g2_o21ai_1 _31129_ (.B1(_08226_),
    .Y(_01352_),
    .A1(_10533_),
    .A2(net4017));
 sg13g2_or2_1 _31130_ (.X(_08227_),
    .B(_08222_),
    .A(_11344_));
 sg13g2_nor2_1 _31131_ (.A(_11331_),
    .B(_08227_),
    .Y(_08228_));
 sg13g2_and2_1 _31132_ (.A(_11331_),
    .B(_08227_),
    .X(_08229_));
 sg13g2_nor3_1 _31133_ (.A(net3681),
    .B(_08228_),
    .C(_08229_),
    .Y(_08230_));
 sg13g2_a21oi_1 _31134_ (.A1(_12616_),
    .A2(_08210_),
    .Y(_08231_),
    .B1(_11332_));
 sg13g2_nor2b_1 _31135_ (.A(_11331_),
    .B_N(_08231_),
    .Y(_08232_));
 sg13g2_xor2_1 _31136_ (.B(_08231_),
    .A(_11331_),
    .X(_08233_));
 sg13g2_o21ai_1 _31137_ (.B1(net3714),
    .Y(_08234_),
    .A1(net2234),
    .A2(net4667));
 sg13g2_a21oi_1 _31138_ (.A1(net4667),
    .A2(_08233_),
    .Y(_08235_),
    .B1(_08234_));
 sg13g2_nor2b_1 _31139_ (.A(net4614),
    .B_N(net1779),
    .Y(_08236_));
 sg13g2_nor4_1 _31140_ (.A(net3947),
    .B(_08230_),
    .C(_08235_),
    .D(_08236_),
    .Y(_08237_));
 sg13g2_a21oi_1 _31141_ (.A1(_10532_),
    .A2(net3941),
    .Y(_01353_),
    .B1(_08237_));
 sg13g2_nand2_1 _31142_ (.Y(_08238_),
    .A(net2234),
    .B(net3947));
 sg13g2_nor3_1 _31143_ (.A(_11330_),
    .B(_11343_),
    .C(_08229_),
    .Y(_08239_));
 sg13g2_o21ai_1 _31144_ (.B1(_11330_),
    .Y(_08240_),
    .A1(_11343_),
    .A2(_08229_));
 sg13g2_nor2_1 _31145_ (.A(net3839),
    .B(_08239_),
    .Y(_08241_));
 sg13g2_a21oi_1 _31146_ (.A1(\u_inv.f_next[50] ),
    .A2(\u_inv.f_reg[50] ),
    .Y(_08242_),
    .B1(_08232_));
 sg13g2_xnor2_1 _31147_ (.Y(_08243_),
    .A(_11330_),
    .B(_08242_));
 sg13g2_nor2_1 _31148_ (.A(\u_inv.f_next[51] ),
    .B(net4668),
    .Y(_08244_));
 sg13g2_a21oi_1 _31149_ (.A1(net4668),
    .A2(_08243_),
    .Y(_08245_),
    .B1(_08244_));
 sg13g2_a221oi_1 _31150_ (.B2(net3839),
    .C1(net4440),
    .B1(_08245_),
    .A1(_08240_),
    .Y(_08246_),
    .A2(_08241_));
 sg13g2_o21ai_1 _31151_ (.B1(net4021),
    .Y(_08247_),
    .A1(net4614),
    .A2(net1838));
 sg13g2_o21ai_1 _31152_ (.B1(_08238_),
    .Y(_01354_),
    .A1(_08246_),
    .A2(_08247_));
 sg13g2_a21oi_1 _31153_ (.A1(_12615_),
    .A2(_08231_),
    .Y(_08248_),
    .B1(_12619_));
 sg13g2_nor2b_1 _31154_ (.A(_11327_),
    .B_N(_08248_),
    .Y(_08249_));
 sg13g2_nand2b_1 _31155_ (.Y(_08250_),
    .B(_11327_),
    .A_N(_08248_));
 sg13g2_nand3b_1 _31156_ (.B(_08250_),
    .C(net4668),
    .Y(_08251_),
    .A_N(_08249_));
 sg13g2_a21oi_1 _31157_ (.A1(net2402),
    .A2(net4546),
    .Y(_08252_),
    .B1(net3703));
 sg13g2_a21oi_1 _31158_ (.A1(_11308_),
    .A2(_11334_),
    .Y(_08253_),
    .B1(_11348_));
 sg13g2_or2_1 _31159_ (.X(_08254_),
    .B(_08253_),
    .A(_11327_));
 sg13g2_xnor2_1 _31160_ (.Y(_08255_),
    .A(_11327_),
    .B(_08253_));
 sg13g2_o21ai_1 _31161_ (.B1(net4021),
    .Y(_08256_),
    .A1(net4614),
    .A2(net1872));
 sg13g2_a221oi_1 _31162_ (.B2(net3694),
    .C1(_08256_),
    .B1(_08255_),
    .A1(_08251_),
    .Y(_08257_),
    .A2(_08252_));
 sg13g2_a21o_1 _31163_ (.A2(net3941),
    .A1(net2702),
    .B1(_08257_),
    .X(_01355_));
 sg13g2_nand2_1 _31164_ (.Y(_08258_),
    .A(net2402),
    .B(net3942));
 sg13g2_nand2_1 _31165_ (.Y(_08259_),
    .A(\u_inv.f_next[53] ),
    .B(net3840));
 sg13g2_o21ai_1 _31166_ (.B1(_08250_),
    .Y(_08260_),
    .A1(_10529_),
    .A2(_10838_));
 sg13g2_xnor2_1 _31167_ (.Y(_08261_),
    .A(_11328_),
    .B(_08260_));
 sg13g2_a22oi_1 _31168_ (.Y(_08262_),
    .B1(_08261_),
    .B2(net4668),
    .A2(_08259_),
    .A1(net3725));
 sg13g2_a21oi_1 _31169_ (.A1(_11340_),
    .A2(_08254_),
    .Y(_08263_),
    .B1(_11328_));
 sg13g2_and3_1 _31170_ (.X(_08264_),
    .A(_11328_),
    .B(_11340_),
    .C(_08254_));
 sg13g2_o21ai_1 _31171_ (.B1(net4380),
    .Y(_08265_),
    .A1(_08263_),
    .A2(_08264_));
 sg13g2_a21oi_1 _31172_ (.A1(net3703),
    .A2(_08265_),
    .Y(_08266_),
    .B1(_08262_));
 sg13g2_o21ai_1 _31173_ (.B1(net4017),
    .Y(_08267_),
    .A1(net4614),
    .A2(net2304));
 sg13g2_o21ai_1 _31174_ (.B1(_08258_),
    .Y(_01356_),
    .A1(_08266_),
    .A2(_08267_));
 sg13g2_o21ai_1 _31175_ (.B1(_11325_),
    .Y(_08268_),
    .A1(_11339_),
    .A2(_08263_));
 sg13g2_or3_1 _31176_ (.A(_11325_),
    .B(_11339_),
    .C(_08263_),
    .X(_08269_));
 sg13g2_nand2_1 _31177_ (.Y(_08270_),
    .A(_08268_),
    .B(_08269_));
 sg13g2_o21ai_1 _31178_ (.B1(_12623_),
    .Y(_08271_),
    .A1(_12613_),
    .A2(_08248_));
 sg13g2_nor2b_1 _31179_ (.A(_11325_),
    .B_N(_08271_),
    .Y(_08272_));
 sg13g2_nand2b_1 _31180_ (.Y(_08273_),
    .B(_11325_),
    .A_N(_08271_));
 sg13g2_nand3b_1 _31181_ (.B(_08273_),
    .C(net4673),
    .Y(_08274_),
    .A_N(_08272_));
 sg13g2_a21oi_1 _31182_ (.A1(\u_inv.f_next[54] ),
    .A2(net4555),
    .Y(_08275_),
    .B1(net3703));
 sg13g2_o21ai_1 _31183_ (.B1(net4021),
    .Y(_08276_),
    .A1(net4614),
    .A2(net1780));
 sg13g2_a221oi_1 _31184_ (.B2(_08275_),
    .C1(_08276_),
    .B1(_08274_),
    .A1(net3694),
    .Y(_08277_),
    .A2(_08270_));
 sg13g2_a21o_1 _31185_ (.A2(net3941),
    .A1(net2857),
    .B1(_08277_),
    .X(_01357_));
 sg13g2_nand2_1 _31186_ (.Y(_08278_),
    .A(net2313),
    .B(net3844));
 sg13g2_a21oi_1 _31187_ (.A1(\u_inv.f_next[54] ),
    .A2(\u_inv.f_reg[54] ),
    .Y(_08279_),
    .B1(_08272_));
 sg13g2_xnor2_1 _31188_ (.Y(_08280_),
    .A(_11324_),
    .B(_08279_));
 sg13g2_a22oi_1 _31189_ (.Y(_08281_),
    .B1(_08280_),
    .B2(net4673),
    .A2(_08278_),
    .A1(net3727));
 sg13g2_o21ai_1 _31190_ (.B1(_08268_),
    .Y(_08282_),
    .A1(_10527_),
    .A2(\u_inv.f_reg[54] ));
 sg13g2_xnor2_1 _31191_ (.Y(_08283_),
    .A(_11324_),
    .B(_08282_));
 sg13g2_o21ai_1 _31192_ (.B1(net4382),
    .Y(_08284_),
    .A1(net3844),
    .A2(_08283_));
 sg13g2_a21oi_1 _31193_ (.A1(net4513),
    .A2(_10966_),
    .Y(_08285_),
    .B1(net3947));
 sg13g2_o21ai_1 _31194_ (.B1(_08285_),
    .Y(_08286_),
    .A1(_08281_),
    .A2(_08284_));
 sg13g2_o21ai_1 _31195_ (.B1(_08286_),
    .Y(_01358_),
    .A1(_10527_),
    .A2(net4021));
 sg13g2_a21o_2 _31196_ (.A2(_08271_),
    .A1(_12612_),
    .B1(_12625_),
    .X(_08287_));
 sg13g2_nand2_1 _31197_ (.Y(_08288_),
    .A(_11321_),
    .B(_08287_));
 sg13g2_nor2_1 _31198_ (.A(_10525_),
    .B(net4673),
    .Y(_08289_));
 sg13g2_o21ai_1 _31199_ (.B1(net4673),
    .Y(_08290_),
    .A1(_11321_),
    .A2(_08287_));
 sg13g2_nor2b_1 _31200_ (.A(_08290_),
    .B_N(_08288_),
    .Y(_08291_));
 sg13g2_o21ai_1 _31201_ (.B1(net3714),
    .Y(_08292_),
    .A1(_08289_),
    .A2(_08291_));
 sg13g2_a21oi_1 _31202_ (.A1(_11308_),
    .A2(_11335_),
    .Y(_08293_),
    .B1(_11352_));
 sg13g2_or2_1 _31203_ (.X(_08294_),
    .B(_08293_),
    .A(_11321_));
 sg13g2_a21oi_1 _31204_ (.A1(_11321_),
    .A2(_08293_),
    .Y(_08295_),
    .B1(net3682));
 sg13g2_a221oi_1 _31205_ (.B2(_08295_),
    .C1(net3948),
    .B1(_08294_),
    .A1(net4513),
    .Y(_08296_),
    .A2(net2184));
 sg13g2_a22oi_1 _31206_ (.Y(_01359_),
    .B1(_08292_),
    .B2(_08296_),
    .A2(net3947),
    .A1(_10526_));
 sg13g2_o21ai_1 _31207_ (.B1(_08288_),
    .Y(_08297_),
    .A1(_10525_),
    .A2(_10834_));
 sg13g2_a21oi_1 _31208_ (.A1(_11317_),
    .A2(_08297_),
    .Y(_08298_),
    .B1(net4555));
 sg13g2_o21ai_1 _31209_ (.B1(_08298_),
    .Y(_08299_),
    .A1(_11317_),
    .A2(_08297_));
 sg13g2_a21oi_1 _31210_ (.A1(\u_inv.f_next[57] ),
    .A2(net4555),
    .Y(_08300_),
    .B1(net3703));
 sg13g2_nand2_1 _31211_ (.Y(_08301_),
    .A(_11362_),
    .B(_08294_));
 sg13g2_nand2b_1 _31212_ (.Y(_08302_),
    .B(_08301_),
    .A_N(_11317_));
 sg13g2_xor2_1 _31213_ (.B(_08301_),
    .A(_11317_),
    .X(_08303_));
 sg13g2_o21ai_1 _31214_ (.B1(net4022),
    .Y(_08304_),
    .A1(net4613),
    .A2(net2104));
 sg13g2_a221oi_1 _31215_ (.B2(net3693),
    .C1(_08304_),
    .B1(_08303_),
    .A1(_08299_),
    .Y(_08305_),
    .A2(_08300_));
 sg13g2_a21o_1 _31216_ (.A2(net3947),
    .A1(net2689),
    .B1(_08305_),
    .X(_01360_));
 sg13g2_a21oi_1 _31217_ (.A1(_12627_),
    .A2(_08287_),
    .Y(_08306_),
    .B1(_12608_));
 sg13g2_xnor2_1 _31218_ (.Y(_08307_),
    .A(_11316_),
    .B(_08306_));
 sg13g2_o21ai_1 _31219_ (.B1(net3843),
    .Y(_08308_),
    .A1(net3248),
    .A2(net4673));
 sg13g2_a21oi_1 _31220_ (.A1(net4673),
    .A2(_08307_),
    .Y(_08309_),
    .B1(_08308_));
 sg13g2_nand2_1 _31221_ (.Y(_08310_),
    .A(_11361_),
    .B(_08302_));
 sg13g2_xnor2_1 _31222_ (.Y(_08311_),
    .A(_11316_),
    .B(_08310_));
 sg13g2_o21ai_1 _31223_ (.B1(net4381),
    .Y(_08312_),
    .A1(net3843),
    .A2(_08311_));
 sg13g2_a21oi_1 _31224_ (.A1(net4513),
    .A2(_10967_),
    .Y(_08313_),
    .B1(net3948));
 sg13g2_o21ai_1 _31225_ (.B1(_08313_),
    .Y(_08314_),
    .A1(_08309_),
    .A2(_08312_));
 sg13g2_o21ai_1 _31226_ (.B1(_08314_),
    .Y(_01361_),
    .A1(_10524_),
    .A2(net4021));
 sg13g2_nand2_1 _31227_ (.Y(_08315_),
    .A(net2655),
    .B(net3843));
 sg13g2_o21ai_1 _31228_ (.B1(_11315_),
    .Y(_08316_),
    .A1(_11316_),
    .A2(_08306_));
 sg13g2_xor2_1 _31229_ (.B(_08316_),
    .A(_11318_),
    .X(_08317_));
 sg13g2_a22oi_1 _31230_ (.Y(_08318_),
    .B1(_08317_),
    .B2(net4673),
    .A2(_08315_),
    .A1(net3727));
 sg13g2_a21oi_1 _31231_ (.A1(_11316_),
    .A2(_08310_),
    .Y(_08319_),
    .B1(_11360_));
 sg13g2_xor2_1 _31232_ (.B(_08319_),
    .A(_11318_),
    .X(_08320_));
 sg13g2_o21ai_1 _31233_ (.B1(net4381),
    .Y(_08321_),
    .A1(net3844),
    .A2(_08320_));
 sg13g2_a21oi_1 _31234_ (.A1(net4513),
    .A2(_10968_),
    .Y(_08322_),
    .B1(net3948));
 sg13g2_o21ai_1 _31235_ (.B1(_08322_),
    .Y(_08323_),
    .A1(_08318_),
    .A2(_08321_));
 sg13g2_o21ai_1 _31236_ (.B1(_08323_),
    .Y(_01362_),
    .A1(_10523_),
    .A2(net4021));
 sg13g2_nand2b_1 _31237_ (.Y(_08324_),
    .B(_12606_),
    .A_N(_08306_));
 sg13g2_nand2b_1 _31238_ (.Y(_08325_),
    .B(_08324_),
    .A_N(_12610_));
 sg13g2_nand2b_1 _31239_ (.Y(_08326_),
    .B(_11313_),
    .A_N(_08325_));
 sg13g2_nor2b_1 _31240_ (.A(_11313_),
    .B_N(_08325_),
    .Y(_08327_));
 sg13g2_nand3b_1 _31241_ (.B(net4673),
    .C(_08326_),
    .Y(_08328_),
    .A_N(_08327_));
 sg13g2_a21oi_1 _31242_ (.A1(\u_inv.f_next[60] ),
    .A2(net4555),
    .Y(_08329_),
    .B1(net3703));
 sg13g2_o21ai_1 _31243_ (.B1(_11364_),
    .Y(_08330_),
    .A1(_11320_),
    .A2(_08294_));
 sg13g2_xnor2_1 _31244_ (.Y(_08331_),
    .A(_11313_),
    .B(_08330_));
 sg13g2_o21ai_1 _31245_ (.B1(net4021),
    .Y(_08332_),
    .A1(net4614),
    .A2(net2046));
 sg13g2_a221oi_1 _31246_ (.B2(net3693),
    .C1(_08332_),
    .B1(_08331_),
    .A1(_08328_),
    .Y(_08333_),
    .A2(_08329_));
 sg13g2_a21o_1 _31247_ (.A2(net3947),
    .A1(net2655),
    .B1(_08333_),
    .X(_01363_));
 sg13g2_a21oi_1 _31248_ (.A1(\u_inv.f_next[60] ),
    .A2(\u_inv.f_reg[60] ),
    .Y(_08334_),
    .B1(_08327_));
 sg13g2_xnor2_1 _31249_ (.Y(_08335_),
    .A(_11312_),
    .B(_08334_));
 sg13g2_o21ai_1 _31250_ (.B1(net3716),
    .Y(_08336_),
    .A1(net2717),
    .A2(net4674));
 sg13g2_a21oi_1 _31251_ (.A1(net4674),
    .A2(_08335_),
    .Y(_08337_),
    .B1(_08336_));
 sg13g2_a21o_1 _31252_ (.A2(_08330_),
    .A1(_11313_),
    .B1(_11354_),
    .X(_08338_));
 sg13g2_and2_1 _31253_ (.A(_11312_),
    .B(_08338_),
    .X(_08339_));
 sg13g2_o21ai_1 _31254_ (.B1(net3693),
    .Y(_08340_),
    .A1(_11312_),
    .A2(_08338_));
 sg13g2_a21oi_1 _31255_ (.A1(net4513),
    .A2(net1919),
    .Y(_08341_),
    .B1(net3950));
 sg13g2_o21ai_1 _31256_ (.B1(_08341_),
    .Y(_08342_),
    .A1(_08339_),
    .A2(_08340_));
 sg13g2_nor2_1 _31257_ (.A(_08337_),
    .B(_08342_),
    .Y(_08343_));
 sg13g2_a21oi_1 _31258_ (.A1(_10521_),
    .A2(net3948),
    .Y(_01364_),
    .B1(_08343_));
 sg13g2_a21oi_1 _31259_ (.A1(_12604_),
    .A2(_08325_),
    .Y(_08344_),
    .B1(_12637_));
 sg13g2_nand2b_1 _31260_ (.Y(_08345_),
    .B(_11310_),
    .A_N(_08344_));
 sg13g2_nand2b_1 _31261_ (.Y(_08346_),
    .B(_08344_),
    .A_N(_11310_));
 sg13g2_nand3_1 _31262_ (.B(_08345_),
    .C(_08346_),
    .A(net4674),
    .Y(_08347_));
 sg13g2_a21oi_1 _31263_ (.A1(net1969),
    .A2(net4555),
    .Y(_08348_),
    .B1(net3704));
 sg13g2_nor2_1 _31264_ (.A(_11353_),
    .B(_08339_),
    .Y(_08349_));
 sg13g2_xnor2_1 _31265_ (.Y(_08350_),
    .A(_11310_),
    .B(_08349_));
 sg13g2_o21ai_1 _31266_ (.B1(net4021),
    .Y(_08351_),
    .A1(net4615),
    .A2(net1764));
 sg13g2_a221oi_1 _31267_ (.B2(net3693),
    .C1(_08351_),
    .B1(_08350_),
    .A1(_08347_),
    .Y(_08352_),
    .A2(_08348_));
 sg13g2_a21o_1 _31268_ (.A2(net3948),
    .A1(net2717),
    .B1(_08352_),
    .X(_01365_));
 sg13g2_nand2_1 _31269_ (.Y(_08353_),
    .A(net1969),
    .B(net3948));
 sg13g2_nand2_1 _31270_ (.Y(_08354_),
    .A(\u_inv.f_next[63] ),
    .B(net3844));
 sg13g2_o21ai_1 _31271_ (.B1(_08345_),
    .Y(_08355_),
    .A1(_10519_),
    .A2(_10828_));
 sg13g2_xnor2_1 _31272_ (.Y(_08356_),
    .A(_11309_),
    .B(_08355_));
 sg13g2_a22oi_1 _31273_ (.Y(_08357_),
    .B1(_08356_),
    .B2(net4674),
    .A2(_08354_),
    .A1(net3727));
 sg13g2_o21ai_1 _31274_ (.B1(_11356_),
    .Y(_08358_),
    .A1(_11310_),
    .A2(_08349_));
 sg13g2_xor2_1 _31275_ (.B(_08358_),
    .A(_11309_),
    .X(_08359_));
 sg13g2_o21ai_1 _31276_ (.B1(net4381),
    .Y(_08360_),
    .A1(net3844),
    .A2(_08359_));
 sg13g2_nor2_1 _31277_ (.A(net4616),
    .B(\u_inv.input_reg[62] ),
    .Y(_08361_));
 sg13g2_o21ai_1 _31278_ (.B1(net4022),
    .Y(_08362_),
    .A1(_08357_),
    .A2(_08360_));
 sg13g2_o21ai_1 _31279_ (.B1(_08353_),
    .Y(_01366_),
    .A1(_08361_),
    .A2(_08362_));
 sg13g2_nand3_1 _31280_ (.B(_11366_),
    .C(_11392_),
    .A(_11337_),
    .Y(_08363_));
 sg13g2_a21oi_1 _31281_ (.A1(_11337_),
    .A2(_11366_),
    .Y(_08364_),
    .B1(_11392_));
 sg13g2_nand3b_1 _31282_ (.B(net3693),
    .C(_08363_),
    .Y(_08365_),
    .A_N(_08364_));
 sg13g2_nand2_1 _31283_ (.Y(_08366_),
    .A(_11392_),
    .B(_12741_));
 sg13g2_xnor2_1 _31284_ (.Y(_08367_),
    .A(_11392_),
    .B(_12741_));
 sg13g2_nor2_1 _31285_ (.A(net2147),
    .B(net4676),
    .Y(_08368_));
 sg13g2_a21oi_1 _31286_ (.A1(net4676),
    .A2(_08367_),
    .Y(_08369_),
    .B1(_08368_));
 sg13g2_a221oi_1 _31287_ (.B2(_08369_),
    .C1(net3947),
    .B1(net3716),
    .A1(net4513),
    .Y(_08370_),
    .A2(net2114));
 sg13g2_a22oi_1 _31288_ (.Y(_01367_),
    .B1(_08365_),
    .B2(_08370_),
    .A2(net3948),
    .A1(_10518_));
 sg13g2_nand2_1 _31289_ (.Y(_08371_),
    .A(net2147),
    .B(net3950));
 sg13g2_nand2_1 _31290_ (.Y(_08372_),
    .A(net2051),
    .B(net3845));
 sg13g2_nand2_1 _31291_ (.Y(_08373_),
    .A(_11391_),
    .B(_08366_));
 sg13g2_xnor2_1 _31292_ (.Y(_08374_),
    .A(_11390_),
    .B(_08373_));
 sg13g2_a22oi_1 _31293_ (.Y(_08375_),
    .B1(_08374_),
    .B2(net4676),
    .A2(_08372_),
    .A1(net3727));
 sg13g2_a21oi_1 _31294_ (.A1(\u_inv.f_next[64] ),
    .A2(_10826_),
    .Y(_08376_),
    .B1(_08364_));
 sg13g2_nor2_1 _31295_ (.A(_11390_),
    .B(_08376_),
    .Y(_08377_));
 sg13g2_a21oi_1 _31296_ (.A1(_11390_),
    .A2(_08376_),
    .Y(_08378_),
    .B1(net3845));
 sg13g2_nor2b_1 _31297_ (.A(_08377_),
    .B_N(_08378_),
    .Y(_08379_));
 sg13g2_nor3_1 _31298_ (.A(net4442),
    .B(_08375_),
    .C(_08379_),
    .Y(_08380_));
 sg13g2_o21ai_1 _31299_ (.B1(net4023),
    .Y(_08381_),
    .A1(net4615),
    .A2(net1798));
 sg13g2_o21ai_1 _31300_ (.B1(_08371_),
    .Y(_01368_),
    .A1(_08380_),
    .A2(_08381_));
 sg13g2_nand2_1 _31301_ (.Y(_08382_),
    .A(net2051),
    .B(net3950));
 sg13g2_nand2b_1 _31302_ (.Y(_08383_),
    .B(_08373_),
    .A_N(_11388_));
 sg13g2_nand2_1 _31303_ (.Y(_08384_),
    .A(_11389_),
    .B(_08383_));
 sg13g2_xnor2_1 _31304_ (.Y(_08385_),
    .A(_11387_),
    .B(_08384_));
 sg13g2_o21ai_1 _31305_ (.B1(net3845),
    .Y(_08386_),
    .A1(\u_inv.f_next[66] ),
    .A2(net4676));
 sg13g2_a21oi_1 _31306_ (.A1(net4676),
    .A2(_08385_),
    .Y(_08387_),
    .B1(_08386_));
 sg13g2_a21oi_1 _31307_ (.A1(\u_inv.f_next[65] ),
    .A2(_10825_),
    .Y(_08388_),
    .B1(_08377_));
 sg13g2_nor2_1 _31308_ (.A(_11387_),
    .B(_08388_),
    .Y(_08389_));
 sg13g2_a21oi_1 _31309_ (.A1(_11387_),
    .A2(_08388_),
    .Y(_08390_),
    .B1(net3845));
 sg13g2_nor2b_1 _31310_ (.A(_08389_),
    .B_N(_08390_),
    .Y(_08391_));
 sg13g2_nor3_1 _31311_ (.A(net4442),
    .B(_08387_),
    .C(_08391_),
    .Y(_08392_));
 sg13g2_o21ai_1 _31312_ (.B1(net4023),
    .Y(_08393_),
    .A1(net4615),
    .A2(net1741));
 sg13g2_o21ai_1 _31313_ (.B1(_08382_),
    .Y(_01369_),
    .A1(_08392_),
    .A2(_08393_));
 sg13g2_a21oi_1 _31314_ (.A1(_11387_),
    .A2(_08384_),
    .Y(_08394_),
    .B1(_11386_));
 sg13g2_xor2_1 _31315_ (.B(_08394_),
    .A(_11385_),
    .X(_08395_));
 sg13g2_nand2_1 _31316_ (.Y(_08396_),
    .A(net2349),
    .B(net3845));
 sg13g2_a22oi_1 _31317_ (.Y(_08397_),
    .B1(_08396_),
    .B2(net3728),
    .A2(_08395_),
    .A1(net4677));
 sg13g2_nor2_1 _31318_ (.A(_11417_),
    .B(_08389_),
    .Y(_08398_));
 sg13g2_xnor2_1 _31319_ (.Y(_08399_),
    .A(_11385_),
    .B(_08398_));
 sg13g2_o21ai_1 _31320_ (.B1(net4381),
    .Y(_08400_),
    .A1(net3846),
    .A2(_08399_));
 sg13g2_a21oi_1 _31321_ (.A1(net4515),
    .A2(_10969_),
    .Y(_08401_),
    .B1(net3950));
 sg13g2_o21ai_1 _31322_ (.B1(_08401_),
    .Y(_08402_),
    .A1(_08397_),
    .A2(_08400_));
 sg13g2_o21ai_1 _31323_ (.B1(_08402_),
    .Y(_01370_),
    .A1(_10515_),
    .A2(net4024));
 sg13g2_o21ai_1 _31324_ (.B1(_12577_),
    .Y(_08403_),
    .A1(_12742_),
    .A2(_08366_));
 sg13g2_a21oi_1 _31325_ (.A1(_11400_),
    .A2(_08403_),
    .Y(_08404_),
    .B1(net4556));
 sg13g2_o21ai_1 _31326_ (.B1(_08404_),
    .Y(_08405_),
    .A1(_11400_),
    .A2(_08403_));
 sg13g2_a21oi_1 _31327_ (.A1(net2060),
    .A2(net4556),
    .Y(_08406_),
    .B1(net3704));
 sg13g2_a21oi_1 _31328_ (.A1(_11367_),
    .A2(_11393_),
    .Y(_08407_),
    .B1(_11422_));
 sg13g2_or2_1 _31329_ (.X(_08408_),
    .B(_08407_),
    .A(_11400_));
 sg13g2_xnor2_1 _31330_ (.Y(_08409_),
    .A(_11400_),
    .B(_08407_));
 sg13g2_o21ai_1 _31331_ (.B1(net4024),
    .Y(_08410_),
    .A1(net4615),
    .A2(net2042));
 sg13g2_a221oi_1 _31332_ (.B2(net3693),
    .C1(_08410_),
    .B1(_08409_),
    .A1(_08405_),
    .Y(_08411_),
    .A2(_08406_));
 sg13g2_a21o_1 _31333_ (.A2(net3951),
    .A1(net2349),
    .B1(_08411_),
    .X(_01371_));
 sg13g2_nand2_1 _31334_ (.Y(_08412_),
    .A(net2060),
    .B(net3959));
 sg13g2_a21oi_1 _31335_ (.A1(_10512_),
    .A2(net4555),
    .Y(_08413_),
    .B1(net3774));
 sg13g2_a21oi_1 _31336_ (.A1(_11400_),
    .A2(_08403_),
    .Y(_08414_),
    .B1(_11399_));
 sg13g2_a21oi_1 _31337_ (.A1(_11398_),
    .A2(_08414_),
    .Y(_08415_),
    .B1(net4556));
 sg13g2_o21ai_1 _31338_ (.B1(_08415_),
    .Y(_08416_),
    .A1(_11398_),
    .A2(_08414_));
 sg13g2_a21oi_1 _31339_ (.A1(_11423_),
    .A2(_08408_),
    .Y(_08417_),
    .B1(_11398_));
 sg13g2_nand3_1 _31340_ (.B(_11423_),
    .C(_08408_),
    .A(_11398_),
    .Y(_08418_));
 sg13g2_nor2b_1 _31341_ (.A(_08417_),
    .B_N(_08418_),
    .Y(_08419_));
 sg13g2_a221oi_1 _31342_ (.B2(net3774),
    .C1(net4443),
    .B1(_08419_),
    .A1(_08413_),
    .Y(_08420_),
    .A2(_08416_));
 sg13g2_o21ai_1 _31343_ (.B1(net4024),
    .Y(_08421_),
    .A1(net4618),
    .A2(net1983));
 sg13g2_o21ai_1 _31344_ (.B1(_08412_),
    .Y(_01372_),
    .A1(_08420_),
    .A2(_08421_));
 sg13g2_nor2_1 _31345_ (.A(_11424_),
    .B(_08417_),
    .Y(_08422_));
 sg13g2_o21ai_1 _31346_ (.B1(_11397_),
    .Y(_08423_),
    .A1(_11424_),
    .A2(_08417_));
 sg13g2_xnor2_1 _31347_ (.Y(_08424_),
    .A(_11397_),
    .B(_08422_));
 sg13g2_o21ai_1 _31348_ (.B1(net4023),
    .Y(_08425_),
    .A1(net4618),
    .A2(net2118));
 sg13g2_a21oi_1 _31349_ (.A1(_12571_),
    .A2(_08403_),
    .Y(_08426_),
    .B1(_12580_));
 sg13g2_xor2_1 _31350_ (.B(_08426_),
    .A(_11397_),
    .X(_08427_));
 sg13g2_o21ai_1 _31351_ (.B1(net3716),
    .Y(_08428_),
    .A1(_10511_),
    .A2(net4676));
 sg13g2_a21oi_1 _31352_ (.A1(net4677),
    .A2(_08427_),
    .Y(_08429_),
    .B1(_08428_));
 sg13g2_nor2_1 _31353_ (.A(_08425_),
    .B(_08429_),
    .Y(_08430_));
 sg13g2_o21ai_1 _31354_ (.B1(_08430_),
    .Y(_08431_),
    .A1(net3682),
    .A2(_08424_));
 sg13g2_o21ai_1 _31355_ (.B1(_08431_),
    .Y(_01373_),
    .A1(_10512_),
    .A2(net4023));
 sg13g2_nand2_1 _31356_ (.Y(_08432_),
    .A(net1539),
    .B(net3951));
 sg13g2_nand2b_1 _31357_ (.Y(_08433_),
    .B(_08423_),
    .A_N(_11428_));
 sg13g2_xnor2_1 _31358_ (.Y(_08434_),
    .A(_11394_),
    .B(_08433_));
 sg13g2_a21oi_1 _31359_ (.A1(_10510_),
    .A2(net4556),
    .Y(_08435_),
    .B1(net3774));
 sg13g2_o21ai_1 _31360_ (.B1(_11396_),
    .Y(_08436_),
    .A1(_11397_),
    .A2(_08426_));
 sg13g2_a21oi_1 _31361_ (.A1(_11395_),
    .A2(_08436_),
    .Y(_08437_),
    .B1(net4556));
 sg13g2_o21ai_1 _31362_ (.B1(_08437_),
    .Y(_08438_),
    .A1(_11395_),
    .A2(_08436_));
 sg13g2_a221oi_1 _31363_ (.B2(_08438_),
    .C1(net4443),
    .B1(_08435_),
    .A1(net3774),
    .Y(_08439_),
    .A2(_08434_));
 sg13g2_o21ai_1 _31364_ (.B1(net4023),
    .Y(_08440_),
    .A1(net4615),
    .A2(\u_inv.input_reg[70] ));
 sg13g2_o21ai_1 _31365_ (.B1(_08432_),
    .Y(_01374_),
    .A1(_08439_),
    .A2(_08440_));
 sg13g2_and3_1 _31366_ (.X(_08441_),
    .A(_11392_),
    .B(_12741_),
    .C(_12743_));
 sg13g2_nor2_1 _31367_ (.A(_12582_),
    .B(_08441_),
    .Y(_08442_));
 sg13g2_nand2b_1 _31368_ (.Y(_08443_),
    .B(_08442_),
    .A_N(_11372_));
 sg13g2_nor2b_1 _31369_ (.A(_08442_),
    .B_N(_11372_),
    .Y(_08444_));
 sg13g2_nand3b_1 _31370_ (.B(net4683),
    .C(_08443_),
    .Y(_08445_),
    .A_N(_08444_));
 sg13g2_o21ai_1 _31371_ (.B1(_08445_),
    .Y(_08446_),
    .A1(_10509_),
    .A2(net4683));
 sg13g2_a21oi_1 _31372_ (.A1(_11367_),
    .A2(_11402_),
    .Y(_08447_),
    .B1(_11430_));
 sg13g2_or2_1 _31373_ (.X(_08448_),
    .B(_08447_),
    .A(_11372_));
 sg13g2_a21oi_1 _31374_ (.A1(_11372_),
    .A2(_08447_),
    .Y(_08449_),
    .B1(net3683));
 sg13g2_nand2_1 _31375_ (.Y(_08450_),
    .A(_08448_),
    .B(_08449_));
 sg13g2_a221oi_1 _31376_ (.B2(_08446_),
    .C1(net3958),
    .B1(net3716),
    .A1(net4514),
    .Y(_08451_),
    .A2(net2265));
 sg13g2_a22oi_1 _31377_ (.Y(_01375_),
    .B1(_08450_),
    .B2(_08451_),
    .A2(net3958),
    .A1(_10510_));
 sg13g2_nand2_1 _31378_ (.Y(_08452_),
    .A(net2067),
    .B(net3958));
 sg13g2_nand2_1 _31379_ (.Y(_08453_),
    .A(\u_inv.f_next[73] ),
    .B(net3851));
 sg13g2_a21oi_1 _31380_ (.A1(\u_inv.f_next[72] ),
    .A2(\u_inv.f_reg[72] ),
    .Y(_08454_),
    .B1(_08444_));
 sg13g2_xor2_1 _31381_ (.B(_08454_),
    .A(_11373_),
    .X(_08455_));
 sg13g2_a22oi_1 _31382_ (.Y(_08456_),
    .B1(_08455_),
    .B2(net4683),
    .A2(_08453_),
    .A1(net3730));
 sg13g2_a21oi_1 _31383_ (.A1(_11410_),
    .A2(_08448_),
    .Y(_08457_),
    .B1(_11373_));
 sg13g2_and3_1 _31384_ (.X(_08458_),
    .A(_11373_),
    .B(_11410_),
    .C(_08448_));
 sg13g2_o21ai_1 _31385_ (.B1(net4383),
    .Y(_08459_),
    .A1(_08457_),
    .A2(_08458_));
 sg13g2_a21oi_1 _31386_ (.A1(net3704),
    .A2(_08459_),
    .Y(_08460_),
    .B1(_08456_));
 sg13g2_o21ai_1 _31387_ (.B1(net4027),
    .Y(_08461_),
    .A1(net4618),
    .A2(net2027));
 sg13g2_o21ai_1 _31388_ (.B1(_08452_),
    .Y(_01376_),
    .A1(_08460_),
    .A2(_08461_));
 sg13g2_nand2_1 _31389_ (.Y(_08462_),
    .A(net2308),
    .B(net3958));
 sg13g2_a21oi_1 _31390_ (.A1(\u_inv.f_next[73] ),
    .A2(_10817_),
    .Y(_08463_),
    .B1(_08457_));
 sg13g2_nor2_1 _31391_ (.A(_11370_),
    .B(_08463_),
    .Y(_08464_));
 sg13g2_a21oi_1 _31392_ (.A1(_11370_),
    .A2(_08463_),
    .Y(_08465_),
    .B1(net3851));
 sg13g2_nor2b_1 _31393_ (.A(_08464_),
    .B_N(_08465_),
    .Y(_08466_));
 sg13g2_o21ai_1 _31394_ (.B1(_12551_),
    .Y(_08467_),
    .A1(_12583_),
    .A2(_08442_));
 sg13g2_xnor2_1 _31395_ (.Y(_08468_),
    .A(_11370_),
    .B(_08467_));
 sg13g2_o21ai_1 _31396_ (.B1(net3852),
    .Y(_08469_),
    .A1(\u_inv.f_next[74] ),
    .A2(net4683));
 sg13g2_a21oi_1 _31397_ (.A1(net4683),
    .A2(_08468_),
    .Y(_08470_),
    .B1(_08469_));
 sg13g2_nor3_1 _31398_ (.A(net4445),
    .B(_08466_),
    .C(_08470_),
    .Y(_08471_));
 sg13g2_o21ai_1 _31399_ (.B1(net4027),
    .Y(_08472_),
    .A1(net4618),
    .A2(net1955));
 sg13g2_o21ai_1 _31400_ (.B1(_08462_),
    .Y(_01377_),
    .A1(_08471_),
    .A2(_08472_));
 sg13g2_nor2_1 _31401_ (.A(_11408_),
    .B(_08464_),
    .Y(_08473_));
 sg13g2_a21oi_1 _31402_ (.A1(_11368_),
    .A2(_08473_),
    .Y(_08474_),
    .B1(net3683));
 sg13g2_o21ai_1 _31403_ (.B1(_08474_),
    .Y(_08475_),
    .A1(_11368_),
    .A2(_08473_));
 sg13g2_a21oi_1 _31404_ (.A1(_11370_),
    .A2(_08467_),
    .Y(_08476_),
    .B1(_11369_));
 sg13g2_xnor2_1 _31405_ (.Y(_08477_),
    .A(_11368_),
    .B(_08476_));
 sg13g2_mux2_1 _31406_ (.A0(net2979),
    .A1(_08477_),
    .S(net4683),
    .X(_08478_));
 sg13g2_a221oi_1 _31407_ (.B2(_08478_),
    .C1(net3958),
    .B1(net3717),
    .A1(net4516),
    .Y(_08479_),
    .A2(net2496));
 sg13g2_a22oi_1 _31408_ (.Y(_01378_),
    .B1(_08475_),
    .B2(_08479_),
    .A2(net3958),
    .A1(_10507_));
 sg13g2_a21oi_2 _31409_ (.B1(_12554_),
    .Y(_08480_),
    .A2(_08467_),
    .A1(_12549_));
 sg13g2_o21ai_1 _31410_ (.B1(net4683),
    .Y(_08481_),
    .A1(_11382_),
    .A2(_08480_));
 sg13g2_a21o_1 _31411_ (.A2(_08480_),
    .A1(_11382_),
    .B1(_08481_),
    .X(_08482_));
 sg13g2_a21oi_1 _31412_ (.A1(net3037),
    .A2(net4569),
    .Y(_08483_),
    .B1(net3704));
 sg13g2_o21ai_1 _31413_ (.B1(_11413_),
    .Y(_08484_),
    .A1(_11374_),
    .A2(_08447_));
 sg13g2_and2_1 _31414_ (.A(_11382_),
    .B(_08484_),
    .X(_08485_));
 sg13g2_xnor2_1 _31415_ (.Y(_08486_),
    .A(_11382_),
    .B(_08484_));
 sg13g2_o21ai_1 _31416_ (.B1(net4028),
    .Y(_08487_),
    .A1(net4618),
    .A2(net1923));
 sg13g2_a221oi_1 _31417_ (.B2(net3695),
    .C1(_08487_),
    .B1(_08486_),
    .A1(_08482_),
    .Y(_08488_),
    .A2(_08483_));
 sg13g2_a21o_1 _31418_ (.A2(net3958),
    .A1(net2979),
    .B1(_08488_),
    .X(_01379_));
 sg13g2_nand2_1 _31419_ (.Y(_08489_),
    .A(net2769),
    .B(net3851));
 sg13g2_o21ai_1 _31420_ (.B1(_11381_),
    .Y(_08490_),
    .A1(_11382_),
    .A2(_08480_));
 sg13g2_xor2_1 _31421_ (.B(_08490_),
    .A(_11380_),
    .X(_08491_));
 sg13g2_a22oi_1 _31422_ (.Y(_08492_),
    .B1(_08491_),
    .B2(net4683),
    .A2(_08489_),
    .A1(net3730));
 sg13g2_o21ai_1 _31423_ (.B1(_11380_),
    .Y(_08493_),
    .A1(_11407_),
    .A2(_08485_));
 sg13g2_or3_1 _31424_ (.A(_11380_),
    .B(_11407_),
    .C(_08485_),
    .X(_08494_));
 sg13g2_nand2_1 _31425_ (.Y(_08495_),
    .A(_08493_),
    .B(_08494_));
 sg13g2_o21ai_1 _31426_ (.B1(net4383),
    .Y(_08496_),
    .A1(net3851),
    .A2(_08495_));
 sg13g2_a21oi_1 _31427_ (.A1(net4516),
    .A2(_10970_),
    .Y(_08497_),
    .B1(net3959));
 sg13g2_o21ai_1 _31428_ (.B1(_08497_),
    .Y(_08498_),
    .A1(_08492_),
    .A2(_08496_));
 sg13g2_o21ai_1 _31429_ (.B1(_08498_),
    .Y(_01380_),
    .A1(_10505_),
    .A2(net4027));
 sg13g2_or3_1 _31430_ (.A(_11380_),
    .B(_11382_),
    .C(_08480_),
    .X(_08499_));
 sg13g2_a21oi_1 _31431_ (.A1(_12558_),
    .A2(_08499_),
    .Y(_08500_),
    .B1(_11378_));
 sg13g2_nand3_1 _31432_ (.B(_12558_),
    .C(_08499_),
    .A(_11378_),
    .Y(_08501_));
 sg13g2_nand3b_1 _31433_ (.B(_08501_),
    .C(net4684),
    .Y(_08502_),
    .A_N(_08500_));
 sg13g2_a21oi_1 _31434_ (.A1(net2271),
    .A2(net4569),
    .Y(_08503_),
    .B1(net3705));
 sg13g2_nand2_1 _31435_ (.Y(_08504_),
    .A(_11406_),
    .B(_08493_));
 sg13g2_xnor2_1 _31436_ (.Y(_08505_),
    .A(_11378_),
    .B(_08504_));
 sg13g2_o21ai_1 _31437_ (.B1(net4027),
    .Y(_08506_),
    .A1(net4618),
    .A2(net1895));
 sg13g2_a221oi_1 _31438_ (.B2(net3695),
    .C1(_08506_),
    .B1(_08505_),
    .A1(_08502_),
    .Y(_08507_),
    .A2(_08503_));
 sg13g2_a21o_1 _31439_ (.A2(net3958),
    .A1(net2769),
    .B1(_08507_),
    .X(_01381_));
 sg13g2_nand2_1 _31440_ (.Y(_08508_),
    .A(net2568),
    .B(net3851));
 sg13g2_nor2_1 _31441_ (.A(_11377_),
    .B(_08500_),
    .Y(_08509_));
 sg13g2_xnor2_1 _31442_ (.Y(_08510_),
    .A(_11376_),
    .B(_08509_));
 sg13g2_a22oi_1 _31443_ (.Y(_08511_),
    .B1(_08510_),
    .B2(net4684),
    .A2(_08508_),
    .A1(net3730));
 sg13g2_a21oi_1 _31444_ (.A1(_11378_),
    .A2(_08504_),
    .Y(_08512_),
    .B1(_11431_));
 sg13g2_xor2_1 _31445_ (.B(_08512_),
    .A(_11376_),
    .X(_08513_));
 sg13g2_o21ai_1 _31446_ (.B1(net4383),
    .Y(_08514_),
    .A1(net3851),
    .A2(_08513_));
 sg13g2_a21oi_1 _31447_ (.A1(net4516),
    .A2(_10971_),
    .Y(_08515_),
    .B1(net3959));
 sg13g2_o21ai_1 _31448_ (.B1(_08515_),
    .Y(_08516_),
    .A1(_08511_),
    .A2(_08514_));
 sg13g2_o21ai_1 _31449_ (.B1(_08516_),
    .Y(_01382_),
    .A1(_10503_),
    .A2(net4028));
 sg13g2_o21ai_1 _31450_ (.B1(_12584_),
    .Y(_08517_),
    .A1(_12582_),
    .A2(_08441_));
 sg13g2_nand3_1 _31451_ (.B(_12561_),
    .C(_08517_),
    .A(_11468_),
    .Y(_08518_));
 sg13g2_a21oi_1 _31452_ (.A1(_12561_),
    .A2(_08517_),
    .Y(_08519_),
    .B1(_11468_));
 sg13g2_nand3b_1 _31453_ (.B(net4684),
    .C(_08518_),
    .Y(_08520_),
    .A_N(_08519_));
 sg13g2_a21oi_1 _31454_ (.A1(net3071),
    .A2(net4569),
    .Y(_08521_),
    .B1(net3705));
 sg13g2_o21ai_1 _31455_ (.B1(_11468_),
    .Y(_08522_),
    .A1(_11405_),
    .A2(_11434_));
 sg13g2_xor2_1 _31456_ (.B(_11468_),
    .A(_11435_),
    .X(_08523_));
 sg13g2_o21ai_1 _31457_ (.B1(net4027),
    .Y(_08524_),
    .A1(net4618),
    .A2(net1847));
 sg13g2_a221oi_1 _31458_ (.B2(net3695),
    .C1(_08524_),
    .B1(_08523_),
    .A1(_08520_),
    .Y(_08525_),
    .A2(_08521_));
 sg13g2_a21o_1 _31459_ (.A2(net3959),
    .A1(net2568),
    .B1(_08525_),
    .X(_01383_));
 sg13g2_nand2_1 _31460_ (.Y(_08526_),
    .A(net2375),
    .B(net3851));
 sg13g2_a21o_1 _31461_ (.A2(\u_inv.f_reg[80] ),
    .A1(\u_inv.f_next[80] ),
    .B1(_08519_),
    .X(_08527_));
 sg13g2_xnor2_1 _31462_ (.Y(_08528_),
    .A(_11471_),
    .B(_08527_));
 sg13g2_a22oi_1 _31463_ (.Y(_08529_),
    .B1(_08528_),
    .B2(net4684),
    .A2(_08526_),
    .A1(net3730));
 sg13g2_a21oi_1 _31464_ (.A1(_11480_),
    .A2(_08522_),
    .Y(_08530_),
    .B1(_11471_));
 sg13g2_nand3_1 _31465_ (.B(_11480_),
    .C(_08522_),
    .A(_11471_),
    .Y(_08531_));
 sg13g2_nand2_1 _31466_ (.Y(_08532_),
    .A(net3822),
    .B(_08531_));
 sg13g2_o21ai_1 _31467_ (.B1(net4383),
    .Y(_08533_),
    .A1(_08530_),
    .A2(_08532_));
 sg13g2_a21oi_1 _31468_ (.A1(net4516),
    .A2(_10972_),
    .Y(_08534_),
    .B1(net3959));
 sg13g2_o21ai_1 _31469_ (.B1(_08534_),
    .Y(_08535_),
    .A1(_08529_),
    .A2(_08533_));
 sg13g2_o21ai_1 _31470_ (.B1(_08535_),
    .Y(_01384_),
    .A1(_10501_),
    .A2(net4027));
 sg13g2_nand2_1 _31471_ (.Y(_08536_),
    .A(_11469_),
    .B(_08527_));
 sg13g2_nand2_1 _31472_ (.Y(_08537_),
    .A(_11470_),
    .B(_08536_));
 sg13g2_inv_1 _31473_ (.Y(_08538_),
    .A(_08537_));
 sg13g2_o21ai_1 _31474_ (.B1(net4687),
    .Y(_08539_),
    .A1(_11466_),
    .A2(_08538_));
 sg13g2_a21o_1 _31475_ (.A2(_08538_),
    .A1(_11466_),
    .B1(_08539_),
    .X(_08540_));
 sg13g2_a21oi_1 _31476_ (.A1(\u_inv.f_next[82] ),
    .A2(net4568),
    .Y(_08541_),
    .B1(net3705));
 sg13g2_o21ai_1 _31477_ (.B1(_11466_),
    .Y(_08542_),
    .A1(_11479_),
    .A2(_08530_));
 sg13g2_or3_1 _31478_ (.A(_11466_),
    .B(_11479_),
    .C(_08530_),
    .X(_08543_));
 sg13g2_nand2_1 _31479_ (.Y(_08544_),
    .A(_08542_),
    .B(_08543_));
 sg13g2_o21ai_1 _31480_ (.B1(net4027),
    .Y(_08545_),
    .A1(net4619),
    .A2(net2099));
 sg13g2_a221oi_1 _31481_ (.B2(net3695),
    .C1(_08545_),
    .B1(_08544_),
    .A1(_08540_),
    .Y(_08546_),
    .A2(_08541_));
 sg13g2_a21o_1 _31482_ (.A2(net3959),
    .A1(net2375),
    .B1(_08546_),
    .X(_01385_));
 sg13g2_o21ai_1 _31483_ (.B1(_11465_),
    .Y(_08547_),
    .A1(_11466_),
    .A2(_08538_));
 sg13g2_xnor2_1 _31484_ (.Y(_08548_),
    .A(_11463_),
    .B(_08547_));
 sg13g2_o21ai_1 _31485_ (.B1(net3717),
    .Y(_08549_),
    .A1(net3084),
    .A2(net4687));
 sg13g2_a21o_1 _31486_ (.A2(_08548_),
    .A1(net4687),
    .B1(_08549_),
    .X(_08550_));
 sg13g2_a21oi_1 _31487_ (.A1(_11478_),
    .A2(_08542_),
    .Y(_08551_),
    .B1(_11463_));
 sg13g2_nand3_1 _31488_ (.B(_11478_),
    .C(_08542_),
    .A(_11463_),
    .Y(_08552_));
 sg13g2_nor2_1 _31489_ (.A(net3683),
    .B(_08551_),
    .Y(_08553_));
 sg13g2_a221oi_1 _31490_ (.B2(_08553_),
    .C1(net3962),
    .B1(_08552_),
    .A1(net4517),
    .Y(_08554_),
    .A2(net2597));
 sg13g2_a22oi_1 _31491_ (.Y(_01386_),
    .B1(_08550_),
    .B2(_08554_),
    .A2(net3962),
    .A1(_10499_));
 sg13g2_a21oi_2 _31492_ (.B1(_12569_),
    .Y(_08555_),
    .A2(_08519_),
    .A1(_12564_));
 sg13g2_inv_1 _31493_ (.Y(_08556_),
    .A(_08555_));
 sg13g2_nand2_1 _31494_ (.Y(_08557_),
    .A(_11459_),
    .B(_08555_));
 sg13g2_nor2_1 _31495_ (.A(_11459_),
    .B(_08555_),
    .Y(_08558_));
 sg13g2_nor2_1 _31496_ (.A(net4568),
    .B(_08558_),
    .Y(_08559_));
 sg13g2_a221oi_1 _31497_ (.B2(_08559_),
    .C1(net3705),
    .B1(_08557_),
    .A1(net3153),
    .Y(_08560_),
    .A2(net4568));
 sg13g2_o21ai_1 _31498_ (.B1(_11484_),
    .Y(_08561_),
    .A1(_11435_),
    .A2(_11472_));
 sg13g2_nand2_1 _31499_ (.Y(_08562_),
    .A(_11459_),
    .B(_08561_));
 sg13g2_or2_1 _31500_ (.X(_08563_),
    .B(_08561_),
    .A(_11459_));
 sg13g2_a21oi_1 _31501_ (.A1(_08562_),
    .A2(_08563_),
    .Y(_08564_),
    .B1(net3683));
 sg13g2_o21ai_1 _31502_ (.B1(net4029),
    .Y(_08565_),
    .A1(net4619),
    .A2(net1858));
 sg13g2_nor3_1 _31503_ (.A(_08560_),
    .B(_08564_),
    .C(_08565_),
    .Y(_08566_));
 sg13g2_a21o_1 _31504_ (.A2(net3962),
    .A1(net3084),
    .B1(_08566_),
    .X(_01387_));
 sg13g2_a21oi_1 _31505_ (.A1(\u_inv.f_next[84] ),
    .A2(net2532),
    .Y(_08567_),
    .B1(_08558_));
 sg13g2_xnor2_1 _31506_ (.Y(_08568_),
    .A(_11461_),
    .B(_08567_));
 sg13g2_o21ai_1 _31507_ (.B1(net3717),
    .Y(_08569_),
    .A1(\u_inv.f_next[85] ),
    .A2(net4687));
 sg13g2_a21o_1 _31508_ (.A2(_08568_),
    .A1(net4687),
    .B1(_08569_),
    .X(_08570_));
 sg13g2_and2_1 _31509_ (.A(_11486_),
    .B(_08562_),
    .X(_08571_));
 sg13g2_or2_1 _31510_ (.X(_08572_),
    .B(_08571_),
    .A(_11460_));
 sg13g2_a21oi_1 _31511_ (.A1(_11460_),
    .A2(_08571_),
    .Y(_08573_),
    .B1(net3683));
 sg13g2_a221oi_1 _31512_ (.B2(_08573_),
    .C1(net3962),
    .B1(_08572_),
    .A1(net4517),
    .Y(_08574_),
    .A2(net2268));
 sg13g2_a22oi_1 _31513_ (.Y(_01388_),
    .B1(_08570_),
    .B2(_08574_),
    .A2(net3962),
    .A1(_10497_));
 sg13g2_a21oi_1 _31514_ (.A1(_12545_),
    .A2(_08556_),
    .Y(_08575_),
    .B1(_12542_));
 sg13g2_a21oi_1 _31515_ (.A1(_11457_),
    .A2(_08575_),
    .Y(_08576_),
    .B1(net4568));
 sg13g2_o21ai_1 _31516_ (.B1(_08576_),
    .Y(_08577_),
    .A1(_11457_),
    .A2(_08575_));
 sg13g2_a21oi_1 _31517_ (.A1(net3227),
    .A2(net4568),
    .Y(_08578_),
    .B1(net3705));
 sg13g2_nand2_1 _31518_ (.Y(_08579_),
    .A(_11485_),
    .B(_08572_));
 sg13g2_and2_1 _31519_ (.A(_11457_),
    .B(_08579_),
    .X(_08580_));
 sg13g2_xnor2_1 _31520_ (.Y(_08581_),
    .A(_11457_),
    .B(_08579_));
 sg13g2_o21ai_1 _31521_ (.B1(net4028),
    .Y(_08582_),
    .A1(net4619),
    .A2(net2025));
 sg13g2_a221oi_1 _31522_ (.B2(net3695),
    .C1(_08582_),
    .B1(_08581_),
    .A1(_08577_),
    .Y(_08583_),
    .A2(_08578_));
 sg13g2_a21o_1 _31523_ (.A2(net3962),
    .A1(net3156),
    .B1(_08583_),
    .X(_01389_));
 sg13g2_o21ai_1 _31524_ (.B1(_11456_),
    .Y(_08584_),
    .A1(_11457_),
    .A2(_08575_));
 sg13g2_or2_1 _31525_ (.X(_08585_),
    .B(_08584_),
    .A(_11455_));
 sg13g2_a21oi_1 _31526_ (.A1(_11455_),
    .A2(_08584_),
    .Y(_08586_),
    .B1(net4569));
 sg13g2_o21ai_1 _31527_ (.B1(net3717),
    .Y(_08587_),
    .A1(net2819),
    .A2(net4684));
 sg13g2_a21o_1 _31528_ (.A2(_08586_),
    .A1(_08585_),
    .B1(_08587_),
    .X(_08588_));
 sg13g2_nor3_1 _31529_ (.A(_11455_),
    .B(_11488_),
    .C(_08580_),
    .Y(_08589_));
 sg13g2_o21ai_1 _31530_ (.B1(_11455_),
    .Y(_08590_),
    .A1(_11488_),
    .A2(_08580_));
 sg13g2_nor2_1 _31531_ (.A(net3683),
    .B(_08589_),
    .Y(_08591_));
 sg13g2_a221oi_1 _31532_ (.B2(_08591_),
    .C1(net3962),
    .B1(_08590_),
    .A1(net4516),
    .Y(_08592_),
    .A2(net2182));
 sg13g2_a22oi_1 _31533_ (.Y(_01390_),
    .B1(_08588_),
    .B2(_08592_),
    .A2(net3959),
    .A1(_10495_));
 sg13g2_o21ai_1 _31534_ (.B1(_12544_),
    .Y(_08593_),
    .A1(_12546_),
    .A2(_08555_));
 sg13g2_o21ai_1 _31535_ (.B1(net4686),
    .Y(_08594_),
    .A1(_11452_),
    .A2(_08593_));
 sg13g2_a21o_1 _31536_ (.A2(_08593_),
    .A1(_11452_),
    .B1(_08594_),
    .X(_08595_));
 sg13g2_a21oi_1 _31537_ (.A1(\u_inv.f_next[88] ),
    .A2(net4568),
    .Y(_08596_),
    .B1(net3705));
 sg13g2_o21ai_1 _31538_ (.B1(_11492_),
    .Y(_08597_),
    .A1(_11435_),
    .A2(_11474_));
 sg13g2_nor2b_1 _31539_ (.A(_11452_),
    .B_N(_08597_),
    .Y(_08598_));
 sg13g2_xor2_1 _31540_ (.B(_08597_),
    .A(_11452_),
    .X(_08599_));
 sg13g2_o21ai_1 _31541_ (.B1(net4029),
    .Y(_08600_),
    .A1(net4618),
    .A2(net1861));
 sg13g2_a221oi_1 _31542_ (.B2(net3696),
    .C1(_08600_),
    .B1(_08599_),
    .A1(_08595_),
    .Y(_08601_),
    .A2(_08596_));
 sg13g2_a21o_1 _31543_ (.A2(net3962),
    .A1(net2819),
    .B1(_08601_),
    .X(_01391_));
 sg13g2_a21oi_1 _31544_ (.A1(_11452_),
    .A2(_08593_),
    .Y(_08602_),
    .B1(_11451_));
 sg13g2_xor2_1 _31545_ (.B(_08602_),
    .A(_11448_),
    .X(_08603_));
 sg13g2_o21ai_1 _31546_ (.B1(net3717),
    .Y(_08604_),
    .A1(net2865),
    .A2(net4686));
 sg13g2_a21o_1 _31547_ (.A2(_08603_),
    .A1(net4686),
    .B1(_08604_),
    .X(_08605_));
 sg13g2_a21oi_1 _31548_ (.A1(\u_inv.f_next[88] ),
    .A2(_10802_),
    .Y(_08606_),
    .B1(_08598_));
 sg13g2_xor2_1 _31549_ (.B(_08606_),
    .A(_11448_),
    .X(_08607_));
 sg13g2_a221oi_1 _31550_ (.B2(_08607_),
    .C1(net3960),
    .B1(net3696),
    .A1(net4516),
    .Y(_08608_),
    .A2(net2204));
 sg13g2_a22oi_1 _31551_ (.Y(_01392_),
    .B1(_08605_),
    .B2(_08608_),
    .A2(net3960),
    .A1(_10493_));
 sg13g2_a21oi_2 _31552_ (.B1(_12591_),
    .Y(_08609_),
    .A2(_08593_),
    .A1(_12538_));
 sg13g2_xnor2_1 _31553_ (.Y(_08610_),
    .A(_11447_),
    .B(_08609_));
 sg13g2_o21ai_1 _31554_ (.B1(net3717),
    .Y(_08611_),
    .A1(net3111),
    .A2(net4686));
 sg13g2_a21oi_1 _31555_ (.A1(net4686),
    .A2(_08610_),
    .Y(_08612_),
    .B1(_08611_));
 sg13g2_o21ai_1 _31556_ (.B1(_11500_),
    .Y(_08613_),
    .A1(_11448_),
    .A2(_08606_));
 sg13g2_and2_1 _31557_ (.A(_11447_),
    .B(_08613_),
    .X(_08614_));
 sg13g2_o21ai_1 _31558_ (.B1(net3695),
    .Y(_08615_),
    .A1(_11447_),
    .A2(_08613_));
 sg13g2_a21oi_1 _31559_ (.A1(net4516),
    .A2(net1886),
    .Y(_08616_),
    .B1(net3960));
 sg13g2_o21ai_1 _31560_ (.B1(_08616_),
    .Y(_08617_),
    .A1(_08614_),
    .A2(_08615_));
 sg13g2_nor2_1 _31561_ (.A(_08612_),
    .B(_08617_),
    .Y(_08618_));
 sg13g2_a21oi_1 _31562_ (.A1(_10492_),
    .A2(net3961),
    .Y(_01393_),
    .B1(_08618_));
 sg13g2_nand2_1 _31563_ (.Y(_08619_),
    .A(net2940),
    .B(net3852));
 sg13g2_o21ai_1 _31564_ (.B1(_11445_),
    .Y(_08620_),
    .A1(_11447_),
    .A2(_08609_));
 sg13g2_xnor2_1 _31565_ (.Y(_08621_),
    .A(_11449_),
    .B(_08620_));
 sg13g2_a22oi_1 _31566_ (.Y(_08622_),
    .B1(_08621_),
    .B2(net4686),
    .A2(_08619_),
    .A1(net3730));
 sg13g2_nor2_1 _31567_ (.A(_11499_),
    .B(_08614_),
    .Y(_08623_));
 sg13g2_xnor2_1 _31568_ (.Y(_08624_),
    .A(_11449_),
    .B(_08623_));
 sg13g2_o21ai_1 _31569_ (.B1(net4383),
    .Y(_08625_),
    .A1(net3852),
    .A2(_08624_));
 sg13g2_a21oi_1 _31570_ (.A1(net4516),
    .A2(_10973_),
    .Y(_08626_),
    .B1(net3960));
 sg13g2_o21ai_1 _31571_ (.B1(_08626_),
    .Y(_08627_),
    .A1(_08622_),
    .A2(_08625_));
 sg13g2_o21ai_1 _31572_ (.B1(_08627_),
    .Y(_01394_),
    .A1(_10491_),
    .A2(net4028));
 sg13g2_o21ai_1 _31573_ (.B1(_12594_),
    .Y(_08628_),
    .A1(_12539_),
    .A2(_08609_));
 sg13g2_a21oi_1 _31574_ (.A1(_11442_),
    .A2(_08628_),
    .Y(_08629_),
    .B1(net4569));
 sg13g2_o21ai_1 _31575_ (.B1(_08629_),
    .Y(_08630_),
    .A1(_11442_),
    .A2(_08628_));
 sg13g2_a21oi_1 _31576_ (.A1(net2353),
    .A2(net4568),
    .Y(_08631_),
    .B1(net3705));
 sg13g2_a21oi_1 _31577_ (.A1(_11450_),
    .A2(_08598_),
    .Y(_08632_),
    .B1(_11504_));
 sg13g2_nor2_1 _31578_ (.A(_11442_),
    .B(_08632_),
    .Y(_08633_));
 sg13g2_xnor2_1 _31579_ (.Y(_08634_),
    .A(_11442_),
    .B(_08632_));
 sg13g2_o21ai_1 _31580_ (.B1(net4028),
    .Y(_08635_),
    .A1(net4619),
    .A2(net1733));
 sg13g2_a221oi_1 _31581_ (.B2(net3695),
    .C1(_08635_),
    .B1(_08634_),
    .A1(_08630_),
    .Y(_08636_),
    .A2(_08631_));
 sg13g2_a21o_1 _31582_ (.A2(net3960),
    .A1(net2940),
    .B1(_08636_),
    .X(_01395_));
 sg13g2_a21oi_1 _31583_ (.A1(_11442_),
    .A2(_08628_),
    .Y(_08637_),
    .B1(_11441_));
 sg13g2_xnor2_1 _31584_ (.Y(_08638_),
    .A(_11440_),
    .B(_08637_));
 sg13g2_nand2_1 _31585_ (.Y(_08639_),
    .A(net4687),
    .B(_08638_));
 sg13g2_a21oi_1 _31586_ (.A1(\u_inv.f_next[93] ),
    .A2(net4568),
    .Y(_08640_),
    .B1(net3705));
 sg13g2_nor2_1 _31587_ (.A(_11494_),
    .B(_08633_),
    .Y(_08641_));
 sg13g2_xnor2_1 _31588_ (.Y(_08642_),
    .A(_11440_),
    .B(_08641_));
 sg13g2_o21ai_1 _31589_ (.B1(net4028),
    .Y(_08643_),
    .A1(net4619),
    .A2(net1920));
 sg13g2_a221oi_1 _31590_ (.B2(net3695),
    .C1(_08643_),
    .B1(_08642_),
    .A1(_08639_),
    .Y(_08644_),
    .A2(_08640_));
 sg13g2_a21o_1 _31591_ (.A2(net3961),
    .A1(net2353),
    .B1(_08644_),
    .X(_01396_));
 sg13g2_a21oi_1 _31592_ (.A1(_12536_),
    .A2(_08628_),
    .Y(_08645_),
    .B1(_12586_));
 sg13g2_xnor2_1 _31593_ (.Y(_08646_),
    .A(_11438_),
    .B(_08645_));
 sg13g2_a21oi_1 _31594_ (.A1(net4686),
    .A2(_08646_),
    .Y(_08647_),
    .B1(net3706));
 sg13g2_o21ai_1 _31595_ (.B1(_08647_),
    .Y(_08648_),
    .A1(net1799),
    .A2(net4686));
 sg13g2_o21ai_1 _31596_ (.B1(_11493_),
    .Y(_08649_),
    .A1(_11440_),
    .A2(_08641_));
 sg13g2_or2_1 _31597_ (.X(_08650_),
    .B(_08649_),
    .A(_11438_));
 sg13g2_and2_1 _31598_ (.A(_11438_),
    .B(_08649_),
    .X(_08651_));
 sg13g2_nor2_1 _31599_ (.A(net3683),
    .B(_08651_),
    .Y(_08652_));
 sg13g2_a221oi_1 _31600_ (.B2(_08652_),
    .C1(net3961),
    .B1(_08650_),
    .A1(net4517),
    .Y(_08653_),
    .A2(net2385));
 sg13g2_a22oi_1 _31601_ (.Y(_01397_),
    .B1(_08648_),
    .B2(_08653_),
    .A2(net3961),
    .A1(_10488_));
 sg13g2_nand2_1 _31602_ (.Y(_08654_),
    .A(net1799),
    .B(net3960));
 sg13g2_o21ai_1 _31603_ (.B1(_11437_),
    .Y(_08655_),
    .A1(_11438_),
    .A2(_08645_));
 sg13g2_nand2_1 _31604_ (.Y(_08656_),
    .A(_11436_),
    .B(_08655_));
 sg13g2_nor2_1 _31605_ (.A(_11436_),
    .B(_08655_),
    .Y(_08657_));
 sg13g2_nor2_1 _31606_ (.A(net4582),
    .B(_08657_),
    .Y(_08658_));
 sg13g2_a221oi_1 _31607_ (.B2(_08658_),
    .C1(net3799),
    .B1(_08656_),
    .A1(_10486_),
    .Y(_08659_),
    .A2(net4582));
 sg13g2_nor2_1 _31608_ (.A(_11497_),
    .B(_08651_),
    .Y(_08660_));
 sg13g2_xor2_1 _31609_ (.B(_08660_),
    .A(_11436_),
    .X(_08661_));
 sg13g2_o21ai_1 _31610_ (.B1(net4383),
    .Y(_08662_),
    .A1(net3855),
    .A2(_08661_));
 sg13g2_nor2_1 _31611_ (.A(_08659_),
    .B(_08662_),
    .Y(_08663_));
 sg13g2_o21ai_1 _31612_ (.B1(net4028),
    .Y(_08664_),
    .A1(net4620),
    .A2(\u_inv.input_reg[94] ));
 sg13g2_o21ai_1 _31613_ (.B1(_08654_),
    .Y(_01398_),
    .A1(_08663_),
    .A2(_08664_));
 sg13g2_o21ai_1 _31614_ (.B1(net3699),
    .Y(_08665_),
    .A1(_11509_),
    .A2(_11567_));
 sg13g2_a21oi_1 _31615_ (.A1(_11509_),
    .A2(_11567_),
    .Y(_08666_),
    .B1(_08665_));
 sg13g2_nand2b_1 _31616_ (.Y(_08667_),
    .B(_12746_),
    .A_N(_11567_));
 sg13g2_xnor2_1 _31617_ (.Y(_08668_),
    .A(_11567_),
    .B(_12745_));
 sg13g2_a21oi_1 _31618_ (.A1(net4703),
    .A2(_08668_),
    .Y(_08669_),
    .B1(net3706));
 sg13g2_o21ai_1 _31619_ (.B1(_08669_),
    .Y(_08670_),
    .A1(net2499),
    .A2(net4695));
 sg13g2_nor2b_1 _31620_ (.A(net4620),
    .B_N(net1637),
    .Y(_08671_));
 sg13g2_nor3_1 _31621_ (.A(net3971),
    .B(_08666_),
    .C(_08671_),
    .Y(_08672_));
 sg13g2_a22oi_1 _31622_ (.Y(_01399_),
    .B1(_08670_),
    .B2(_08672_),
    .A2(net3971),
    .A1(_10486_));
 sg13g2_a21oi_1 _31623_ (.A1(_11509_),
    .A2(_11567_),
    .Y(_08673_),
    .B1(_11602_));
 sg13g2_or2_1 _31624_ (.X(_08674_),
    .B(_08673_),
    .A(_11569_));
 sg13g2_a21oi_1 _31625_ (.A1(_11569_),
    .A2(_08673_),
    .Y(_08675_),
    .B1(net3684));
 sg13g2_o21ai_1 _31626_ (.B1(_08667_),
    .Y(_08676_),
    .A1(_10485_),
    .A2(_10794_));
 sg13g2_nor2_1 _31627_ (.A(_10484_),
    .B(net4696),
    .Y(_08677_));
 sg13g2_o21ai_1 _31628_ (.B1(net4704),
    .Y(_08678_),
    .A1(_11569_),
    .A2(_08676_));
 sg13g2_a21oi_1 _31629_ (.A1(_11569_),
    .A2(_08676_),
    .Y(_08679_),
    .B1(_08678_));
 sg13g2_o21ai_1 _31630_ (.B1(net3717),
    .Y(_08680_),
    .A1(_08677_),
    .A2(_08679_));
 sg13g2_a221oi_1 _31631_ (.B2(_08675_),
    .C1(net3972),
    .B1(_08674_),
    .A1(net4518),
    .Y(_08681_),
    .A2(net2398));
 sg13g2_a22oi_1 _31632_ (.Y(_01400_),
    .B1(_08680_),
    .B2(_08681_),
    .A2(net3980),
    .A1(_10485_));
 sg13g2_nand2_1 _31633_ (.Y(_08682_),
    .A(_11601_),
    .B(_08674_));
 sg13g2_and2_1 _31634_ (.A(_11565_),
    .B(_08682_),
    .X(_08683_));
 sg13g2_nor2_1 _31635_ (.A(net3684),
    .B(_08683_),
    .Y(_08684_));
 sg13g2_o21ai_1 _31636_ (.B1(_08684_),
    .Y(_08685_),
    .A1(_11565_),
    .A2(_08682_));
 sg13g2_a21oi_1 _31637_ (.A1(_12468_),
    .A2(_08667_),
    .Y(_08686_),
    .B1(_11568_));
 sg13g2_nor2b_1 _31638_ (.A(_11565_),
    .B_N(_08686_),
    .Y(_08687_));
 sg13g2_xor2_1 _31639_ (.B(_08686_),
    .A(_11565_),
    .X(_08688_));
 sg13g2_nor2_1 _31640_ (.A(net2086),
    .B(net4696),
    .Y(_08689_));
 sg13g2_a21oi_1 _31641_ (.A1(net4696),
    .A2(_08688_),
    .Y(_08690_),
    .B1(_08689_));
 sg13g2_a221oi_1 _31642_ (.B2(_08690_),
    .C1(net3972),
    .B1(net3717),
    .A1(net4518),
    .Y(_08691_),
    .A2(net2541));
 sg13g2_a22oi_1 _31643_ (.Y(_01401_),
    .B1(_08685_),
    .B2(_08691_),
    .A2(net3973),
    .A1(_10484_));
 sg13g2_nand2_1 _31644_ (.Y(_08692_),
    .A(net2086),
    .B(net3973));
 sg13g2_nor2_1 _31645_ (.A(_11606_),
    .B(_08683_),
    .Y(_08693_));
 sg13g2_xor2_1 _31646_ (.B(_08693_),
    .A(_11566_),
    .X(_08694_));
 sg13g2_nor2_1 _31647_ (.A(net3863),
    .B(_08694_),
    .Y(_08695_));
 sg13g2_nand2_1 _31648_ (.Y(_08696_),
    .A(net1761),
    .B(net3860));
 sg13g2_a21oi_1 _31649_ (.A1(\u_inv.f_next[98] ),
    .A2(\u_inv.f_reg[98] ),
    .Y(_08697_),
    .B1(_08687_));
 sg13g2_xnor2_1 _31650_ (.Y(_08698_),
    .A(_11566_),
    .B(_08697_));
 sg13g2_a22oi_1 _31651_ (.Y(_08699_),
    .B1(_08698_),
    .B2(net4704),
    .A2(_08696_),
    .A1(net3735));
 sg13g2_nor3_1 _31652_ (.A(net4448),
    .B(_08695_),
    .C(_08699_),
    .Y(_08700_));
 sg13g2_o21ai_1 _31653_ (.B1(net4031),
    .Y(_08701_),
    .A1(net4623),
    .A2(net1929));
 sg13g2_o21ai_1 _31654_ (.B1(_08692_),
    .Y(_01402_),
    .A1(_08700_),
    .A2(_08701_));
 sg13g2_nand2_1 _31655_ (.Y(_08702_),
    .A(net1761),
    .B(net3980));
 sg13g2_a21oi_1 _31656_ (.A1(_11509_),
    .A2(_11571_),
    .Y(_08703_),
    .B1(_11608_));
 sg13g2_or2_1 _31657_ (.X(_08704_),
    .B(_08703_),
    .A(_11575_));
 sg13g2_a21oi_1 _31658_ (.A1(_11575_),
    .A2(_08703_),
    .Y(_08705_),
    .B1(net3860));
 sg13g2_o21ai_1 _31659_ (.B1(_12472_),
    .Y(_08706_),
    .A1(_12747_),
    .A2(_08667_));
 sg13g2_xnor2_1 _31660_ (.Y(_08707_),
    .A(_11575_),
    .B(_08706_));
 sg13g2_nor2_1 _31661_ (.A(\u_inv.f_next[100] ),
    .B(net4703),
    .Y(_08708_));
 sg13g2_a21oi_1 _31662_ (.A1(net4703),
    .A2(_08707_),
    .Y(_08709_),
    .B1(_08708_));
 sg13g2_a221oi_1 _31663_ (.B2(net3860),
    .C1(net4448),
    .B1(_08709_),
    .A1(_08704_),
    .Y(_08710_),
    .A2(_08705_));
 sg13g2_o21ai_1 _31664_ (.B1(net4032),
    .Y(_08711_),
    .A1(net4623),
    .A2(\u_inv.input_reg[99] ));
 sg13g2_o21ai_1 _31665_ (.B1(_08702_),
    .Y(_01403_),
    .A1(_08710_),
    .A2(_08711_));
 sg13g2_nand2_1 _31666_ (.Y(_08712_),
    .A(_11609_),
    .B(_08704_));
 sg13g2_a21oi_1 _31667_ (.A1(_11609_),
    .A2(_08704_),
    .Y(_08713_),
    .B1(_11573_));
 sg13g2_o21ai_1 _31668_ (.B1(net3699),
    .Y(_08714_),
    .A1(_11572_),
    .A2(_08712_));
 sg13g2_a21oi_1 _31669_ (.A1(_11575_),
    .A2(_08706_),
    .Y(_08715_),
    .B1(_11574_));
 sg13g2_xnor2_1 _31670_ (.Y(_08716_),
    .A(_11572_),
    .B(_08715_));
 sg13g2_o21ai_1 _31671_ (.B1(net3720),
    .Y(_08717_),
    .A1(net2018),
    .A2(net4703));
 sg13g2_a21oi_1 _31672_ (.A1(net4703),
    .A2(_08716_),
    .Y(_08718_),
    .B1(_08717_));
 sg13g2_a21oi_1 _31673_ (.A1(net4518),
    .A2(net1980),
    .Y(_08719_),
    .B1(net3973));
 sg13g2_o21ai_1 _31674_ (.B1(_08719_),
    .Y(_08720_),
    .A1(_08713_),
    .A2(_08714_));
 sg13g2_nor2_1 _31675_ (.A(_08718_),
    .B(_08720_),
    .Y(_08721_));
 sg13g2_a21oi_1 _31676_ (.A1(_10481_),
    .A2(net3980),
    .Y(_01404_),
    .B1(_08721_));
 sg13g2_nand2_1 _31677_ (.Y(_08722_),
    .A(net2018),
    .B(net3980));
 sg13g2_or2_1 _31678_ (.X(_08723_),
    .B(_08713_),
    .A(_11610_));
 sg13g2_nor2_1 _31679_ (.A(_11580_),
    .B(_08723_),
    .Y(_08724_));
 sg13g2_and2_1 _31680_ (.A(_11580_),
    .B(_08723_),
    .X(_08725_));
 sg13g2_nor3_1 _31681_ (.A(net3860),
    .B(_08724_),
    .C(_08725_),
    .Y(_08726_));
 sg13g2_a21oi_1 _31682_ (.A1(_12465_),
    .A2(_08706_),
    .Y(_08727_),
    .B1(_12476_));
 sg13g2_xnor2_1 _31683_ (.Y(_08728_),
    .A(_11580_),
    .B(_08727_));
 sg13g2_o21ai_1 _31684_ (.B1(net3863),
    .Y(_08729_),
    .A1(\u_inv.f_next[102] ),
    .A2(net4703));
 sg13g2_a21oi_1 _31685_ (.A1(net4703),
    .A2(_08728_),
    .Y(_08730_),
    .B1(_08729_));
 sg13g2_nor3_1 _31686_ (.A(net4448),
    .B(_08726_),
    .C(_08730_),
    .Y(_08731_));
 sg13g2_o21ai_1 _31687_ (.B1(net4035),
    .Y(_08732_),
    .A1(net4623),
    .A2(net1876));
 sg13g2_o21ai_1 _31688_ (.B1(_08722_),
    .Y(_01405_),
    .A1(_08731_),
    .A2(_08732_));
 sg13g2_o21ai_1 _31689_ (.B1(_11579_),
    .Y(_08733_),
    .A1(_11580_),
    .A2(_08727_));
 sg13g2_a21oi_1 _31690_ (.A1(_11577_),
    .A2(_08733_),
    .Y(_08734_),
    .B1(net4591));
 sg13g2_o21ai_1 _31691_ (.B1(_08734_),
    .Y(_08735_),
    .A1(_11577_),
    .A2(_08733_));
 sg13g2_o21ai_1 _31692_ (.B1(_08735_),
    .Y(_08736_),
    .A1(_10478_),
    .A2(net4703));
 sg13g2_a21oi_1 _31693_ (.A1(net3860),
    .A2(_08736_),
    .Y(_08737_),
    .B1(net4448));
 sg13g2_nor2_1 _31694_ (.A(_11614_),
    .B(_08725_),
    .Y(_08738_));
 sg13g2_a21oi_1 _31695_ (.A1(_11577_),
    .A2(_08738_),
    .Y(_08739_),
    .B1(net3860));
 sg13g2_o21ai_1 _31696_ (.B1(_08739_),
    .Y(_08740_),
    .A1(_11577_),
    .A2(_08738_));
 sg13g2_o21ai_1 _31697_ (.B1(net4035),
    .Y(_08741_),
    .A1(net4623),
    .A2(net2075));
 sg13g2_a21o_1 _31698_ (.A2(_08740_),
    .A1(_08737_),
    .B1(_08741_),
    .X(_08742_));
 sg13g2_o21ai_1 _31699_ (.B1(_08742_),
    .Y(_01406_),
    .A1(_10479_),
    .A2(net4035));
 sg13g2_nand2_1 _31700_ (.Y(_08743_),
    .A(net2328),
    .B(net3981));
 sg13g2_a21oi_1 _31701_ (.A1(_11509_),
    .A2(_11581_),
    .Y(_08744_),
    .B1(_11616_));
 sg13g2_or2_1 _31702_ (.X(_08745_),
    .B(_08744_),
    .A(_11557_));
 sg13g2_a21oi_1 _31703_ (.A1(_11557_),
    .A2(_08744_),
    .Y(_08746_),
    .B1(net3861));
 sg13g2_nor3_1 _31704_ (.A(_11567_),
    .B(_12745_),
    .C(_12748_),
    .Y(_08747_));
 sg13g2_nor2b_2 _31705_ (.A(_08747_),
    .B_N(_12478_),
    .Y(_08748_));
 sg13g2_nor2b_1 _31706_ (.A(_08748_),
    .B_N(_11557_),
    .Y(_08749_));
 sg13g2_xor2_1 _31707_ (.B(_08748_),
    .A(_11557_),
    .X(_08750_));
 sg13g2_nor2_1 _31708_ (.A(\u_inv.f_next[104] ),
    .B(net4708),
    .Y(_08751_));
 sg13g2_a21oi_1 _31709_ (.A1(net4708),
    .A2(_08750_),
    .Y(_08752_),
    .B1(_08751_));
 sg13g2_a221oi_1 _31710_ (.B2(net3861),
    .C1(net4448),
    .B1(_08752_),
    .A1(_08745_),
    .Y(_08753_),
    .A2(_08746_));
 sg13g2_o21ai_1 _31711_ (.B1(net4038),
    .Y(_08754_),
    .A1(net4623),
    .A2(net2289));
 sg13g2_o21ai_1 _31712_ (.B1(_08743_),
    .Y(_01407_),
    .A1(_08753_),
    .A2(_08754_));
 sg13g2_nand3_1 _31713_ (.B(_11627_),
    .C(_08745_),
    .A(_11558_),
    .Y(_08755_));
 sg13g2_a21oi_1 _31714_ (.A1(_11627_),
    .A2(_08745_),
    .Y(_08756_),
    .B1(_11558_));
 sg13g2_nor2_1 _31715_ (.A(net3687),
    .B(_08756_),
    .Y(_08757_));
 sg13g2_a21oi_1 _31716_ (.A1(\u_inv.f_next[104] ),
    .A2(net2595),
    .Y(_08758_),
    .B1(_08749_));
 sg13g2_xnor2_1 _31717_ (.Y(_08759_),
    .A(_11559_),
    .B(_08758_));
 sg13g2_o21ai_1 _31718_ (.B1(net3720),
    .Y(_08760_),
    .A1(\u_inv.f_next[105] ),
    .A2(net4707));
 sg13g2_a21o_1 _31719_ (.A2(_08759_),
    .A1(net4707),
    .B1(_08760_),
    .X(_08761_));
 sg13g2_a221oi_1 _31720_ (.B2(_08757_),
    .C1(net3982),
    .B1(_08755_),
    .A1(net4521),
    .Y(_08762_),
    .A2(net2443));
 sg13g2_a22oi_1 _31721_ (.Y(_01408_),
    .B1(_08761_),
    .B2(_08762_),
    .A2(net3982),
    .A1(_10477_));
 sg13g2_a21o_1 _31722_ (.A2(_10785_),
    .A1(net4957),
    .B1(_08756_),
    .X(_08763_));
 sg13g2_and2_1 _31723_ (.A(_11561_),
    .B(_08763_),
    .X(_08764_));
 sg13g2_nor2_1 _31724_ (.A(net3687),
    .B(_08764_),
    .Y(_08765_));
 sg13g2_o21ai_1 _31725_ (.B1(_08765_),
    .Y(_08766_),
    .A1(_11561_),
    .A2(_08763_));
 sg13g2_o21ai_1 _31726_ (.B1(_12523_),
    .Y(_08767_),
    .A1(_12498_),
    .A2(_08748_));
 sg13g2_nor2b_1 _31727_ (.A(_11561_),
    .B_N(_08767_),
    .Y(_08768_));
 sg13g2_xor2_1 _31728_ (.B(_08767_),
    .A(_11561_),
    .X(_08769_));
 sg13g2_nor2_1 _31729_ (.A(net3284),
    .B(net4707),
    .Y(_08770_));
 sg13g2_a21oi_1 _31730_ (.A1(net4707),
    .A2(_08769_),
    .Y(_08771_),
    .B1(_08770_));
 sg13g2_a221oi_1 _31731_ (.B2(_08771_),
    .C1(net3982),
    .B1(net3720),
    .A1(net4521),
    .Y(_08772_),
    .A2(net1998));
 sg13g2_a22oi_1 _31732_ (.Y(_01409_),
    .B1(_08766_),
    .B2(_08772_),
    .A2(net3982),
    .A1(_10476_));
 sg13g2_o21ai_1 _31733_ (.B1(_11560_),
    .Y(_08773_),
    .A1(_11625_),
    .A2(_08764_));
 sg13g2_or3_1 _31734_ (.A(_11560_),
    .B(_11625_),
    .C(_08764_),
    .X(_08774_));
 sg13g2_nand3_1 _31735_ (.B(_08773_),
    .C(_08774_),
    .A(net3699),
    .Y(_08775_));
 sg13g2_a21oi_1 _31736_ (.A1(\u_inv.f_next[106] ),
    .A2(\u_inv.f_reg[106] ),
    .Y(_08776_),
    .B1(_08768_));
 sg13g2_xnor2_1 _31737_ (.Y(_08777_),
    .A(_11560_),
    .B(_08776_));
 sg13g2_o21ai_1 _31738_ (.B1(net3720),
    .Y(_08778_),
    .A1(net2585),
    .A2(net4707));
 sg13g2_a21oi_1 _31739_ (.A1(net4707),
    .A2(_08777_),
    .Y(_08779_),
    .B1(_08778_));
 sg13g2_a21oi_1 _31740_ (.A1(net4521),
    .A2(net1951),
    .Y(_08780_),
    .B1(net3982));
 sg13g2_nor2b_1 _31741_ (.A(_08779_),
    .B_N(_08780_),
    .Y(_08781_));
 sg13g2_a22oi_1 _31742_ (.Y(_01410_),
    .B1(_08775_),
    .B2(_08781_),
    .A2(net3982),
    .A1(_10475_));
 sg13g2_a21o_2 _31743_ (.A2(_08767_),
    .A1(_12497_),
    .B1(_12526_),
    .X(_08782_));
 sg13g2_nor2b_1 _31744_ (.A(_11555_),
    .B_N(_08782_),
    .Y(_08783_));
 sg13g2_xnor2_1 _31745_ (.Y(_08784_),
    .A(_11555_),
    .B(_08782_));
 sg13g2_o21ai_1 _31746_ (.B1(net3720),
    .Y(_08785_),
    .A1(_10473_),
    .A2(net4706));
 sg13g2_a21oi_1 _31747_ (.A1(net4706),
    .A2(_08784_),
    .Y(_08786_),
    .B1(_08785_));
 sg13g2_o21ai_1 _31748_ (.B1(_11629_),
    .Y(_08787_),
    .A1(_11563_),
    .A2(_08745_));
 sg13g2_and2_1 _31749_ (.A(_11555_),
    .B(_08787_),
    .X(_08788_));
 sg13g2_xor2_1 _31750_ (.B(_08787_),
    .A(_11555_),
    .X(_08789_));
 sg13g2_o21ai_1 _31751_ (.B1(net4036),
    .Y(_08790_),
    .A1(net4624),
    .A2(net2085));
 sg13g2_nor2_1 _31752_ (.A(_08786_),
    .B(_08790_),
    .Y(_08791_));
 sg13g2_o21ai_1 _31753_ (.B1(_08791_),
    .Y(_08792_),
    .A1(net3687),
    .A2(_08789_));
 sg13g2_o21ai_1 _31754_ (.B1(_08792_),
    .Y(_01411_),
    .A1(_10474_),
    .A2(net4036));
 sg13g2_nand2_1 _31755_ (.Y(_08793_),
    .A(net2526),
    .B(net3861));
 sg13g2_a21oi_1 _31756_ (.A1(\u_inv.f_next[108] ),
    .A2(\u_inv.f_reg[108] ),
    .Y(_08794_),
    .B1(_08783_));
 sg13g2_xnor2_1 _31757_ (.Y(_08795_),
    .A(_11554_),
    .B(_08794_));
 sg13g2_a22oi_1 _31758_ (.Y(_08796_),
    .B1(_08795_),
    .B2(net4706),
    .A2(_08793_),
    .A1(net3735));
 sg13g2_o21ai_1 _31759_ (.B1(_11554_),
    .Y(_08797_),
    .A1(_11619_),
    .A2(_08788_));
 sg13g2_or3_1 _31760_ (.A(_11554_),
    .B(_11619_),
    .C(_08788_),
    .X(_08798_));
 sg13g2_nand2_1 _31761_ (.Y(_08799_),
    .A(_08797_),
    .B(_08798_));
 sg13g2_o21ai_1 _31762_ (.B1(net4386),
    .Y(_08800_),
    .A1(net3861),
    .A2(_08799_));
 sg13g2_a21oi_1 _31763_ (.A1(net4521),
    .A2(_10974_),
    .Y(_08801_),
    .B1(net3983));
 sg13g2_o21ai_1 _31764_ (.B1(_08801_),
    .Y(_08802_),
    .A1(_08796_),
    .A2(_08800_));
 sg13g2_o21ai_1 _31765_ (.B1(_08802_),
    .Y(_01412_),
    .A1(_10473_),
    .A2(net4036));
 sg13g2_a21oi_1 _31766_ (.A1(_11618_),
    .A2(_08797_),
    .Y(_08803_),
    .B1(_11552_));
 sg13g2_nand3_1 _31767_ (.B(_11618_),
    .C(_08797_),
    .A(_11552_),
    .Y(_08804_));
 sg13g2_nand2b_1 _31768_ (.Y(_08805_),
    .B(_08804_),
    .A_N(_08803_));
 sg13g2_o21ai_1 _31769_ (.B1(net4036),
    .Y(_08806_),
    .A1(net4628),
    .A2(net2117));
 sg13g2_a21oi_1 _31770_ (.A1(_12494_),
    .A2(_08782_),
    .Y(_08807_),
    .B1(_12530_));
 sg13g2_nand2b_1 _31771_ (.Y(_08808_),
    .B(_08807_),
    .A_N(_11552_));
 sg13g2_nand2b_1 _31772_ (.Y(_08809_),
    .B(_11552_),
    .A_N(_08807_));
 sg13g2_nand3_1 _31773_ (.B(_08808_),
    .C(_08809_),
    .A(net4706),
    .Y(_08810_));
 sg13g2_a21oi_1 _31774_ (.A1(net2100),
    .A2(net4593),
    .Y(_08811_),
    .B1(net3709));
 sg13g2_a221oi_1 _31775_ (.B2(_08811_),
    .C1(_08806_),
    .B1(_08810_),
    .A1(net3699),
    .Y(_08812_),
    .A2(_08805_));
 sg13g2_a21o_1 _31776_ (.A2(net3983),
    .A1(net2526),
    .B1(_08812_),
    .X(_01413_));
 sg13g2_nand2_1 _31777_ (.Y(_08813_),
    .A(net2100),
    .B(net3983));
 sg13g2_a21oi_1 _31778_ (.A1(\u_inv.f_next[110] ),
    .A2(_10780_),
    .Y(_08814_),
    .B1(_08803_));
 sg13g2_xnor2_1 _31779_ (.Y(_08815_),
    .A(_11550_),
    .B(_08814_));
 sg13g2_and2_1 _31780_ (.A(_11551_),
    .B(_08809_),
    .X(_08816_));
 sg13g2_xor2_1 _31781_ (.B(_08816_),
    .A(_11550_),
    .X(_08817_));
 sg13g2_nand2_1 _31782_ (.Y(_08818_),
    .A(\u_inv.f_next[111] ),
    .B(net3861));
 sg13g2_a22oi_1 _31783_ (.Y(_08819_),
    .B1(_08818_),
    .B2(net3735),
    .A2(_08817_),
    .A1(net4706));
 sg13g2_o21ai_1 _31784_ (.B1(net4385),
    .Y(_08820_),
    .A1(net3862),
    .A2(_08815_));
 sg13g2_nor2_1 _31785_ (.A(_08819_),
    .B(_08820_),
    .Y(_08821_));
 sg13g2_o21ai_1 _31786_ (.B1(net4037),
    .Y(_08822_),
    .A1(net4628),
    .A2(\u_inv.input_reg[110] ));
 sg13g2_o21ai_1 _31787_ (.B1(_08813_),
    .Y(_01414_),
    .A1(_08821_),
    .A2(_08822_));
 sg13g2_o21ai_1 _31788_ (.B1(_12531_),
    .Y(_08823_),
    .A1(_12499_),
    .A2(_08748_));
 sg13g2_xor2_1 _31789_ (.B(_08823_),
    .A(_11534_),
    .X(_08824_));
 sg13g2_o21ai_1 _31790_ (.B1(net3718),
    .Y(_08825_),
    .A1(_10469_),
    .A2(net4715));
 sg13g2_a21oi_1 _31791_ (.A1(net4715),
    .A2(_08824_),
    .Y(_08826_),
    .B1(_08825_));
 sg13g2_a21oi_2 _31792_ (.B1(_11632_),
    .Y(_08827_),
    .A2(_11582_),
    .A1(_11509_));
 sg13g2_or2_1 _31793_ (.X(_08828_),
    .B(_08827_),
    .A(_11534_));
 sg13g2_xor2_1 _31794_ (.B(_08827_),
    .A(_11534_),
    .X(_08829_));
 sg13g2_o21ai_1 _31795_ (.B1(net4044),
    .Y(_08830_),
    .A1(net4628),
    .A2(net2621));
 sg13g2_nor2_1 _31796_ (.A(_08826_),
    .B(_08830_),
    .Y(_08831_));
 sg13g2_o21ai_1 _31797_ (.B1(_08831_),
    .Y(_08832_),
    .A1(net3685),
    .A2(_08829_));
 sg13g2_o21ai_1 _31798_ (.B1(_08832_),
    .Y(_01415_),
    .A1(_10470_),
    .A2(net4036));
 sg13g2_nand2_1 _31799_ (.Y(_08833_),
    .A(net1527),
    .B(net3992));
 sg13g2_nand2_1 _31800_ (.Y(_08834_),
    .A(\u_inv.f_next[113] ),
    .B(net3869));
 sg13g2_a21oi_1 _31801_ (.A1(_11534_),
    .A2(_08823_),
    .Y(_08835_),
    .B1(_11533_));
 sg13g2_xor2_1 _31802_ (.B(_08835_),
    .A(_11535_),
    .X(_08836_));
 sg13g2_a22oi_1 _31803_ (.Y(_08837_),
    .B1(_08836_),
    .B2(net4716),
    .A2(_08834_),
    .A1(net3733));
 sg13g2_a21oi_1 _31804_ (.A1(_11590_),
    .A2(_08828_),
    .Y(_08838_),
    .B1(_11535_));
 sg13g2_and3_1 _31805_ (.X(_08839_),
    .A(_11535_),
    .B(_11590_),
    .C(_08828_));
 sg13g2_o21ai_1 _31806_ (.B1(net4385),
    .Y(_08840_),
    .A1(_08838_),
    .A2(_08839_));
 sg13g2_a21oi_1 _31807_ (.A1(net3707),
    .A2(_08840_),
    .Y(_08841_),
    .B1(_08837_));
 sg13g2_o21ai_1 _31808_ (.B1(net4045),
    .Y(_08842_),
    .A1(net4628),
    .A2(\u_inv.input_reg[112] ));
 sg13g2_o21ai_1 _31809_ (.B1(_08833_),
    .Y(_01416_),
    .A1(_08841_),
    .A2(_08842_));
 sg13g2_nor2_1 _31810_ (.A(_11589_),
    .B(_08838_),
    .Y(_08843_));
 sg13g2_xnor2_1 _31811_ (.Y(_08844_),
    .A(_11532_),
    .B(_08843_));
 sg13g2_o21ai_1 _31812_ (.B1(net4045),
    .Y(_08845_),
    .A1(net4629),
    .A2(net1793));
 sg13g2_a21oi_2 _31813_ (.B1(_12501_),
    .Y(_08846_),
    .A2(_08823_),
    .A1(_12488_));
 sg13g2_a21oi_1 _31814_ (.A1(_11531_),
    .A2(_08846_),
    .Y(_08847_),
    .B1(net4599));
 sg13g2_o21ai_1 _31815_ (.B1(_08847_),
    .Y(_08848_),
    .A1(_11531_),
    .A2(_08846_));
 sg13g2_a21oi_1 _31816_ (.A1(net2404),
    .A2(net4599),
    .Y(_08849_),
    .B1(net3707));
 sg13g2_a221oi_1 _31817_ (.B2(_08849_),
    .C1(_08845_),
    .B1(_08848_),
    .A1(net3698),
    .Y(_08850_),
    .A2(_08844_));
 sg13g2_a21o_1 _31818_ (.A2(net3992),
    .A1(net2661),
    .B1(_08850_),
    .X(_01417_));
 sg13g2_o21ai_1 _31819_ (.B1(_11588_),
    .Y(_08851_),
    .A1(_11532_),
    .A2(_08843_));
 sg13g2_xor2_1 _31820_ (.B(_08851_),
    .A(_11529_),
    .X(_08852_));
 sg13g2_nand2_1 _31821_ (.Y(_08853_),
    .A(net2997),
    .B(net3870));
 sg13g2_o21ai_1 _31822_ (.B1(_11530_),
    .Y(_08854_),
    .A1(_11531_),
    .A2(_08846_));
 sg13g2_xnor2_1 _31823_ (.Y(_08855_),
    .A(_11529_),
    .B(_08854_));
 sg13g2_a22oi_1 _31824_ (.Y(_08856_),
    .B1(_08855_),
    .B2(net4716),
    .A2(_08853_),
    .A1(net3733));
 sg13g2_o21ai_1 _31825_ (.B1(net4385),
    .Y(_08857_),
    .A1(net3872),
    .A2(_08852_));
 sg13g2_a21oi_1 _31826_ (.A1(net4519),
    .A2(_10975_),
    .Y(_08858_),
    .B1(net3991));
 sg13g2_o21ai_1 _31827_ (.B1(_08858_),
    .Y(_08859_),
    .A1(_08856_),
    .A2(_08857_));
 sg13g2_o21ai_1 _31828_ (.B1(_08859_),
    .Y(_01418_),
    .A1(_10467_),
    .A2(net4045));
 sg13g2_o21ai_1 _31829_ (.B1(_12504_),
    .Y(_08860_),
    .A1(_12487_),
    .A2(_08846_));
 sg13g2_a21oi_1 _31830_ (.A1(_11543_),
    .A2(_08860_),
    .Y(_08861_),
    .B1(net4597));
 sg13g2_o21ai_1 _31831_ (.B1(_08861_),
    .Y(_08862_),
    .A1(_11543_),
    .A2(_08860_));
 sg13g2_a21oi_1 _31832_ (.A1(net2223),
    .A2(net4598),
    .Y(_08863_),
    .B1(net3707));
 sg13g2_o21ai_1 _31833_ (.B1(_11594_),
    .Y(_08864_),
    .A1(_11536_),
    .A2(_08827_));
 sg13g2_and2_1 _31834_ (.A(_11544_),
    .B(_08864_),
    .X(_08865_));
 sg13g2_xnor2_1 _31835_ (.Y(_08866_),
    .A(_11544_),
    .B(_08864_));
 sg13g2_o21ai_1 _31836_ (.B1(net4049),
    .Y(_08867_),
    .A1(net4631),
    .A2(net2286));
 sg13g2_a221oi_1 _31837_ (.B2(net3698),
    .C1(_08867_),
    .B1(_08866_),
    .A1(_08862_),
    .Y(_08868_),
    .A2(_08863_));
 sg13g2_a21o_1 _31838_ (.A2(net3993),
    .A1(net2997),
    .B1(_08868_),
    .X(_01419_));
 sg13g2_nand2_1 _31839_ (.Y(_08869_),
    .A(net2989),
    .B(net3871));
 sg13g2_a21oi_1 _31840_ (.A1(_11543_),
    .A2(_08860_),
    .Y(_08870_),
    .B1(_11542_));
 sg13g2_xnor2_1 _31841_ (.Y(_08871_),
    .A(_11541_),
    .B(_08870_));
 sg13g2_a22oi_1 _31842_ (.Y(_08872_),
    .B1(_08871_),
    .B2(net4720),
    .A2(_08869_),
    .A1(net3732));
 sg13g2_o21ai_1 _31843_ (.B1(_11541_),
    .Y(_08873_),
    .A1(_11587_),
    .A2(_08865_));
 sg13g2_or3_1 _31844_ (.A(_11541_),
    .B(_11587_),
    .C(_08865_),
    .X(_08874_));
 sg13g2_nand2_1 _31845_ (.Y(_08875_),
    .A(_08873_),
    .B(_08874_));
 sg13g2_o21ai_1 _31846_ (.B1(net4384),
    .Y(_08876_),
    .A1(net3871),
    .A2(_08875_));
 sg13g2_a21oi_1 _31847_ (.A1(net4519),
    .A2(_10976_),
    .Y(_08877_),
    .B1(net3993));
 sg13g2_o21ai_1 _31848_ (.B1(_08877_),
    .Y(_08878_),
    .A1(_08872_),
    .A2(_08876_));
 sg13g2_o21ai_1 _31849_ (.B1(_08878_),
    .Y(_01420_),
    .A1(_10465_),
    .A2(net4049));
 sg13g2_a21oi_1 _31850_ (.A1(_12486_),
    .A2(_08860_),
    .Y(_08879_),
    .B1(_12509_));
 sg13g2_a21oi_1 _31851_ (.A1(_11539_),
    .A2(_08879_),
    .Y(_08880_),
    .B1(net4598));
 sg13g2_o21ai_1 _31852_ (.B1(_08880_),
    .Y(_08881_),
    .A1(_11539_),
    .A2(_08879_));
 sg13g2_a21oi_1 _31853_ (.A1(\u_inv.f_next[118] ),
    .A2(net4598),
    .Y(_08882_),
    .B1(net3707));
 sg13g2_nand2_1 _31854_ (.Y(_08883_),
    .A(_11586_),
    .B(_08873_));
 sg13g2_xnor2_1 _31855_ (.Y(_08884_),
    .A(_11539_),
    .B(_08883_));
 sg13g2_o21ai_1 _31856_ (.B1(net4049),
    .Y(_08885_),
    .A1(net4631),
    .A2(net2179));
 sg13g2_a221oi_1 _31857_ (.B2(net3698),
    .C1(_08885_),
    .B1(_08884_),
    .A1(_08881_),
    .Y(_08886_),
    .A2(_08882_));
 sg13g2_a21o_1 _31858_ (.A2(net3993),
    .A1(net2989),
    .B1(_08886_),
    .X(_01421_));
 sg13g2_nand2_1 _31859_ (.Y(_08887_),
    .A(net2767),
    .B(net3871));
 sg13g2_o21ai_1 _31860_ (.B1(_11538_),
    .Y(_08888_),
    .A1(_11539_),
    .A2(_08879_));
 sg13g2_xor2_1 _31861_ (.B(_08888_),
    .A(_11537_),
    .X(_08889_));
 sg13g2_a22oi_1 _31862_ (.Y(_08890_),
    .B1(_08889_),
    .B2(net4720),
    .A2(_08887_),
    .A1(net3732));
 sg13g2_a21oi_1 _31863_ (.A1(_11539_),
    .A2(_08883_),
    .Y(_08891_),
    .B1(_11598_));
 sg13g2_xor2_1 _31864_ (.B(_08891_),
    .A(_11537_),
    .X(_08892_));
 sg13g2_o21ai_1 _31865_ (.B1(net4384),
    .Y(_08893_),
    .A1(net3871),
    .A2(_08892_));
 sg13g2_a21oi_1 _31866_ (.A1(net4520),
    .A2(_10977_),
    .Y(_08894_),
    .B1(net3994));
 sg13g2_o21ai_1 _31867_ (.B1(_08894_),
    .Y(_08895_),
    .A1(_08890_),
    .A2(_08893_));
 sg13g2_o21ai_1 _31868_ (.B1(_08895_),
    .Y(_01422_),
    .A1(_10463_),
    .A2(net4049));
 sg13g2_a21oi_1 _31869_ (.A1(_12490_),
    .A2(_08823_),
    .Y(_08896_),
    .B1(_12511_));
 sg13g2_nand2_1 _31870_ (.Y(_08897_),
    .A(_11514_),
    .B(_08896_));
 sg13g2_nor2_1 _31871_ (.A(_11514_),
    .B(_08896_),
    .Y(_08898_));
 sg13g2_nand3b_1 _31872_ (.B(net4721),
    .C(_08897_),
    .Y(_08899_),
    .A_N(_08898_));
 sg13g2_a21oi_1 _31873_ (.A1(\u_inv.f_next[120] ),
    .A2(net4598),
    .Y(_08900_),
    .B1(net3707));
 sg13g2_o21ai_1 _31874_ (.B1(_11600_),
    .Y(_08901_),
    .A1(_11546_),
    .A2(_08827_));
 sg13g2_xnor2_1 _31875_ (.Y(_08902_),
    .A(_11514_),
    .B(_08901_));
 sg13g2_o21ai_1 _31876_ (.B1(net4049),
    .Y(_08903_),
    .A1(net4630),
    .A2(net2451));
 sg13g2_a221oi_1 _31877_ (.B2(net3698),
    .C1(_08903_),
    .B1(_08902_),
    .A1(_08899_),
    .Y(_08904_),
    .A2(_08900_));
 sg13g2_a21o_1 _31878_ (.A2(net3993),
    .A1(net2767),
    .B1(_08904_),
    .X(_01423_));
 sg13g2_a21oi_1 _31879_ (.A1(\u_inv.f_next[120] ),
    .A2(\u_inv.f_reg[120] ),
    .Y(_08905_),
    .B1(_08898_));
 sg13g2_o21ai_1 _31880_ (.B1(net4721),
    .Y(_08906_),
    .A1(_11517_),
    .A2(_08905_));
 sg13g2_a21oi_1 _31881_ (.A1(_11517_),
    .A2(_08905_),
    .Y(_08907_),
    .B1(_08906_));
 sg13g2_a21oi_1 _31882_ (.A1(_10460_),
    .A2(net4597),
    .Y(_08908_),
    .B1(_08907_));
 sg13g2_a21oi_1 _31883_ (.A1(_11514_),
    .A2(_08901_),
    .Y(_08909_),
    .B1(_11636_));
 sg13g2_a21oi_1 _31884_ (.A1(_11517_),
    .A2(_08909_),
    .Y(_08910_),
    .B1(net3685));
 sg13g2_o21ai_1 _31885_ (.B1(_08910_),
    .Y(_08911_),
    .A1(_11517_),
    .A2(_08909_));
 sg13g2_a221oi_1 _31886_ (.B2(_08908_),
    .C1(net3994),
    .B1(net3719),
    .A1(net4519),
    .Y(_08912_),
    .A2(net2252));
 sg13g2_a22oi_1 _31887_ (.Y(_01424_),
    .B1(_08911_),
    .B2(_08912_),
    .A2(net3994),
    .A1(_10461_));
 sg13g2_a21oi_1 _31888_ (.A1(_11515_),
    .A2(_08905_),
    .Y(_08913_),
    .B1(_11516_));
 sg13g2_nor2b_1 _31889_ (.A(_11512_),
    .B_N(_08913_),
    .Y(_08914_));
 sg13g2_xnor2_1 _31890_ (.Y(_08915_),
    .A(_11512_),
    .B(_08913_));
 sg13g2_nand2_1 _31891_ (.Y(_08916_),
    .A(net4721),
    .B(_08915_));
 sg13g2_a21oi_1 _31892_ (.A1(net2164),
    .A2(net4597),
    .Y(_08917_),
    .B1(net3707));
 sg13g2_o21ai_1 _31893_ (.B1(_11635_),
    .Y(_08918_),
    .A1(_11517_),
    .A2(_08909_));
 sg13g2_xnor2_1 _31894_ (.Y(_08919_),
    .A(_11512_),
    .B(_08918_));
 sg13g2_a221oi_1 _31895_ (.B2(net3698),
    .C1(net3994),
    .B1(_08919_),
    .A1(_08916_),
    .Y(_08920_),
    .A2(_08917_));
 sg13g2_o21ai_1 _31896_ (.B1(_08920_),
    .Y(_08921_),
    .A1(net4631),
    .A2(net2667));
 sg13g2_o21ai_1 _31897_ (.B1(_08921_),
    .Y(_01425_),
    .A1(_10460_),
    .A2(net4050));
 sg13g2_nand2_1 _31898_ (.Y(_08922_),
    .A(net2164),
    .B(net3994));
 sg13g2_a21oi_1 _31899_ (.A1(net2164),
    .A2(\u_inv.f_reg[122] ),
    .Y(_08923_),
    .B1(_08914_));
 sg13g2_xnor2_1 _31900_ (.Y(_08924_),
    .A(_11510_),
    .B(_08923_));
 sg13g2_o21ai_1 _31901_ (.B1(net3718),
    .Y(_08925_),
    .A1(_10458_),
    .A2(net4721));
 sg13g2_a21oi_1 _31902_ (.A1(net4721),
    .A2(_08924_),
    .Y(_08926_),
    .B1(_08925_));
 sg13g2_a21oi_1 _31903_ (.A1(_11512_),
    .A2(_08918_),
    .Y(_08927_),
    .B1(_11634_));
 sg13g2_a21oi_1 _31904_ (.A1(_11511_),
    .A2(_08927_),
    .Y(_08928_),
    .B1(net3685));
 sg13g2_o21ai_1 _31905_ (.B1(_08928_),
    .Y(_08929_),
    .A1(_11511_),
    .A2(_08927_));
 sg13g2_o21ai_1 _31906_ (.B1(net4049),
    .Y(_08930_),
    .A1(net4631),
    .A2(\u_inv.input_reg[122] ));
 sg13g2_nand2b_1 _31907_ (.Y(_08931_),
    .B(_08929_),
    .A_N(_08930_));
 sg13g2_o21ai_1 _31908_ (.B1(_08922_),
    .Y(_01426_),
    .A1(_08926_),
    .A2(_08931_));
 sg13g2_nand2b_1 _31909_ (.Y(_08932_),
    .B(_08898_),
    .A_N(_12483_));
 sg13g2_nand2_2 _31910_ (.Y(_08933_),
    .A(_12515_),
    .B(_08932_));
 sg13g2_xor2_1 _31911_ (.B(_08933_),
    .A(_11526_),
    .X(_08934_));
 sg13g2_o21ai_1 _31912_ (.B1(net3718),
    .Y(_08935_),
    .A1(_10457_),
    .A2(net4720));
 sg13g2_a21oi_1 _31913_ (.A1(net4720),
    .A2(_08934_),
    .Y(_08936_),
    .B1(_08935_));
 sg13g2_a21oi_1 _31914_ (.A1(_11519_),
    .A2(_08901_),
    .Y(_08937_),
    .B1(_11640_));
 sg13g2_or2_1 _31915_ (.X(_08938_),
    .B(_08937_),
    .A(_11526_));
 sg13g2_xor2_1 _31916_ (.B(_08937_),
    .A(_11526_),
    .X(_08939_));
 sg13g2_o21ai_1 _31917_ (.B1(net4048),
    .Y(_08940_),
    .A1(net4630),
    .A2(net1904));
 sg13g2_nor2_1 _31918_ (.A(_08936_),
    .B(_08940_),
    .Y(_08941_));
 sg13g2_o21ai_1 _31919_ (.B1(_08941_),
    .Y(_08942_),
    .A1(net3686),
    .A2(_08939_));
 sg13g2_o21ai_1 _31920_ (.B1(_08942_),
    .Y(_01427_),
    .A1(_10458_),
    .A2(net4050));
 sg13g2_nand2_1 _31921_ (.Y(_08943_),
    .A(net1558),
    .B(net3993));
 sg13g2_nand2_1 _31922_ (.Y(_08944_),
    .A(\u_inv.f_next[125] ),
    .B(net3871));
 sg13g2_a21oi_1 _31923_ (.A1(_11526_),
    .A2(_08933_),
    .Y(_08945_),
    .B1(_11525_));
 sg13g2_xor2_1 _31924_ (.B(_08945_),
    .A(_11524_),
    .X(_08946_));
 sg13g2_a22oi_1 _31925_ (.Y(_08947_),
    .B1(_08946_),
    .B2(net4720),
    .A2(_08944_),
    .A1(net3732));
 sg13g2_a21oi_1 _31926_ (.A1(_11641_),
    .A2(_08938_),
    .Y(_08948_),
    .B1(_11524_));
 sg13g2_and3_1 _31927_ (.X(_08949_),
    .A(_11524_),
    .B(_11641_),
    .C(_08938_));
 sg13g2_o21ai_1 _31928_ (.B1(net4385),
    .Y(_08950_),
    .A1(_08948_),
    .A2(_08949_));
 sg13g2_a21oi_1 _31929_ (.A1(net3707),
    .A2(_08950_),
    .Y(_08951_),
    .B1(_08947_));
 sg13g2_o21ai_1 _31930_ (.B1(net4049),
    .Y(_08952_),
    .A1(net4631),
    .A2(\u_inv.input_reg[124] ));
 sg13g2_o21ai_1 _31931_ (.B1(_08943_),
    .Y(_01428_),
    .A1(_08951_),
    .A2(_08952_));
 sg13g2_o21ai_1 _31932_ (.B1(_11522_),
    .Y(_08953_),
    .A1(_11642_),
    .A2(_08948_));
 sg13g2_nor3_1 _31933_ (.A(_11522_),
    .B(_11642_),
    .C(_08948_),
    .Y(_08954_));
 sg13g2_nor2_1 _31934_ (.A(net3686),
    .B(_08954_),
    .Y(_08955_));
 sg13g2_a21oi_1 _31935_ (.A1(_12480_),
    .A2(_08933_),
    .Y(_08956_),
    .B1(_12518_));
 sg13g2_xnor2_1 _31936_ (.Y(_08957_),
    .A(_11522_),
    .B(_08956_));
 sg13g2_a21oi_1 _31937_ (.A1(net4720),
    .A2(_08957_),
    .Y(_08958_),
    .B1(net3707));
 sg13g2_o21ai_1 _31938_ (.B1(_08958_),
    .Y(_08959_),
    .A1(net2821),
    .A2(net4720));
 sg13g2_a221oi_1 _31939_ (.B2(_08955_),
    .C1(net3993),
    .B1(_08953_),
    .A1(net4519),
    .Y(_08960_),
    .A2(net2079));
 sg13g2_a22oi_1 _31940_ (.Y(_01429_),
    .B1(_08959_),
    .B2(_08960_),
    .A2(net3993),
    .A1(_10456_));
 sg13g2_nand2_1 _31941_ (.Y(_08961_),
    .A(net2545),
    .B(net3871));
 sg13g2_o21ai_1 _31942_ (.B1(_11521_),
    .Y(_08962_),
    .A1(_11522_),
    .A2(_08956_));
 sg13g2_xor2_1 _31943_ (.B(_08962_),
    .A(_11520_),
    .X(_08963_));
 sg13g2_a22oi_1 _31944_ (.Y(_08964_),
    .B1(_08963_),
    .B2(net4720),
    .A2(_08961_),
    .A1(net3733));
 sg13g2_nand2b_1 _31945_ (.Y(_08965_),
    .B(_08953_),
    .A_N(_11645_));
 sg13g2_xnor2_1 _31946_ (.Y(_08966_),
    .A(_11520_),
    .B(_08965_));
 sg13g2_o21ai_1 _31947_ (.B1(net4384),
    .Y(_08967_),
    .A1(net3871),
    .A2(_08966_));
 sg13g2_a21oi_1 _31948_ (.A1(net4519),
    .A2(_10978_),
    .Y(_08968_),
    .B1(net3993));
 sg13g2_o21ai_1 _31949_ (.B1(_08968_),
    .Y(_08969_),
    .A1(_08964_),
    .A2(_08967_));
 sg13g2_o21ai_1 _31950_ (.B1(_08969_),
    .Y(_01430_),
    .A1(_10455_),
    .A2(net4049));
 sg13g2_nor3_1 _31951_ (.A(_11585_),
    .B(_11649_),
    .C(_11724_),
    .Y(_08970_));
 sg13g2_o21ai_1 _31952_ (.B1(_11724_),
    .Y(_08971_),
    .A1(_11585_),
    .A2(_11649_));
 sg13g2_nand3b_1 _31953_ (.B(_08971_),
    .C(net3698),
    .Y(_08972_),
    .A_N(_08970_));
 sg13g2_a21oi_1 _31954_ (.A1(net4519),
    .A2(net2323),
    .Y(_08973_),
    .B1(net3992));
 sg13g2_xnor2_1 _31955_ (.Y(_08974_),
    .A(_11724_),
    .B(_12750_));
 sg13g2_o21ai_1 _31956_ (.B1(net3718),
    .Y(_08975_),
    .A1(net2561),
    .A2(net4716));
 sg13g2_a21oi_1 _31957_ (.A1(net4716),
    .A2(_08974_),
    .Y(_08976_),
    .B1(_08975_));
 sg13g2_nor2b_1 _31958_ (.A(_08976_),
    .B_N(_08973_),
    .Y(_08977_));
 sg13g2_a22oi_1 _31959_ (.Y(_01431_),
    .B1(_08972_),
    .B2(_08977_),
    .A2(net3992),
    .A1(_10454_));
 sg13g2_nand2_1 _31960_ (.Y(_08978_),
    .A(net2561),
    .B(net3992));
 sg13g2_nand2_1 _31961_ (.Y(_08979_),
    .A(_11841_),
    .B(_08971_));
 sg13g2_and2_1 _31962_ (.A(_11725_),
    .B(_08979_),
    .X(_08980_));
 sg13g2_o21ai_1 _31963_ (.B1(net3820),
    .Y(_08981_),
    .A1(_11725_),
    .A2(_08979_));
 sg13g2_nor2_1 _31964_ (.A(_08980_),
    .B(_08981_),
    .Y(_08982_));
 sg13g2_nand2_1 _31965_ (.Y(_08983_),
    .A(net1878),
    .B(net3870));
 sg13g2_o21ai_1 _31966_ (.B1(_11723_),
    .Y(_08984_),
    .A1(_11724_),
    .A2(_12750_));
 sg13g2_xor2_1 _31967_ (.B(_08984_),
    .A(_11725_),
    .X(_08985_));
 sg13g2_a22oi_1 _31968_ (.Y(_08986_),
    .B1(_08985_),
    .B2(net4719),
    .A2(_08983_),
    .A1(net3732));
 sg13g2_nor3_1 _31969_ (.A(net4447),
    .B(_08982_),
    .C(_08986_),
    .Y(_08987_));
 sg13g2_o21ai_1 _31970_ (.B1(net4046),
    .Y(_08988_),
    .A1(net4630),
    .A2(net2020));
 sg13g2_o21ai_1 _31971_ (.B1(_08978_),
    .Y(_01432_),
    .A1(_08987_),
    .A2(_08988_));
 sg13g2_nand2_1 _31972_ (.Y(_08989_),
    .A(net1878),
    .B(net3992));
 sg13g2_nor3_1 _31973_ (.A(_11722_),
    .B(_11840_),
    .C(_08980_),
    .Y(_08990_));
 sg13g2_o21ai_1 _31974_ (.B1(_11722_),
    .Y(_08991_),
    .A1(_11840_),
    .A2(_08980_));
 sg13g2_nand2_1 _31975_ (.Y(_08992_),
    .A(net3820),
    .B(_08991_));
 sg13g2_nor2_1 _31976_ (.A(_08990_),
    .B(_08992_),
    .Y(_08993_));
 sg13g2_nor3_1 _31977_ (.A(_11724_),
    .B(_11725_),
    .C(_12750_),
    .Y(_08994_));
 sg13g2_nor2_1 _31978_ (.A(_12408_),
    .B(_08994_),
    .Y(_08995_));
 sg13g2_nor2_1 _31979_ (.A(_11722_),
    .B(_08995_),
    .Y(_08996_));
 sg13g2_xnor2_1 _31980_ (.Y(_08997_),
    .A(_11722_),
    .B(_08995_));
 sg13g2_o21ai_1 _31981_ (.B1(net3870),
    .Y(_08998_),
    .A1(\u_inv.f_next[130] ),
    .A2(net4719));
 sg13g2_a21oi_1 _31982_ (.A1(net4719),
    .A2(_08997_),
    .Y(_08999_),
    .B1(_08998_));
 sg13g2_nor3_1 _31983_ (.A(net4446),
    .B(_08993_),
    .C(_08999_),
    .Y(_09000_));
 sg13g2_o21ai_1 _31984_ (.B1(net4046),
    .Y(_09001_),
    .A1(net4625),
    .A2(net1853));
 sg13g2_o21ai_1 _31985_ (.B1(_08989_),
    .Y(_01433_),
    .A1(_09000_),
    .A2(_09001_));
 sg13g2_nand2_1 _31986_ (.Y(_09002_),
    .A(_11839_),
    .B(_08991_));
 sg13g2_xnor2_1 _31987_ (.Y(_09003_),
    .A(_11719_),
    .B(_09002_));
 sg13g2_nand2_1 _31988_ (.Y(_09004_),
    .A(\u_inv.f_next[131] ),
    .B(net3866));
 sg13g2_a21oi_1 _31989_ (.A1(\u_inv.f_next[130] ),
    .A2(\u_inv.f_reg[130] ),
    .Y(_09005_),
    .B1(_08996_));
 sg13g2_xnor2_1 _31990_ (.Y(_09006_),
    .A(_11720_),
    .B(_09005_));
 sg13g2_a22oi_1 _31991_ (.Y(_09007_),
    .B1(_09006_),
    .B2(net4719),
    .A2(_09004_),
    .A1(net3732));
 sg13g2_a21oi_1 _31992_ (.A1(net3821),
    .A2(_09003_),
    .Y(_09008_),
    .B1(_09007_));
 sg13g2_o21ai_1 _31993_ (.B1(net4043),
    .Y(_09009_),
    .A1(net4625),
    .A2(net1817));
 sg13g2_a21o_1 _31994_ (.A2(_09008_),
    .A1(net4384),
    .B1(_09009_),
    .X(_09010_));
 sg13g2_o21ai_1 _31995_ (.B1(_09010_),
    .Y(_01434_),
    .A1(_10451_),
    .A2(net4043));
 sg13g2_nand2_1 _31996_ (.Y(_09011_),
    .A(net2720),
    .B(net3988));
 sg13g2_o21ai_1 _31997_ (.B1(_11845_),
    .Y(_09012_),
    .A1(_11650_),
    .A2(_11726_));
 sg13g2_and2_1 _31998_ (.A(_11715_),
    .B(_09012_),
    .X(_09013_));
 sg13g2_o21ai_1 _31999_ (.B1(net3818),
    .Y(_09014_),
    .A1(_11715_),
    .A2(_09012_));
 sg13g2_nor2_1 _32000_ (.A(_09013_),
    .B(_09014_),
    .Y(_09015_));
 sg13g2_o21ai_1 _32001_ (.B1(_12410_),
    .Y(_09016_),
    .A1(_12750_),
    .A2(_12752_));
 sg13g2_nor2b_1 _32002_ (.A(_11715_),
    .B_N(_09016_),
    .Y(_09017_));
 sg13g2_xor2_1 _32003_ (.B(_09016_),
    .A(_11715_),
    .X(_09018_));
 sg13g2_o21ai_1 _32004_ (.B1(net3865),
    .Y(_09019_),
    .A1(net2097),
    .A2(net4709));
 sg13g2_a21oi_1 _32005_ (.A1(net4709),
    .A2(_09018_),
    .Y(_09020_),
    .B1(_09019_));
 sg13g2_nor3_1 _32006_ (.A(net4446),
    .B(_09015_),
    .C(_09020_),
    .Y(_09021_));
 sg13g2_o21ai_1 _32007_ (.B1(net4040),
    .Y(_09022_),
    .A1(net4625),
    .A2(net2054));
 sg13g2_o21ai_1 _32008_ (.B1(_09011_),
    .Y(_01435_),
    .A1(_09021_),
    .A2(_09022_));
 sg13g2_nand2_1 _32009_ (.Y(_09023_),
    .A(net2097),
    .B(net3986));
 sg13g2_nor2_1 _32010_ (.A(_11847_),
    .B(_09013_),
    .Y(_09024_));
 sg13g2_nor2_1 _32011_ (.A(_11716_),
    .B(_09024_),
    .Y(_09025_));
 sg13g2_a21oi_1 _32012_ (.A1(_11716_),
    .A2(_09024_),
    .Y(_09026_),
    .B1(net3865));
 sg13g2_nor2b_1 _32013_ (.A(_09025_),
    .B_N(_09026_),
    .Y(_09027_));
 sg13g2_nand2_1 _32014_ (.Y(_09028_),
    .A(\u_inv.f_next[133] ),
    .B(net3865));
 sg13g2_a21oi_1 _32015_ (.A1(\u_inv.f_next[132] ),
    .A2(\u_inv.f_reg[132] ),
    .Y(_09029_),
    .B1(_09017_));
 sg13g2_xnor2_1 _32016_ (.Y(_09030_),
    .A(_11717_),
    .B(_09029_));
 sg13g2_a22oi_1 _32017_ (.Y(_09031_),
    .B1(_09030_),
    .B2(net4709),
    .A2(_09028_),
    .A1(net3734));
 sg13g2_nor3_1 _32018_ (.A(net4446),
    .B(_09027_),
    .C(_09031_),
    .Y(_09032_));
 sg13g2_o21ai_1 _32019_ (.B1(net4039),
    .Y(_09033_),
    .A1(net4626),
    .A2(net2008));
 sg13g2_o21ai_1 _32020_ (.B1(_09023_),
    .Y(_01436_),
    .A1(_09032_),
    .A2(_09033_));
 sg13g2_nand2_1 _32021_ (.Y(_09034_),
    .A(net2400),
    .B(net3986));
 sg13g2_nor2_1 _32022_ (.A(_11846_),
    .B(_09025_),
    .Y(_09035_));
 sg13g2_nor2_1 _32023_ (.A(_11713_),
    .B(_09035_),
    .Y(_09036_));
 sg13g2_a21oi_1 _32024_ (.A1(_11713_),
    .A2(_09035_),
    .Y(_09037_),
    .B1(net3865));
 sg13g2_nor2b_1 _32025_ (.A(_09036_),
    .B_N(_09037_),
    .Y(_09038_));
 sg13g2_a21oi_1 _32026_ (.A1(_12403_),
    .A2(_09016_),
    .Y(_09039_),
    .B1(_12400_));
 sg13g2_xnor2_1 _32027_ (.Y(_09040_),
    .A(_11714_),
    .B(_09039_));
 sg13g2_o21ai_1 _32028_ (.B1(net3865),
    .Y(_09041_),
    .A1(\u_inv.f_next[134] ),
    .A2(net4709));
 sg13g2_a21oi_1 _32029_ (.A1(net4709),
    .A2(_09040_),
    .Y(_09042_),
    .B1(_09041_));
 sg13g2_nor3_1 _32030_ (.A(net4446),
    .B(_09038_),
    .C(_09042_),
    .Y(_09043_));
 sg13g2_o21ai_1 _32031_ (.B1(net4039),
    .Y(_09044_),
    .A1(net4626),
    .A2(net1934));
 sg13g2_o21ai_1 _32032_ (.B1(_09034_),
    .Y(_01437_),
    .A1(_09043_),
    .A2(_09044_));
 sg13g2_nand2_1 _32033_ (.Y(_09045_),
    .A(net2618),
    .B(net3988));
 sg13g2_a21oi_1 _32034_ (.A1(\u_inv.f_next[134] ),
    .A2(_10756_),
    .Y(_09046_),
    .B1(_09036_));
 sg13g2_o21ai_1 _32035_ (.B1(net3818),
    .Y(_09047_),
    .A1(_11710_),
    .A2(_09046_));
 sg13g2_a21oi_1 _32036_ (.A1(_11710_),
    .A2(_09046_),
    .Y(_09048_),
    .B1(_09047_));
 sg13g2_nand2_1 _32037_ (.Y(_09049_),
    .A(\u_inv.f_next[135] ),
    .B(net3865));
 sg13g2_o21ai_1 _32038_ (.B1(_11712_),
    .Y(_09050_),
    .A1(_11714_),
    .A2(_09039_));
 sg13g2_xnor2_1 _32039_ (.Y(_09051_),
    .A(_11710_),
    .B(_09050_));
 sg13g2_a22oi_1 _32040_ (.Y(_09052_),
    .B1(_09051_),
    .B2(net4709),
    .A2(_09049_),
    .A1(net3734));
 sg13g2_nor3_1 _32041_ (.A(net4446),
    .B(_09048_),
    .C(_09052_),
    .Y(_09053_));
 sg13g2_o21ai_1 _32042_ (.B1(net4043),
    .Y(_09054_),
    .A1(net4626),
    .A2(net1938));
 sg13g2_o21ai_1 _32043_ (.B1(_09045_),
    .Y(_01438_),
    .A1(_09053_),
    .A2(_09054_));
 sg13g2_a21o_2 _32044_ (.A2(_09016_),
    .A1(_12404_),
    .B1(_12402_),
    .X(_09055_));
 sg13g2_nor2b_1 _32045_ (.A(_11703_),
    .B_N(_09055_),
    .Y(_09056_));
 sg13g2_nand2b_1 _32046_ (.Y(_09057_),
    .B(_11703_),
    .A_N(_09055_));
 sg13g2_nand3b_1 _32047_ (.B(_09057_),
    .C(net4710),
    .Y(_09058_),
    .A_N(_09056_));
 sg13g2_a21oi_1 _32048_ (.A1(\u_inv.f_next[136] ),
    .A2(net4596),
    .Y(_09059_),
    .B1(net3708));
 sg13g2_o21ai_1 _32049_ (.B1(_11853_),
    .Y(_09060_),
    .A1(_11650_),
    .A2(_11727_));
 sg13g2_xnor2_1 _32050_ (.Y(_09061_),
    .A(_11703_),
    .B(_09060_));
 sg13g2_a221oi_1 _32051_ (.B2(net3697),
    .C1(net3989),
    .B1(_09061_),
    .A1(_09058_),
    .Y(_09062_),
    .A2(_09059_));
 sg13g2_o21ai_1 _32052_ (.B1(_09062_),
    .Y(_09063_),
    .A1(net4626),
    .A2(net2062));
 sg13g2_o21ai_1 _32053_ (.B1(_09063_),
    .Y(_01439_),
    .A1(_10446_),
    .A2(net4040));
 sg13g2_a21oi_1 _32054_ (.A1(_11703_),
    .A2(_09060_),
    .Y(_09064_),
    .B1(_11863_));
 sg13g2_nand2_1 _32055_ (.Y(_09065_),
    .A(_11705_),
    .B(_09064_));
 sg13g2_or2_1 _32056_ (.X(_09066_),
    .B(_09064_),
    .A(_11705_));
 sg13g2_nand3_1 _32057_ (.B(_09065_),
    .C(_09066_),
    .A(net3697),
    .Y(_09067_));
 sg13g2_a21oi_1 _32058_ (.A1(\u_inv.f_next[136] ),
    .A2(\u_inv.f_reg[136] ),
    .Y(_09068_),
    .B1(_09056_));
 sg13g2_xnor2_1 _32059_ (.Y(_09069_),
    .A(_11706_),
    .B(_09068_));
 sg13g2_o21ai_1 _32060_ (.B1(net3719),
    .Y(_09070_),
    .A1(net2332),
    .A2(net4710));
 sg13g2_a21oi_1 _32061_ (.A1(net4710),
    .A2(_09069_),
    .Y(_09071_),
    .B1(_09070_));
 sg13g2_a21oi_1 _32062_ (.A1(net4520),
    .A2(net1787),
    .Y(_09072_),
    .B1(net3988));
 sg13g2_nor2b_1 _32063_ (.A(_09071_),
    .B_N(_09072_),
    .Y(_09073_));
 sg13g2_a22oi_1 _32064_ (.Y(_01440_),
    .B1(_09067_),
    .B2(_09073_),
    .A2(net3989),
    .A1(_10445_));
 sg13g2_nand2_1 _32065_ (.Y(_09074_),
    .A(net2332),
    .B(net3988));
 sg13g2_nand2_1 _32066_ (.Y(_09075_),
    .A(_11862_),
    .B(_09066_));
 sg13g2_and2_1 _32067_ (.A(_11702_),
    .B(_09075_),
    .X(_09076_));
 sg13g2_o21ai_1 _32068_ (.B1(net3819),
    .Y(_09077_),
    .A1(_11702_),
    .A2(_09075_));
 sg13g2_nor2_1 _32069_ (.A(_09076_),
    .B(_09077_),
    .Y(_09078_));
 sg13g2_a21oi_2 _32070_ (.B1(_12389_),
    .Y(_09079_),
    .A2(_09055_),
    .A1(_12413_));
 sg13g2_inv_1 _32071_ (.Y(_09080_),
    .A(_09079_));
 sg13g2_xnor2_1 _32072_ (.Y(_09081_),
    .A(_11702_),
    .B(_09079_));
 sg13g2_o21ai_1 _32073_ (.B1(net3867),
    .Y(_09082_),
    .A1(\u_inv.f_next[138] ),
    .A2(net4711));
 sg13g2_a21oi_1 _32074_ (.A1(net4711),
    .A2(_09081_),
    .Y(_09083_),
    .B1(_09082_));
 sg13g2_nor3_1 _32075_ (.A(net4446),
    .B(_09078_),
    .C(_09083_),
    .Y(_09084_));
 sg13g2_o21ai_1 _32076_ (.B1(net4040),
    .Y(_09085_),
    .A1(net4626),
    .A2(net1751));
 sg13g2_o21ai_1 _32077_ (.B1(_09074_),
    .Y(_01441_),
    .A1(_09084_),
    .A2(_09085_));
 sg13g2_nor2_1 _32078_ (.A(net2542),
    .B(net4039),
    .Y(_09086_));
 sg13g2_nor3_1 _32079_ (.A(_11699_),
    .B(_11861_),
    .C(_09076_),
    .Y(_09087_));
 sg13g2_o21ai_1 _32080_ (.B1(_11699_),
    .Y(_09088_),
    .A1(_11861_),
    .A2(_09076_));
 sg13g2_nor2_1 _32081_ (.A(net3685),
    .B(_09087_),
    .Y(_09089_));
 sg13g2_o21ai_1 _32082_ (.B1(_11701_),
    .Y(_09090_),
    .A1(_11702_),
    .A2(_09079_));
 sg13g2_xnor2_1 _32083_ (.Y(_09091_),
    .A(_11700_),
    .B(_09090_));
 sg13g2_o21ai_1 _32084_ (.B1(net3719),
    .Y(_09092_),
    .A1(\u_inv.f_next[139] ),
    .A2(net4710));
 sg13g2_a21oi_1 _32085_ (.A1(net4710),
    .A2(_09091_),
    .Y(_09093_),
    .B1(_09092_));
 sg13g2_a221oi_1 _32086_ (.B2(_09089_),
    .C1(_09093_),
    .B1(_09088_),
    .A1(net4520),
    .Y(_09094_),
    .A2(net2319));
 sg13g2_a21oi_1 _32087_ (.A1(net4039),
    .A2(_09094_),
    .Y(_01442_),
    .B1(_09086_));
 sg13g2_a21oi_1 _32088_ (.A1(_12386_),
    .A2(_09080_),
    .Y(_09095_),
    .B1(_12392_));
 sg13g2_nand2b_1 _32089_ (.Y(_09096_),
    .B(_11696_),
    .A_N(_09095_));
 sg13g2_xnor2_1 _32090_ (.Y(_09097_),
    .A(_11696_),
    .B(_09095_));
 sg13g2_o21ai_1 _32091_ (.B1(net3719),
    .Y(_09098_),
    .A1(_10441_),
    .A2(net4710));
 sg13g2_a21oi_1 _32092_ (.A1(net4710),
    .A2(_09097_),
    .Y(_09099_),
    .B1(_09098_));
 sg13g2_a21oi_1 _32093_ (.A1(_11707_),
    .A2(_09060_),
    .Y(_09100_),
    .B1(_11867_));
 sg13g2_or2_1 _32094_ (.X(_09101_),
    .B(_09100_),
    .A(_11696_));
 sg13g2_xor2_1 _32095_ (.B(_09100_),
    .A(_11696_),
    .X(_09102_));
 sg13g2_o21ai_1 _32096_ (.B1(net4041),
    .Y(_09103_),
    .A1(net4626),
    .A2(net2026));
 sg13g2_nor2_1 _32097_ (.A(_09099_),
    .B(_09103_),
    .Y(_09104_));
 sg13g2_o21ai_1 _32098_ (.B1(_09104_),
    .Y(_09105_),
    .A1(net3685),
    .A2(_09102_));
 sg13g2_o21ai_1 _32099_ (.B1(_09105_),
    .Y(_01443_),
    .A1(_10442_),
    .A2(net4042));
 sg13g2_nand2_1 _32100_ (.Y(_09106_),
    .A(net1728),
    .B(net3989));
 sg13g2_nand2_1 _32101_ (.Y(_09107_),
    .A(\u_inv.f_next[141] ),
    .B(net3866));
 sg13g2_o21ai_1 _32102_ (.B1(_09096_),
    .Y(_09108_),
    .A1(_10441_),
    .A2(_10750_));
 sg13g2_xnor2_1 _32103_ (.Y(_09109_),
    .A(_11695_),
    .B(_09108_));
 sg13g2_a22oi_1 _32104_ (.Y(_09110_),
    .B1(_09109_),
    .B2(net4710),
    .A2(_09107_),
    .A1(net3734));
 sg13g2_a21oi_1 _32105_ (.A1(_11856_),
    .A2(_09101_),
    .Y(_09111_),
    .B1(_11695_));
 sg13g2_and3_1 _32106_ (.X(_09112_),
    .A(_11695_),
    .B(_11856_),
    .C(_09101_));
 sg13g2_nor3_1 _32107_ (.A(net3867),
    .B(_09111_),
    .C(_09112_),
    .Y(_09113_));
 sg13g2_nor3_1 _32108_ (.A(net4446),
    .B(_09110_),
    .C(_09113_),
    .Y(_09114_));
 sg13g2_o21ai_1 _32109_ (.B1(net4039),
    .Y(_09115_),
    .A1(net4626),
    .A2(\u_inv.input_reg[140] ));
 sg13g2_o21ai_1 _32110_ (.B1(_09106_),
    .Y(_01444_),
    .A1(_09114_),
    .A2(_09115_));
 sg13g2_nor2_1 _32111_ (.A(_12383_),
    .B(_09095_),
    .Y(_09116_));
 sg13g2_nor2_1 _32112_ (.A(_12395_),
    .B(_09116_),
    .Y(_09117_));
 sg13g2_xnor2_1 _32113_ (.Y(_09118_),
    .A(_11693_),
    .B(_09117_));
 sg13g2_a21oi_1 _32114_ (.A1(net2799),
    .A2(net4596),
    .Y(_09119_),
    .B1(net3708));
 sg13g2_o21ai_1 _32115_ (.B1(_09119_),
    .Y(_09120_),
    .A1(net4596),
    .A2(_09118_));
 sg13g2_nor3_1 _32116_ (.A(_11693_),
    .B(_11855_),
    .C(_09111_),
    .Y(_09121_));
 sg13g2_o21ai_1 _32117_ (.B1(_11693_),
    .Y(_09122_),
    .A1(_11855_),
    .A2(_09111_));
 sg13g2_nand2b_1 _32118_ (.Y(_09123_),
    .B(_09122_),
    .A_N(_09121_));
 sg13g2_o21ai_1 _32119_ (.B1(net4040),
    .Y(_09124_),
    .A1(net4626),
    .A2(net2225));
 sg13g2_a21oi_1 _32120_ (.A1(net3697),
    .A2(_09123_),
    .Y(_09125_),
    .B1(_09124_));
 sg13g2_nand2_1 _32121_ (.Y(_09126_),
    .A(_09120_),
    .B(_09125_));
 sg13g2_o21ai_1 _32122_ (.B1(_09126_),
    .Y(_01445_),
    .A1(_10440_),
    .A2(net4040));
 sg13g2_nand2_1 _32123_ (.Y(_09127_),
    .A(net2419),
    .B(net3867));
 sg13g2_o21ai_1 _32124_ (.B1(_11692_),
    .Y(_09128_),
    .A1(_11693_),
    .A2(_09117_));
 sg13g2_xnor2_1 _32125_ (.Y(_09129_),
    .A(_11691_),
    .B(_09128_));
 sg13g2_a22oi_1 _32126_ (.Y(_09130_),
    .B1(_09129_),
    .B2(net4711),
    .A2(_09127_),
    .A1(net3734));
 sg13g2_nand2_1 _32127_ (.Y(_09131_),
    .A(_11859_),
    .B(_09122_));
 sg13g2_xor2_1 _32128_ (.B(_09131_),
    .A(_11691_),
    .X(_09132_));
 sg13g2_o21ai_1 _32129_ (.B1(net4384),
    .Y(_09133_),
    .A1(net3867),
    .A2(_09132_));
 sg13g2_a21oi_1 _32130_ (.A1(net4520),
    .A2(_10979_),
    .Y(_09134_),
    .B1(net3989));
 sg13g2_o21ai_1 _32131_ (.B1(_09134_),
    .Y(_09135_),
    .A1(_09130_),
    .A2(_09133_));
 sg13g2_o21ai_1 _32132_ (.B1(_09135_),
    .Y(_01446_),
    .A1(_10439_),
    .A2(net4041));
 sg13g2_a21oi_1 _32133_ (.A1(_12414_),
    .A2(_09055_),
    .Y(_09136_),
    .B1(_12397_));
 sg13g2_a21o_2 _32134_ (.A2(_09055_),
    .A1(_12414_),
    .B1(_12397_),
    .X(_09137_));
 sg13g2_o21ai_1 _32135_ (.B1(net4711),
    .Y(_09138_),
    .A1(_11671_),
    .A2(_09136_));
 sg13g2_a21o_1 _32136_ (.A2(_09136_),
    .A1(_11671_),
    .B1(_09138_),
    .X(_09139_));
 sg13g2_a21oi_1 _32137_ (.A1(net2073),
    .A2(net4596),
    .Y(_09140_),
    .B1(net3708));
 sg13g2_o21ai_1 _32138_ (.B1(_11871_),
    .Y(_09141_),
    .A1(_11650_),
    .A2(_11728_));
 sg13g2_and2_1 _32139_ (.A(_11671_),
    .B(_09141_),
    .X(_09142_));
 sg13g2_xnor2_1 _32140_ (.Y(_09143_),
    .A(_11671_),
    .B(_09141_));
 sg13g2_o21ai_1 _32141_ (.B1(net4040),
    .Y(_09144_),
    .A1(net4625),
    .A2(net1939));
 sg13g2_a221oi_1 _32142_ (.B2(net3697),
    .C1(_09144_),
    .B1(_09143_),
    .A1(_09139_),
    .Y(_09145_),
    .A2(_09140_));
 sg13g2_a21o_1 _32143_ (.A2(net3989),
    .A1(net2419),
    .B1(_09145_),
    .X(_01447_));
 sg13g2_nand2_1 _32144_ (.Y(_09146_),
    .A(net2073),
    .B(net3988));
 sg13g2_o21ai_1 _32145_ (.B1(_11670_),
    .Y(_09147_),
    .A1(_11671_),
    .A2(_09136_));
 sg13g2_xor2_1 _32146_ (.B(_09147_),
    .A(_11674_),
    .X(_09148_));
 sg13g2_nor2_1 _32147_ (.A(\u_inv.f_next[145] ),
    .B(net4712),
    .Y(_09149_));
 sg13g2_a21oi_1 _32148_ (.A1(net4712),
    .A2(_09148_),
    .Y(_09150_),
    .B1(_09149_));
 sg13g2_or2_1 _32149_ (.X(_09151_),
    .B(_09142_),
    .A(_11816_));
 sg13g2_or2_1 _32150_ (.X(_09152_),
    .B(_09151_),
    .A(_11674_));
 sg13g2_a21oi_1 _32151_ (.A1(_11674_),
    .A2(_09151_),
    .Y(_09153_),
    .B1(net3866));
 sg13g2_a221oi_1 _32152_ (.B2(_09153_),
    .C1(net4447),
    .B1(_09152_),
    .A1(net3866),
    .Y(_09154_),
    .A2(_09150_));
 sg13g2_o21ai_1 _32153_ (.B1(net4040),
    .Y(_09155_),
    .A1(net4625),
    .A2(net1925));
 sg13g2_o21ai_1 _32154_ (.B1(_09146_),
    .Y(_01448_),
    .A1(_09154_),
    .A2(_09155_));
 sg13g2_a21oi_2 _32155_ (.B1(_12440_),
    .Y(_09156_),
    .A2(_09137_),
    .A1(_12426_));
 sg13g2_o21ai_1 _32156_ (.B1(net4711),
    .Y(_09157_),
    .A1(_11669_),
    .A2(_09156_));
 sg13g2_a21o_1 _32157_ (.A2(_09156_),
    .A1(_11669_),
    .B1(_09157_),
    .X(_09158_));
 sg13g2_a21oi_1 _32158_ (.A1(\u_inv.f_next[146] ),
    .A2(net4596),
    .Y(_09159_),
    .B1(net3708));
 sg13g2_a21oi_1 _32159_ (.A1(_11674_),
    .A2(_09142_),
    .Y(_09160_),
    .B1(_11818_));
 sg13g2_xnor2_1 _32160_ (.Y(_09161_),
    .A(_11668_),
    .B(_09160_));
 sg13g2_o21ai_1 _32161_ (.B1(net4040),
    .Y(_09162_),
    .A1(net4625),
    .A2(net1928));
 sg13g2_a221oi_1 _32162_ (.B2(net3697),
    .C1(_09162_),
    .B1(_09161_),
    .A1(_09158_),
    .Y(_09163_),
    .A2(_09159_));
 sg13g2_a21o_1 _32163_ (.A2(net3988),
    .A1(net2738),
    .B1(_09163_),
    .X(_01449_));
 sg13g2_o21ai_1 _32164_ (.B1(_11667_),
    .Y(_09164_),
    .A1(_11669_),
    .A2(_09156_));
 sg13g2_xnor2_1 _32165_ (.Y(_09165_),
    .A(_11672_),
    .B(_09164_));
 sg13g2_o21ai_1 _32166_ (.B1(net3719),
    .Y(_09166_),
    .A1(net3018),
    .A2(net4711));
 sg13g2_a21o_1 _32167_ (.A2(_09165_),
    .A1(net4711),
    .B1(_09166_),
    .X(_09167_));
 sg13g2_o21ai_1 _32168_ (.B1(_11820_),
    .Y(_09168_),
    .A1(_11668_),
    .A2(_09160_));
 sg13g2_xnor2_1 _32169_ (.Y(_09169_),
    .A(_11672_),
    .B(_09168_));
 sg13g2_a221oi_1 _32170_ (.B2(_09169_),
    .C1(net3988),
    .B1(net3697),
    .A1(net4520),
    .Y(_09170_),
    .A2(net2534));
 sg13g2_a22oi_1 _32171_ (.Y(_01450_),
    .B1(_09167_),
    .B2(_09170_),
    .A2(net3988),
    .A1(_10435_));
 sg13g2_o21ai_1 _32172_ (.B1(_12444_),
    .Y(_09171_),
    .A1(_12425_),
    .A2(_09156_));
 sg13g2_nand2_1 _32173_ (.Y(_09172_),
    .A(_11663_),
    .B(_09171_));
 sg13g2_xnor2_1 _32174_ (.Y(_09173_),
    .A(_11663_),
    .B(_09171_));
 sg13g2_a21oi_1 _32175_ (.A1(net3242),
    .A2(net4597),
    .Y(_09174_),
    .B1(net3708));
 sg13g2_o21ai_1 _32176_ (.B1(_09174_),
    .Y(_09175_),
    .A1(net4597),
    .A2(_09173_));
 sg13g2_nor2b_2 _32177_ (.A(_11675_),
    .B_N(_09141_),
    .Y(_09176_));
 sg13g2_nor2_1 _32178_ (.A(_11822_),
    .B(_09176_),
    .Y(_09177_));
 sg13g2_o21ai_1 _32179_ (.B1(_11664_),
    .Y(_09178_),
    .A1(_11822_),
    .A2(_09176_));
 sg13g2_xnor2_1 _32180_ (.Y(_09179_),
    .A(_11663_),
    .B(_09177_));
 sg13g2_o21ai_1 _32181_ (.B1(net4041),
    .Y(_09180_),
    .A1(net4625),
    .A2(net1981));
 sg13g2_a21oi_1 _32182_ (.A1(net3697),
    .A2(_09179_),
    .Y(_09181_),
    .B1(_09180_));
 sg13g2_nand2_1 _32183_ (.Y(_09182_),
    .A(_09175_),
    .B(_09181_));
 sg13g2_o21ai_1 _32184_ (.B1(_09182_),
    .Y(_01451_),
    .A1(_10434_),
    .A2(net4041));
 sg13g2_o21ai_1 _32185_ (.B1(_09172_),
    .Y(_09183_),
    .A1(_10433_),
    .A2(_10742_));
 sg13g2_xor2_1 _32186_ (.B(_09183_),
    .A(_11659_),
    .X(_09184_));
 sg13g2_o21ai_1 _32187_ (.B1(net3719),
    .Y(_09185_),
    .A1(_10432_),
    .A2(net4717));
 sg13g2_a21oi_1 _32188_ (.A1(net4717),
    .A2(_09184_),
    .Y(_09186_),
    .B1(_09185_));
 sg13g2_and3_1 _32189_ (.X(_09187_),
    .A(_11659_),
    .B(_11815_),
    .C(_09178_));
 sg13g2_a21oi_1 _32190_ (.A1(_11815_),
    .A2(_09178_),
    .Y(_09188_),
    .B1(_11659_));
 sg13g2_nor2_1 _32191_ (.A(_09187_),
    .B(_09188_),
    .Y(_09189_));
 sg13g2_o21ai_1 _32192_ (.B1(net4041),
    .Y(_09190_),
    .A1(net4627),
    .A2(net2135));
 sg13g2_nor2_1 _32193_ (.A(_09186_),
    .B(_09190_),
    .Y(_09191_));
 sg13g2_o21ai_1 _32194_ (.B1(_09191_),
    .Y(_09192_),
    .A1(net3685),
    .A2(_09189_));
 sg13g2_o21ai_1 _32195_ (.B1(_09192_),
    .Y(_01452_),
    .A1(_10433_),
    .A2(net4041));
 sg13g2_a21oi_1 _32196_ (.A1(_12424_),
    .A2(_09171_),
    .Y(_09193_),
    .B1(_12447_));
 sg13g2_xnor2_1 _32197_ (.Y(_09194_),
    .A(_11662_),
    .B(_09193_));
 sg13g2_a21oi_1 _32198_ (.A1(net3093),
    .A2(net4597),
    .Y(_09195_),
    .B1(net3708));
 sg13g2_o21ai_1 _32199_ (.B1(_09195_),
    .Y(_09196_),
    .A1(net4597),
    .A2(_09194_));
 sg13g2_nor2_1 _32200_ (.A(_11825_),
    .B(_09188_),
    .Y(_09197_));
 sg13g2_nor2_1 _32201_ (.A(_11661_),
    .B(_09197_),
    .Y(_09198_));
 sg13g2_xnor2_1 _32202_ (.Y(_09199_),
    .A(_11661_),
    .B(_09197_));
 sg13g2_o21ai_1 _32203_ (.B1(net4047),
    .Y(_09200_),
    .A1(net4627),
    .A2(net2433));
 sg13g2_a21oi_1 _32204_ (.A1(net3697),
    .A2(_09199_),
    .Y(_09201_),
    .B1(_09200_));
 sg13g2_nand2_1 _32205_ (.Y(_09202_),
    .A(_09196_),
    .B(_09201_));
 sg13g2_o21ai_1 _32206_ (.B1(_09202_),
    .Y(_01453_),
    .A1(_10432_),
    .A2(net4047));
 sg13g2_nand2_1 _32207_ (.Y(_09203_),
    .A(net3042),
    .B(net3870));
 sg13g2_o21ai_1 _32208_ (.B1(_11660_),
    .Y(_09204_),
    .A1(_11662_),
    .A2(_09193_));
 sg13g2_xnor2_1 _32209_ (.Y(_09205_),
    .A(_11665_),
    .B(_09204_));
 sg13g2_a22oi_1 _32210_ (.Y(_09206_),
    .B1(_09205_),
    .B2(net4717),
    .A2(_09203_),
    .A1(net3732));
 sg13g2_or2_1 _32211_ (.X(_09207_),
    .B(_09198_),
    .A(_11824_));
 sg13g2_xor2_1 _32212_ (.B(_09207_),
    .A(_11665_),
    .X(_09208_));
 sg13g2_o21ai_1 _32213_ (.B1(net4384),
    .Y(_09209_),
    .A1(net3870),
    .A2(_09208_));
 sg13g2_a21oi_1 _32214_ (.A1(net4520),
    .A2(_10980_),
    .Y(_09210_),
    .B1(net3995));
 sg13g2_o21ai_1 _32215_ (.B1(_09210_),
    .Y(_09211_),
    .A1(_09206_),
    .A2(_09209_));
 sg13g2_o21ai_1 _32216_ (.B1(_09211_),
    .Y(_01454_),
    .A1(_10431_),
    .A2(net4047));
 sg13g2_a21oi_2 _32217_ (.B1(_12452_),
    .Y(_09212_),
    .A2(_09137_),
    .A1(_12428_));
 sg13g2_nand2b_1 _32218_ (.Y(_09213_),
    .B(_11651_),
    .A_N(_09212_));
 sg13g2_xnor2_1 _32219_ (.Y(_09214_),
    .A(_11651_),
    .B(_09212_));
 sg13g2_o21ai_1 _32220_ (.B1(net3719),
    .Y(_09215_),
    .A1(_10429_),
    .A2(net4717));
 sg13g2_a21oi_1 _32221_ (.A1(net4717),
    .A2(_09214_),
    .Y(_09216_),
    .B1(_09215_));
 sg13g2_a21oi_2 _32222_ (.B1(_11829_),
    .Y(_09217_),
    .A2(_09176_),
    .A1(_11666_));
 sg13g2_nor2_1 _32223_ (.A(_11651_),
    .B(_09217_),
    .Y(_09218_));
 sg13g2_xor2_1 _32224_ (.B(_09217_),
    .A(_11651_),
    .X(_09219_));
 sg13g2_o21ai_1 _32225_ (.B1(net4047),
    .Y(_09220_),
    .A1(net4625),
    .A2(net1989));
 sg13g2_nor2_1 _32226_ (.A(_09216_),
    .B(_09220_),
    .Y(_09221_));
 sg13g2_o21ai_1 _32227_ (.B1(_09221_),
    .Y(_09222_),
    .A1(net3685),
    .A2(_09219_));
 sg13g2_o21ai_1 _32228_ (.B1(_09222_),
    .Y(_01455_),
    .A1(_10430_),
    .A2(net4047));
 sg13g2_nand2_1 _32229_ (.Y(_09223_),
    .A(net2878),
    .B(net3870));
 sg13g2_o21ai_1 _32230_ (.B1(_09213_),
    .Y(_09224_),
    .A1(_10429_),
    .A2(_10738_));
 sg13g2_xnor2_1 _32231_ (.Y(_09225_),
    .A(_11652_),
    .B(_09224_));
 sg13g2_a22oi_1 _32232_ (.Y(_09226_),
    .B1(_09225_),
    .B2(net4717),
    .A2(_09223_),
    .A1(net3732));
 sg13g2_nor2_1 _32233_ (.A(_11808_),
    .B(_09218_),
    .Y(_09227_));
 sg13g2_or2_1 _32234_ (.X(_09228_),
    .B(_09227_),
    .A(_11652_));
 sg13g2_xnor2_1 _32235_ (.Y(_09229_),
    .A(_11652_),
    .B(_09227_));
 sg13g2_o21ai_1 _32236_ (.B1(net4384),
    .Y(_09230_),
    .A1(net3870),
    .A2(_09229_));
 sg13g2_a21oi_1 _32237_ (.A1(net4520),
    .A2(_10981_),
    .Y(_09231_),
    .B1(net3995));
 sg13g2_o21ai_1 _32238_ (.B1(_09231_),
    .Y(_09232_),
    .A1(_09226_),
    .A2(_09230_));
 sg13g2_o21ai_1 _32239_ (.B1(_09232_),
    .Y(_01456_),
    .A1(_10429_),
    .A2(net4047));
 sg13g2_and3_1 _32240_ (.X(_09233_),
    .A(_11654_),
    .B(_11807_),
    .C(_09228_));
 sg13g2_a21oi_1 _32241_ (.A1(_11807_),
    .A2(_09228_),
    .Y(_09234_),
    .B1(_11654_));
 sg13g2_nor2_1 _32242_ (.A(_09233_),
    .B(_09234_),
    .Y(_09235_));
 sg13g2_o21ai_1 _32243_ (.B1(net4047),
    .Y(_09236_),
    .A1(net4630),
    .A2(net1819));
 sg13g2_nor2_1 _32244_ (.A(_12420_),
    .B(_09212_),
    .Y(_09237_));
 sg13g2_nor2_1 _32245_ (.A(_12434_),
    .B(_09237_),
    .Y(_09238_));
 sg13g2_nor2b_1 _32246_ (.A(_09238_),
    .B_N(_11654_),
    .Y(_09239_));
 sg13g2_xnor2_1 _32247_ (.Y(_09240_),
    .A(_11654_),
    .B(_09238_));
 sg13g2_o21ai_1 _32248_ (.B1(net3718),
    .Y(_09241_),
    .A1(_10427_),
    .A2(net4718));
 sg13g2_a21oi_1 _32249_ (.A1(net4718),
    .A2(_09240_),
    .Y(_09242_),
    .B1(_09241_));
 sg13g2_nor2_1 _32250_ (.A(_09236_),
    .B(_09242_),
    .Y(_09243_));
 sg13g2_o21ai_1 _32251_ (.B1(_09243_),
    .Y(_09244_),
    .A1(net3686),
    .A2(_09235_));
 sg13g2_o21ai_1 _32252_ (.B1(_09244_),
    .Y(_01457_),
    .A1(_10428_),
    .A2(net4048));
 sg13g2_nor2_1 _32253_ (.A(_11806_),
    .B(_09234_),
    .Y(_09245_));
 sg13g2_xnor2_1 _32254_ (.Y(_09246_),
    .A(_11656_),
    .B(_09245_));
 sg13g2_nor2_1 _32255_ (.A(_11653_),
    .B(_09239_),
    .Y(_09247_));
 sg13g2_xnor2_1 _32256_ (.Y(_09248_),
    .A(_11656_),
    .B(_09247_));
 sg13g2_o21ai_1 _32257_ (.B1(net3718),
    .Y(_09249_),
    .A1(net3199),
    .A2(net4718));
 sg13g2_a21o_1 _32258_ (.A2(_09248_),
    .A1(net4718),
    .B1(_09249_),
    .X(_09250_));
 sg13g2_a221oi_1 _32259_ (.B2(_09246_),
    .C1(net3995),
    .B1(net3698),
    .A1(net4519),
    .Y(_09251_),
    .A2(net2698));
 sg13g2_a22oi_1 _32260_ (.Y(_01458_),
    .B1(_09250_),
    .B2(_09251_),
    .A2(net3995),
    .A1(_10427_));
 sg13g2_nor2_1 _32261_ (.A(_10426_),
    .B(net4048),
    .Y(_09252_));
 sg13g2_a21o_2 _32262_ (.A2(_09237_),
    .A1(_12419_),
    .B1(_12438_),
    .X(_09253_));
 sg13g2_nor2b_1 _32263_ (.A(_11684_),
    .B_N(_09253_),
    .Y(_09254_));
 sg13g2_xnor2_1 _32264_ (.Y(_09255_),
    .A(_11684_),
    .B(_09253_));
 sg13g2_o21ai_1 _32265_ (.B1(net3718),
    .Y(_09256_),
    .A1(_10425_),
    .A2(net4717));
 sg13g2_a21oi_1 _32266_ (.A1(net4718),
    .A2(_09255_),
    .Y(_09257_),
    .B1(_09256_));
 sg13g2_o21ai_1 _32267_ (.B1(_11813_),
    .Y(_09258_),
    .A1(_11658_),
    .A2(_09217_));
 sg13g2_xnor2_1 _32268_ (.Y(_09259_),
    .A(_11684_),
    .B(_09258_));
 sg13g2_nand2_1 _32269_ (.Y(_09260_),
    .A(net3698),
    .B(_09259_));
 sg13g2_o21ai_1 _32270_ (.B1(net4047),
    .Y(_09261_),
    .A1(net4630),
    .A2(net2550));
 sg13g2_nor2_1 _32271_ (.A(_09257_),
    .B(_09261_),
    .Y(_09262_));
 sg13g2_a21o_1 _32272_ (.A2(_09262_),
    .A1(_09260_),
    .B1(_09252_),
    .X(_01459_));
 sg13g2_nand2_1 _32273_ (.Y(_09263_),
    .A(net1748),
    .B(net3995));
 sg13g2_nand2_1 _32274_ (.Y(_09264_),
    .A(\u_inv.f_next[157] ),
    .B(net3870));
 sg13g2_a21oi_1 _32275_ (.A1(\u_inv.f_next[156] ),
    .A2(\u_inv.f_reg[156] ),
    .Y(_09265_),
    .B1(_09254_));
 sg13g2_xnor2_1 _32276_ (.Y(_09266_),
    .A(_11683_),
    .B(_09265_));
 sg13g2_a22oi_1 _32277_ (.Y(_09267_),
    .B1(_09266_),
    .B2(net4717),
    .A2(_09264_),
    .A1(net3732));
 sg13g2_a21o_1 _32278_ (.A2(_09258_),
    .A1(_11684_),
    .B1(_11834_),
    .X(_09268_));
 sg13g2_nand2_1 _32279_ (.Y(_09269_),
    .A(_11683_),
    .B(_09268_));
 sg13g2_inv_1 _32280_ (.Y(_09270_),
    .A(_09269_));
 sg13g2_nor2_1 _32281_ (.A(_11683_),
    .B(_09268_),
    .Y(_09271_));
 sg13g2_o21ai_1 _32282_ (.B1(net4384),
    .Y(_09272_),
    .A1(_09270_),
    .A2(_09271_));
 sg13g2_a21oi_1 _32283_ (.A1(net3708),
    .A2(_09272_),
    .Y(_09273_),
    .B1(_09267_));
 sg13g2_o21ai_1 _32284_ (.B1(net4048),
    .Y(_09274_),
    .A1(net4630),
    .A2(\u_inv.input_reg[156] ));
 sg13g2_o21ai_1 _32285_ (.B1(_09263_),
    .Y(_01460_),
    .A1(_09273_),
    .A2(_09274_));
 sg13g2_nand2_1 _32286_ (.Y(_09275_),
    .A(_11833_),
    .B(_09269_));
 sg13g2_xnor2_1 _32287_ (.Y(_09276_),
    .A(_11680_),
    .B(_09275_));
 sg13g2_a22oi_1 _32288_ (.Y(_09277_),
    .B1(_09253_),
    .B2(_12417_),
    .A2(_12430_),
    .A1(_11682_));
 sg13g2_xnor2_1 _32289_ (.Y(_09278_),
    .A(_11680_),
    .B(_09277_));
 sg13g2_o21ai_1 _32290_ (.B1(net3720),
    .Y(_09279_),
    .A1(_10423_),
    .A2(net4719));
 sg13g2_a21oi_1 _32291_ (.A1(net4719),
    .A2(_09278_),
    .Y(_09280_),
    .B1(_09279_));
 sg13g2_o21ai_1 _32292_ (.B1(net4048),
    .Y(_09281_),
    .A1(net4630),
    .A2(net2239));
 sg13g2_nor2_1 _32293_ (.A(_09280_),
    .B(_09281_),
    .Y(_09282_));
 sg13g2_o21ai_1 _32294_ (.B1(_09282_),
    .Y(_09283_),
    .A1(net3686),
    .A2(_09276_));
 sg13g2_o21ai_1 _32295_ (.B1(_09283_),
    .Y(_01461_),
    .A1(_10424_),
    .A2(net4048));
 sg13g2_nand2_1 _32296_ (.Y(_09284_),
    .A(net1475),
    .B(net3995));
 sg13g2_a21oi_1 _32297_ (.A1(_11681_),
    .A2(_09275_),
    .Y(_09285_),
    .B1(_11832_));
 sg13g2_xnor2_1 _32298_ (.Y(_09286_),
    .A(_11678_),
    .B(_09285_));
 sg13g2_a21oi_1 _32299_ (.A1(_10422_),
    .A2(net4597),
    .Y(_09287_),
    .B1(net3821));
 sg13g2_o21ai_1 _32300_ (.B1(_11679_),
    .Y(_09288_),
    .A1(_11681_),
    .A2(_09277_));
 sg13g2_o21ai_1 _32301_ (.B1(net4719),
    .Y(_09289_),
    .A1(_11678_),
    .A2(_09288_));
 sg13g2_a21o_1 _32302_ (.A2(_09288_),
    .A1(_11678_),
    .B1(_09289_),
    .X(_09290_));
 sg13g2_a221oi_1 _32303_ (.B2(_09290_),
    .C1(net4449),
    .B1(_09287_),
    .A1(net3821),
    .Y(_09291_),
    .A2(_09286_));
 sg13g2_o21ai_1 _32304_ (.B1(net4048),
    .Y(_09292_),
    .A1(net4630),
    .A2(\u_inv.input_reg[158] ));
 sg13g2_o21ai_1 _32305_ (.B1(_09284_),
    .Y(_01462_),
    .A1(_09291_),
    .A2(_09292_));
 sg13g2_o21ai_1 _32306_ (.B1(_11729_),
    .Y(_09293_),
    .A1(_11585_),
    .A2(_11649_));
 sg13g2_nand2_2 _32307_ (.Y(_09294_),
    .A(_11873_),
    .B(_09293_));
 sg13g2_nor2_1 _32308_ (.A(net4432),
    .B(_09294_),
    .Y(_09295_));
 sg13g2_and2_1 _32309_ (.A(net4432),
    .B(_09294_),
    .X(_09296_));
 sg13g2_nor3_1 _32310_ (.A(net3685),
    .B(_09295_),
    .C(_09296_),
    .Y(_09297_));
 sg13g2_nand2_1 _32311_ (.Y(_09298_),
    .A(net4519),
    .B(net1219));
 sg13g2_a21oi_2 _32312_ (.B1(_12457_),
    .Y(_09299_),
    .A2(_12753_),
    .A1(_12751_));
 sg13g2_nor2_1 _32313_ (.A(net4432),
    .B(_09299_),
    .Y(_09300_));
 sg13g2_xnor2_1 _32314_ (.Y(_09301_),
    .A(net4432),
    .B(_09299_));
 sg13g2_o21ai_1 _32315_ (.B1(net3718),
    .Y(_09302_),
    .A1(\u_inv.f_next[160] ),
    .A2(net4714));
 sg13g2_a21oi_1 _32316_ (.A1(net4714),
    .A2(_09301_),
    .Y(_09303_),
    .B1(_09302_));
 sg13g2_nor3_2 _32317_ (.A(net3991),
    .B(_09297_),
    .C(_09303_),
    .Y(_09304_));
 sg13g2_a22oi_1 _32318_ (.Y(_01463_),
    .B1(_09298_),
    .B2(_09304_),
    .A2(net3992),
    .A1(_10422_));
 sg13g2_o21ai_1 _32319_ (.B1(_11793_),
    .Y(_09305_),
    .A1(_11881_),
    .A2(_09296_));
 sg13g2_nor3_1 _32320_ (.A(_11793_),
    .B(_11881_),
    .C(_09296_),
    .Y(_09306_));
 sg13g2_o21ai_1 _32321_ (.B1(net4044),
    .Y(_09307_),
    .A1(net4628),
    .A2(net1947));
 sg13g2_a21oi_1 _32322_ (.A1(\u_inv.f_next[160] ),
    .A2(\u_inv.f_reg[160] ),
    .Y(_09308_),
    .B1(_09300_));
 sg13g2_nor2_1 _32323_ (.A(net3869),
    .B(_09306_),
    .Y(_09309_));
 sg13g2_nand2_1 _32324_ (.Y(_09310_),
    .A(\u_inv.f_next[161] ),
    .B(net3869));
 sg13g2_xnor2_1 _32325_ (.Y(_09311_),
    .A(_11793_),
    .B(_09308_));
 sg13g2_a22oi_1 _32326_ (.Y(_09312_),
    .B1(_09311_),
    .B2(net4714),
    .A2(_09310_),
    .A1(net3733));
 sg13g2_a21oi_1 _32327_ (.A1(_09305_),
    .A2(_09309_),
    .Y(_09313_),
    .B1(_09312_));
 sg13g2_a21o_1 _32328_ (.A2(_09313_),
    .A1(net4385),
    .B1(_09307_),
    .X(_09314_));
 sg13g2_o21ai_1 _32329_ (.B1(_09314_),
    .Y(_01464_),
    .A1(_10421_),
    .A2(net4044));
 sg13g2_nand2_1 _32330_ (.Y(_09315_),
    .A(net2140),
    .B(net3991));
 sg13g2_and2_1 _32331_ (.A(_11880_),
    .B(_09305_),
    .X(_09316_));
 sg13g2_nor2_1 _32332_ (.A(_11791_),
    .B(_09316_),
    .Y(_09317_));
 sg13g2_a21oi_1 _32333_ (.A1(_11791_),
    .A2(_09316_),
    .Y(_09318_),
    .B1(net3869));
 sg13g2_nor2b_1 _32334_ (.A(_09317_),
    .B_N(_09318_),
    .Y(_09319_));
 sg13g2_nor3_1 _32335_ (.A(net4432),
    .B(_11793_),
    .C(_09299_),
    .Y(_09320_));
 sg13g2_nor2_1 _32336_ (.A(_12360_),
    .B(_09320_),
    .Y(_09321_));
 sg13g2_xnor2_1 _32337_ (.Y(_09322_),
    .A(_11790_),
    .B(_09321_));
 sg13g2_o21ai_1 _32338_ (.B1(net3872),
    .Y(_09323_),
    .A1(net1772),
    .A2(net4715));
 sg13g2_a21oi_1 _32339_ (.A1(net4715),
    .A2(_09322_),
    .Y(_09324_),
    .B1(_09323_));
 sg13g2_nor3_1 _32340_ (.A(net4447),
    .B(_09319_),
    .C(_09324_),
    .Y(_09325_));
 sg13g2_o21ai_1 _32341_ (.B1(net4044),
    .Y(_09326_),
    .A1(net4629),
    .A2(net1887));
 sg13g2_o21ai_1 _32342_ (.B1(_09315_),
    .Y(_01465_),
    .A1(_09325_),
    .A2(_09326_));
 sg13g2_nand2_1 _32343_ (.Y(_09327_),
    .A(net1772),
    .B(net3991));
 sg13g2_or2_1 _32344_ (.X(_09328_),
    .B(_09317_),
    .A(_11879_));
 sg13g2_o21ai_1 _32345_ (.B1(net3820),
    .Y(_09329_),
    .A1(_11788_),
    .A2(_09328_));
 sg13g2_a21oi_1 _32346_ (.A1(_11788_),
    .A2(_09328_),
    .Y(_09330_),
    .B1(_09329_));
 sg13g2_nand2_1 _32347_ (.Y(_09331_),
    .A(\u_inv.f_next[163] ),
    .B(net3869));
 sg13g2_o21ai_1 _32348_ (.B1(_11789_),
    .Y(_09332_),
    .A1(_11790_),
    .A2(_09321_));
 sg13g2_xor2_1 _32349_ (.B(_09332_),
    .A(_11788_),
    .X(_09333_));
 sg13g2_a22oi_1 _32350_ (.Y(_09334_),
    .B1(_09333_),
    .B2(net4714),
    .A2(_09331_),
    .A1(net3733));
 sg13g2_nor3_1 _32351_ (.A(net4447),
    .B(_09330_),
    .C(_09334_),
    .Y(_09335_));
 sg13g2_o21ai_1 _32352_ (.B1(net4044),
    .Y(_09336_),
    .A1(net4629),
    .A2(\u_inv.input_reg[162] ));
 sg13g2_o21ai_1 _32353_ (.B1(_09327_),
    .Y(_01466_),
    .A1(_09335_),
    .A2(_09336_));
 sg13g2_nand2_1 _32354_ (.Y(_09337_),
    .A(net1908),
    .B(net3991));
 sg13g2_a21oi_1 _32355_ (.A1(_11794_),
    .A2(_09294_),
    .Y(_09338_),
    .B1(_11885_));
 sg13g2_o21ai_1 _32356_ (.B1(net3820),
    .Y(_09339_),
    .A1(_11798_),
    .A2(_09338_));
 sg13g2_a21oi_1 _32357_ (.A1(_11798_),
    .A2(_09338_),
    .Y(_09340_),
    .B1(_09339_));
 sg13g2_nor3_1 _32358_ (.A(_11792_),
    .B(_12458_),
    .C(_09299_),
    .Y(_09341_));
 sg13g2_nand2b_2 _32359_ (.Y(_09342_),
    .B(_12362_),
    .A_N(_09341_));
 sg13g2_nand2_1 _32360_ (.Y(_09343_),
    .A(_11798_),
    .B(_09342_));
 sg13g2_xnor2_1 _32361_ (.Y(_09344_),
    .A(_11798_),
    .B(_09342_));
 sg13g2_o21ai_1 _32362_ (.B1(net3869),
    .Y(_09345_),
    .A1(\u_inv.f_next[164] ),
    .A2(net4714));
 sg13g2_a21oi_1 _32363_ (.A1(net4714),
    .A2(_09344_),
    .Y(_09346_),
    .B1(_09345_));
 sg13g2_nor3_1 _32364_ (.A(net4447),
    .B(_09340_),
    .C(_09346_),
    .Y(_09347_));
 sg13g2_o21ai_1 _32365_ (.B1(net4044),
    .Y(_09348_),
    .A1(net4628),
    .A2(net1818));
 sg13g2_o21ai_1 _32366_ (.B1(_09337_),
    .Y(_01467_),
    .A1(_09347_),
    .A2(_09348_));
 sg13g2_nand2_1 _32367_ (.Y(_09349_),
    .A(net2256),
    .B(net3991));
 sg13g2_o21ai_1 _32368_ (.B1(_11877_),
    .Y(_09350_),
    .A1(_11798_),
    .A2(_09338_));
 sg13g2_nand2_1 _32369_ (.Y(_09351_),
    .A(_11800_),
    .B(_09350_));
 sg13g2_o21ai_1 _32370_ (.B1(net3820),
    .Y(_09352_),
    .A1(_11800_),
    .A2(_09350_));
 sg13g2_nor2b_1 _32371_ (.A(_09352_),
    .B_N(_09351_),
    .Y(_09353_));
 sg13g2_o21ai_1 _32372_ (.B1(_09343_),
    .Y(_09354_),
    .A1(_10417_),
    .A2(_10726_));
 sg13g2_xnor2_1 _32373_ (.Y(_09355_),
    .A(_11799_),
    .B(_09354_));
 sg13g2_nand2_1 _32374_ (.Y(_09356_),
    .A(\u_inv.f_next[165] ),
    .B(net3869));
 sg13g2_a22oi_1 _32375_ (.Y(_09357_),
    .B1(_09356_),
    .B2(net3733),
    .A2(_09355_),
    .A1(net4715));
 sg13g2_nor3_1 _32376_ (.A(net4447),
    .B(_09353_),
    .C(_09357_),
    .Y(_09358_));
 sg13g2_o21ai_1 _32377_ (.B1(net4046),
    .Y(_09359_),
    .A1(net4629),
    .A2(net1896));
 sg13g2_o21ai_1 _32378_ (.B1(_09349_),
    .Y(_01468_),
    .A1(_09358_),
    .A2(_09359_));
 sg13g2_nand2_1 _32379_ (.Y(_09360_),
    .A(net2854),
    .B(net3991));
 sg13g2_nand2_1 _32380_ (.Y(_09361_),
    .A(_11876_),
    .B(_09351_));
 sg13g2_o21ai_1 _32381_ (.B1(net3820),
    .Y(_09362_),
    .A1(_11797_),
    .A2(_09361_));
 sg13g2_a21oi_1 _32382_ (.A1(_11797_),
    .A2(_09361_),
    .Y(_09363_),
    .B1(_09362_));
 sg13g2_a21oi_1 _32383_ (.A1(_12356_),
    .A2(_09342_),
    .Y(_09364_),
    .B1(_12365_));
 sg13g2_xnor2_1 _32384_ (.Y(_09365_),
    .A(_11797_),
    .B(_09364_));
 sg13g2_o21ai_1 _32385_ (.B1(net3869),
    .Y(_09366_),
    .A1(net2021),
    .A2(net4715));
 sg13g2_a21oi_1 _32386_ (.A1(net4715),
    .A2(_09365_),
    .Y(_09367_),
    .B1(_09366_));
 sg13g2_nor3_1 _32387_ (.A(net4447),
    .B(_09363_),
    .C(_09367_),
    .Y(_09368_));
 sg13g2_o21ai_1 _32388_ (.B1(net4044),
    .Y(_09369_),
    .A1(net4628),
    .A2(net1882));
 sg13g2_o21ai_1 _32389_ (.B1(_09360_),
    .Y(_01469_),
    .A1(_09368_),
    .A2(_09369_));
 sg13g2_nand2_1 _32390_ (.Y(_09370_),
    .A(net2021),
    .B(net3991));
 sg13g2_a21oi_1 _32391_ (.A1(_11797_),
    .A2(_09361_),
    .Y(_09371_),
    .B1(_11875_));
 sg13g2_xnor2_1 _32392_ (.Y(_09372_),
    .A(_11795_),
    .B(_09371_));
 sg13g2_o21ai_1 _32393_ (.B1(_11796_),
    .Y(_09373_),
    .A1(_11797_),
    .A2(_09364_));
 sg13g2_o21ai_1 _32394_ (.B1(net4714),
    .Y(_09374_),
    .A1(_11795_),
    .A2(_09373_));
 sg13g2_a21o_1 _32395_ (.A2(_09373_),
    .A1(_11795_),
    .B1(_09374_),
    .X(_09375_));
 sg13g2_o21ai_1 _32396_ (.B1(_09375_),
    .Y(_09376_),
    .A1(\u_inv.f_next[167] ),
    .A2(net4714));
 sg13g2_o21ai_1 _32397_ (.B1(net4385),
    .Y(_09377_),
    .A1(net3820),
    .A2(_09376_));
 sg13g2_a21oi_1 _32398_ (.A1(net3820),
    .A2(_09372_),
    .Y(_09378_),
    .B1(_09377_));
 sg13g2_o21ai_1 _32399_ (.B1(net4044),
    .Y(_09379_),
    .A1(net4628),
    .A2(net2000));
 sg13g2_o21ai_1 _32400_ (.B1(_09370_),
    .Y(_01470_),
    .A1(_09378_),
    .A2(_09379_));
 sg13g2_a21oi_2 _32401_ (.B1(_11888_),
    .Y(_09380_),
    .A2(_09294_),
    .A1(_11803_));
 sg13g2_or2_1 _32402_ (.X(_09381_),
    .B(_09380_),
    .A(_11783_));
 sg13g2_a21oi_1 _32403_ (.A1(_11783_),
    .A2(_09380_),
    .Y(_09382_),
    .B1(net3861));
 sg13g2_a21oi_2 _32404_ (.B1(_12367_),
    .Y(_09383_),
    .A2(_09300_),
    .A1(_12459_));
 sg13g2_xnor2_1 _32405_ (.Y(_09384_),
    .A(_11784_),
    .B(_09383_));
 sg13g2_o21ai_1 _32406_ (.B1(net3861),
    .Y(_09385_),
    .A1(\u_inv.f_next[168] ),
    .A2(net4706));
 sg13g2_a21oi_1 _32407_ (.A1(net4706),
    .A2(_09384_),
    .Y(_09386_),
    .B1(_09385_));
 sg13g2_a21oi_1 _32408_ (.A1(_09381_),
    .A2(_09382_),
    .Y(_09387_),
    .B1(_09386_));
 sg13g2_o21ai_1 _32409_ (.B1(net4037),
    .Y(_09388_),
    .A1(net4629),
    .A2(net1885));
 sg13g2_a21o_1 _32410_ (.A2(_09387_),
    .A1(net4386),
    .B1(_09388_),
    .X(_09389_));
 sg13g2_o21ai_1 _32411_ (.B1(_09389_),
    .Y(_01471_),
    .A1(_10414_),
    .A2(net4036));
 sg13g2_nand2_1 _32412_ (.Y(_09390_),
    .A(net2818),
    .B(net3983));
 sg13g2_o21ai_1 _32413_ (.B1(_09381_),
    .Y(_09391_),
    .A1(_10413_),
    .A2(\u_inv.f_reg[168] ));
 sg13g2_and2_1 _32414_ (.A(_11785_),
    .B(_09391_),
    .X(_09392_));
 sg13g2_o21ai_1 _32415_ (.B1(net3815),
    .Y(_09393_),
    .A1(_11785_),
    .A2(_09391_));
 sg13g2_nor2_1 _32416_ (.A(_09392_),
    .B(_09393_),
    .Y(_09394_));
 sg13g2_nand2_1 _32417_ (.Y(_09395_),
    .A(net2083),
    .B(net3861));
 sg13g2_o21ai_1 _32418_ (.B1(_11782_),
    .Y(_09396_),
    .A1(_11784_),
    .A2(_09383_));
 sg13g2_xor2_1 _32419_ (.B(_09396_),
    .A(_11785_),
    .X(_09397_));
 sg13g2_a22oi_1 _32420_ (.Y(_09398_),
    .B1(_09397_),
    .B2(net4706),
    .A2(_09395_),
    .A1(net3735));
 sg13g2_nor3_1 _32421_ (.A(net4448),
    .B(_09394_),
    .C(_09398_),
    .Y(_09399_));
 sg13g2_o21ai_1 _32422_ (.B1(net4037),
    .Y(_09400_),
    .A1(net4623),
    .A2(net1851));
 sg13g2_o21ai_1 _32423_ (.B1(_09390_),
    .Y(_01472_),
    .A1(_09399_),
    .A2(_09400_));
 sg13g2_nand2_1 _32424_ (.Y(_09401_),
    .A(net2083),
    .B(net3983));
 sg13g2_a21o_1 _32425_ (.A2(_10721_),
    .A1(\u_inv.f_next[169] ),
    .B1(_09392_),
    .X(_09402_));
 sg13g2_nand2_1 _32426_ (.Y(_09403_),
    .A(_11780_),
    .B(_09402_));
 sg13g2_o21ai_1 _32427_ (.B1(net3815),
    .Y(_09404_),
    .A1(_11780_),
    .A2(_09402_));
 sg13g2_nor2b_1 _32428_ (.A(_09404_),
    .B_N(_09403_),
    .Y(_09405_));
 sg13g2_o21ai_1 _32429_ (.B1(_12375_),
    .Y(_09406_),
    .A1(_12352_),
    .A2(_09383_));
 sg13g2_xnor2_1 _32430_ (.Y(_09407_),
    .A(_11779_),
    .B(_09406_));
 sg13g2_o21ai_1 _32431_ (.B1(net3862),
    .Y(_09408_),
    .A1(\u_inv.f_next[170] ),
    .A2(net4707));
 sg13g2_a21oi_1 _32432_ (.A1(net4707),
    .A2(_09407_),
    .Y(_09409_),
    .B1(_09408_));
 sg13g2_nor3_1 _32433_ (.A(net4448),
    .B(_09405_),
    .C(_09409_),
    .Y(_09410_));
 sg13g2_o21ai_1 _32434_ (.B1(net4036),
    .Y(_09411_),
    .A1(net4624),
    .A2(net1975));
 sg13g2_o21ai_1 _32435_ (.B1(_09401_),
    .Y(_01473_),
    .A1(_09410_),
    .A2(_09411_));
 sg13g2_nand2b_1 _32436_ (.Y(_09412_),
    .B(_09403_),
    .A_N(_11890_));
 sg13g2_a21oi_1 _32437_ (.A1(_11777_),
    .A2(_09412_),
    .Y(_09413_),
    .B1(net3687));
 sg13g2_o21ai_1 _32438_ (.B1(_09413_),
    .Y(_09414_),
    .A1(_11777_),
    .A2(_09412_));
 sg13g2_a21oi_1 _32439_ (.A1(_11779_),
    .A2(_09406_),
    .Y(_09415_),
    .B1(_11778_));
 sg13g2_or2_1 _32440_ (.X(_09416_),
    .B(_09415_),
    .A(_11776_));
 sg13g2_a21oi_1 _32441_ (.A1(_11776_),
    .A2(_09415_),
    .Y(_09417_),
    .B1(net4592));
 sg13g2_a221oi_1 _32442_ (.B2(_09417_),
    .C1(net3709),
    .B1(_09416_),
    .A1(_10410_),
    .Y(_09418_),
    .A2(net4592));
 sg13g2_a21oi_1 _32443_ (.A1(net4521),
    .A2(net2426),
    .Y(_09419_),
    .B1(net3982));
 sg13g2_nor2b_1 _32444_ (.A(_09418_),
    .B_N(_09419_),
    .Y(_09420_));
 sg13g2_a22oi_1 _32445_ (.Y(_01474_),
    .B1(_09414_),
    .B2(_09420_),
    .A2(net3982),
    .A1(_10411_));
 sg13g2_a21oi_2 _32446_ (.B1(_12378_),
    .Y(_09421_),
    .A2(_09406_),
    .A1(_12353_));
 sg13g2_xnor2_1 _32447_ (.Y(_09422_),
    .A(_11774_),
    .B(_09421_));
 sg13g2_a21oi_1 _32448_ (.A1(net2429),
    .A2(net4592),
    .Y(_09423_),
    .B1(net3709));
 sg13g2_o21ai_1 _32449_ (.B1(_09423_),
    .Y(_09424_),
    .A1(net4593),
    .A2(_09422_));
 sg13g2_o21ai_1 _32450_ (.B1(_11893_),
    .Y(_09425_),
    .A1(_11786_),
    .A2(_09380_));
 sg13g2_and2_1 _32451_ (.A(_11774_),
    .B(_09425_),
    .X(_09426_));
 sg13g2_xnor2_1 _32452_ (.Y(_09427_),
    .A(_11774_),
    .B(_09425_));
 sg13g2_o21ai_1 _32453_ (.B1(net4035),
    .Y(_09428_),
    .A1(net4624),
    .A2(net1848));
 sg13g2_a21oi_1 _32454_ (.A1(net3699),
    .A2(_09427_),
    .Y(_09429_),
    .B1(_09428_));
 sg13g2_nand2_1 _32455_ (.Y(_09430_),
    .A(_09424_),
    .B(_09429_));
 sg13g2_o21ai_1 _32456_ (.B1(_09430_),
    .Y(_01475_),
    .A1(_10410_),
    .A2(net4036));
 sg13g2_nand2_1 _32457_ (.Y(_09431_),
    .A(net2429),
    .B(net3980));
 sg13g2_o21ai_1 _32458_ (.B1(_11773_),
    .Y(_09432_),
    .A1(_11774_),
    .A2(_09421_));
 sg13g2_or2_1 _32459_ (.X(_09433_),
    .B(_09432_),
    .A(_11772_));
 sg13g2_a21oi_1 _32460_ (.A1(_11772_),
    .A2(_09432_),
    .Y(_09434_),
    .B1(net4591));
 sg13g2_a221oi_1 _32461_ (.B2(_09434_),
    .C1(net3815),
    .B1(_09433_),
    .A1(_10408_),
    .Y(_09435_),
    .A2(net4591));
 sg13g2_nor3_1 _32462_ (.A(_11772_),
    .B(_11894_),
    .C(_09426_),
    .Y(_09436_));
 sg13g2_and2_1 _32463_ (.A(_11772_),
    .B(_09426_),
    .X(_09437_));
 sg13g2_nand2_1 _32464_ (.Y(_09438_),
    .A(_11895_),
    .B(net3815));
 sg13g2_nor3_1 _32465_ (.A(_09436_),
    .B(_09437_),
    .C(_09438_),
    .Y(_09439_));
 sg13g2_nor3_1 _32466_ (.A(net4448),
    .B(_09435_),
    .C(_09439_),
    .Y(_09440_));
 sg13g2_o21ai_1 _32467_ (.B1(net4035),
    .Y(_09441_),
    .A1(net4624),
    .A2(net2056));
 sg13g2_o21ai_1 _32468_ (.B1(_09431_),
    .Y(_01476_),
    .A1(_09440_),
    .A2(_09441_));
 sg13g2_nor2_1 _32469_ (.A(_11896_),
    .B(_09437_),
    .Y(_09442_));
 sg13g2_or2_1 _32470_ (.X(_09443_),
    .B(_09442_),
    .A(_11770_));
 sg13g2_xnor2_1 _32471_ (.Y(_09444_),
    .A(_11770_),
    .B(_09442_));
 sg13g2_o21ai_1 _32472_ (.B1(_12369_),
    .Y(_09445_),
    .A1(_12350_),
    .A2(_09421_));
 sg13g2_a21oi_1 _32473_ (.A1(_11770_),
    .A2(_09445_),
    .Y(_09446_),
    .B1(net4591));
 sg13g2_o21ai_1 _32474_ (.B1(_09446_),
    .Y(_09447_),
    .A1(_11770_),
    .A2(_09445_));
 sg13g2_a21oi_1 _32475_ (.A1(net2630),
    .A2(net4591),
    .Y(_09448_),
    .B1(net3709));
 sg13g2_o21ai_1 _32476_ (.B1(net4035),
    .Y(_09449_),
    .A1(net4623),
    .A2(net2173));
 sg13g2_a221oi_1 _32477_ (.B2(_09448_),
    .C1(_09449_),
    .B1(_09447_),
    .A1(net3699),
    .Y(_09450_),
    .A2(_09444_));
 sg13g2_a21o_1 _32478_ (.A2(net3981),
    .A1(net2202),
    .B1(_09450_),
    .X(_01477_));
 sg13g2_a21oi_1 _32479_ (.A1(_11897_),
    .A2(_09443_),
    .Y(_09451_),
    .B1(_11768_));
 sg13g2_nand3_1 _32480_ (.B(_11897_),
    .C(_09443_),
    .A(_11768_),
    .Y(_09452_));
 sg13g2_nor2_1 _32481_ (.A(net3687),
    .B(_09451_),
    .Y(_09453_));
 sg13g2_a21oi_1 _32482_ (.A1(_11770_),
    .A2(_09445_),
    .Y(_09454_),
    .B1(_11769_));
 sg13g2_xor2_1 _32483_ (.B(_09454_),
    .A(_11768_),
    .X(_09455_));
 sg13g2_o21ai_1 _32484_ (.B1(net3720),
    .Y(_09456_),
    .A1(net2191),
    .A2(net4704));
 sg13g2_a21o_1 _32485_ (.A2(_09455_),
    .A1(net4704),
    .B1(_09456_),
    .X(_09457_));
 sg13g2_a221oi_1 _32486_ (.B2(_09453_),
    .C1(net3980),
    .B1(_09452_),
    .A1(net4521),
    .Y(_09458_),
    .A2(net2461));
 sg13g2_a22oi_1 _32487_ (.Y(_01478_),
    .B1(_09457_),
    .B2(_09458_),
    .A2(net3980),
    .A1(_10407_));
 sg13g2_nand2_1 _32488_ (.Y(_09459_),
    .A(net2191),
    .B(net3980));
 sg13g2_a21oi_2 _32489_ (.B1(_11804_),
    .Y(_09460_),
    .A2(_09293_),
    .A1(_11873_));
 sg13g2_nor2_1 _32490_ (.A(_11902_),
    .B(_09460_),
    .Y(_09461_));
 sg13g2_or2_1 _32491_ (.X(_09462_),
    .B(_09461_),
    .A(_11759_));
 sg13g2_a21oi_1 _32492_ (.A1(_11759_),
    .A2(_09461_),
    .Y(_09463_),
    .B1(net3856));
 sg13g2_nor3_1 _32493_ (.A(net4432),
    .B(_12460_),
    .C(_09299_),
    .Y(_09464_));
 sg13g2_nand2b_2 _32494_ (.Y(_09465_),
    .B(_12381_),
    .A_N(_09464_));
 sg13g2_nand2_1 _32495_ (.Y(_09466_),
    .A(_11759_),
    .B(_09465_));
 sg13g2_xnor2_1 _32496_ (.Y(_09467_),
    .A(_11759_),
    .B(_09465_));
 sg13g2_nor2_1 _32497_ (.A(\u_inv.f_next[176] ),
    .B(net4695),
    .Y(_09468_));
 sg13g2_a21oi_1 _32498_ (.A1(net4695),
    .A2(_09467_),
    .Y(_09469_),
    .B1(_09468_));
 sg13g2_a221oi_1 _32499_ (.B2(net3856),
    .C1(net4445),
    .B1(_09469_),
    .A1(_09462_),
    .Y(_09470_),
    .A2(_09463_));
 sg13g2_o21ai_1 _32500_ (.B1(net4035),
    .Y(_09471_),
    .A1(net4623),
    .A2(net1898));
 sg13g2_o21ai_1 _32501_ (.B1(_09459_),
    .Y(_01479_),
    .A1(_09470_),
    .A2(_09471_));
 sg13g2_nand2_1 _32502_ (.Y(_09472_),
    .A(net2044),
    .B(net3972));
 sg13g2_o21ai_1 _32503_ (.B1(_09466_),
    .Y(_09473_),
    .A1(_10405_),
    .A2(_10714_));
 sg13g2_xnor2_1 _32504_ (.Y(_09474_),
    .A(_11760_),
    .B(_09473_));
 sg13g2_nor2_1 _32505_ (.A(\u_inv.f_next[177] ),
    .B(net4695),
    .Y(_09475_));
 sg13g2_a21oi_1 _32506_ (.A1(net4695),
    .A2(_09474_),
    .Y(_09476_),
    .B1(_09475_));
 sg13g2_and2_1 _32507_ (.A(_11760_),
    .B(_11922_),
    .X(_09477_));
 sg13g2_nor2_1 _32508_ (.A(_11760_),
    .B(_09462_),
    .Y(_09478_));
 sg13g2_a21oi_1 _32509_ (.A1(_09462_),
    .A2(_09477_),
    .Y(_09479_),
    .B1(net3856));
 sg13g2_a21o_1 _32510_ (.A2(_09462_),
    .A1(_11922_),
    .B1(_11760_),
    .X(_09480_));
 sg13g2_a221oi_1 _32511_ (.B2(_09480_),
    .C1(net4449),
    .B1(_09479_),
    .A1(net3856),
    .Y(_09481_),
    .A2(_09476_));
 sg13g2_o21ai_1 _32512_ (.B1(net4031),
    .Y(_09482_),
    .A1(net4621),
    .A2(net1995));
 sg13g2_o21ai_1 _32513_ (.B1(_09472_),
    .Y(_01480_),
    .A1(_09481_),
    .A2(_09482_));
 sg13g2_nand2_1 _32514_ (.Y(_09483_),
    .A(net2231),
    .B(net3972));
 sg13g2_or2_1 _32515_ (.X(_09484_),
    .B(_09478_),
    .A(_11923_));
 sg13g2_o21ai_1 _32516_ (.B1(net3802),
    .Y(_09485_),
    .A1(net4433),
    .A2(_09484_));
 sg13g2_a21oi_1 _32517_ (.A1(net4433),
    .A2(_09484_),
    .Y(_09486_),
    .B1(_09485_));
 sg13g2_a21oi_2 _32518_ (.B1(_12323_),
    .Y(_09487_),
    .A2(_09465_),
    .A1(_12346_));
 sg13g2_xnor2_1 _32519_ (.Y(_09488_),
    .A(net4433),
    .B(_09487_));
 sg13g2_o21ai_1 _32520_ (.B1(net3856),
    .Y(_09489_),
    .A1(\u_inv.f_next[178] ),
    .A2(net4695));
 sg13g2_a21oi_1 _32521_ (.A1(net4695),
    .A2(_09488_),
    .Y(_09490_),
    .B1(_09489_));
 sg13g2_nor3_1 _32522_ (.A(net4449),
    .B(_09486_),
    .C(_09490_),
    .Y(_09491_));
 sg13g2_o21ai_1 _32523_ (.B1(net4032),
    .Y(_09492_),
    .A1(net4621),
    .A2(\u_inv.input_reg[177] ));
 sg13g2_o21ai_1 _32524_ (.B1(_09483_),
    .Y(_01481_),
    .A1(_09491_),
    .A2(_09492_));
 sg13g2_a21oi_1 _32525_ (.A1(_11763_),
    .A2(_09484_),
    .Y(_09493_),
    .B1(_11920_));
 sg13g2_xor2_1 _32526_ (.B(_09493_),
    .A(_11764_),
    .X(_09494_));
 sg13g2_nand2_1 _32527_ (.Y(_09495_),
    .A(net2671),
    .B(net3856));
 sg13g2_o21ai_1 _32528_ (.B1(_11762_),
    .Y(_09496_),
    .A1(net4433),
    .A2(_09487_));
 sg13g2_xor2_1 _32529_ (.B(_09496_),
    .A(_11764_),
    .X(_09497_));
 sg13g2_a22oi_1 _32530_ (.Y(_09498_),
    .B1(_09497_),
    .B2(net4695),
    .A2(_09495_),
    .A1(net3731));
 sg13g2_o21ai_1 _32531_ (.B1(net4383),
    .Y(_09499_),
    .A1(net3856),
    .A2(_09494_));
 sg13g2_a21oi_1 _32532_ (.A1(net4518),
    .A2(_10982_),
    .Y(_09500_),
    .B1(net3973));
 sg13g2_o21ai_1 _32533_ (.B1(_09500_),
    .Y(_09501_),
    .A1(_09498_),
    .A2(_09499_));
 sg13g2_o21ai_1 _32534_ (.B1(_09501_),
    .Y(_01482_),
    .A1(_10403_),
    .A2(net4031));
 sg13g2_o21ai_1 _32535_ (.B1(_12326_),
    .Y(_09502_),
    .A1(_12321_),
    .A2(_09487_));
 sg13g2_a21oi_1 _32536_ (.A1(_11755_),
    .A2(_09502_),
    .Y(_09503_),
    .B1(net4581));
 sg13g2_o21ai_1 _32537_ (.B1(_09503_),
    .Y(_09504_),
    .A1(_11755_),
    .A2(_09502_));
 sg13g2_a21oi_1 _32538_ (.A1(net2497),
    .A2(net4581),
    .Y(_09505_),
    .B1(net3706));
 sg13g2_o21ai_1 _32539_ (.B1(_11765_),
    .Y(_09506_),
    .A1(_11902_),
    .A2(_09460_));
 sg13g2_nand2_1 _32540_ (.Y(_09507_),
    .A(_11925_),
    .B(_09506_));
 sg13g2_a21oi_1 _32541_ (.A1(_11925_),
    .A2(_09506_),
    .Y(_09508_),
    .B1(_11755_));
 sg13g2_xnor2_1 _32542_ (.Y(_09509_),
    .A(_11756_),
    .B(_09507_));
 sg13g2_o21ai_1 _32543_ (.B1(net4031),
    .Y(_09510_),
    .A1(net4621),
    .A2(net2023));
 sg13g2_a221oi_1 _32544_ (.B2(net3696),
    .C1(_09510_),
    .B1(_09509_),
    .A1(_09504_),
    .Y(_09511_),
    .A2(_09505_));
 sg13g2_a21o_1 _32545_ (.A2(net3972),
    .A1(net2671),
    .B1(_09511_),
    .X(_01483_));
 sg13g2_a21oi_1 _32546_ (.A1(_11755_),
    .A2(_09502_),
    .Y(_09512_),
    .B1(_11754_));
 sg13g2_xnor2_1 _32547_ (.Y(_09513_),
    .A(_11757_),
    .B(_09512_));
 sg13g2_a21oi_1 _32548_ (.A1(net2616),
    .A2(net4581),
    .Y(_09514_),
    .B1(net3706));
 sg13g2_o21ai_1 _32549_ (.B1(_09514_),
    .Y(_09515_),
    .A1(net4581),
    .A2(_09513_));
 sg13g2_o21ai_1 _32550_ (.B1(_11757_),
    .Y(_09516_),
    .A1(_11928_),
    .A2(_09508_));
 sg13g2_or3_1 _32551_ (.A(_11757_),
    .B(_11928_),
    .C(_09508_),
    .X(_09517_));
 sg13g2_nand2_1 _32552_ (.Y(_09518_),
    .A(_09516_),
    .B(_09517_));
 sg13g2_o21ai_1 _32553_ (.B1(net4031),
    .Y(_09519_),
    .A1(net4621),
    .A2(net1953));
 sg13g2_a21oi_1 _32554_ (.A1(net3696),
    .A2(_09518_),
    .Y(_09520_),
    .B1(_09519_));
 sg13g2_nand2_1 _32555_ (.Y(_09521_),
    .A(_09515_),
    .B(_09520_));
 sg13g2_o21ai_1 _32556_ (.B1(_09521_),
    .Y(_01484_),
    .A1(_10401_),
    .A2(net4031));
 sg13g2_nand3_1 _32557_ (.B(_11927_),
    .C(_09516_),
    .A(_11752_),
    .Y(_09522_));
 sg13g2_a21o_1 _32558_ (.A2(_09516_),
    .A1(_11927_),
    .B1(_11752_),
    .X(_09523_));
 sg13g2_nand3_1 _32559_ (.B(_09522_),
    .C(_09523_),
    .A(net3802),
    .Y(_09524_));
 sg13g2_a21oi_1 _32560_ (.A1(_12319_),
    .A2(_09502_),
    .Y(_09525_),
    .B1(_12331_));
 sg13g2_xnor2_1 _32561_ (.Y(_09526_),
    .A(_11753_),
    .B(_09525_));
 sg13g2_a21oi_1 _32562_ (.A1(net4697),
    .A2(_09526_),
    .Y(_09527_),
    .B1(net3802));
 sg13g2_o21ai_1 _32563_ (.B1(_09527_),
    .Y(_09528_),
    .A1(\u_inv.f_next[182] ),
    .A2(net4697));
 sg13g2_nand3_1 _32564_ (.B(_09524_),
    .C(_09528_),
    .A(net4383),
    .Y(_09529_));
 sg13g2_o21ai_1 _32565_ (.B1(_09529_),
    .Y(_09530_),
    .A1(net4621),
    .A2(net2076));
 sg13g2_nor2_1 _32566_ (.A(net2616),
    .B(net4031),
    .Y(_09531_));
 sg13g2_a21oi_1 _32567_ (.A1(net4030),
    .A2(_09530_),
    .Y(_01485_),
    .B1(_09531_));
 sg13g2_a21oi_1 _32568_ (.A1(_11930_),
    .A2(_09523_),
    .Y(_09532_),
    .B1(_11749_));
 sg13g2_nand3_1 _32569_ (.B(_11930_),
    .C(_09523_),
    .A(_11749_),
    .Y(_09533_));
 sg13g2_nor2_1 _32570_ (.A(net3684),
    .B(_09532_),
    .Y(_09534_));
 sg13g2_o21ai_1 _32571_ (.B1(_11751_),
    .Y(_09535_),
    .A1(_11753_),
    .A2(_09525_));
 sg13g2_xnor2_1 _32572_ (.Y(_09536_),
    .A(_11749_),
    .B(_09535_));
 sg13g2_o21ai_1 _32573_ (.B1(net3721),
    .Y(_09537_),
    .A1(net2366),
    .A2(net4697));
 sg13g2_a21o_1 _32574_ (.A2(_09536_),
    .A1(net4697),
    .B1(_09537_),
    .X(_09538_));
 sg13g2_a221oi_1 _32575_ (.B2(_09534_),
    .C1(net3972),
    .B1(_09533_),
    .A1(net4518),
    .Y(_09539_),
    .A2(net2651));
 sg13g2_a22oi_1 _32576_ (.Y(_01486_),
    .B1(_09538_),
    .B2(_09539_),
    .A2(net3972),
    .A1(_10399_));
 sg13g2_nand2_1 _32577_ (.Y(_09540_),
    .A(net2366),
    .B(net3972));
 sg13g2_o21ai_1 _32578_ (.B1(_11934_),
    .Y(_09541_),
    .A1(_11758_),
    .A2(_09506_));
 sg13g2_nor2_1 _32579_ (.A(_11744_),
    .B(_09541_),
    .Y(_09542_));
 sg13g2_nand2_1 _32580_ (.Y(_09543_),
    .A(_11744_),
    .B(_09541_));
 sg13g2_nor2_1 _32581_ (.A(net3855),
    .B(_09542_),
    .Y(_09544_));
 sg13g2_a21oi_2 _32582_ (.B1(_12334_),
    .Y(_09545_),
    .A2(_09465_),
    .A1(_12347_));
 sg13g2_nor2_1 _32583_ (.A(_11744_),
    .B(_09545_),
    .Y(_09546_));
 sg13g2_xnor2_1 _32584_ (.Y(_09547_),
    .A(_11744_),
    .B(_09545_));
 sg13g2_nand2_1 _32585_ (.Y(_09548_),
    .A(_10397_),
    .B(net4582));
 sg13g2_a21oi_1 _32586_ (.A1(net4693),
    .A2(_09547_),
    .Y(_09549_),
    .B1(net3799));
 sg13g2_a221oi_1 _32587_ (.B2(_09549_),
    .C1(net4445),
    .B1(_09548_),
    .A1(_09543_),
    .Y(_09550_),
    .A2(_09544_));
 sg13g2_o21ai_1 _32588_ (.B1(net4031),
    .Y(_09551_),
    .A1(net4621),
    .A2(net2189));
 sg13g2_o21ai_1 _32589_ (.B1(_09540_),
    .Y(_01487_),
    .A1(_09550_),
    .A2(_09551_));
 sg13g2_nand2_1 _32590_ (.Y(_09552_),
    .A(net2151),
    .B(net3971));
 sg13g2_a21o_1 _32591_ (.A2(_09543_),
    .A1(_11906_),
    .B1(_11745_),
    .X(_09553_));
 sg13g2_nand3_1 _32592_ (.B(_11906_),
    .C(_09543_),
    .A(_11745_),
    .Y(_09554_));
 sg13g2_o21ai_1 _32593_ (.B1(net4030),
    .Y(_09555_),
    .A1(net4620),
    .A2(net1891));
 sg13g2_a21oi_1 _32594_ (.A1(\u_inv.f_next[184] ),
    .A2(\u_inv.f_reg[184] ),
    .Y(_09556_),
    .B1(_09546_));
 sg13g2_and3_1 _32595_ (.X(_09557_),
    .A(net3799),
    .B(_09553_),
    .C(_09554_));
 sg13g2_nand2_1 _32596_ (.Y(_09558_),
    .A(\u_inv.f_next[185] ),
    .B(net3855));
 sg13g2_xor2_1 _32597_ (.B(_09556_),
    .A(_11745_),
    .X(_09559_));
 sg13g2_a22oi_1 _32598_ (.Y(_09560_),
    .B1(_09559_),
    .B2(net4693),
    .A2(_09558_),
    .A1(net3730));
 sg13g2_nor3_1 _32599_ (.A(net4445),
    .B(_09557_),
    .C(_09560_),
    .Y(_09561_));
 sg13g2_o21ai_1 _32600_ (.B1(_09552_),
    .Y(_01488_),
    .A1(_09555_),
    .A2(_09561_));
 sg13g2_nand2_1 _32601_ (.Y(_09562_),
    .A(net2175),
    .B(net3971));
 sg13g2_nand2_1 _32602_ (.Y(_09563_),
    .A(_11905_),
    .B(_09553_));
 sg13g2_and2_1 _32603_ (.A(_11743_),
    .B(_09563_),
    .X(_09564_));
 sg13g2_o21ai_1 _32604_ (.B1(net3799),
    .Y(_09565_),
    .A1(_11743_),
    .A2(_09563_));
 sg13g2_a21oi_1 _32605_ (.A1(_11745_),
    .A2(_09546_),
    .Y(_09566_),
    .B1(_12336_));
 sg13g2_xnor2_1 _32606_ (.Y(_09567_),
    .A(_11743_),
    .B(_09566_));
 sg13g2_o21ai_1 _32607_ (.B1(net3855),
    .Y(_09568_),
    .A1(\u_inv.f_next[186] ),
    .A2(net4694));
 sg13g2_a21oi_1 _32608_ (.A1(net4694),
    .A2(_09567_),
    .Y(_09569_),
    .B1(_09568_));
 sg13g2_o21ai_1 _32609_ (.B1(net4386),
    .Y(_09570_),
    .A1(_09564_),
    .A2(_09565_));
 sg13g2_nor2_1 _32610_ (.A(_09569_),
    .B(_09570_),
    .Y(_09571_));
 sg13g2_o21ai_1 _32611_ (.B1(net4030),
    .Y(_09572_),
    .A1(net4620),
    .A2(net1790));
 sg13g2_o21ai_1 _32612_ (.B1(_09562_),
    .Y(_01489_),
    .A1(_09571_),
    .A2(_09572_));
 sg13g2_nor2_1 _32613_ (.A(_11904_),
    .B(_09564_),
    .Y(_09573_));
 sg13g2_a21oi_1 _32614_ (.A1(_11740_),
    .A2(_09573_),
    .Y(_09574_),
    .B1(net3684));
 sg13g2_o21ai_1 _32615_ (.B1(_09574_),
    .Y(_09575_),
    .A1(_11740_),
    .A2(_09573_));
 sg13g2_o21ai_1 _32616_ (.B1(_11742_),
    .Y(_09576_),
    .A1(_11743_),
    .A2(_09566_));
 sg13g2_xnor2_1 _32617_ (.Y(_09577_),
    .A(_11740_),
    .B(_09576_));
 sg13g2_o21ai_1 _32618_ (.B1(net3721),
    .Y(_09578_),
    .A1(net2984),
    .A2(net4694));
 sg13g2_a21oi_1 _32619_ (.A1(net4694),
    .A2(_09577_),
    .Y(_09579_),
    .B1(_09578_));
 sg13g2_a21oi_1 _32620_ (.A1(net4518),
    .A2(net1930),
    .Y(_09580_),
    .B1(net3975));
 sg13g2_nor2b_1 _32621_ (.A(_09579_),
    .B_N(_09580_),
    .Y(_09581_));
 sg13g2_a22oi_1 _32622_ (.Y(_01490_),
    .B1(_09575_),
    .B2(_09581_),
    .A2(net3971),
    .A1(_10395_));
 sg13g2_a21o_1 _32623_ (.A2(_09541_),
    .A1(_11747_),
    .B1(_11909_),
    .X(_09582_));
 sg13g2_and2_1 _32624_ (.A(_11737_),
    .B(_09582_),
    .X(_09583_));
 sg13g2_o21ai_1 _32625_ (.B1(net3799),
    .Y(_09584_),
    .A1(_11737_),
    .A2(_09582_));
 sg13g2_nor3_1 _32626_ (.A(_11744_),
    .B(_12313_),
    .C(_09545_),
    .Y(_09585_));
 sg13g2_nand2b_2 _32627_ (.Y(_09586_),
    .B(_12338_),
    .A_N(_09585_));
 sg13g2_xnor2_1 _32628_ (.Y(_09587_),
    .A(_11736_),
    .B(_09586_));
 sg13g2_o21ai_1 _32629_ (.B1(net3855),
    .Y(_09588_),
    .A1(net2188),
    .A2(net4693));
 sg13g2_a21oi_1 _32630_ (.A1(net4693),
    .A2(_09587_),
    .Y(_09589_),
    .B1(_09588_));
 sg13g2_o21ai_1 _32631_ (.B1(net4386),
    .Y(_09590_),
    .A1(_09583_),
    .A2(_09584_));
 sg13g2_or2_1 _32632_ (.X(_09591_),
    .B(net1716),
    .A(net4620));
 sg13g2_o21ai_1 _32633_ (.B1(_09591_),
    .Y(_09592_),
    .A1(_09589_),
    .A2(_09590_));
 sg13g2_nor2_1 _32634_ (.A(net2984),
    .B(net4030),
    .Y(_09593_));
 sg13g2_a21oi_1 _32635_ (.A1(net4030),
    .A2(_09592_),
    .Y(_01491_),
    .B1(_09593_));
 sg13g2_nand2_1 _32636_ (.Y(_09594_),
    .A(net2188),
    .B(net3971));
 sg13g2_nand2_1 _32637_ (.Y(_09595_),
    .A(net2129),
    .B(net3855));
 sg13g2_a21oi_1 _32638_ (.A1(_11736_),
    .A2(_09586_),
    .Y(_09596_),
    .B1(_11735_));
 sg13g2_xnor2_1 _32639_ (.Y(_09597_),
    .A(_11734_),
    .B(_09596_));
 sg13g2_a22oi_1 _32640_ (.Y(_09598_),
    .B1(_09597_),
    .B2(net4693),
    .A2(_09595_),
    .A1(net3731));
 sg13g2_nor3_1 _32641_ (.A(_11734_),
    .B(_11913_),
    .C(_09583_),
    .Y(_09599_));
 sg13g2_nand2_1 _32642_ (.Y(_09600_),
    .A(_11734_),
    .B(_09583_));
 sg13g2_inv_1 _32643_ (.Y(_09601_),
    .A(_09600_));
 sg13g2_nor4_1 _32644_ (.A(_11914_),
    .B(net3855),
    .C(_09599_),
    .D(_09601_),
    .Y(_09602_));
 sg13g2_nor3_1 _32645_ (.A(net4445),
    .B(_09598_),
    .C(_09602_),
    .Y(_09603_));
 sg13g2_o21ai_1 _32646_ (.B1(net4033),
    .Y(_09604_),
    .A1(net4620),
    .A2(net1868));
 sg13g2_o21ai_1 _32647_ (.B1(_09594_),
    .Y(_01492_),
    .A1(_09603_),
    .A2(_09604_));
 sg13g2_nand2_1 _32648_ (.Y(_09605_),
    .A(net2129),
    .B(net3971));
 sg13g2_nand2_1 _32649_ (.Y(_09606_),
    .A(_11915_),
    .B(_09600_));
 sg13g2_o21ai_1 _32650_ (.B1(net3799),
    .Y(_09607_),
    .A1(_11733_),
    .A2(_09606_));
 sg13g2_a21oi_1 _32651_ (.A1(_11733_),
    .A2(_09606_),
    .Y(_09608_),
    .B1(_09607_));
 sg13g2_a21oi_1 _32652_ (.A1(_12315_),
    .A2(_09586_),
    .Y(_09609_),
    .B1(_12340_));
 sg13g2_xnor2_1 _32653_ (.Y(_09610_),
    .A(_11733_),
    .B(_09609_));
 sg13g2_o21ai_1 _32654_ (.B1(net3855),
    .Y(_09611_),
    .A1(\u_inv.f_next[190] ),
    .A2(net4693));
 sg13g2_a21oi_1 _32655_ (.A1(net4693),
    .A2(_09610_),
    .Y(_09612_),
    .B1(_09611_));
 sg13g2_nor3_1 _32656_ (.A(net4445),
    .B(_09608_),
    .C(_09612_),
    .Y(_09613_));
 sg13g2_o21ai_1 _32657_ (.B1(net4030),
    .Y(_09614_),
    .A1(net4620),
    .A2(net1844));
 sg13g2_o21ai_1 _32658_ (.B1(_09605_),
    .Y(_01493_),
    .A1(_09613_),
    .A2(_09614_));
 sg13g2_nand2_1 _32659_ (.Y(_09615_),
    .A(net2316),
    .B(net3971));
 sg13g2_a21oi_1 _32660_ (.A1(_11733_),
    .A2(_09606_),
    .Y(_09616_),
    .B1(_11912_));
 sg13g2_xor2_1 _32661_ (.B(_09616_),
    .A(_11730_),
    .X(_09617_));
 sg13g2_a21oi_1 _32662_ (.A1(_10390_),
    .A2(net4582),
    .Y(_09618_),
    .B1(net3799));
 sg13g2_o21ai_1 _32663_ (.B1(_11731_),
    .Y(_09619_),
    .A1(_11733_),
    .A2(_09609_));
 sg13g2_xnor2_1 _32664_ (.Y(_09620_),
    .A(_11730_),
    .B(_09619_));
 sg13g2_nand2_1 _32665_ (.Y(_09621_),
    .A(net4693),
    .B(_09620_));
 sg13g2_a221oi_1 _32666_ (.B2(_09621_),
    .C1(net4445),
    .B1(_09618_),
    .A1(net3803),
    .Y(_09622_),
    .A2(_09617_));
 sg13g2_o21ai_1 _32667_ (.B1(net4033),
    .Y(_09623_),
    .A1(net4620),
    .A2(net1982));
 sg13g2_o21ai_1 _32668_ (.B1(_09615_),
    .Y(_01494_),
    .A1(_09622_),
    .A2(_09623_));
 sg13g2_a21oi_1 _32669_ (.A1(_11939_),
    .A2(_12000_),
    .Y(_09624_),
    .B1(net3683));
 sg13g2_o21ai_1 _32670_ (.B1(_09624_),
    .Y(_09625_),
    .A1(_11939_),
    .A2(_12000_));
 sg13g2_a21oi_1 _32671_ (.A1(net4517),
    .A2(net2121),
    .Y(_09626_),
    .B1(net3960));
 sg13g2_nand2_1 _32672_ (.Y(_09627_),
    .A(_11999_),
    .B(_12755_));
 sg13g2_xnor2_1 _32673_ (.Y(_09628_),
    .A(_11999_),
    .B(_12755_));
 sg13g2_o21ai_1 _32674_ (.B1(net3716),
    .Y(_09629_),
    .A1(net2242),
    .A2(net4676));
 sg13g2_a21oi_2 _32675_ (.B1(_09629_),
    .Y(_09630_),
    .A2(_09628_),
    .A1(net4676));
 sg13g2_nor2b_1 _32676_ (.A(_09630_),
    .B_N(_09626_),
    .Y(_09631_));
 sg13g2_a22oi_1 _32677_ (.Y(_01495_),
    .B1(_09625_),
    .B2(_09631_),
    .A2(net3960),
    .A1(_10390_));
 sg13g2_nand2_1 _32678_ (.Y(_09632_),
    .A(net2242),
    .B(net3951));
 sg13g2_a21oi_1 _32679_ (.A1(_11939_),
    .A2(_12000_),
    .Y(_09633_),
    .B1(_12020_));
 sg13g2_o21ai_1 _32680_ (.B1(net3775),
    .Y(_09634_),
    .A1(_12001_),
    .A2(_09633_));
 sg13g2_a21oi_1 _32681_ (.A1(_12001_),
    .A2(_09633_),
    .Y(_09635_),
    .B1(_09634_));
 sg13g2_nand2_1 _32682_ (.Y(_09636_),
    .A(\u_inv.f_next[193] ),
    .B(net3845));
 sg13g2_o21ai_1 _32683_ (.B1(_09627_),
    .Y(_09637_),
    .A1(_10389_),
    .A2(_10698_));
 sg13g2_xnor2_1 _32684_ (.Y(_09638_),
    .A(_12001_),
    .B(_09637_));
 sg13g2_a22oi_1 _32685_ (.Y(_09639_),
    .B1(_09638_),
    .B2(net4677),
    .A2(_09636_),
    .A1(net3727));
 sg13g2_nor3_1 _32686_ (.A(net4443),
    .B(_09635_),
    .C(_09639_),
    .Y(_09640_));
 sg13g2_o21ai_1 _32687_ (.B1(net4023),
    .Y(_09641_),
    .A1(net4615),
    .A2(net2238));
 sg13g2_o21ai_1 _32688_ (.B1(_09632_),
    .Y(_01496_),
    .A1(_09640_),
    .A2(_09641_));
 sg13g2_o21ai_1 _32689_ (.B1(_12019_),
    .Y(_09642_),
    .A1(_12001_),
    .A2(_09633_));
 sg13g2_xor2_1 _32690_ (.B(_09642_),
    .A(_11997_),
    .X(_09643_));
 sg13g2_nand2_1 _32691_ (.Y(_09644_),
    .A(net3693),
    .B(_09643_));
 sg13g2_a21oi_2 _32692_ (.B1(_12259_),
    .Y(_09645_),
    .A2(_12756_),
    .A1(_12755_));
 sg13g2_a21oi_1 _32693_ (.A1(_11997_),
    .A2(_09645_),
    .Y(_09646_),
    .B1(net4556));
 sg13g2_o21ai_1 _32694_ (.B1(_09646_),
    .Y(_09647_),
    .A1(_11997_),
    .A2(_09645_));
 sg13g2_o21ai_1 _32695_ (.B1(_09647_),
    .Y(_09648_),
    .A1(_10387_),
    .A2(net4677));
 sg13g2_a221oi_1 _32696_ (.B2(_09648_),
    .C1(net3950),
    .B1(net3716),
    .A1(net4513),
    .Y(_09649_),
    .A2(net2305));
 sg13g2_a22oi_1 _32697_ (.Y(_01497_),
    .B1(_09644_),
    .B2(_09649_),
    .A2(net3950),
    .A1(_10388_));
 sg13g2_o21ai_1 _32698_ (.B1(_11996_),
    .Y(_09650_),
    .A1(_11997_),
    .A2(_09645_));
 sg13g2_xnor2_1 _32699_ (.Y(_09651_),
    .A(_11995_),
    .B(_09650_));
 sg13g2_o21ai_1 _32700_ (.B1(net4381),
    .Y(_09652_),
    .A1(_10386_),
    .A2(net4677));
 sg13g2_a21oi_1 _32701_ (.A1(net4677),
    .A2(_09651_),
    .Y(_09653_),
    .B1(_09652_));
 sg13g2_a21o_1 _32702_ (.A2(_09642_),
    .A1(_11997_),
    .B1(_12018_),
    .X(_09654_));
 sg13g2_a21oi_1 _32703_ (.A1(_11995_),
    .A2(_09654_),
    .Y(_09655_),
    .B1(net3845));
 sg13g2_o21ai_1 _32704_ (.B1(_09655_),
    .Y(_09656_),
    .A1(_11995_),
    .A2(_09654_));
 sg13g2_o21ai_1 _32705_ (.B1(_09656_),
    .Y(_09657_),
    .A1(net3700),
    .A2(_09653_));
 sg13g2_o21ai_1 _32706_ (.B1(net4023),
    .Y(_09658_),
    .A1(net4615),
    .A2(net2462));
 sg13g2_nand2b_1 _32707_ (.Y(_09659_),
    .B(_09657_),
    .A_N(_09658_));
 sg13g2_o21ai_1 _32708_ (.B1(_09659_),
    .Y(_01498_),
    .A1(_10387_),
    .A2(net4023));
 sg13g2_nor2_1 _32709_ (.A(_12257_),
    .B(_09645_),
    .Y(_09660_));
 sg13g2_nor2_1 _32710_ (.A(_12262_),
    .B(_09660_),
    .Y(_09661_));
 sg13g2_inv_2 _32711_ (.Y(_09662_),
    .A(_09661_));
 sg13g2_a21oi_1 _32712_ (.A1(_12011_),
    .A2(_09662_),
    .Y(_09663_),
    .B1(net4555));
 sg13g2_o21ai_1 _32713_ (.B1(_09663_),
    .Y(_09664_),
    .A1(_12011_),
    .A2(_09662_));
 sg13g2_a21oi_1 _32714_ (.A1(net1770),
    .A2(net4555),
    .Y(_09665_),
    .B1(net3704));
 sg13g2_a21oi_1 _32715_ (.A1(_11939_),
    .A2(_12002_),
    .Y(_09666_),
    .B1(_12025_));
 sg13g2_or2_1 _32716_ (.X(_09667_),
    .B(_09666_),
    .A(_12011_));
 sg13g2_xnor2_1 _32717_ (.Y(_09668_),
    .A(_12011_),
    .B(_09666_));
 sg13g2_o21ai_1 _32718_ (.B1(net4022),
    .Y(_09669_),
    .A1(net4615),
    .A2(net2201));
 sg13g2_a221oi_1 _32719_ (.B2(net3693),
    .C1(_09669_),
    .B1(_09668_),
    .A1(_09664_),
    .Y(_09670_),
    .A2(_09665_));
 sg13g2_a21o_1 _32720_ (.A2(net3950),
    .A1(net2440),
    .B1(_09670_),
    .X(_01499_));
 sg13g2_nand2_1 _32721_ (.Y(_09671_),
    .A(net1770),
    .B(net3949));
 sg13g2_nand2_1 _32722_ (.Y(_09672_),
    .A(net1704),
    .B(net3843));
 sg13g2_a21oi_1 _32723_ (.A1(_12011_),
    .A2(_09662_),
    .Y(_09673_),
    .B1(_12010_));
 sg13g2_xor2_1 _32724_ (.B(_09673_),
    .A(_12009_),
    .X(_09674_));
 sg13g2_a22oi_1 _32725_ (.Y(_09675_),
    .B1(_09674_),
    .B2(net4675),
    .A2(_09672_),
    .A1(net3727));
 sg13g2_a21oi_1 _32726_ (.A1(_12017_),
    .A2(_09667_),
    .Y(_09676_),
    .B1(_12009_));
 sg13g2_and3_1 _32727_ (.X(_09677_),
    .A(_12009_),
    .B(_12017_),
    .C(_09667_));
 sg13g2_nor3_1 _32728_ (.A(net3843),
    .B(_09676_),
    .C(_09677_),
    .Y(_09678_));
 sg13g2_nor3_1 _32729_ (.A(net4442),
    .B(_09675_),
    .C(_09678_),
    .Y(_09679_));
 sg13g2_o21ai_1 _32730_ (.B1(net4022),
    .Y(_09680_),
    .A1(net4613),
    .A2(\u_inv.input_reg[196] ));
 sg13g2_o21ai_1 _32731_ (.B1(_09671_),
    .Y(_01500_),
    .A1(_09679_),
    .A2(_09680_));
 sg13g2_nand2_1 _32732_ (.Y(_09681_),
    .A(net1704),
    .B(net3949));
 sg13g2_or2_1 _32733_ (.X(_09682_),
    .B(_09676_),
    .A(_12016_));
 sg13g2_o21ai_1 _32734_ (.B1(net3774),
    .Y(_09683_),
    .A1(_12007_),
    .A2(_09682_));
 sg13g2_a21oi_1 _32735_ (.A1(_12007_),
    .A2(_09682_),
    .Y(_09684_),
    .B1(_09683_));
 sg13g2_a21oi_1 _32736_ (.A1(_12255_),
    .A2(_09662_),
    .Y(_09685_),
    .B1(_12266_));
 sg13g2_nor2_1 _32737_ (.A(_12007_),
    .B(_09685_),
    .Y(_09686_));
 sg13g2_xnor2_1 _32738_ (.Y(_09687_),
    .A(_12007_),
    .B(_09685_));
 sg13g2_o21ai_1 _32739_ (.B1(net3843),
    .Y(_09688_),
    .A1(net1627),
    .A2(net4675));
 sg13g2_a21oi_1 _32740_ (.A1(net4675),
    .A2(_09687_),
    .Y(_09689_),
    .B1(_09688_));
 sg13g2_nor3_1 _32741_ (.A(net4442),
    .B(_09684_),
    .C(_09689_),
    .Y(_09690_));
 sg13g2_o21ai_1 _32742_ (.B1(net4020),
    .Y(_09691_),
    .A1(net4613),
    .A2(\u_inv.input_reg[197] ));
 sg13g2_o21ai_1 _32743_ (.B1(_09681_),
    .Y(_01501_),
    .A1(_09690_),
    .A2(_09691_));
 sg13g2_nand2_1 _32744_ (.Y(_09692_),
    .A(net1627),
    .B(net3949));
 sg13g2_a21oi_1 _32745_ (.A1(_12007_),
    .A2(_09682_),
    .Y(_09693_),
    .B1(_12029_));
 sg13g2_o21ai_1 _32746_ (.B1(net3774),
    .Y(_09694_),
    .A1(_12004_),
    .A2(_09693_));
 sg13g2_a21oi_1 _32747_ (.A1(_12004_),
    .A2(_09693_),
    .Y(_09695_),
    .B1(_09694_));
 sg13g2_nand2_1 _32748_ (.Y(_09696_),
    .A(\u_inv.f_next[199] ),
    .B(net3843));
 sg13g2_nor2_1 _32749_ (.A(_12006_),
    .B(_09686_),
    .Y(_09697_));
 sg13g2_xnor2_1 _32750_ (.Y(_09698_),
    .A(_12005_),
    .B(_09697_));
 sg13g2_a22oi_1 _32751_ (.Y(_09699_),
    .B1(_09698_),
    .B2(net4675),
    .A2(_09696_),
    .A1(net3727));
 sg13g2_nor3_1 _32752_ (.A(net4442),
    .B(_09695_),
    .C(_09699_),
    .Y(_09700_));
 sg13g2_o21ai_1 _32753_ (.B1(net4020),
    .Y(_09701_),
    .A1(net4613),
    .A2(\u_inv.input_reg[198] ));
 sg13g2_o21ai_1 _32754_ (.B1(_09692_),
    .Y(_01502_),
    .A1(_09700_),
    .A2(_09701_));
 sg13g2_a21oi_1 _32755_ (.A1(_11939_),
    .A2(_12013_),
    .Y(_09702_),
    .B1(_12031_));
 sg13g2_nand2_1 _32756_ (.Y(_09703_),
    .A(_11991_),
    .B(_09702_));
 sg13g2_nor2_1 _32757_ (.A(_11991_),
    .B(_09702_),
    .Y(_09704_));
 sg13g2_nor2_1 _32758_ (.A(net3681),
    .B(_09704_),
    .Y(_09705_));
 sg13g2_a21oi_1 _32759_ (.A1(_12755_),
    .A2(_12758_),
    .Y(_09706_),
    .B1(_12268_));
 sg13g2_xnor2_1 _32760_ (.Y(_09707_),
    .A(_11992_),
    .B(_09706_));
 sg13g2_o21ai_1 _32761_ (.B1(net3716),
    .Y(_09708_),
    .A1(net2509),
    .A2(net4675));
 sg13g2_a21o_1 _32762_ (.A2(_09707_),
    .A1(net4675),
    .B1(_09708_),
    .X(_09709_));
 sg13g2_a221oi_1 _32763_ (.B2(_09705_),
    .C1(net3949),
    .B1(_09703_),
    .A1(net4513),
    .Y(_09710_),
    .A2(net1915));
 sg13g2_a22oi_1 _32764_ (.Y(_01503_),
    .B1(_09709_),
    .B2(_09710_),
    .A2(net3949),
    .A1(_10382_));
 sg13g2_nand2_1 _32765_ (.Y(_09711_),
    .A(net2509),
    .B(net3949));
 sg13g2_a21o_1 _32766_ (.A2(_10690_),
    .A1(\u_inv.f_next[200] ),
    .B1(_09704_),
    .X(_09712_));
 sg13g2_nand2_1 _32767_ (.Y(_09713_),
    .A(_11979_),
    .B(_09712_));
 sg13g2_o21ai_1 _32768_ (.B1(net3774),
    .Y(_09714_),
    .A1(_11979_),
    .A2(_09712_));
 sg13g2_nor2b_1 _32769_ (.A(_09714_),
    .B_N(_09713_),
    .Y(_09715_));
 sg13g2_nand2_1 _32770_ (.Y(_09716_),
    .A(net1992),
    .B(net3843));
 sg13g2_o21ai_1 _32771_ (.B1(_11990_),
    .Y(_09717_),
    .A1(_11992_),
    .A2(_09706_));
 sg13g2_xor2_1 _32772_ (.B(_09717_),
    .A(_11979_),
    .X(_09718_));
 sg13g2_a22oi_1 _32773_ (.Y(_09719_),
    .B1(_09718_),
    .B2(net4675),
    .A2(_09716_),
    .A1(net3727));
 sg13g2_nor3_1 _32774_ (.A(net4442),
    .B(_09715_),
    .C(_09719_),
    .Y(_09720_));
 sg13g2_o21ai_1 _32775_ (.B1(net4020),
    .Y(_09721_),
    .A1(net4613),
    .A2(net1913));
 sg13g2_o21ai_1 _32776_ (.B1(_09711_),
    .Y(_01504_),
    .A1(_09720_),
    .A2(_09721_));
 sg13g2_nand2_1 _32777_ (.Y(_09722_),
    .A(net1992),
    .B(net3949));
 sg13g2_nand2_1 _32778_ (.Y(_09723_),
    .A(_12033_),
    .B(_09713_));
 sg13g2_o21ai_1 _32779_ (.B1(net3774),
    .Y(_09724_),
    .A1(_11978_),
    .A2(_09723_));
 sg13g2_a21oi_1 _32780_ (.A1(_11978_),
    .A2(_09723_),
    .Y(_09725_),
    .B1(_09724_));
 sg13g2_or2_1 _32781_ (.X(_09726_),
    .B(_09706_),
    .A(_12273_));
 sg13g2_and2_1 _32782_ (.A(_12281_),
    .B(_09726_),
    .X(_09727_));
 sg13g2_nor2_1 _32783_ (.A(_11978_),
    .B(_09727_),
    .Y(_09728_));
 sg13g2_xnor2_1 _32784_ (.Y(_09729_),
    .A(_11978_),
    .B(_09727_));
 sg13g2_o21ai_1 _32785_ (.B1(net3839),
    .Y(_09730_),
    .A1(net1959),
    .A2(net4665));
 sg13g2_a21oi_1 _32786_ (.A1(net4665),
    .A2(_09729_),
    .Y(_09731_),
    .B1(_09730_));
 sg13g2_nor3_1 _32787_ (.A(net4442),
    .B(_09725_),
    .C(_09731_),
    .Y(_09732_));
 sg13g2_o21ai_1 _32788_ (.B1(net4020),
    .Y(_09733_),
    .A1(net4617),
    .A2(net1810));
 sg13g2_o21ai_1 _32789_ (.B1(_09722_),
    .Y(_01505_),
    .A1(_09732_),
    .A2(_09733_));
 sg13g2_nand2_1 _32790_ (.Y(_09734_),
    .A(net1959),
    .B(net3940));
 sg13g2_a21oi_1 _32791_ (.A1(_11978_),
    .A2(_09723_),
    .Y(_09735_),
    .B1(_12032_));
 sg13g2_xnor2_1 _32792_ (.Y(_09736_),
    .A(_11981_),
    .B(_09735_));
 sg13g2_a21oi_1 _32793_ (.A1(\u_inv.f_next[202] ),
    .A2(\u_inv.f_reg[202] ),
    .Y(_09737_),
    .B1(_09728_));
 sg13g2_a21oi_1 _32794_ (.A1(_11980_),
    .A2(_09737_),
    .Y(_09738_),
    .B1(net4546));
 sg13g2_o21ai_1 _32795_ (.B1(_09738_),
    .Y(_09739_),
    .A1(_11980_),
    .A2(_09737_));
 sg13g2_o21ai_1 _32796_ (.B1(_09739_),
    .Y(_09740_),
    .A1(\u_inv.f_next[203] ),
    .A2(net4665));
 sg13g2_o21ai_1 _32797_ (.B1(net4381),
    .Y(_09741_),
    .A1(net3763),
    .A2(_09740_));
 sg13g2_a21oi_1 _32798_ (.A1(net3763),
    .A2(_09736_),
    .Y(_09742_),
    .B1(_09741_));
 sg13g2_o21ai_1 _32799_ (.B1(net4020),
    .Y(_09743_),
    .A1(net4617),
    .A2(\u_inv.input_reg[202] ));
 sg13g2_o21ai_1 _32800_ (.B1(_09734_),
    .Y(_01506_),
    .A1(_09742_),
    .A2(_09743_));
 sg13g2_o21ai_1 _32801_ (.B1(_12038_),
    .Y(_09744_),
    .A1(_11993_),
    .A2(_09702_));
 sg13g2_and2_1 _32802_ (.A(_11984_),
    .B(_09744_),
    .X(_09745_));
 sg13g2_xor2_1 _32803_ (.B(_09744_),
    .A(_11984_),
    .X(_09746_));
 sg13g2_nor2_1 _32804_ (.A(_12272_),
    .B(_09727_),
    .Y(_09747_));
 sg13g2_nor2_1 _32805_ (.A(_12284_),
    .B(_09747_),
    .Y(_09748_));
 sg13g2_or2_1 _32806_ (.X(_09749_),
    .B(_09747_),
    .A(_12284_));
 sg13g2_xnor2_1 _32807_ (.Y(_09750_),
    .A(_11984_),
    .B(_09749_));
 sg13g2_o21ai_1 _32808_ (.B1(net3714),
    .Y(_09751_),
    .A1(_10377_),
    .A2(net4665));
 sg13g2_a21oi_1 _32809_ (.A1(net4665),
    .A2(_09750_),
    .Y(_09752_),
    .B1(_09751_));
 sg13g2_o21ai_1 _32810_ (.B1(net4020),
    .Y(_09753_),
    .A1(net4613),
    .A2(net1987));
 sg13g2_nor2_1 _32811_ (.A(_09752_),
    .B(_09753_),
    .Y(_09754_));
 sg13g2_o21ai_1 _32812_ (.B1(_09754_),
    .Y(_09755_),
    .A1(net3681),
    .A2(_09746_));
 sg13g2_o21ai_1 _32813_ (.B1(_09755_),
    .Y(_01507_),
    .A1(_10378_),
    .A2(net4017));
 sg13g2_o21ai_1 _32814_ (.B1(_11982_),
    .Y(_09756_),
    .A1(_12039_),
    .A2(_09745_));
 sg13g2_or3_1 _32815_ (.A(_11982_),
    .B(_12039_),
    .C(_09745_),
    .X(_09757_));
 sg13g2_nand3_1 _32816_ (.B(_09756_),
    .C(_09757_),
    .A(net3763),
    .Y(_09758_));
 sg13g2_nand2_1 _32817_ (.Y(_09759_),
    .A(\u_inv.f_next[205] ),
    .B(net3839));
 sg13g2_o21ai_1 _32818_ (.B1(_11983_),
    .Y(_09760_),
    .A1(_11984_),
    .A2(_09748_));
 sg13g2_xor2_1 _32819_ (.B(_09760_),
    .A(_11982_),
    .X(_09761_));
 sg13g2_a22oi_1 _32820_ (.Y(_09762_),
    .B1(_09761_),
    .B2(net4665),
    .A2(_09759_),
    .A1(net3726));
 sg13g2_nor2_1 _32821_ (.A(net4442),
    .B(_09762_),
    .Y(_09763_));
 sg13g2_o21ai_1 _32822_ (.B1(net4020),
    .Y(_09764_),
    .A1(net4613),
    .A2(net1911));
 sg13g2_a21o_1 _32823_ (.A2(_09763_),
    .A1(_09758_),
    .B1(_09764_),
    .X(_09765_));
 sg13g2_o21ai_1 _32824_ (.B1(_09765_),
    .Y(_01508_),
    .A1(_10377_),
    .A2(net4017));
 sg13g2_and3_1 _32825_ (.X(_09766_),
    .A(_11989_),
    .B(_12040_),
    .C(_09756_));
 sg13g2_a21oi_1 _32826_ (.A1(_12040_),
    .A2(_09756_),
    .Y(_09767_),
    .B1(_11989_));
 sg13g2_nor2_1 _32827_ (.A(_09766_),
    .B(_09767_),
    .Y(_09768_));
 sg13g2_o21ai_1 _32828_ (.B1(net4017),
    .Y(_09769_),
    .A1(net4611),
    .A2(net1943));
 sg13g2_a21oi_1 _32829_ (.A1(_12269_),
    .A2(_09749_),
    .Y(_09770_),
    .B1(_12276_));
 sg13g2_xnor2_1 _32830_ (.Y(_09771_),
    .A(_11989_),
    .B(_09770_));
 sg13g2_o21ai_1 _32831_ (.B1(net3715),
    .Y(_09772_),
    .A1(_10375_),
    .A2(net4666));
 sg13g2_a21oi_1 _32832_ (.A1(net4665),
    .A2(_09771_),
    .Y(_09773_),
    .B1(_09772_));
 sg13g2_nor2_1 _32833_ (.A(_09769_),
    .B(_09773_),
    .Y(_09774_));
 sg13g2_o21ai_1 _32834_ (.B1(_09774_),
    .Y(_09775_),
    .A1(net3681),
    .A2(_09768_));
 sg13g2_o21ai_1 _32835_ (.B1(_09775_),
    .Y(_01509_),
    .A1(_10376_),
    .A2(net4017));
 sg13g2_nand2_1 _32836_ (.Y(_09776_),
    .A(net2664),
    .B(net3940));
 sg13g2_a21oi_1 _32837_ (.A1(\u_inv.f_next[206] ),
    .A2(_10684_),
    .Y(_09777_),
    .B1(_09767_));
 sg13g2_o21ai_1 _32838_ (.B1(net3763),
    .Y(_09778_),
    .A1(_11986_),
    .A2(_09777_));
 sg13g2_a21oi_1 _32839_ (.A1(_11986_),
    .A2(_09777_),
    .Y(_09779_),
    .B1(_09778_));
 sg13g2_nand2_1 _32840_ (.Y(_09780_),
    .A(net2177),
    .B(net3839));
 sg13g2_o21ai_1 _32841_ (.B1(_11987_),
    .Y(_09781_),
    .A1(_11988_),
    .A2(_09770_));
 sg13g2_xnor2_1 _32842_ (.Y(_09782_),
    .A(_11986_),
    .B(_09781_));
 sg13g2_a22oi_1 _32843_ (.Y(_09783_),
    .B1(_09782_),
    .B2(net4666),
    .A2(_09780_),
    .A1(net3726));
 sg13g2_nor3_1 _32844_ (.A(net4440),
    .B(_09779_),
    .C(_09783_),
    .Y(_09784_));
 sg13g2_o21ai_1 _32845_ (.B1(net4020),
    .Y(_09785_),
    .A1(net4613),
    .A2(net1781));
 sg13g2_o21ai_1 _32846_ (.B1(_09776_),
    .Y(_01510_),
    .A1(_09784_),
    .A2(_09785_));
 sg13g2_nand2_1 _32847_ (.Y(_09786_),
    .A(net2177),
    .B(net3940));
 sg13g2_a21oi_2 _32848_ (.B1(_12046_),
    .Y(_09787_),
    .A2(_12014_),
    .A1(_11939_));
 sg13g2_o21ai_1 _32849_ (.B1(net3763),
    .Y(_09788_),
    .A1(_11963_),
    .A2(_09787_));
 sg13g2_a21oi_1 _32850_ (.A1(_11963_),
    .A2(_09787_),
    .Y(_09789_),
    .B1(_09788_));
 sg13g2_a21o_2 _32851_ (.A2(_12759_),
    .A1(_12755_),
    .B1(_12288_),
    .X(_09790_));
 sg13g2_xnor2_1 _32852_ (.Y(_09791_),
    .A(_11963_),
    .B(_09790_));
 sg13g2_o21ai_1 _32853_ (.B1(net3839),
    .Y(_09792_),
    .A1(\u_inv.f_next[208] ),
    .A2(net4664));
 sg13g2_a21oi_1 _32854_ (.A1(net4665),
    .A2(_09791_),
    .Y(_09793_),
    .B1(_09792_));
 sg13g2_nor3_1 _32855_ (.A(net4441),
    .B(_09789_),
    .C(_09793_),
    .Y(_09794_));
 sg13g2_o21ai_1 _32856_ (.B1(net4017),
    .Y(_09795_),
    .A1(net4611),
    .A2(net1823));
 sg13g2_o21ai_1 _32857_ (.B1(_09786_),
    .Y(_01511_),
    .A1(_09794_),
    .A2(_09795_));
 sg13g2_o21ai_1 _32858_ (.B1(_12056_),
    .Y(_09796_),
    .A1(_11963_),
    .A2(_09787_));
 sg13g2_nand2_1 _32859_ (.Y(_09797_),
    .A(_11965_),
    .B(_09796_));
 sg13g2_o21ai_1 _32860_ (.B1(net3694),
    .Y(_09798_),
    .A1(_11965_),
    .A2(_09796_));
 sg13g2_nand2b_1 _32861_ (.Y(_09799_),
    .B(_09797_),
    .A_N(_09798_));
 sg13g2_a21oi_1 _32862_ (.A1(_11963_),
    .A2(_09790_),
    .Y(_09800_),
    .B1(_11962_));
 sg13g2_xnor2_1 _32863_ (.Y(_09801_),
    .A(_11965_),
    .B(_09800_));
 sg13g2_o21ai_1 _32864_ (.B1(net3715),
    .Y(_09802_),
    .A1(net2549),
    .A2(net4664));
 sg13g2_a21oi_1 _32865_ (.A1(net4664),
    .A2(_09801_),
    .Y(_09803_),
    .B1(_09802_));
 sg13g2_a21oi_1 _32866_ (.A1(net4514),
    .A2(net2053),
    .Y(_09804_),
    .B1(net3939));
 sg13g2_nor2b_1 _32867_ (.A(_09803_),
    .B_N(_09804_),
    .Y(_09805_));
 sg13g2_a22oi_1 _32868_ (.Y(_01512_),
    .B1(_09799_),
    .B2(_09805_),
    .A2(net3939),
    .A1(_10373_));
 sg13g2_nand2_1 _32869_ (.Y(_09806_),
    .A(net2549),
    .B(net3939));
 sg13g2_nand2_1 _32870_ (.Y(_09807_),
    .A(_12055_),
    .B(_09797_));
 sg13g2_and2_1 _32871_ (.A(_11960_),
    .B(_09807_),
    .X(_09808_));
 sg13g2_o21ai_1 _32872_ (.B1(net3763),
    .Y(_09809_),
    .A1(_11960_),
    .A2(_09807_));
 sg13g2_nor2_1 _32873_ (.A(_09808_),
    .B(_09809_),
    .Y(_09810_));
 sg13g2_nand2b_1 _32874_ (.Y(_09811_),
    .B(_09790_),
    .A_N(_12250_));
 sg13g2_and2_1 _32875_ (.A(_12300_),
    .B(_09811_),
    .X(_09812_));
 sg13g2_xnor2_1 _32876_ (.Y(_09813_),
    .A(_11960_),
    .B(_09812_));
 sg13g2_o21ai_1 _32877_ (.B1(net3839),
    .Y(_09814_),
    .A1(net2206),
    .A2(net4664));
 sg13g2_a21oi_1 _32878_ (.A1(net4664),
    .A2(_09813_),
    .Y(_09815_),
    .B1(_09814_));
 sg13g2_nor3_1 _32879_ (.A(net4441),
    .B(_09810_),
    .C(_09815_),
    .Y(_09816_));
 sg13g2_o21ai_1 _32880_ (.B1(net4014),
    .Y(_09817_),
    .A1(net4609),
    .A2(net1797));
 sg13g2_o21ai_1 _32881_ (.B1(_09806_),
    .Y(_01513_),
    .A1(_09816_),
    .A2(_09817_));
 sg13g2_nand2_1 _32882_ (.Y(_09818_),
    .A(net2206),
    .B(net3939));
 sg13g2_nor2_1 _32883_ (.A(_12054_),
    .B(_09808_),
    .Y(_09819_));
 sg13g2_xnor2_1 _32884_ (.Y(_09820_),
    .A(_11958_),
    .B(_09819_));
 sg13g2_o21ai_1 _32885_ (.B1(_11959_),
    .Y(_09821_),
    .A1(_11960_),
    .A2(_09812_));
 sg13g2_a21oi_1 _32886_ (.A1(_10370_),
    .A2(net4547),
    .Y(_09822_),
    .B1(net3763));
 sg13g2_o21ai_1 _32887_ (.B1(net4664),
    .Y(_09823_),
    .A1(_11958_),
    .A2(_09821_));
 sg13g2_a21o_1 _32888_ (.A2(_09821_),
    .A1(_11958_),
    .B1(_09823_),
    .X(_09824_));
 sg13g2_a221oi_1 _32889_ (.B2(_09824_),
    .C1(net4441),
    .B1(_09822_),
    .A1(net3763),
    .Y(_09825_),
    .A2(_09820_));
 sg13g2_o21ai_1 _32890_ (.B1(net4014),
    .Y(_09826_),
    .A1(net4612),
    .A2(net1866));
 sg13g2_o21ai_1 _32891_ (.B1(_09818_),
    .Y(_01514_),
    .A1(_09825_),
    .A2(_09826_));
 sg13g2_o21ai_1 _32892_ (.B1(_12058_),
    .Y(_09827_),
    .A1(_11966_),
    .A2(_09787_));
 sg13g2_xnor2_1 _32893_ (.Y(_09828_),
    .A(_11974_),
    .B(_09827_));
 sg13g2_a21oi_1 _32894_ (.A1(_12300_),
    .A2(_09811_),
    .Y(_09829_),
    .B1(_12251_));
 sg13g2_nor2_2 _32895_ (.A(_12303_),
    .B(_09829_),
    .Y(_09830_));
 sg13g2_inv_1 _32896_ (.Y(_09831_),
    .A(_09830_));
 sg13g2_o21ai_1 _32897_ (.B1(net4664),
    .Y(_09832_),
    .A1(_11974_),
    .A2(_09830_));
 sg13g2_a21o_1 _32898_ (.A2(_09830_),
    .A1(_11974_),
    .B1(_09832_),
    .X(_09833_));
 sg13g2_a21oi_1 _32899_ (.A1(net2983),
    .A2(net4547),
    .Y(_09834_),
    .B1(net3703));
 sg13g2_a221oi_1 _32900_ (.B2(_09834_),
    .C1(net3940),
    .B1(_09833_),
    .A1(net3694),
    .Y(_09835_),
    .A2(_09828_));
 sg13g2_o21ai_1 _32901_ (.B1(_09835_),
    .Y(_09836_),
    .A1(net4612),
    .A2(net1966));
 sg13g2_o21ai_1 _32902_ (.B1(_09836_),
    .Y(_01515_),
    .A1(_10370_),
    .A2(net4016));
 sg13g2_o21ai_1 _32903_ (.B1(_11973_),
    .Y(_09837_),
    .A1(_11974_),
    .A2(_09830_));
 sg13g2_xnor2_1 _32904_ (.Y(_09838_),
    .A(_11972_),
    .B(_09837_));
 sg13g2_o21ai_1 _32905_ (.B1(net3714),
    .Y(_09839_),
    .A1(net2477),
    .A2(net4664));
 sg13g2_a21oi_1 _32906_ (.A1(net4666),
    .A2(_09838_),
    .Y(_09840_),
    .B1(_09839_));
 sg13g2_a21oi_1 _32907_ (.A1(_11974_),
    .A2(_09827_),
    .Y(_09841_),
    .B1(_12051_));
 sg13g2_nor2_1 _32908_ (.A(_11972_),
    .B(_09841_),
    .Y(_09842_));
 sg13g2_a21oi_1 _32909_ (.A1(_11972_),
    .A2(_09841_),
    .Y(_09843_),
    .B1(net3681));
 sg13g2_nor2b_1 _32910_ (.A(_09842_),
    .B_N(_09843_),
    .Y(_09844_));
 sg13g2_nor2b_1 _32911_ (.A(net4611),
    .B_N(net2128),
    .Y(_09845_));
 sg13g2_nor4_1 _32912_ (.A(net3939),
    .B(_09840_),
    .C(_09844_),
    .D(_09845_),
    .Y(_09846_));
 sg13g2_a21oi_1 _32913_ (.A1(_10369_),
    .A2(net3939),
    .Y(_01516_),
    .B1(_09846_));
 sg13g2_or2_1 _32914_ (.X(_09847_),
    .B(_09842_),
    .A(_12050_));
 sg13g2_a21oi_1 _32915_ (.A1(_11969_),
    .A2(_09847_),
    .Y(_09848_),
    .B1(net3681));
 sg13g2_o21ai_1 _32916_ (.B1(_09848_),
    .Y(_09849_),
    .A1(_11969_),
    .A2(_09847_));
 sg13g2_a21oi_1 _32917_ (.A1(_12248_),
    .A2(_09831_),
    .Y(_09850_),
    .B1(_12307_));
 sg13g2_xnor2_1 _32918_ (.Y(_09851_),
    .A(_11969_),
    .B(_09850_));
 sg13g2_nor2_1 _32919_ (.A(net1696),
    .B(net4661),
    .Y(_09852_));
 sg13g2_a21oi_1 _32920_ (.A1(net4661),
    .A2(_09851_),
    .Y(_09853_),
    .B1(_09852_));
 sg13g2_a221oi_1 _32921_ (.B2(_09853_),
    .C1(net3939),
    .B1(net3715),
    .A1(net4514),
    .Y(_09854_),
    .A2(net2220));
 sg13g2_a22oi_1 _32922_ (.Y(_01517_),
    .B1(_09849_),
    .B2(_09854_),
    .A2(net3939),
    .A1(_10368_));
 sg13g2_nand2_1 _32923_ (.Y(_09855_),
    .A(net1696),
    .B(net3938));
 sg13g2_o21ai_1 _32924_ (.B1(_11968_),
    .Y(_09856_),
    .A1(_11969_),
    .A2(_09850_));
 sg13g2_xor2_1 _32925_ (.B(_09856_),
    .A(_11967_),
    .X(_09857_));
 sg13g2_nand2_1 _32926_ (.Y(_09858_),
    .A(net4661),
    .B(_09857_));
 sg13g2_a21oi_1 _32927_ (.A1(_10366_),
    .A2(net4546),
    .Y(_09859_),
    .B1(net3762));
 sg13g2_a21oi_1 _32928_ (.A1(_11969_),
    .A2(_09847_),
    .Y(_09860_),
    .B1(_12047_));
 sg13g2_xnor2_1 _32929_ (.Y(_09861_),
    .A(_11967_),
    .B(_09860_));
 sg13g2_a221oi_1 _32930_ (.B2(net3762),
    .C1(net4440),
    .B1(_09861_),
    .A1(_09858_),
    .Y(_09862_),
    .A2(_09859_));
 sg13g2_o21ai_1 _32931_ (.B1(net4017),
    .Y(_09863_),
    .A1(net4609),
    .A2(\u_inv.input_reg[214] ));
 sg13g2_o21ai_1 _32932_ (.B1(_09855_),
    .Y(_01518_),
    .A1(_09862_),
    .A2(_09863_));
 sg13g2_nand2_1 _32933_ (.Y(_09864_),
    .A(net2124),
    .B(net3938));
 sg13g2_o21ai_1 _32934_ (.B1(_12061_),
    .Y(_09865_),
    .A1(_11976_),
    .A2(_09787_));
 sg13g2_o21ai_1 _32935_ (.B1(net3762),
    .Y(_09866_),
    .A1(_11944_),
    .A2(_09865_));
 sg13g2_a21oi_1 _32936_ (.A1(_11944_),
    .A2(_09865_),
    .Y(_09867_),
    .B1(_09866_));
 sg13g2_a21oi_1 _32937_ (.A1(_12252_),
    .A2(_09790_),
    .Y(_09868_),
    .B1(_12309_));
 sg13g2_nor2_1 _32938_ (.A(_11944_),
    .B(_09868_),
    .Y(_09869_));
 sg13g2_xnor2_1 _32939_ (.Y(_09870_),
    .A(_11944_),
    .B(_09868_));
 sg13g2_o21ai_1 _32940_ (.B1(net3838),
    .Y(_09871_),
    .A1(\u_inv.f_next[216] ),
    .A2(net4661));
 sg13g2_a21oi_1 _32941_ (.A1(net4661),
    .A2(_09870_),
    .Y(_09872_),
    .B1(_09871_));
 sg13g2_nor3_1 _32942_ (.A(net4440),
    .B(_09867_),
    .C(_09872_),
    .Y(_09873_));
 sg13g2_o21ai_1 _32943_ (.B1(net4014),
    .Y(_09874_),
    .A1(net4609),
    .A2(net1796));
 sg13g2_o21ai_1 _32944_ (.B1(_09864_),
    .Y(_01519_),
    .A1(_09873_),
    .A2(_09874_));
 sg13g2_nand2_1 _32945_ (.Y(_09875_),
    .A(net2195),
    .B(net3938));
 sg13g2_a21oi_1 _32946_ (.A1(_11944_),
    .A2(_09865_),
    .Y(_09876_),
    .B1(_12063_));
 sg13g2_nor2_1 _32947_ (.A(_11945_),
    .B(_09876_),
    .Y(_09877_));
 sg13g2_a21oi_1 _32948_ (.A1(_11945_),
    .A2(_09876_),
    .Y(_09878_),
    .B1(net3837));
 sg13g2_nor2b_1 _32949_ (.A(_09877_),
    .B_N(_09878_),
    .Y(_09879_));
 sg13g2_nand2_1 _32950_ (.Y(_09880_),
    .A(\u_inv.f_next[217] ),
    .B(net3837));
 sg13g2_a21oi_1 _32951_ (.A1(\u_inv.f_next[216] ),
    .A2(\u_inv.f_reg[216] ),
    .Y(_09881_),
    .B1(_09869_));
 sg13g2_xor2_1 _32952_ (.B(_09881_),
    .A(_11945_),
    .X(_09882_));
 sg13g2_a22oi_1 _32953_ (.Y(_09883_),
    .B1(_09882_),
    .B2(net4660),
    .A2(_09880_),
    .A1(net3725));
 sg13g2_nor3_1 _32954_ (.A(net4441),
    .B(_09879_),
    .C(_09883_),
    .Y(_09884_));
 sg13g2_o21ai_1 _32955_ (.B1(net4014),
    .Y(_09885_),
    .A1(net4609),
    .A2(net2040));
 sg13g2_o21ai_1 _32956_ (.B1(_09875_),
    .Y(_01520_),
    .A1(_09884_),
    .A2(_09885_));
 sg13g2_nand2_1 _32957_ (.Y(_09886_),
    .A(net2258),
    .B(net3938));
 sg13g2_a21oi_1 _32958_ (.A1(\u_inv.f_next[217] ),
    .A2(_10673_),
    .Y(_09887_),
    .B1(_09877_));
 sg13g2_nor2_1 _32959_ (.A(_11942_),
    .B(_09887_),
    .Y(_09888_));
 sg13g2_a21oi_1 _32960_ (.A1(_11942_),
    .A2(_09887_),
    .Y(_09889_),
    .B1(net3837));
 sg13g2_nor2b_1 _32961_ (.A(_09888_),
    .B_N(_09889_),
    .Y(_09890_));
 sg13g2_a21o_1 _32962_ (.A2(_09869_),
    .A1(_11945_),
    .B1(_12290_),
    .X(_09891_));
 sg13g2_xnor2_1 _32963_ (.Y(_09892_),
    .A(_11942_),
    .B(_09891_));
 sg13g2_o21ai_1 _32964_ (.B1(net3837),
    .Y(_09893_),
    .A1(net2109),
    .A2(net4660));
 sg13g2_a21oi_1 _32965_ (.A1(net4660),
    .A2(_09892_),
    .Y(_09894_),
    .B1(_09893_));
 sg13g2_nor3_1 _32966_ (.A(net4441),
    .B(_09890_),
    .C(_09894_),
    .Y(_09895_));
 sg13g2_o21ai_1 _32967_ (.B1(net4014),
    .Y(_09896_),
    .A1(net4609),
    .A2(net1988));
 sg13g2_o21ai_1 _32968_ (.B1(_09886_),
    .Y(_01521_),
    .A1(_09895_),
    .A2(_09896_));
 sg13g2_nand2_1 _32969_ (.Y(_09897_),
    .A(net2109),
    .B(net3938));
 sg13g2_a21oi_1 _32970_ (.A1(_11942_),
    .A2(_09891_),
    .Y(_09898_),
    .B1(_11941_));
 sg13g2_xnor2_1 _32971_ (.Y(_09899_),
    .A(_11940_),
    .B(_09898_));
 sg13g2_nor2_1 _32972_ (.A(\u_inv.f_next[219] ),
    .B(net4660),
    .Y(_09900_));
 sg13g2_a21oi_1 _32973_ (.A1(net4660),
    .A2(_09899_),
    .Y(_09901_),
    .B1(_09900_));
 sg13g2_o21ai_1 _32974_ (.B1(_11940_),
    .Y(_09902_),
    .A1(_12062_),
    .A2(_09888_));
 sg13g2_nor3_1 _32975_ (.A(_11940_),
    .B(_12062_),
    .C(_09888_),
    .Y(_09903_));
 sg13g2_nor2_1 _32976_ (.A(net3837),
    .B(_09903_),
    .Y(_09904_));
 sg13g2_a221oi_1 _32977_ (.B2(_09904_),
    .C1(net4441),
    .B1(_09902_),
    .A1(net3837),
    .Y(_09905_),
    .A2(_09901_));
 sg13g2_o21ai_1 _32978_ (.B1(net4014),
    .Y(_09906_),
    .A1(net4609),
    .A2(net1824));
 sg13g2_o21ai_1 _32979_ (.B1(_09897_),
    .Y(_01522_),
    .A1(_09905_),
    .A2(_09906_));
 sg13g2_nand2_1 _32980_ (.Y(_09907_),
    .A(net2236),
    .B(net3938));
 sg13g2_a21oi_1 _32981_ (.A1(_11947_),
    .A2(_09865_),
    .Y(_09908_),
    .B1(_12068_));
 sg13g2_o21ai_1 _32982_ (.B1(net3762),
    .Y(_09909_),
    .A1(_11955_),
    .A2(_09908_));
 sg13g2_a21oi_1 _32983_ (.A1(_11955_),
    .A2(_09908_),
    .Y(_09910_),
    .B1(_09909_));
 sg13g2_nand2b_1 _32984_ (.Y(_09911_),
    .B(_09869_),
    .A_N(_12245_));
 sg13g2_nand2_2 _32985_ (.Y(_09912_),
    .A(_12293_),
    .B(_09911_));
 sg13g2_xnor2_1 _32986_ (.Y(_09913_),
    .A(_11955_),
    .B(_09912_));
 sg13g2_o21ai_1 _32987_ (.B1(net3837),
    .Y(_09914_),
    .A1(net1709),
    .A2(net4660));
 sg13g2_a21oi_1 _32988_ (.A1(net4660),
    .A2(_09913_),
    .Y(_09915_),
    .B1(_09914_));
 sg13g2_nor3_1 _32989_ (.A(net4440),
    .B(_09910_),
    .C(_09915_),
    .Y(_09916_));
 sg13g2_o21ai_1 _32990_ (.B1(net4014),
    .Y(_09917_),
    .A1(net4609),
    .A2(net1792));
 sg13g2_o21ai_1 _32991_ (.B1(_09907_),
    .Y(_01523_),
    .A1(_09916_),
    .A2(_09917_));
 sg13g2_nand2_1 _32992_ (.Y(_09918_),
    .A(net1709),
    .B(net3938));
 sg13g2_o21ai_1 _32993_ (.B1(_12069_),
    .Y(_09919_),
    .A1(_11955_),
    .A2(_09908_));
 sg13g2_and2_1 _32994_ (.A(_11953_),
    .B(_09919_),
    .X(_09920_));
 sg13g2_o21ai_1 _32995_ (.B1(net3762),
    .Y(_09921_),
    .A1(_11953_),
    .A2(_09919_));
 sg13g2_nor2_1 _32996_ (.A(_09920_),
    .B(_09921_),
    .Y(_09922_));
 sg13g2_nand2_1 _32997_ (.Y(_09923_),
    .A(\u_inv.f_next[221] ),
    .B(net3837));
 sg13g2_a21oi_1 _32998_ (.A1(_11955_),
    .A2(_09912_),
    .Y(_09924_),
    .B1(_11954_));
 sg13g2_xnor2_1 _32999_ (.Y(_09925_),
    .A(_11953_),
    .B(_09924_));
 sg13g2_a22oi_1 _33000_ (.Y(_09926_),
    .B1(_09925_),
    .B2(net4660),
    .A2(_09923_),
    .A1(net3725));
 sg13g2_nor3_1 _33001_ (.A(net4440),
    .B(_09922_),
    .C(_09926_),
    .Y(_09927_));
 sg13g2_o21ai_1 _33002_ (.B1(net4016),
    .Y(_09928_),
    .A1(net4609),
    .A2(\u_inv.input_reg[220] ));
 sg13g2_o21ai_1 _33003_ (.B1(_09918_),
    .Y(_01524_),
    .A1(_09927_),
    .A2(_09928_));
 sg13g2_nand2_1 _33004_ (.Y(_09929_),
    .A(net2277),
    .B(net3929));
 sg13g2_nor3_1 _33005_ (.A(_11950_),
    .B(_12070_),
    .C(_09920_),
    .Y(_09930_));
 sg13g2_o21ai_1 _33006_ (.B1(_11950_),
    .Y(_09931_),
    .A1(_12070_),
    .A2(_09920_));
 sg13g2_nor2_1 _33007_ (.A(net3838),
    .B(_09930_),
    .Y(_09932_));
 sg13g2_a21oi_1 _33008_ (.A1(_12242_),
    .A2(_09912_),
    .Y(_09933_),
    .B1(_12295_));
 sg13g2_xnor2_1 _33009_ (.Y(_09934_),
    .A(_11950_),
    .B(_09933_));
 sg13g2_nand2_1 _33010_ (.Y(_09935_),
    .A(_10359_),
    .B(net4538));
 sg13g2_a21oi_1 _33011_ (.A1(net4661),
    .A2(_09934_),
    .Y(_09936_),
    .B1(net3762));
 sg13g2_a221oi_1 _33012_ (.B2(_09936_),
    .C1(net4440),
    .B1(_09935_),
    .A1(_09931_),
    .Y(_09937_),
    .A2(_09932_));
 sg13g2_o21ai_1 _33013_ (.B1(net4012),
    .Y(_09938_),
    .A1(net4605),
    .A2(net2081));
 sg13g2_o21ai_1 _33014_ (.B1(_09929_),
    .Y(_01525_),
    .A1(_09937_),
    .A2(_09938_));
 sg13g2_nand2_1 _33015_ (.Y(_09939_),
    .A(net1463),
    .B(net3929));
 sg13g2_nand2b_1 _33016_ (.Y(_09940_),
    .B(_09931_),
    .A_N(_12073_));
 sg13g2_xor2_1 _33017_ (.B(_09940_),
    .A(_11948_),
    .X(_09941_));
 sg13g2_a21oi_1 _33018_ (.A1(_10358_),
    .A2(net4538),
    .Y(_09942_),
    .B1(net3754));
 sg13g2_o21ai_1 _33019_ (.B1(_11949_),
    .Y(_09943_),
    .A1(_11950_),
    .A2(_09933_));
 sg13g2_o21ai_1 _33020_ (.B1(net4661),
    .Y(_09944_),
    .A1(_11948_),
    .A2(_09943_));
 sg13g2_a21o_1 _33021_ (.A2(_09943_),
    .A1(_11948_),
    .B1(_09944_),
    .X(_09945_));
 sg13g2_a221oi_1 _33022_ (.B2(_09945_),
    .C1(net4438),
    .B1(_09942_),
    .A1(net3754),
    .Y(_09946_),
    .A2(_09941_));
 sg13g2_o21ai_1 _33023_ (.B1(net4012),
    .Y(_09947_),
    .A1(net4607),
    .A2(\u_inv.input_reg[222] ));
 sg13g2_o21ai_1 _33024_ (.B1(_09939_),
    .Y(_01526_),
    .A1(_09946_),
    .A2(_09947_));
 sg13g2_nand2_1 _33025_ (.Y(_09948_),
    .A(_12079_),
    .B(_12086_));
 sg13g2_a21oi_1 _33026_ (.A1(_12079_),
    .A2(_12086_),
    .Y(_09949_),
    .B1(net3679));
 sg13g2_o21ai_1 _33027_ (.B1(_09949_),
    .Y(_09950_),
    .A1(_12079_),
    .A2(_12086_));
 sg13g2_nor2_1 _33028_ (.A(_12086_),
    .B(_12761_),
    .Y(_09951_));
 sg13g2_nand2_1 _33029_ (.Y(_09952_),
    .A(_12086_),
    .B(_12761_));
 sg13g2_nand3b_1 _33030_ (.B(_09952_),
    .C(net4654),
    .Y(_09953_),
    .A_N(_09951_));
 sg13g2_o21ai_1 _33031_ (.B1(_09953_),
    .Y(_09954_),
    .A1(_10357_),
    .A2(net4654));
 sg13g2_a221oi_1 _33032_ (.B2(_09954_),
    .C1(net3929),
    .B1(net3713),
    .A1(net4515),
    .Y(_09955_),
    .A2(net2113));
 sg13g2_a22oi_1 _33033_ (.Y(_01527_),
    .B1(_09950_),
    .B2(_09955_),
    .A2(net3929),
    .A1(_10358_));
 sg13g2_nand2_1 _33034_ (.Y(_09956_),
    .A(net2049),
    .B(net3929));
 sg13g2_a21oi_1 _33035_ (.A1(\u_inv.f_next[224] ),
    .A2(\u_inv.f_reg[224] ),
    .Y(_09957_),
    .B1(_09951_));
 sg13g2_xnor2_1 _33036_ (.Y(_09958_),
    .A(_12087_),
    .B(_09957_));
 sg13g2_mux2_1 _33037_ (.A0(net4967),
    .A1(_09958_),
    .S(net4654),
    .X(_09959_));
 sg13g2_and2_1 _33038_ (.A(_12126_),
    .B(_09948_),
    .X(_09960_));
 sg13g2_nor2_1 _33039_ (.A(_12087_),
    .B(_09960_),
    .Y(_09961_));
 sg13g2_nand2_1 _33040_ (.Y(_09962_),
    .A(_12087_),
    .B(_09960_));
 sg13g2_nor2_1 _33041_ (.A(net3833),
    .B(_09961_),
    .Y(_09963_));
 sg13g2_a221oi_1 _33042_ (.B2(_09963_),
    .C1(net4439),
    .B1(_09962_),
    .A1(net3833),
    .Y(_09964_),
    .A2(_09959_));
 sg13g2_o21ai_1 _33043_ (.B1(net4012),
    .Y(_09965_),
    .A1(net4605),
    .A2(net1835));
 sg13g2_o21ai_1 _33044_ (.B1(_09956_),
    .Y(_01528_),
    .A1(_09964_),
    .A2(_09965_));
 sg13g2_nand2_1 _33045_ (.Y(_09966_),
    .A(net2266),
    .B(net3929));
 sg13g2_a21oi_1 _33046_ (.A1(\u_inv.f_next[225] ),
    .A2(_10665_),
    .Y(_09967_),
    .B1(_09961_));
 sg13g2_nor2_1 _33047_ (.A(_12081_),
    .B(_09967_),
    .Y(_09968_));
 sg13g2_a21oi_1 _33048_ (.A1(_12081_),
    .A2(_09967_),
    .Y(_09969_),
    .B1(net3831));
 sg13g2_nor2b_1 _33049_ (.A(_09968_),
    .B_N(_09969_),
    .Y(_09970_));
 sg13g2_a21oi_1 _33050_ (.A1(_12087_),
    .A2(_09951_),
    .Y(_09971_),
    .B1(_12777_));
 sg13g2_xnor2_1 _33051_ (.Y(_09972_),
    .A(_12082_),
    .B(_09971_));
 sg13g2_o21ai_1 _33052_ (.B1(net3831),
    .Y(_09973_),
    .A1(\u_inv.f_next[226] ),
    .A2(net4649));
 sg13g2_a21oi_1 _33053_ (.A1(net4649),
    .A2(_09972_),
    .Y(_09974_),
    .B1(_09973_));
 sg13g2_nor3_1 _33054_ (.A(net4438),
    .B(_09970_),
    .C(_09974_),
    .Y(_09975_));
 sg13g2_o21ai_1 _33055_ (.B1(net4012),
    .Y(_09976_),
    .A1(net4607),
    .A2(net1884));
 sg13g2_o21ai_1 _33056_ (.B1(_09966_),
    .Y(_01529_),
    .A1(_09975_),
    .A2(_09976_));
 sg13g2_nor2_1 _33057_ (.A(net2700),
    .B(net4006),
    .Y(_09977_));
 sg13g2_nor3_1 _33058_ (.A(_12084_),
    .B(_12124_),
    .C(_09968_),
    .Y(_09978_));
 sg13g2_o21ai_1 _33059_ (.B1(_12084_),
    .Y(_09979_),
    .A1(_12124_),
    .A2(_09968_));
 sg13g2_nor2_1 _33060_ (.A(net3680),
    .B(_09978_),
    .Y(_09980_));
 sg13g2_o21ai_1 _33061_ (.B1(_12080_),
    .Y(_09981_),
    .A1(_12082_),
    .A2(_09971_));
 sg13g2_xnor2_1 _33062_ (.Y(_09982_),
    .A(_12083_),
    .B(_09981_));
 sg13g2_o21ai_1 _33063_ (.B1(net3712),
    .Y(_09983_),
    .A1(\u_inv.f_next[227] ),
    .A2(net4649));
 sg13g2_a21oi_1 _33064_ (.A1(net4649),
    .A2(_09982_),
    .Y(_09984_),
    .B1(_09983_));
 sg13g2_a221oi_1 _33065_ (.B2(_09980_),
    .C1(_09984_),
    .B1(_09979_),
    .A1(net4515),
    .Y(_09985_),
    .A2(net2093));
 sg13g2_a21oi_1 _33066_ (.A1(net4006),
    .A2(_09985_),
    .Y(_01530_),
    .B1(_09977_));
 sg13g2_o21ai_1 _33067_ (.B1(_12779_),
    .Y(_09986_),
    .A1(_12761_),
    .A2(_12774_));
 sg13g2_nand2_1 _33068_ (.Y(_09987_),
    .A(_12095_),
    .B(_09986_));
 sg13g2_xnor2_1 _33069_ (.Y(_09988_),
    .A(_12095_),
    .B(_09986_));
 sg13g2_o21ai_1 _33070_ (.B1(net3712),
    .Y(_09989_),
    .A1(net3277),
    .A2(net4649));
 sg13g2_a21o_1 _33071_ (.A2(_09988_),
    .A1(net4649),
    .B1(_09989_),
    .X(_09990_));
 sg13g2_a21oi_1 _33072_ (.A1(_12079_),
    .A2(_12088_),
    .Y(_09991_),
    .B1(_12129_));
 sg13g2_xnor2_1 _33073_ (.Y(_09992_),
    .A(_12096_),
    .B(_09991_));
 sg13g2_a221oi_1 _33074_ (.B2(_09992_),
    .C1(net3926),
    .B1(net3691),
    .A1(net4512),
    .Y(_09993_),
    .A2(net2494));
 sg13g2_a22oi_1 _33075_ (.Y(_01531_),
    .B1(_09990_),
    .B2(_09993_),
    .A2(net3926),
    .A1(_10354_));
 sg13g2_nand2_1 _33076_ (.Y(_09994_),
    .A(net2212),
    .B(net3831));
 sg13g2_o21ai_1 _33077_ (.B1(_09987_),
    .Y(_09995_),
    .A1(_10353_),
    .A2(_10662_));
 sg13g2_xnor2_1 _33078_ (.Y(_09996_),
    .A(_12093_),
    .B(_09995_));
 sg13g2_a22oi_1 _33079_ (.Y(_09997_),
    .B1(_09996_),
    .B2(net4649),
    .A2(_09994_),
    .A1(net3724));
 sg13g2_o21ai_1 _33080_ (.B1(_12122_),
    .Y(_09998_),
    .A1(_12095_),
    .A2(_09991_));
 sg13g2_and2_1 _33081_ (.A(_12094_),
    .B(_09998_),
    .X(_09999_));
 sg13g2_o21ai_1 _33082_ (.B1(net3752),
    .Y(_10000_),
    .A1(_12094_),
    .A2(_09998_));
 sg13g2_o21ai_1 _33083_ (.B1(net4378),
    .Y(_10001_),
    .A1(_09999_),
    .A2(_10000_));
 sg13g2_a21oi_1 _33084_ (.A1(net4515),
    .A2(_10983_),
    .Y(_10002_),
    .B1(net3926));
 sg13g2_o21ai_1 _33085_ (.B1(_10002_),
    .Y(_10003_),
    .A1(_09997_),
    .A2(_10001_));
 sg13g2_o21ai_1 _33086_ (.B1(_10003_),
    .Y(_01532_),
    .A1(_10353_),
    .A2(net4007));
 sg13g2_nand2_1 _33087_ (.Y(_10004_),
    .A(net2212),
    .B(net3928));
 sg13g2_nor3_1 _33088_ (.A(_12092_),
    .B(_12121_),
    .C(_09999_),
    .Y(_10005_));
 sg13g2_o21ai_1 _33089_ (.B1(_12092_),
    .Y(_10006_),
    .A1(_12121_),
    .A2(_09999_));
 sg13g2_nor2_1 _33090_ (.A(net3832),
    .B(_10005_),
    .Y(_10007_));
 sg13g2_a21oi_1 _33091_ (.A1(_12763_),
    .A2(_09986_),
    .Y(_10008_),
    .B1(_12787_));
 sg13g2_xnor2_1 _33092_ (.Y(_10009_),
    .A(_12092_),
    .B(_10008_));
 sg13g2_nand2_1 _33093_ (.Y(_10010_),
    .A(_10351_),
    .B(net4536));
 sg13g2_a21oi_1 _33094_ (.A1(net4649),
    .A2(_10009_),
    .Y(_10011_),
    .B1(net3753));
 sg13g2_a221oi_1 _33095_ (.B2(_10011_),
    .C1(net4438),
    .B1(_10010_),
    .A1(_10006_),
    .Y(_10012_),
    .A2(_10007_));
 sg13g2_o21ai_1 _33096_ (.B1(net4007),
    .Y(_10013_),
    .A1(net4604),
    .A2(\u_inv.input_reg[229] ));
 sg13g2_o21ai_1 _33097_ (.B1(_10004_),
    .Y(_01533_),
    .A1(_10012_),
    .A2(_10013_));
 sg13g2_nand2_1 _33098_ (.Y(_10014_),
    .A(_12134_),
    .B(_10006_));
 sg13g2_xnor2_1 _33099_ (.Y(_10015_),
    .A(_12089_),
    .B(_10014_));
 sg13g2_nand2_1 _33100_ (.Y(_10016_),
    .A(\u_inv.f_next[231] ),
    .B(net3831));
 sg13g2_o21ai_1 _33101_ (.B1(_12090_),
    .Y(_10017_),
    .A1(_12092_),
    .A2(_10008_));
 sg13g2_xnor2_1 _33102_ (.Y(_10018_),
    .A(_12089_),
    .B(_10017_));
 sg13g2_a22oi_1 _33103_ (.Y(_10019_),
    .B1(_10018_),
    .B2(net4648),
    .A2(_10016_),
    .A1(net3724));
 sg13g2_a21oi_1 _33104_ (.A1(net3752),
    .A2(_10015_),
    .Y(_10020_),
    .B1(_10019_));
 sg13g2_o21ai_1 _33105_ (.B1(net4007),
    .Y(_10021_),
    .A1(net4604),
    .A2(net2448));
 sg13g2_a21o_1 _33106_ (.A2(_10020_),
    .A1(net4378),
    .B1(_10021_),
    .X(_10022_));
 sg13g2_o21ai_1 _33107_ (.B1(_10022_),
    .Y(_01534_),
    .A1(_10351_),
    .A2(net4006));
 sg13g2_nand2b_1 _33108_ (.Y(_10023_),
    .B(_09986_),
    .A_N(_12764_));
 sg13g2_and2_1 _33109_ (.A(_12789_),
    .B(_10023_),
    .X(_10024_));
 sg13g2_nand2_1 _33110_ (.Y(_10025_),
    .A(_12789_),
    .B(_10023_));
 sg13g2_xnor2_1 _33111_ (.Y(_10026_),
    .A(_12103_),
    .B(_10024_));
 sg13g2_a21oi_1 _33112_ (.A1(net2947),
    .A2(net4537),
    .Y(_10027_),
    .B1(net3702));
 sg13g2_o21ai_1 _33113_ (.B1(_10027_),
    .Y(_10028_),
    .A1(net4537),
    .A2(_10026_));
 sg13g2_and3_1 _33114_ (.X(_10029_),
    .A(_12079_),
    .B(_12088_),
    .C(_12097_));
 sg13g2_or2_1 _33115_ (.X(_10030_),
    .B(_10029_),
    .A(_12136_));
 sg13g2_nand2_1 _33116_ (.Y(_10031_),
    .A(_12103_),
    .B(_10030_));
 sg13g2_xnor2_1 _33117_ (.Y(_10032_),
    .A(_12103_),
    .B(_10030_));
 sg13g2_o21ai_1 _33118_ (.B1(net4007),
    .Y(_10033_),
    .A1(net4604),
    .A2(net2327));
 sg13g2_a21oi_1 _33119_ (.A1(net3692),
    .A2(_10032_),
    .Y(_10034_),
    .B1(_10033_));
 sg13g2_nand2_1 _33120_ (.Y(_10035_),
    .A(_10028_),
    .B(_10034_));
 sg13g2_o21ai_1 _33121_ (.B1(_10035_),
    .Y(_01535_),
    .A1(_10350_),
    .A2(net4006));
 sg13g2_a21oi_1 _33122_ (.A1(_10348_),
    .A2(net4537),
    .Y(_10036_),
    .B1(net3752));
 sg13g2_o21ai_1 _33123_ (.B1(_12102_),
    .Y(_10037_),
    .A1(_12103_),
    .A2(_10024_));
 sg13g2_xnor2_1 _33124_ (.Y(_10038_),
    .A(_12105_),
    .B(_10037_));
 sg13g2_o21ai_1 _33125_ (.B1(_10036_),
    .Y(_10039_),
    .A1(net4537),
    .A2(_10038_));
 sg13g2_a21oi_1 _33126_ (.A1(_12147_),
    .A2(_10031_),
    .Y(_10040_),
    .B1(_12104_));
 sg13g2_nand3_1 _33127_ (.B(_12147_),
    .C(_10031_),
    .A(_12104_),
    .Y(_10041_));
 sg13g2_nor2_1 _33128_ (.A(net3832),
    .B(_10040_),
    .Y(_10042_));
 sg13g2_a21oi_1 _33129_ (.A1(_10041_),
    .A2(_10042_),
    .Y(_10043_),
    .B1(net4438));
 sg13g2_a21oi_1 _33130_ (.A1(_10039_),
    .A2(_10043_),
    .Y(_10044_),
    .B1(net3926));
 sg13g2_o21ai_1 _33131_ (.B1(_10044_),
    .Y(_10045_),
    .A1(net4607),
    .A2(net2185));
 sg13g2_o21ai_1 _33132_ (.B1(_10045_),
    .Y(_01536_),
    .A1(_10349_),
    .A2(net4007));
 sg13g2_nand2_1 _33133_ (.Y(_10046_),
    .A(net2193),
    .B(net3928));
 sg13g2_nor3_1 _33134_ (.A(_12100_),
    .B(_12146_),
    .C(_10040_),
    .Y(_10047_));
 sg13g2_o21ai_1 _33135_ (.B1(_12100_),
    .Y(_10048_),
    .A1(_12146_),
    .A2(_10040_));
 sg13g2_nor2_1 _33136_ (.A(net3831),
    .B(_10047_),
    .Y(_10049_));
 sg13g2_a21oi_1 _33137_ (.A1(_12769_),
    .A2(_10025_),
    .Y(_10050_),
    .B1(_12782_));
 sg13g2_xnor2_1 _33138_ (.Y(_10051_),
    .A(_12100_),
    .B(_10050_));
 sg13g2_nand2_1 _33139_ (.Y(_10052_),
    .A(_10347_),
    .B(net4537));
 sg13g2_a21oi_1 _33140_ (.A1(net4648),
    .A2(_10051_),
    .Y(_10053_),
    .B1(net3752));
 sg13g2_a221oi_1 _33141_ (.B2(_10053_),
    .C1(net4439),
    .B1(_10052_),
    .A1(_10048_),
    .Y(_10054_),
    .A2(_10049_));
 sg13g2_o21ai_1 _33142_ (.B1(net4013),
    .Y(_10055_),
    .A1(net4607),
    .A2(net1897));
 sg13g2_o21ai_1 _33143_ (.B1(_10046_),
    .Y(_01537_),
    .A1(_10054_),
    .A2(_10055_));
 sg13g2_nand2_1 _33144_ (.Y(_10056_),
    .A(net1412),
    .B(net3926));
 sg13g2_nor2b_1 _33145_ (.A(_12145_),
    .B_N(_10048_),
    .Y(_10057_));
 sg13g2_xnor2_1 _33146_ (.Y(_10058_),
    .A(_12098_),
    .B(_10057_));
 sg13g2_a21oi_1 _33147_ (.A1(_10346_),
    .A2(net4537),
    .Y(_10059_),
    .B1(net3752));
 sg13g2_o21ai_1 _33148_ (.B1(_12099_),
    .Y(_10060_),
    .A1(_12100_),
    .A2(_10050_));
 sg13g2_o21ai_1 _33149_ (.B1(net4648),
    .Y(_10061_),
    .A1(_12098_),
    .A2(_10060_));
 sg13g2_a21o_1 _33150_ (.A2(_10060_),
    .A1(_12098_),
    .B1(_10061_),
    .X(_10062_));
 sg13g2_a221oi_1 _33151_ (.B2(_10062_),
    .C1(net4439),
    .B1(_10059_),
    .A1(net3752),
    .Y(_10063_),
    .A2(_10058_));
 sg13g2_o21ai_1 _33152_ (.B1(net4006),
    .Y(_10064_),
    .A1(net4607),
    .A2(\u_inv.input_reg[234] ));
 sg13g2_o21ai_1 _33153_ (.B1(_10056_),
    .Y(_01538_),
    .A1(_10063_),
    .A2(_10064_));
 sg13g2_o21ai_1 _33154_ (.B1(_12784_),
    .Y(_10065_),
    .A1(_12771_),
    .A2(_10024_));
 sg13g2_xnor2_1 _33155_ (.Y(_10066_),
    .A(_12110_),
    .B(_10065_));
 sg13g2_o21ai_1 _33156_ (.B1(net3711),
    .Y(_10067_),
    .A1(_10345_),
    .A2(net4648));
 sg13g2_a21oi_1 _33157_ (.A1(net4648),
    .A2(_10066_),
    .Y(_10068_),
    .B1(_10067_));
 sg13g2_o21ai_1 _33158_ (.B1(_12107_),
    .Y(_10069_),
    .A1(_12136_),
    .A2(_10029_));
 sg13g2_nand2_1 _33159_ (.Y(_10070_),
    .A(_12150_),
    .B(_10069_));
 sg13g2_xnor2_1 _33160_ (.Y(_10071_),
    .A(_12111_),
    .B(_10070_));
 sg13g2_nor2_1 _33161_ (.A(net3679),
    .B(_10071_),
    .Y(_10072_));
 sg13g2_o21ai_1 _33162_ (.B1(net4006),
    .Y(_10073_),
    .A1(net4607),
    .A2(net2096));
 sg13g2_or3_1 _33163_ (.A(_10068_),
    .B(_10072_),
    .C(_10073_),
    .X(_10074_));
 sg13g2_o21ai_1 _33164_ (.B1(_10074_),
    .Y(_01539_),
    .A1(_10346_),
    .A2(net4006));
 sg13g2_nand2_1 _33165_ (.Y(_10075_),
    .A(net1625),
    .B(net3926));
 sg13g2_a21oi_1 _33166_ (.A1(_12111_),
    .A2(_10065_),
    .Y(_10076_),
    .B1(_12109_));
 sg13g2_xnor2_1 _33167_ (.Y(_10077_),
    .A(_12112_),
    .B(_10076_));
 sg13g2_a21oi_1 _33168_ (.A1(\u_inv.f_next[237] ),
    .A2(net4537),
    .Y(_10078_),
    .B1(net4438));
 sg13g2_o21ai_1 _33169_ (.B1(_10078_),
    .Y(_10079_),
    .A1(net4537),
    .A2(_10077_));
 sg13g2_a21o_1 _33170_ (.A2(_10070_),
    .A1(_12110_),
    .B1(_12137_),
    .X(_10080_));
 sg13g2_a21oi_1 _33171_ (.A1(_12150_),
    .A2(_10069_),
    .Y(_10081_),
    .B1(_12113_));
 sg13g2_o21ai_1 _33172_ (.B1(net3752),
    .Y(_10082_),
    .A1(_12112_),
    .A2(_10080_));
 sg13g2_a21oi_1 _33173_ (.A1(_12112_),
    .A2(_10080_),
    .Y(_10083_),
    .B1(_10082_));
 sg13g2_a21oi_1 _33174_ (.A1(net3679),
    .A2(_10079_),
    .Y(_10084_),
    .B1(_10083_));
 sg13g2_o21ai_1 _33175_ (.B1(net4013),
    .Y(_10085_),
    .A1(net4607),
    .A2(\u_inv.input_reg[236] ));
 sg13g2_o21ai_1 _33176_ (.B1(_10075_),
    .Y(_01540_),
    .A1(_10084_),
    .A2(_10085_));
 sg13g2_nand2_1 _33177_ (.Y(_10086_),
    .A(net1967),
    .B(net3926));
 sg13g2_a21oi_1 _33178_ (.A1(_12766_),
    .A2(_10065_),
    .Y(_10087_),
    .B1(_12792_));
 sg13g2_xnor2_1 _33179_ (.Y(_10088_),
    .A(_12116_),
    .B(_10087_));
 sg13g2_nor2_1 _33180_ (.A(\u_inv.f_next[238] ),
    .B(net4648),
    .Y(_10089_));
 sg13g2_a21oi_1 _33181_ (.A1(net4648),
    .A2(_10088_),
    .Y(_10090_),
    .B1(_10089_));
 sg13g2_or3_1 _33182_ (.A(_12116_),
    .B(_12139_),
    .C(_10081_),
    .X(_10091_));
 sg13g2_o21ai_1 _33183_ (.B1(_12116_),
    .Y(_10092_),
    .A1(_12139_),
    .A2(_10081_));
 sg13g2_a21o_1 _33184_ (.A2(_10092_),
    .A1(_10091_),
    .B1(net4438),
    .X(_10093_));
 sg13g2_a22oi_1 _33185_ (.Y(_10094_),
    .B1(_10093_),
    .B2(net3701),
    .A2(_10090_),
    .A1(net3831));
 sg13g2_o21ai_1 _33186_ (.B1(net4004),
    .Y(_10095_),
    .A1(net4604),
    .A2(\u_inv.input_reg[237] ));
 sg13g2_o21ai_1 _33187_ (.B1(_10086_),
    .Y(_01541_),
    .A1(_10094_),
    .A2(_10095_));
 sg13g2_nand2_1 _33188_ (.Y(_10096_),
    .A(net2764),
    .B(net3831));
 sg13g2_o21ai_1 _33189_ (.B1(_12115_),
    .Y(_10097_),
    .A1(_12116_),
    .A2(_10087_));
 sg13g2_xnor2_1 _33190_ (.Y(_10098_),
    .A(_12114_),
    .B(_10097_));
 sg13g2_a22oi_1 _33191_ (.Y(_10099_),
    .B1(_10098_),
    .B2(net4648),
    .A2(_10096_),
    .A1(net3724));
 sg13g2_nand2b_1 _33192_ (.Y(_10100_),
    .B(_10092_),
    .A_N(_12140_));
 sg13g2_xor2_1 _33193_ (.B(_10100_),
    .A(_12114_),
    .X(_10101_));
 sg13g2_o21ai_1 _33194_ (.B1(net4378),
    .Y(_10102_),
    .A1(net3831),
    .A2(_10101_));
 sg13g2_a21oi_1 _33195_ (.A1(net4511),
    .A2(_10984_),
    .Y(_10103_),
    .B1(net3926));
 sg13g2_o21ai_1 _33196_ (.B1(_10103_),
    .Y(_10104_),
    .A1(_10099_),
    .A2(_10102_));
 sg13g2_o21ai_1 _33197_ (.B1(_10104_),
    .Y(_01542_),
    .A1(_10343_),
    .A2(net4006));
 sg13g2_xnor2_1 _33198_ (.Y(_10105_),
    .A(_12152_),
    .B(_12158_));
 sg13g2_a21oi_1 _33199_ (.A1(net4511),
    .A2(net2205),
    .Y(_10106_),
    .B1(net3919));
 sg13g2_nand2_2 _33200_ (.Y(_10107_),
    .A(_12157_),
    .B(_12798_));
 sg13g2_nor2_1 _33201_ (.A(_12157_),
    .B(_12798_),
    .Y(_10108_));
 sg13g2_nor2_1 _33202_ (.A(net4526),
    .B(_10108_),
    .Y(_10109_));
 sg13g2_a22oi_1 _33203_ (.Y(_10110_),
    .B1(_10107_),
    .B2(_10109_),
    .A2(net4526),
    .A1(\u_inv.f_next[240] ));
 sg13g2_a21oi_1 _33204_ (.A1(net3825),
    .A2(_10110_),
    .Y(_10111_),
    .B1(net4434));
 sg13g2_o21ai_1 _33205_ (.B1(_10111_),
    .Y(_10112_),
    .A1(net3825),
    .A2(_10105_));
 sg13g2_a22oi_1 _33206_ (.Y(_01543_),
    .B1(_10106_),
    .B2(_10112_),
    .A2(net3919),
    .A1(_10342_));
 sg13g2_nand2_1 _33207_ (.Y(_10113_),
    .A(net2696),
    .B(net3915));
 sg13g2_o21ai_1 _33208_ (.B1(_12175_),
    .Y(_10114_),
    .A1(_12152_),
    .A2(_12157_));
 sg13g2_nand2_1 _33209_ (.Y(_10115_),
    .A(_12160_),
    .B(_10114_));
 sg13g2_o21ai_1 _33210_ (.B1(net3742),
    .Y(_10116_),
    .A1(_12160_),
    .A2(_10114_));
 sg13g2_nor2b_1 _33211_ (.A(_10116_),
    .B_N(_10115_),
    .Y(_10117_));
 sg13g2_nand2_1 _33212_ (.Y(_10118_),
    .A(\u_inv.f_next[241] ),
    .B(net3825));
 sg13g2_o21ai_1 _33213_ (.B1(_10107_),
    .Y(_10119_),
    .A1(_10341_),
    .A2(_10650_));
 sg13g2_xnor2_1 _33214_ (.Y(_10120_),
    .A(_12159_),
    .B(_10119_));
 sg13g2_a22oi_1 _33215_ (.Y(_10121_),
    .B1(_10120_),
    .B2(net4636),
    .A2(_10118_),
    .A1(net3722));
 sg13g2_nor3_1 _33216_ (.A(net4434),
    .B(_10117_),
    .C(_10121_),
    .Y(_10122_));
 sg13g2_o21ai_1 _33217_ (.B1(net4005),
    .Y(_10123_),
    .A1(net4603),
    .A2(net2004));
 sg13g2_o21ai_1 _33218_ (.B1(_10113_),
    .Y(_01544_),
    .A1(_10122_),
    .A2(_10123_));
 sg13g2_nand3_1 _33219_ (.B(_12174_),
    .C(_10115_),
    .A(_12155_),
    .Y(_10124_));
 sg13g2_a21o_1 _33220_ (.A2(_10115_),
    .A1(_12174_),
    .B1(_12155_),
    .X(_10125_));
 sg13g2_nand3_1 _33221_ (.B(_10124_),
    .C(_10125_),
    .A(net3690),
    .Y(_10126_));
 sg13g2_o21ai_1 _33222_ (.B1(_12231_),
    .Y(_10127_),
    .A1(_12160_),
    .A2(_10107_));
 sg13g2_xnor2_1 _33223_ (.Y(_10128_),
    .A(_12155_),
    .B(_10127_));
 sg13g2_o21ai_1 _33224_ (.B1(net3711),
    .Y(_10129_),
    .A1(net1826),
    .A2(net4637));
 sg13g2_a21oi_1 _33225_ (.A1(net4637),
    .A2(_10128_),
    .Y(_10130_),
    .B1(_10129_));
 sg13g2_a21oi_1 _33226_ (.A1(net4511),
    .A2(net2126),
    .Y(_10131_),
    .B1(net3916));
 sg13g2_nor2b_1 _33227_ (.A(_10130_),
    .B_N(_10131_),
    .Y(_10132_));
 sg13g2_a22oi_1 _33228_ (.Y(_01545_),
    .B1(_10126_),
    .B2(_10132_),
    .A2(net3916),
    .A1(_10340_));
 sg13g2_nand2_1 _33229_ (.Y(_10133_),
    .A(net1826),
    .B(net3916));
 sg13g2_a21oi_1 _33230_ (.A1(_12155_),
    .A2(_10127_),
    .Y(_10134_),
    .B1(_12154_));
 sg13g2_xor2_1 _33231_ (.B(_10134_),
    .A(_12153_),
    .X(_10135_));
 sg13g2_a21oi_1 _33232_ (.A1(\u_inv.f_next[243] ),
    .A2(net4526),
    .Y(_10136_),
    .B1(net4435));
 sg13g2_o21ai_1 _33233_ (.B1(_10136_),
    .Y(_10137_),
    .A1(net4528),
    .A2(_10135_));
 sg13g2_a21oi_1 _33234_ (.A1(_12173_),
    .A2(_10125_),
    .Y(_10138_),
    .B1(_12153_));
 sg13g2_nand3_1 _33235_ (.B(_12173_),
    .C(_10125_),
    .A(_12153_),
    .Y(_10139_));
 sg13g2_nor2_1 _33236_ (.A(net3827),
    .B(_10138_),
    .Y(_10140_));
 sg13g2_a22oi_1 _33237_ (.Y(_10141_),
    .B1(_10139_),
    .B2(_10140_),
    .A2(_10137_),
    .A1(net3679));
 sg13g2_o21ai_1 _33238_ (.B1(net4000),
    .Y(_10142_),
    .A1(net4603),
    .A2(\u_inv.input_reg[242] ));
 sg13g2_o21ai_1 _33239_ (.B1(_10133_),
    .Y(_01546_),
    .A1(_10141_),
    .A2(_10142_));
 sg13g2_nand2_1 _33240_ (.Y(_10143_),
    .A(net2181),
    .B(net3915));
 sg13g2_nor3_1 _33241_ (.A(_12160_),
    .B(_12229_),
    .C(_10107_),
    .Y(_10144_));
 sg13g2_nand2b_2 _33242_ (.Y(_10145_),
    .B(_12235_),
    .A_N(_10144_));
 sg13g2_xnor2_1 _33243_ (.Y(_10146_),
    .A(_12164_),
    .B(_10145_));
 sg13g2_nand2_1 _33244_ (.Y(_10147_),
    .A(_10337_),
    .B(net4526));
 sg13g2_a21oi_1 _33245_ (.A1(net4636),
    .A2(_10146_),
    .Y(_10148_),
    .B1(net3742));
 sg13g2_o21ai_1 _33246_ (.B1(_12178_),
    .Y(_10149_),
    .A1(_12152_),
    .A2(_12161_));
 sg13g2_xnor2_1 _33247_ (.Y(_10150_),
    .A(_12164_),
    .B(_10149_));
 sg13g2_a221oi_1 _33248_ (.B2(net3742),
    .C1(net4437),
    .B1(_10150_),
    .A1(_10147_),
    .Y(_10151_),
    .A2(_10148_));
 sg13g2_o21ai_1 _33249_ (.B1(net4005),
    .Y(_10152_),
    .A1(net4603),
    .A2(net1932));
 sg13g2_o21ai_1 _33250_ (.B1(_10143_),
    .Y(_01547_),
    .A1(_10151_),
    .A2(_10152_));
 sg13g2_nand2_1 _33251_ (.Y(_10153_),
    .A(net1439),
    .B(net3915));
 sg13g2_nand2_1 _33252_ (.Y(_10154_),
    .A(\u_inv.f_next[245] ),
    .B(net3826));
 sg13g2_a21oi_1 _33253_ (.A1(_12164_),
    .A2(_10145_),
    .Y(_10155_),
    .B1(_12163_));
 sg13g2_xor2_1 _33254_ (.B(_10155_),
    .A(_12162_),
    .X(_10156_));
 sg13g2_a22oi_1 _33255_ (.Y(_10157_),
    .B1(_10156_),
    .B2(net4636),
    .A2(_10154_),
    .A1(net3722));
 sg13g2_a21oi_1 _33256_ (.A1(_12165_),
    .A2(_10149_),
    .Y(_10158_),
    .B1(_12172_));
 sg13g2_nor2_1 _33257_ (.A(_12162_),
    .B(_10158_),
    .Y(_10159_));
 sg13g2_a21oi_1 _33258_ (.A1(_12162_),
    .A2(_10158_),
    .Y(_10160_),
    .B1(net3826));
 sg13g2_nor2b_1 _33259_ (.A(_10159_),
    .B_N(_10160_),
    .Y(_10161_));
 sg13g2_nor3_1 _33260_ (.A(net4437),
    .B(_10157_),
    .C(_10161_),
    .Y(_10162_));
 sg13g2_o21ai_1 _33261_ (.B1(net4005),
    .Y(_10163_),
    .A1(net4603),
    .A2(\u_inv.input_reg[244] ));
 sg13g2_o21ai_1 _33262_ (.B1(_10153_),
    .Y(_01548_),
    .A1(_10162_),
    .A2(_10163_));
 sg13g2_nand2_1 _33263_ (.Y(_10164_),
    .A(net2197),
    .B(net3915));
 sg13g2_o21ai_1 _33264_ (.B1(_12171_),
    .Y(_10165_),
    .A1(_12162_),
    .A2(_10158_));
 sg13g2_nor2_1 _33265_ (.A(_12168_),
    .B(_10165_),
    .Y(_10166_));
 sg13g2_nand2_1 _33266_ (.Y(_10167_),
    .A(_12168_),
    .B(_10165_));
 sg13g2_nor2_1 _33267_ (.A(net3826),
    .B(_10166_),
    .Y(_10168_));
 sg13g2_a21oi_1 _33268_ (.A1(_12227_),
    .A2(_10145_),
    .Y(_10169_),
    .B1(_12237_));
 sg13g2_xnor2_1 _33269_ (.Y(_10170_),
    .A(_12168_),
    .B(_10169_));
 sg13g2_nand2_1 _33270_ (.Y(_10171_),
    .A(_10335_),
    .B(net4526));
 sg13g2_a21oi_1 _33271_ (.A1(net4636),
    .A2(_10170_),
    .Y(_10172_),
    .B1(net3742));
 sg13g2_a221oi_1 _33272_ (.B2(_10172_),
    .C1(net4437),
    .B1(_10171_),
    .A1(_10167_),
    .Y(_10173_),
    .A2(_10168_));
 sg13g2_o21ai_1 _33273_ (.B1(net4005),
    .Y(_10174_),
    .A1(net4603),
    .A2(net1852));
 sg13g2_o21ai_1 _33274_ (.B1(_10164_),
    .Y(_01549_),
    .A1(_10173_),
    .A2(_10174_));
 sg13g2_nand2_1 _33275_ (.Y(_10175_),
    .A(net1661),
    .B(net3915));
 sg13g2_a21oi_1 _33276_ (.A1(_12168_),
    .A2(_10165_),
    .Y(_10176_),
    .B1(_12183_));
 sg13g2_xor2_1 _33277_ (.B(_10176_),
    .A(_12166_),
    .X(_10177_));
 sg13g2_nor2_1 _33278_ (.A(net3826),
    .B(_10177_),
    .Y(_10178_));
 sg13g2_nand2_1 _33279_ (.Y(_10179_),
    .A(\u_inv.f_next[247] ),
    .B(net3826));
 sg13g2_o21ai_1 _33280_ (.B1(_12167_),
    .Y(_10180_),
    .A1(_12168_),
    .A2(_10169_));
 sg13g2_xor2_1 _33281_ (.B(_10180_),
    .A(_12166_),
    .X(_10181_));
 sg13g2_a22oi_1 _33282_ (.Y(_10182_),
    .B1(_10181_),
    .B2(net4636),
    .A2(_10179_),
    .A1(net3722));
 sg13g2_nor3_1 _33283_ (.A(net4434),
    .B(_10178_),
    .C(_10182_),
    .Y(_10183_));
 sg13g2_o21ai_1 _33284_ (.B1(net4005),
    .Y(_10184_),
    .A1(net4603),
    .A2(\u_inv.input_reg[246] ));
 sg13g2_o21ai_1 _33285_ (.B1(_10175_),
    .Y(_01550_),
    .A1(_10183_),
    .A2(_10184_));
 sg13g2_nand2_1 _33286_ (.Y(_10185_),
    .A(net2336),
    .B(net3915));
 sg13g2_o21ai_1 _33287_ (.B1(net3742),
    .Y(_10186_),
    .A1(_12186_),
    .A2(_12188_));
 sg13g2_a21oi_1 _33288_ (.A1(_12186_),
    .A2(_12188_),
    .Y(_10187_),
    .B1(_10186_));
 sg13g2_xnor2_1 _33289_ (.Y(_10188_),
    .A(_12188_),
    .B(_12800_));
 sg13g2_o21ai_1 _33290_ (.B1(net3825),
    .Y(_10189_),
    .A1(\u_inv.f_next[248] ),
    .A2(net4636));
 sg13g2_a21oi_1 _33291_ (.A1(net4636),
    .A2(_10188_),
    .Y(_10190_),
    .B1(_10189_));
 sg13g2_nor3_1 _33292_ (.A(net4434),
    .B(_10187_),
    .C(_10190_),
    .Y(_10191_));
 sg13g2_o21ai_1 _33293_ (.B1(net4000),
    .Y(_10192_),
    .A1(net4603),
    .A2(net1965));
 sg13g2_o21ai_1 _33294_ (.B1(_10185_),
    .Y(_01551_),
    .A1(_10191_),
    .A2(_10192_));
 sg13g2_nand2_1 _33295_ (.Y(_10193_),
    .A(net2890),
    .B(net3915));
 sg13g2_a21oi_1 _33296_ (.A1(_12186_),
    .A2(_12188_),
    .Y(_10194_),
    .B1(_12197_));
 sg13g2_and2_1 _33297_ (.A(_12190_),
    .B(_10194_),
    .X(_10195_));
 sg13g2_nor2_1 _33298_ (.A(_12190_),
    .B(_10194_),
    .Y(_10196_));
 sg13g2_nor3_1 _33299_ (.A(net3825),
    .B(_10195_),
    .C(_10196_),
    .Y(_10197_));
 sg13g2_nand2_1 _33300_ (.Y(_10198_),
    .A(\u_inv.f_next[249] ),
    .B(net3825));
 sg13g2_o21ai_1 _33301_ (.B1(_12187_),
    .Y(_10199_),
    .A1(_12188_),
    .A2(_12800_));
 sg13g2_xnor2_1 _33302_ (.Y(_10200_),
    .A(_12190_),
    .B(_10199_));
 sg13g2_a22oi_1 _33303_ (.Y(_10201_),
    .B1(_10200_),
    .B2(net4637),
    .A2(_10198_),
    .A1(net3722));
 sg13g2_nor3_1 _33304_ (.A(net4434),
    .B(_10197_),
    .C(_10201_),
    .Y(_10202_));
 sg13g2_o21ai_1 _33305_ (.B1(net4000),
    .Y(_10203_),
    .A1(net4601),
    .A2(net2180));
 sg13g2_o21ai_1 _33306_ (.B1(_10193_),
    .Y(_01552_),
    .A1(_10202_),
    .A2(_10203_));
 sg13g2_nand2_1 _33307_ (.Y(_10204_),
    .A(net3171),
    .B(net3916));
 sg13g2_o21ai_1 _33308_ (.B1(_12193_),
    .Y(_10205_),
    .A1(_12196_),
    .A2(_10196_));
 sg13g2_nor3_1 _33309_ (.A(_12193_),
    .B(_12196_),
    .C(_10196_),
    .Y(_10206_));
 sg13g2_nor2_1 _33310_ (.A(net3826),
    .B(_10206_),
    .Y(_10207_));
 sg13g2_nor2b_1 _33311_ (.A(_12800_),
    .B_N(_12802_),
    .Y(_10208_));
 sg13g2_nor2_1 _33312_ (.A(_12806_),
    .B(_10208_),
    .Y(_10209_));
 sg13g2_xnor2_1 _33313_ (.Y(_10210_),
    .A(_12193_),
    .B(_10209_));
 sg13g2_nand2_1 _33314_ (.Y(_10211_),
    .A(_10331_),
    .B(net4526));
 sg13g2_a21oi_1 _33315_ (.A1(net4637),
    .A2(_10210_),
    .Y(_10212_),
    .B1(net3742));
 sg13g2_a221oi_1 _33316_ (.B2(_10212_),
    .C1(net4434),
    .B1(_10211_),
    .A1(_10205_),
    .Y(_10213_),
    .A2(_10207_));
 sg13g2_o21ai_1 _33317_ (.B1(net4001),
    .Y(_10214_),
    .A1(net4601),
    .A2(net1946));
 sg13g2_o21ai_1 _33318_ (.B1(_10204_),
    .Y(_01553_),
    .A1(_10213_),
    .A2(_10214_));
 sg13g2_nand2_1 _33319_ (.Y(_10215_),
    .A(_12195_),
    .B(_10205_));
 sg13g2_o21ai_1 _33320_ (.B1(net3689),
    .Y(_10216_),
    .A1(_12189_),
    .A2(_10215_));
 sg13g2_a21o_1 _33321_ (.A2(_10215_),
    .A1(_12189_),
    .B1(_10216_),
    .X(_10217_));
 sg13g2_o21ai_1 _33322_ (.B1(_12192_),
    .Y(_10218_),
    .A1(_12193_),
    .A2(_10209_));
 sg13g2_o21ai_1 _33323_ (.B1(net4638),
    .Y(_10219_),
    .A1(_12189_),
    .A2(_10218_));
 sg13g2_a21oi_1 _33324_ (.A1(_12189_),
    .A2(_10218_),
    .Y(_10220_),
    .B1(_10219_));
 sg13g2_o21ai_1 _33325_ (.B1(net3713),
    .Y(_10221_),
    .A1(\u_inv.f_next[251] ),
    .A2(net4639));
 sg13g2_nand2_1 _33326_ (.Y(_10222_),
    .A(net4512),
    .B(net1723));
 sg13g2_o21ai_1 _33327_ (.B1(_10222_),
    .Y(_10223_),
    .A1(_10220_),
    .A2(_10221_));
 sg13g2_nor2_1 _33328_ (.A(net3916),
    .B(_10223_),
    .Y(_10224_));
 sg13g2_a22oi_1 _33329_ (.Y(_01554_),
    .B1(_10217_),
    .B2(_10224_),
    .A2(net3916),
    .A1(_10331_));
 sg13g2_nand2b_1 _33330_ (.Y(_10225_),
    .B(_12206_),
    .A_N(_12202_));
 sg13g2_a21oi_1 _33331_ (.A1(_12202_),
    .A2(_12205_),
    .Y(_10226_),
    .B1(net3827));
 sg13g2_nand2_1 _33332_ (.Y(_10227_),
    .A(_12205_),
    .B(_12808_));
 sg13g2_xnor2_1 _33333_ (.Y(_10228_),
    .A(_12205_),
    .B(_12808_));
 sg13g2_o21ai_1 _33334_ (.B1(net3827),
    .Y(_10229_),
    .A1(\u_inv.f_next[252] ),
    .A2(net4638));
 sg13g2_a21oi_1 _33335_ (.A1(net4638),
    .A2(_10228_),
    .Y(_10230_),
    .B1(_10229_));
 sg13g2_a21oi_1 _33336_ (.A1(_10225_),
    .A2(_10226_),
    .Y(_10231_),
    .B1(_10230_));
 sg13g2_o21ai_1 _33337_ (.B1(net4001),
    .Y(_10232_),
    .A1(net4601),
    .A2(net1756));
 sg13g2_a21o_1 _33338_ (.A2(_10231_),
    .A1(net4379),
    .B1(_10232_),
    .X(_10233_));
 sg13g2_o21ai_1 _33339_ (.B1(_10233_),
    .Y(_01555_),
    .A1(_10330_),
    .A2(net4000));
 sg13g2_nand2_1 _33340_ (.Y(_10234_),
    .A(net2244),
    .B(net3916));
 sg13g2_nand2_1 _33341_ (.Y(_10235_),
    .A(_12204_),
    .B(_10227_));
 sg13g2_xor2_1 _33342_ (.B(_10235_),
    .A(_12203_),
    .X(_10236_));
 sg13g2_nand2_1 _33343_ (.Y(_10237_),
    .A(\u_inv.f_next[253] ),
    .B(net3827));
 sg13g2_a22oi_1 _33344_ (.Y(_10238_),
    .B1(_10237_),
    .B2(net3722),
    .A2(_10236_),
    .A1(net4638));
 sg13g2_nand2b_1 _33345_ (.Y(_10239_),
    .B(_10225_),
    .A_N(_12209_));
 sg13g2_nor2_1 _33346_ (.A(_12203_),
    .B(_10239_),
    .Y(_10240_));
 sg13g2_a21o_1 _33347_ (.A2(_10239_),
    .A1(_12203_),
    .B1(net3827),
    .X(_10241_));
 sg13g2_o21ai_1 _33348_ (.B1(net4379),
    .Y(_10242_),
    .A1(_10240_),
    .A2(_10241_));
 sg13g2_nor2_1 _33349_ (.A(net4601),
    .B(net1948),
    .Y(_10243_));
 sg13g2_o21ai_1 _33350_ (.B1(net4000),
    .Y(_10244_),
    .A1(_10238_),
    .A2(_10242_));
 sg13g2_o21ai_1 _33351_ (.B1(_10234_),
    .Y(_01556_),
    .A1(_10243_),
    .A2(_10244_));
 sg13g2_nand2_1 _33352_ (.Y(_10245_),
    .A(_11077_),
    .B(_12211_));
 sg13g2_o21ai_1 _33353_ (.B1(net3742),
    .Y(_10246_),
    .A1(_11077_),
    .A2(_12211_));
 sg13g2_nand2b_1 _33354_ (.Y(_10247_),
    .B(_10245_),
    .A_N(_10246_));
 sg13g2_xnor2_1 _33355_ (.Y(_10248_),
    .A(_11077_),
    .B(_12811_));
 sg13g2_o21ai_1 _33356_ (.B1(net3827),
    .Y(_10249_),
    .A1(\u_inv.f_next[254] ),
    .A2(net4638));
 sg13g2_a21oi_1 _33357_ (.A1(net4638),
    .A2(_10248_),
    .Y(_10250_),
    .B1(_10249_));
 sg13g2_nor2_1 _33358_ (.A(net4435),
    .B(_10250_),
    .Y(_10251_));
 sg13g2_o21ai_1 _33359_ (.B1(net4001),
    .Y(_10252_),
    .A1(net4601),
    .A2(net1952));
 sg13g2_a21o_1 _33360_ (.A2(_10251_),
    .A1(_10247_),
    .B1(_10252_),
    .X(_10253_));
 sg13g2_o21ai_1 _33361_ (.B1(_10253_),
    .Y(_01557_),
    .A1(_10328_),
    .A2(net4000));
 sg13g2_nand2_1 _33362_ (.Y(_10254_),
    .A(net2535),
    .B(net3917));
 sg13g2_nand2_1 _33363_ (.Y(_10255_),
    .A(net2560),
    .B(net3827));
 sg13g2_o21ai_1 _33364_ (.B1(_11076_),
    .Y(_10256_),
    .A1(_11077_),
    .A2(_12811_));
 sg13g2_xnor2_1 _33365_ (.Y(_10257_),
    .A(_11072_),
    .B(_10256_));
 sg13g2_a22oi_1 _33366_ (.Y(_10258_),
    .B1(_10257_),
    .B2(net4638),
    .A2(_10255_),
    .A1(net3722));
 sg13g2_and3_1 _33367_ (.X(_10259_),
    .A(_11072_),
    .B(_11073_),
    .C(_10245_));
 sg13g2_a21oi_1 _33368_ (.A1(_11073_),
    .A2(_10245_),
    .Y(_10260_),
    .B1(_11072_));
 sg13g2_nor3_1 _33369_ (.A(net3828),
    .B(_10259_),
    .C(_10260_),
    .Y(_10261_));
 sg13g2_nor3_1 _33370_ (.A(net4435),
    .B(_10258_),
    .C(_10261_),
    .Y(_10262_));
 sg13g2_o21ai_1 _33371_ (.B1(net4001),
    .Y(_10263_),
    .A1(net4601),
    .A2(net2010));
 sg13g2_o21ai_1 _33372_ (.B1(_10254_),
    .Y(_01558_),
    .A1(_10262_),
    .A2(_10263_));
 sg13g2_nand2_1 _33373_ (.Y(_10264_),
    .A(net2530),
    .B(net3917));
 sg13g2_nor2_1 _33374_ (.A(_11070_),
    .B(_12212_),
    .Y(_10265_));
 sg13g2_nor2b_1 _33375_ (.A(_10265_),
    .B_N(_12223_),
    .Y(_10266_));
 sg13g2_nand2_1 _33376_ (.Y(_10267_),
    .A(\u_inv.f_next[256] ),
    .B(net3825));
 sg13g2_nand3_1 _33377_ (.B(_11071_),
    .C(_12813_),
    .A(_11070_),
    .Y(_10268_));
 sg13g2_nor2_1 _33378_ (.A(net4526),
    .B(_12814_),
    .Y(_10269_));
 sg13g2_a22oi_1 _33379_ (.Y(_10270_),
    .B1(_10268_),
    .B2(_10269_),
    .A2(_10267_),
    .A1(net3722));
 sg13g2_nor3_1 _33380_ (.A(net4434),
    .B(_10266_),
    .C(_10270_),
    .Y(_10271_));
 sg13g2_o21ai_1 _33381_ (.B1(net4001),
    .Y(_10272_),
    .A1(net4602),
    .A2(net2037));
 sg13g2_o21ai_1 _33382_ (.B1(_10264_),
    .Y(_01559_),
    .A1(_10271_),
    .A2(_10272_));
 sg13g2_nor2_1 _33383_ (.A(net1857),
    .B(net1227),
    .Y(_10273_));
 sg13g2_nor4_1 _33384_ (.A(net1562),
    .B(net1088),
    .C(_13579_),
    .D(_13592_),
    .Y(_10274_));
 sg13g2_and4_1 _33385_ (.A(net2119),
    .B(net1067),
    .C(_10273_),
    .D(_10274_),
    .X(_10275_));
 sg13g2_o21ai_1 _33386_ (.B1(net4965),
    .Y(_01560_),
    .A1(net4435),
    .A2(_10275_));
 sg13g2_nand2_1 _33387_ (.Y(_10276_),
    .A(net4379),
    .B(_10275_));
 sg13g2_o21ai_1 _33388_ (.B1(_10276_),
    .Y(_01561_),
    .A1(_11043_),
    .A2(_11046_));
 sg13g2_nor3_1 _33389_ (.A(\u_inv.input_valid ),
    .B(_10632_),
    .C(\u_inv.load_input ),
    .Y(_10277_));
 sg13g2_nor2_1 _33390_ (.A(\u_inv.input_reg[0] ),
    .B(net4245),
    .Y(_10278_));
 sg13g2_a21oi_1 _33391_ (.A1(_10988_),
    .A2(net4245),
    .Y(_01562_),
    .B1(_10278_));
 sg13g2_nor2_1 _33392_ (.A(net1529),
    .B(net4243),
    .Y(_10279_));
 sg13g2_a21oi_1 _33393_ (.A1(_10989_),
    .A2(net4243),
    .Y(_01563_),
    .B1(_10279_));
 sg13g2_nor2_1 _33394_ (.A(net1621),
    .B(net4243),
    .Y(_10280_));
 sg13g2_a21oi_1 _33395_ (.A1(_10990_),
    .A2(net4243),
    .Y(_01564_),
    .B1(_10280_));
 sg13g2_nor2_1 _33396_ (.A(net1267),
    .B(net4243),
    .Y(_10281_));
 sg13g2_a21oi_1 _33397_ (.A1(_10991_),
    .A2(net4243),
    .Y(_01565_),
    .B1(_10281_));
 sg13g2_nor2_1 _33398_ (.A(net1214),
    .B(net4243),
    .Y(_10282_));
 sg13g2_a21oi_1 _33399_ (.A1(_10992_),
    .A2(net4244),
    .Y(_01566_),
    .B1(_10282_));
 sg13g2_nor2_1 _33400_ (.A(net1300),
    .B(net4244),
    .Y(_10283_));
 sg13g2_a21oi_1 _33401_ (.A1(_10993_),
    .A2(net4244),
    .Y(_01567_),
    .B1(_10283_));
 sg13g2_nor2_1 _33402_ (.A(\u_inv.input_reg[6] ),
    .B(net4244),
    .Y(_10284_));
 sg13g2_a21oi_1 _33403_ (.A1(_10994_),
    .A2(net4243),
    .Y(_01568_),
    .B1(_10284_));
 sg13g2_nor2_1 _33404_ (.A(net1670),
    .B(net4245),
    .Y(_10285_));
 sg13g2_a21oi_1 _33405_ (.A1(_10995_),
    .A2(net4245),
    .Y(_01569_),
    .B1(_10285_));
 sg13g2_mux2_1 _33406_ (.A0(net2059),
    .A1(net1446),
    .S(net4245),
    .X(_01570_));
 sg13g2_mux2_1 _33407_ (.A0(net1815),
    .A1(net1249),
    .S(net4244),
    .X(_01571_));
 sg13g2_mux2_1 _33408_ (.A0(net1999),
    .A1(net1593),
    .S(net4244),
    .X(_01572_));
 sg13g2_mux2_1 _33409_ (.A0(net1963),
    .A1(net1241),
    .S(net4244),
    .X(_01573_));
 sg13g2_mux2_1 _33410_ (.A0(net1862),
    .A1(net1212),
    .S(net4251),
    .X(_01574_));
 sg13g2_mux2_1 _33411_ (.A0(net1875),
    .A1(net1143),
    .S(net4251),
    .X(_01575_));
 sg13g2_mux2_1 _33412_ (.A0(net1811),
    .A1(\shift_reg[14] ),
    .S(net4251),
    .X(_01576_));
 sg13g2_mux2_1 _33413_ (.A0(net1785),
    .A1(\shift_reg[15] ),
    .S(net4251),
    .X(_01577_));
 sg13g2_mux2_1 _33414_ (.A0(net1683),
    .A1(\shift_reg[16] ),
    .S(net4251),
    .X(_01578_));
 sg13g2_mux2_1 _33415_ (.A0(net1845),
    .A1(\shift_reg[17] ),
    .S(net4251),
    .X(_01579_));
 sg13g2_mux2_1 _33416_ (.A0(net1619),
    .A1(\shift_reg[18] ),
    .S(net4251),
    .X(_01580_));
 sg13g2_mux2_1 _33417_ (.A0(net1855),
    .A1(\shift_reg[19] ),
    .S(net4251),
    .X(_01581_));
 sg13g2_mux2_1 _33418_ (.A0(net2065),
    .A1(net1419),
    .S(net4253),
    .X(_01582_));
 sg13g2_mux2_1 _33419_ (.A0(net1962),
    .A1(net1251),
    .S(net4252),
    .X(_01583_));
 sg13g2_mux2_1 _33420_ (.A0(net1937),
    .A1(net1359),
    .S(net4252),
    .X(_01584_));
 sg13g2_mux2_1 _33421_ (.A0(net1912),
    .A1(net1487),
    .S(net4252),
    .X(_01585_));
 sg13g2_mux2_1 _33422_ (.A0(net2009),
    .A1(net1633),
    .S(net4252),
    .X(_01586_));
 sg13g2_mux2_1 _33423_ (.A0(net1737),
    .A1(net1230),
    .S(net4252),
    .X(_01587_));
 sg13g2_mux2_1 _33424_ (.A0(net1758),
    .A1(net1210),
    .S(net4252),
    .X(_01588_));
 sg13g2_mux2_1 _33425_ (.A0(net1837),
    .A1(net1584),
    .S(net4253),
    .X(_01589_));
 sg13g2_mux2_1 _33426_ (.A0(net1784),
    .A1(net1160),
    .S(net4252),
    .X(_01590_));
 sg13g2_mux2_1 _33427_ (.A0(net1747),
    .A1(net1461),
    .S(net4252),
    .X(_01591_));
 sg13g2_mux2_1 _33428_ (.A0(net1722),
    .A1(net1155),
    .S(net4256),
    .X(_01592_));
 sg13g2_mux2_1 _33429_ (.A0(net1663),
    .A1(net1148),
    .S(net4256),
    .X(_01593_));
 sg13g2_mux2_1 _33430_ (.A0(net1694),
    .A1(net1384),
    .S(net4256),
    .X(_01594_));
 sg13g2_mux2_1 _33431_ (.A0(net1717),
    .A1(net1132),
    .S(net4256),
    .X(_01595_));
 sg13g2_mux2_1 _33432_ (.A0(net1695),
    .A1(net1388),
    .S(net4256),
    .X(_01596_));
 sg13g2_mux2_1 _33433_ (.A0(net1795),
    .A1(net1162),
    .S(net4256),
    .X(_01597_));
 sg13g2_mux2_1 _33434_ (.A0(net1940),
    .A1(net1429),
    .S(net4256),
    .X(_01598_));
 sg13g2_mux2_1 _33435_ (.A0(net1802),
    .A1(net1355),
    .S(net4257),
    .X(_01599_));
 sg13g2_mux2_1 _33436_ (.A0(net1814),
    .A1(net1261),
    .S(net4257),
    .X(_01600_));
 sg13g2_mux2_1 _33437_ (.A0(net1993),
    .A1(net1479),
    .S(net4256),
    .X(_01601_));
 sg13g2_mux2_1 _33438_ (.A0(net1767),
    .A1(net1336),
    .S(net4258),
    .X(_01602_));
 sg13g2_mux2_1 _33439_ (.A0(net1902),
    .A1(net1310),
    .S(net4258),
    .X(_01603_));
 sg13g2_mux2_1 _33440_ (.A0(net1860),
    .A1(net1274),
    .S(net4257),
    .X(_01604_));
 sg13g2_mux2_1 _33441_ (.A0(net1863),
    .A1(net1483),
    .S(net4259),
    .X(_01605_));
 sg13g2_mux2_1 _33442_ (.A0(net2015),
    .A1(net1151),
    .S(net4258),
    .X(_01606_));
 sg13g2_mux2_1 _33443_ (.A0(net1978),
    .A1(\shift_reg[45] ),
    .S(net4258),
    .X(_01607_));
 sg13g2_mux2_1 _33444_ (.A0(net1720),
    .A1(\shift_reg[46] ),
    .S(net4258),
    .X(_01608_));
 sg13g2_mux2_1 _33445_ (.A0(net1803),
    .A1(net1711),
    .S(net4258),
    .X(_01609_));
 sg13g2_mux2_1 _33446_ (.A0(net1718),
    .A1(\shift_reg[48] ),
    .S(net4264),
    .X(_01610_));
 sg13g2_mux2_1 _33447_ (.A0(net1779),
    .A1(net1420),
    .S(net4261),
    .X(_01611_));
 sg13g2_mux2_1 _33448_ (.A0(net1838),
    .A1(net1198),
    .S(net4261),
    .X(_01612_));
 sg13g2_mux2_1 _33449_ (.A0(net1872),
    .A1(net1123),
    .S(net4261),
    .X(_01613_));
 sg13g2_mux2_1 _33450_ (.A0(net2304),
    .A1(net1278),
    .S(net4264),
    .X(_01614_));
 sg13g2_mux2_1 _33451_ (.A0(net1780),
    .A1(net1541),
    .S(net4264),
    .X(_01615_));
 sg13g2_mux2_1 _33452_ (.A0(net1750),
    .A1(net1284),
    .S(net4263),
    .X(_01616_));
 sg13g2_mux2_1 _33453_ (.A0(net2184),
    .A1(net1232),
    .S(net4261),
    .X(_01617_));
 sg13g2_mux2_1 _33454_ (.A0(net2104),
    .A1(net1350),
    .S(net4262),
    .X(_01618_));
 sg13g2_mux2_1 _33455_ (.A0(net1725),
    .A1(net1650),
    .S(net4261),
    .X(_01619_));
 sg13g2_mux2_1 _33456_ (.A0(net1801),
    .A1(net1572),
    .S(net4262),
    .X(_01620_));
 sg13g2_mux2_1 _33457_ (.A0(net2046),
    .A1(net1383),
    .S(net4262),
    .X(_01621_));
 sg13g2_mux2_1 _33458_ (.A0(net1919),
    .A1(net1589),
    .S(net4262),
    .X(_01622_));
 sg13g2_mux2_1 _33459_ (.A0(net1764),
    .A1(\shift_reg[61] ),
    .S(net4262),
    .X(_01623_));
 sg13g2_mux2_1 _33460_ (.A0(net2453),
    .A1(net1332),
    .S(net4263),
    .X(_01624_));
 sg13g2_mux2_1 _33461_ (.A0(net2114),
    .A1(net1519),
    .S(net4262),
    .X(_01625_));
 sg13g2_mux2_1 _33462_ (.A0(net1798),
    .A1(net1579),
    .S(net4262),
    .X(_01626_));
 sg13g2_mux2_1 _33463_ (.A0(net1741),
    .A1(net1473),
    .S(net4262),
    .X(_01627_));
 sg13g2_mux2_1 _33464_ (.A0(net1813),
    .A1(net1485),
    .S(net4270),
    .X(_01628_));
 sg13g2_mux2_1 _33465_ (.A0(net2042),
    .A1(net1386),
    .S(net4270),
    .X(_01629_));
 sg13g2_mux2_1 _33466_ (.A0(net1983),
    .A1(net1286),
    .S(net4267),
    .X(_01630_));
 sg13g2_mux2_1 _33467_ (.A0(net2118),
    .A1(net1157),
    .S(net4270),
    .X(_01631_));
 sg13g2_mux2_1 _33468_ (.A0(net2111),
    .A1(net1408),
    .S(net4267),
    .X(_01632_));
 sg13g2_mux2_1 _33469_ (.A0(net2265),
    .A1(net1257),
    .S(net4267),
    .X(_01633_));
 sg13g2_mux2_1 _33470_ (.A0(net2027),
    .A1(net1208),
    .S(net4267),
    .X(_01634_));
 sg13g2_mux2_1 _33471_ (.A0(net1955),
    .A1(net1570),
    .S(net4267),
    .X(_01635_));
 sg13g2_mux2_1 _33472_ (.A0(net2496),
    .A1(net1238),
    .S(net4269),
    .X(_01636_));
 sg13g2_mux2_1 _33473_ (.A0(net1923),
    .A1(net1402),
    .S(net4267),
    .X(_01637_));
 sg13g2_mux2_1 _33474_ (.A0(net1715),
    .A1(net1459),
    .S(net4267),
    .X(_01638_));
 sg13g2_mux2_1 _33475_ (.A0(net1895),
    .A1(net1477),
    .S(net4268),
    .X(_01639_));
 sg13g2_mux2_1 _33476_ (.A0(net1708),
    .A1(net1380),
    .S(net4267),
    .X(_01640_));
 sg13g2_mux2_1 _33477_ (.A0(net1847),
    .A1(net1317),
    .S(net4268),
    .X(_01641_));
 sg13g2_mux2_1 _33478_ (.A0(net1974),
    .A1(net1339),
    .S(net4268),
    .X(_01642_));
 sg13g2_mux2_1 _33479_ (.A0(net2099),
    .A1(net1282),
    .S(net4268),
    .X(_01643_));
 sg13g2_mux2_1 _33480_ (.A0(net2597),
    .A1(net1465),
    .S(net4269),
    .X(_01644_));
 sg13g2_mux2_1 _33481_ (.A0(net1858),
    .A1(net1343),
    .S(net4268),
    .X(_01645_));
 sg13g2_mux2_1 _33482_ (.A0(net2268),
    .A1(net1471),
    .S(net4268),
    .X(_01646_));
 sg13g2_mux2_1 _33483_ (.A0(net2025),
    .A1(net1253),
    .S(net4268),
    .X(_01647_));
 sg13g2_mux2_1 _33484_ (.A0(net2182),
    .A1(net1444),
    .S(net4268),
    .X(_01648_));
 sg13g2_mux2_1 _33485_ (.A0(net1861),
    .A1(net1247),
    .S(net4269),
    .X(_01649_));
 sg13g2_mux2_1 _33486_ (.A0(net2204),
    .A1(net1291),
    .S(net4272),
    .X(_01650_));
 sg13g2_mux2_1 _33487_ (.A0(net1886),
    .A1(net1328),
    .S(net4271),
    .X(_01651_));
 sg13g2_mux2_1 _33488_ (.A0(net1682),
    .A1(net1378),
    .S(net4271),
    .X(_01652_));
 sg13g2_mux2_1 _33489_ (.A0(net1733),
    .A1(net1615),
    .S(net4271),
    .X(_01653_));
 sg13g2_mux2_1 _33490_ (.A0(net1920),
    .A1(net1481),
    .S(net4271),
    .X(_01654_));
 sg13g2_mux2_1 _33491_ (.A0(net2385),
    .A1(net1204),
    .S(net4271),
    .X(_01655_));
 sg13g2_mux2_1 _33492_ (.A0(net2071),
    .A1(net1330),
    .S(net4272),
    .X(_01656_));
 sg13g2_mux2_1 _33493_ (.A0(net1637),
    .A1(\shift_reg[95] ),
    .S(net4271),
    .X(_01657_));
 sg13g2_mux2_1 _33494_ (.A0(net2398),
    .A1(net1731),
    .S(net4275),
    .X(_01658_));
 sg13g2_mux2_1 _33495_ (.A0(net2541),
    .A1(net1361),
    .S(net4273),
    .X(_01659_));
 sg13g2_mux2_1 _33496_ (.A0(net1929),
    .A1(net1899),
    .S(net4275),
    .X(_01660_));
 sg13g2_mux2_1 _33497_ (.A0(net2157),
    .A1(net1469),
    .S(net4274),
    .X(_01661_));
 sg13g2_mux2_1 _33498_ (.A0(net1980),
    .A1(net1766),
    .S(net4275),
    .X(_01662_));
 sg13g2_mux2_1 _33499_ (.A0(net1876),
    .A1(\shift_reg[101] ),
    .S(net4287),
    .X(_01663_));
 sg13g2_mux2_1 _33500_ (.A0(net2075),
    .A1(net1991),
    .S(net4275),
    .X(_01664_));
 sg13g2_mux2_1 _33501_ (.A0(net2289),
    .A1(net2183),
    .S(net4275),
    .X(_01665_));
 sg13g2_mux2_1 _33502_ (.A0(net2443),
    .A1(net1736),
    .S(net4276),
    .X(_01666_));
 sg13g2_mux2_1 _33503_ (.A0(net1998),
    .A1(net1173),
    .S(net4276),
    .X(_01667_));
 sg13g2_mux2_1 _33504_ (.A0(net1951),
    .A1(net1396),
    .S(net4276),
    .X(_01668_));
 sg13g2_mux2_1 _33505_ (.A0(net2085),
    .A1(net1404),
    .S(net4277),
    .X(_01669_));
 sg13g2_mux2_1 _33506_ (.A0(net1888),
    .A1(net1196),
    .S(net4282),
    .X(_01670_));
 sg13g2_mux2_1 _33507_ (.A0(net2117),
    .A1(net1864),
    .S(net4286),
    .X(_01671_));
 sg13g2_mux2_1 _33508_ (.A0(net2408),
    .A1(net1776),
    .S(net4277),
    .X(_01672_));
 sg13g2_mux2_1 _33509_ (.A0(net2621),
    .A1(net2161),
    .S(net4277),
    .X(_01673_));
 sg13g2_mux2_1 _33510_ (.A0(net2557),
    .A1(net1353),
    .S(net4276),
    .X(_01674_));
 sg13g2_mux2_1 _33511_ (.A0(net1793),
    .A1(net1629),
    .S(net4284),
    .X(_01675_));
 sg13g2_mux2_1 _33512_ (.A0(net2031),
    .A1(net1107),
    .S(net4277),
    .X(_01676_));
 sg13g2_mux2_1 _33513_ (.A0(net2286),
    .A1(net1922),
    .S(net4285),
    .X(_01677_));
 sg13g2_mux2_1 _33514_ (.A0(net1894),
    .A1(net1635),
    .S(net4284),
    .X(_01678_));
 sg13g2_mux2_1 _33515_ (.A0(net2179),
    .A1(net1259),
    .S(net4285),
    .X(_01679_));
 sg13g2_mux2_1 _33516_ (.A0(net2654),
    .A1(net1961),
    .S(net4285),
    .X(_01680_));
 sg13g2_mux2_1 _33517_ (.A0(net2451),
    .A1(net1774),
    .S(net4285),
    .X(_01681_));
 sg13g2_mux2_1 _33518_ (.A0(net2252),
    .A1(net1889),
    .S(net4284),
    .X(_01682_));
 sg13g2_mux2_1 _33519_ (.A0(net2667),
    .A1(net1500),
    .S(net4284),
    .X(_01683_));
 sg13g2_mux2_1 _33520_ (.A0(net2299),
    .A1(net1417),
    .S(net4284),
    .X(_01684_));
 sg13g2_mux2_1 _33521_ (.A0(net1904),
    .A1(net1698),
    .S(net4283),
    .X(_01685_));
 sg13g2_mux2_1 _33522_ (.A0(net2105),
    .A1(net1180),
    .S(net4283),
    .X(_01686_));
 sg13g2_mux2_1 _33523_ (.A0(net2079),
    .A1(net1986),
    .S(net4284),
    .X(_01687_));
 sg13g2_mux2_1 _33524_ (.A0(net1740),
    .A1(net1530),
    .S(net4284),
    .X(_01688_));
 sg13g2_mux2_1 _33525_ (.A0(net2323),
    .A1(net1112),
    .S(net4283),
    .X(_01689_));
 sg13g2_mux2_1 _33526_ (.A0(net2020),
    .A1(net1326),
    .S(net4281),
    .X(_01690_));
 sg13g2_mux2_1 _33527_ (.A0(net1853),
    .A1(net1555),
    .S(net4281),
    .X(_01691_));
 sg13g2_mux2_1 _33528_ (.A0(net1817),
    .A1(net1606),
    .S(net4281),
    .X(_01692_));
 sg13g2_mux2_1 _33529_ (.A0(net2054),
    .A1(net1288),
    .S(net4281),
    .X(_01693_));
 sg13g2_mux2_1 _33530_ (.A0(net2008),
    .A1(net1218),
    .S(net4279),
    .X(_01694_));
 sg13g2_mux2_1 _33531_ (.A0(net1934),
    .A1(net1265),
    .S(net4278),
    .X(_01695_));
 sg13g2_mux2_1 _33532_ (.A0(net1938),
    .A1(net1414),
    .S(net4279),
    .X(_01696_));
 sg13g2_mux2_1 _33533_ (.A0(net2062),
    .A1(net1394),
    .S(net4278),
    .X(_01697_));
 sg13g2_mux2_1 _33534_ (.A0(net1787),
    .A1(net1221),
    .S(net4278),
    .X(_01698_));
 sg13g2_mux2_1 _33535_ (.A0(net1751),
    .A1(\shift_reg[137] ),
    .S(net4278),
    .X(_01699_));
 sg13g2_mux2_1 _33536_ (.A0(net2319),
    .A1(net1178),
    .S(net4278),
    .X(_01700_));
 sg13g2_mux2_1 _33537_ (.A0(net2026),
    .A1(net1234),
    .S(net4278),
    .X(_01701_));
 sg13g2_mux2_1 _33538_ (.A0(net1958),
    .A1(net1364),
    .S(net4278),
    .X(_01702_));
 sg13g2_mux2_1 _33539_ (.A0(net2225),
    .A1(net1517),
    .S(net4279),
    .X(_01703_));
 sg13g2_mux2_1 _33540_ (.A0(net2463),
    .A1(net1592),
    .S(net4279),
    .X(_01704_));
 sg13g2_mux2_1 _33541_ (.A0(net1939),
    .A1(net1648),
    .S(net4278),
    .X(_01705_));
 sg13g2_mux2_1 _33542_ (.A0(net1925),
    .A1(net1536),
    .S(net4280),
    .X(_01706_));
 sg13g2_mux2_1 _33543_ (.A0(net1928),
    .A1(net1489),
    .S(net4280),
    .X(_01707_));
 sg13g2_mux2_1 _33544_ (.A0(net2534),
    .A1(net1869),
    .S(net4280),
    .X(_01708_));
 sg13g2_mux2_1 _33545_ (.A0(net1981),
    .A1(net1612),
    .S(net4280),
    .X(_01709_));
 sg13g2_mux2_1 _33546_ (.A0(net2135),
    .A1(net1496),
    .S(net4280),
    .X(_01710_));
 sg13g2_mux2_1 _33547_ (.A0(net2433),
    .A1(net1524),
    .S(net4281),
    .X(_01711_));
 sg13g2_mux2_1 _33548_ (.A0(net2016),
    .A1(net1917),
    .S(net4280),
    .X(_01712_));
 sg13g2_mux2_1 _33549_ (.A0(net1989),
    .A1(net1600),
    .S(net4280),
    .X(_01713_));
 sg13g2_mux2_1 _33550_ (.A0(net2488),
    .A1(net2439),
    .S(net4280),
    .X(_01714_));
 sg13g2_mux2_1 _33551_ (.A0(net1819),
    .A1(\shift_reg[153] ),
    .S(net4285),
    .X(_01715_));
 sg13g2_mux2_1 _33552_ (.A0(net2698),
    .A1(net1657),
    .S(net4283),
    .X(_01716_));
 sg13g2_mux2_1 _33553_ (.A0(net2550),
    .A1(net1644),
    .S(net4283),
    .X(_01717_));
 sg13g2_mux2_1 _33554_ (.A0(net1831),
    .A1(\shift_reg[156] ),
    .S(net4285),
    .X(_01718_));
 sg13g2_mux2_1 _33555_ (.A0(net2239),
    .A1(net1545),
    .S(net4283),
    .X(_01719_));
 sg13g2_mux2_1 _33556_ (.A0(net2216),
    .A1(net1673),
    .S(net4283),
    .X(_01720_));
 sg13g2_mux2_1 _33557_ (.A0(net1219),
    .A1(net1679),
    .S(net4283),
    .X(_01721_));
 sg13g2_mux2_1 _33558_ (.A0(net1947),
    .A1(net1276),
    .S(net4284),
    .X(_01722_));
 sg13g2_mux2_1 _33559_ (.A0(net1887),
    .A1(net1365),
    .S(net4282),
    .X(_01723_));
 sg13g2_mux2_1 _33560_ (.A0(net1972),
    .A1(net1312),
    .S(net4286),
    .X(_01724_));
 sg13g2_mux2_1 _33561_ (.A0(net1818),
    .A1(net1702),
    .S(net4282),
    .X(_01725_));
 sg13g2_mux2_1 _33562_ (.A0(net1896),
    .A1(net1243),
    .S(net4282),
    .X(_01726_));
 sg13g2_mux2_1 _33563_ (.A0(net1882),
    .A1(net1651),
    .S(net4282),
    .X(_01727_));
 sg13g2_mux2_1 _33564_ (.A0(net2000),
    .A1(net1269),
    .S(net4282),
    .X(_01728_));
 sg13g2_mux2_1 _33565_ (.A0(net1885),
    .A1(net1435),
    .S(net4282),
    .X(_01729_));
 sg13g2_mux2_1 _33566_ (.A0(net1851),
    .A1(net1554),
    .S(net4282),
    .X(_01730_));
 sg13g2_mux2_1 _33567_ (.A0(net1975),
    .A1(net1441),
    .S(net4277),
    .X(_01731_));
 sg13g2_mux2_1 _33568_ (.A0(net2426),
    .A1(net1333),
    .S(net4277),
    .X(_01732_));
 sg13g2_mux2_1 _33569_ (.A0(net1848),
    .A1(net1406),
    .S(net4276),
    .X(_01733_));
 sg13g2_mux2_1 _33570_ (.A0(net2056),
    .A1(net1726),
    .S(net4276),
    .X(_01734_));
 sg13g2_mux2_1 _33571_ (.A0(net2173),
    .A1(net1498),
    .S(net4276),
    .X(_01735_));
 sg13g2_mux2_1 _33572_ (.A0(net2461),
    .A1(net1727),
    .S(net4276),
    .X(_01736_));
 sg13g2_mux2_1 _33573_ (.A0(net1898),
    .A1(net1304),
    .S(net4275),
    .X(_01737_));
 sg13g2_mux2_1 _33574_ (.A0(net1995),
    .A1(net1503),
    .S(net4274),
    .X(_01738_));
 sg13g2_mux2_1 _33575_ (.A0(net2368),
    .A1(net1272),
    .S(net4275),
    .X(_01739_));
 sg13g2_mux2_1 _33576_ (.A0(net2006),
    .A1(net1809),
    .S(net4275),
    .X(_01740_));
 sg13g2_mux2_1 _33577_ (.A0(net2023),
    .A1(net1675),
    .S(net4273),
    .X(_01741_));
 sg13g2_mux2_1 _33578_ (.A0(net1953),
    .A1(net1616),
    .S(net4273),
    .X(_01742_));
 sg13g2_mux2_1 _33579_ (.A0(net2076),
    .A1(net1422),
    .S(net4273),
    .X(_01743_));
 sg13g2_mux2_1 _33580_ (.A0(net2651),
    .A1(net1596),
    .S(net4273),
    .X(_01744_));
 sg13g2_mux2_1 _33581_ (.A0(net2189),
    .A1(net1167),
    .S(net4273),
    .X(_01745_));
 sg13g2_mux2_1 _33582_ (.A0(net1891),
    .A1(\shift_reg[184] ),
    .S(net4273),
    .X(_01746_));
 sg13g2_mux2_1 _33583_ (.A0(net1790),
    .A1(\shift_reg[185] ),
    .S(net4273),
    .X(_01747_));
 sg13g2_mux2_1 _33584_ (.A0(net1930),
    .A1(net1687),
    .S(net4271),
    .X(_01748_));
 sg13g2_mux2_1 _33585_ (.A0(net1716),
    .A1(net1714),
    .S(net4271),
    .X(_01749_));
 sg13g2_mux2_1 _33586_ (.A0(net1868),
    .A1(net1513),
    .S(net4272),
    .X(_01750_));
 sg13g2_mux2_1 _33587_ (.A0(net1844),
    .A1(net1841),
    .S(net4272),
    .X(_01751_));
 sg13g2_mux2_1 _33588_ (.A0(net1982),
    .A1(net1843),
    .S(net4272),
    .X(_01752_));
 sg13g2_mux2_1 _33589_ (.A0(net2121),
    .A1(net1345),
    .S(net4269),
    .X(_01753_));
 sg13g2_mux2_1 _33590_ (.A0(net2238),
    .A1(net1659),
    .S(net4263),
    .X(_01754_));
 sg13g2_mux2_1 _33591_ (.A0(net2305),
    .A1(net1280),
    .S(net4263),
    .X(_01755_));
 sg13g2_mux2_1 _33592_ (.A0(net2462),
    .A1(net1398),
    .S(net4265),
    .X(_01756_));
 sg13g2_mux2_1 _33593_ (.A0(net2201),
    .A1(net1763),
    .S(net4260),
    .X(_01757_));
 sg13g2_mux2_1 _33594_ (.A0(net1990),
    .A1(net1854),
    .S(net4263),
    .X(_01758_));
 sg13g2_mux2_1 _33595_ (.A0(net1833),
    .A1(\shift_reg[197] ),
    .S(net4261),
    .X(_01759_));
 sg13g2_mux2_1 _33596_ (.A0(net1839),
    .A1(\shift_reg[198] ),
    .S(net4261),
    .X(_01760_));
 sg13g2_mux2_1 _33597_ (.A0(net1915),
    .A1(\shift_reg[199] ),
    .S(net4261),
    .X(_01761_));
 sg13g2_mux2_1 _33598_ (.A0(net1913),
    .A1(net1808),
    .S(net4260),
    .X(_01762_));
 sg13g2_mux2_1 _33599_ (.A0(net1810),
    .A1(net1567),
    .S(net4260),
    .X(_01763_));
 sg13g2_mux2_1 _33600_ (.A0(net2041),
    .A1(net1357),
    .S(net4260),
    .X(_01764_));
 sg13g2_mux2_1 _33601_ (.A0(net1987),
    .A1(net1200),
    .S(net4260),
    .X(_01765_));
 sg13g2_mux2_1 _33602_ (.A0(net1911),
    .A1(net1315),
    .S(net4260),
    .X(_01766_));
 sg13g2_mux2_1 _33603_ (.A0(net1943),
    .A1(net1424),
    .S(net4260),
    .X(_01767_));
 sg13g2_mux2_1 _33604_ (.A0(net1781),
    .A1(\shift_reg[206] ),
    .S(net4260),
    .X(_01768_));
 sg13g2_mux2_1 _33605_ (.A0(net1823),
    .A1(net1323),
    .S(net4255),
    .X(_01769_));
 sg13g2_mux2_1 _33606_ (.A0(net2053),
    .A1(net1371),
    .S(net4255),
    .X(_01770_));
 sg13g2_mux2_1 _33607_ (.A0(net1797),
    .A1(net1164),
    .S(net4254),
    .X(_01771_));
 sg13g2_mux2_1 _33608_ (.A0(net1866),
    .A1(net1557),
    .S(net4254),
    .X(_01772_));
 sg13g2_mux2_1 _33609_ (.A0(net1966),
    .A1(net1494),
    .S(net4255),
    .X(_01773_));
 sg13g2_mux2_1 _33610_ (.A0(net2128),
    .A1(net1618),
    .S(net4255),
    .X(_01774_));
 sg13g2_mux2_1 _33611_ (.A0(net2220),
    .A1(net1182),
    .S(net4258),
    .X(_01775_));
 sg13g2_mux2_1 _33612_ (.A0(net2131),
    .A1(net1306),
    .S(net4255),
    .X(_01776_));
 sg13g2_mux2_1 _33613_ (.A0(net1796),
    .A1(net1136),
    .S(net4254),
    .X(_01777_));
 sg13g2_mux2_1 _33614_ (.A0(net2040),
    .A1(net1125),
    .S(net4254),
    .X(_01778_));
 sg13g2_mux2_1 _33615_ (.A0(net1988),
    .A1(net1443),
    .S(net4254),
    .X(_01779_));
 sg13g2_mux2_1 _33616_ (.A0(net1824),
    .A1(net1642),
    .S(net4254),
    .X(_01780_));
 sg13g2_mux2_1 _33617_ (.A0(net1792),
    .A1(net1587),
    .S(net4254),
    .X(_01781_));
 sg13g2_mux2_1 _33618_ (.A0(net1807),
    .A1(net1730),
    .S(net4254),
    .X(_01782_));
 sg13g2_mux2_1 _33619_ (.A0(net2081),
    .A1(\shift_reg[221] ),
    .S(net4253),
    .X(_01783_));
 sg13g2_mux2_1 _33620_ (.A0(net1825),
    .A1(net1602),
    .S(net4250),
    .X(_01784_));
 sg13g2_mux2_1 _33621_ (.A0(net2113),
    .A1(net1090),
    .S(net4250),
    .X(_01785_));
 sg13g2_mux2_1 _33622_ (.A0(net1835),
    .A1(\shift_reg[224] ),
    .S(net4250),
    .X(_01786_));
 sg13g2_mux2_1 _33623_ (.A0(net1884),
    .A1(net1544),
    .S(net4250),
    .X(_01787_));
 sg13g2_mux2_1 _33624_ (.A0(net2093),
    .A1(net1927),
    .S(net4250),
    .X(_01788_));
 sg13g2_mux2_1 _33625_ (.A0(net2494),
    .A1(net1146),
    .S(net4248),
    .X(_01789_));
 sg13g2_mux2_1 _33626_ (.A0(net1742),
    .A1(net1685),
    .S(net4249),
    .X(_01790_));
 sg13g2_mux2_1 _33627_ (.A0(net2294),
    .A1(net1192),
    .S(net4249),
    .X(_01791_));
 sg13g2_mux2_1 _33628_ (.A0(net2448),
    .A1(net1202),
    .S(net4249),
    .X(_01792_));
 sg13g2_mux2_1 _33629_ (.A0(net2327),
    .A1(net1512),
    .S(net4248),
    .X(_01793_));
 sg13g2_mux2_1 _33630_ (.A0(net2185),
    .A1(net1188),
    .S(net4249),
    .X(_01794_));
 sg13g2_mux2_1 _33631_ (.A0(net1897),
    .A1(net1319),
    .S(net4248),
    .X(_01795_));
 sg13g2_mux2_1 _33632_ (.A0(net1973),
    .A1(net1129),
    .S(net4248),
    .X(_01796_));
 sg13g2_mux2_1 _33633_ (.A0(net2096),
    .A1(net1340),
    .S(net4248),
    .X(_01797_));
 sg13g2_mux2_1 _33634_ (.A0(net1828),
    .A1(net1194),
    .S(net4248),
    .X(_01798_));
 sg13g2_mux2_1 _33635_ (.A0(net2160),
    .A1(net1118),
    .S(net4248),
    .X(_01799_));
 sg13g2_mux2_1 _33636_ (.A0(net1732),
    .A1(net1302),
    .S(net4248),
    .X(_01800_));
 sg13g2_mux2_1 _33637_ (.A0(net2205),
    .A1(net1105),
    .S(net4247),
    .X(_01801_));
 sg13g2_mux2_1 _33638_ (.A0(net2004),
    .A1(\shift_reg[240] ),
    .S(net4242),
    .X(_01802_));
 sg13g2_mux2_1 _33639_ (.A0(net2126),
    .A1(net1138),
    .S(net4242),
    .X(_01803_));
 sg13g2_mux2_1 _33640_ (.A0(net1849),
    .A1(net1549),
    .S(net4242),
    .X(_01804_));
 sg13g2_mux2_1 _33641_ (.A0(net1932),
    .A1(\shift_reg[243] ),
    .S(net4242),
    .X(_01805_));
 sg13g2_mux2_1 _33642_ (.A0(net1788),
    .A1(\shift_reg[244] ),
    .S(net4242),
    .X(_01806_));
 sg13g2_mux2_1 _33643_ (.A0(net1852),
    .A1(net1639),
    .S(net4242),
    .X(_01807_));
 sg13g2_mux2_1 _33644_ (.A0(net1783),
    .A1(net1564),
    .S(net4242),
    .X(_01808_));
 sg13g2_mux2_1 _33645_ (.A0(net1965),
    .A1(net1706),
    .S(net4242),
    .X(_01809_));
 sg13g2_mux2_1 _33646_ (.A0(net2180),
    .A1(net1127),
    .S(net4246),
    .X(_01810_));
 sg13g2_mux2_1 _33647_ (.A0(net1946),
    .A1(net1097),
    .S(net4246),
    .X(_01811_));
 sg13g2_mux2_1 _33648_ (.A0(net1723),
    .A1(net1086),
    .S(net4246),
    .X(_01812_));
 sg13g2_mux2_1 _33649_ (.A0(net1756),
    .A1(net1115),
    .S(net4246),
    .X(_01813_));
 sg13g2_mux2_1 _33650_ (.A0(net1948),
    .A1(net1153),
    .S(net4246),
    .X(_01814_));
 sg13g2_mux2_1 _33651_ (.A0(net1952),
    .A1(net1121),
    .S(net4246),
    .X(_01815_));
 sg13g2_mux2_1 _33652_ (.A0(net2010),
    .A1(net1099),
    .S(net4246),
    .X(_01816_));
 sg13g2_mux2_1 _33653_ (.A0(net2037),
    .A1(net1109),
    .S(net4246),
    .X(_01817_));
 sg13g2_nor2_1 _33654_ (.A(net1599),
    .B(net4039),
    .Y(_10286_));
 sg13g2_a21oi_1 _33655_ (.A1(net1599),
    .A2(net3907),
    .Y(_01818_),
    .B1(_10286_));
 sg13g2_and2_1 _33656_ (.A(net1599),
    .B(net1603),
    .X(_10287_));
 sg13g2_a21o_1 _33657_ (.A2(_10287_),
    .A1(_12214_),
    .B1(net4446),
    .X(_10288_));
 sg13g2_nand3_1 _33658_ (.B(_12214_),
    .C(net3908),
    .A(net1599),
    .Y(_10289_));
 sg13g2_a22oi_1 _33659_ (.Y(_01819_),
    .B1(_10289_),
    .B2(_10628_),
    .A2(_10288_),
    .A1(net4039));
 sg13g2_o21ai_1 _33660_ (.B1(net1603),
    .Y(_10290_),
    .A1(net1599),
    .A2(_12220_));
 sg13g2_xnor2_1 _33661_ (.Y(_10291_),
    .A(net2841),
    .B(_10290_));
 sg13g2_a22oi_1 _33662_ (.Y(_10292_),
    .B1(net3908),
    .B2(_10291_),
    .A2(net3986),
    .A1(net2841));
 sg13g2_inv_1 _33663_ (.Y(_01820_),
    .A(_10292_));
 sg13g2_a21oi_1 _33664_ (.A1(\u_inv.delta_reg[2] ),
    .A2(_10287_),
    .Y(_10293_),
    .B1(net2467));
 sg13g2_nand3_1 _33665_ (.B(\u_inv.delta_reg[2] ),
    .C(_10287_),
    .A(\u_inv.delta_reg[3] ),
    .Y(_10294_));
 sg13g2_nand2_1 _33666_ (.Y(_10295_),
    .A(net3865),
    .B(_10294_));
 sg13g2_o21ai_1 _33667_ (.B1(net2467),
    .Y(_10296_),
    .A1(net1603),
    .A2(\u_inv.delta_reg[2] ));
 sg13g2_nand3_1 _33668_ (.B(net3819),
    .C(_10296_),
    .A(_12215_),
    .Y(_10297_));
 sg13g2_o21ai_1 _33669_ (.B1(_10297_),
    .Y(_10298_),
    .A1(_10293_),
    .A2(_10295_));
 sg13g2_a22oi_1 _33670_ (.Y(_10299_),
    .B1(net3907),
    .B2(_10298_),
    .A2(net3986),
    .A1(net2467));
 sg13g2_inv_1 _33671_ (.Y(_01821_),
    .A(net2468));
 sg13g2_nand2_1 _33672_ (.Y(_10300_),
    .A(_12215_),
    .B(_10295_));
 sg13g2_xnor2_1 _33673_ (.Y(_10301_),
    .A(net2600),
    .B(_10300_));
 sg13g2_a22oi_1 _33674_ (.Y(_10302_),
    .B1(net3907),
    .B2(_10301_),
    .A2(net3986),
    .A1(net2600));
 sg13g2_inv_1 _33675_ (.Y(_01822_),
    .A(_10302_));
 sg13g2_nor2_1 _33676_ (.A(_10629_),
    .B(_10294_),
    .Y(_10303_));
 sg13g2_a21oi_1 _33677_ (.A1(_12216_),
    .A2(net3818),
    .Y(_10304_),
    .B1(_10303_));
 sg13g2_xnor2_1 _33678_ (.Y(_10305_),
    .A(net2953),
    .B(_10304_));
 sg13g2_a22oi_1 _33679_ (.Y(_10306_),
    .B1(net3908),
    .B2(_10305_),
    .A2(net3987),
    .A1(net2953));
 sg13g2_inv_1 _33680_ (.Y(_01823_),
    .A(net2954));
 sg13g2_nand2_1 _33681_ (.Y(_10307_),
    .A(net1521),
    .B(net3987));
 sg13g2_o21ai_1 _33682_ (.B1(net1521),
    .Y(_10308_),
    .A1(\u_inv.delta_reg[5] ),
    .A2(_12216_));
 sg13g2_nor2_1 _33683_ (.A(_12214_),
    .B(_12217_),
    .Y(_10309_));
 sg13g2_a21oi_1 _33684_ (.A1(\u_inv.delta_reg[5] ),
    .A2(_10303_),
    .Y(_10310_),
    .B1(net1521));
 sg13g2_nand3_1 _33685_ (.B(net1521),
    .C(_10303_),
    .A(\u_inv.delta_reg[5] ),
    .Y(_10311_));
 sg13g2_nor2b_1 _33686_ (.A(_10310_),
    .B_N(_10311_),
    .Y(_10312_));
 sg13g2_a22oi_1 _33687_ (.Y(_10313_),
    .B1(_10312_),
    .B2(net3866),
    .A2(_10309_),
    .A1(_10308_));
 sg13g2_o21ai_1 _33688_ (.B1(_10307_),
    .Y(_01824_),
    .A1(net4239),
    .A2(_10313_));
 sg13g2_nand2b_1 _33689_ (.Y(_10314_),
    .B(_10311_),
    .A_N(_10309_));
 sg13g2_xnor2_1 _33690_ (.Y(_10315_),
    .A(_10630_),
    .B(_10314_));
 sg13g2_a22oi_1 _33691_ (.Y(_10316_),
    .B1(net3907),
    .B2(_10315_),
    .A2(net3987),
    .A1(net1680));
 sg13g2_inv_1 _33692_ (.Y(_01825_),
    .A(net1681));
 sg13g2_nand2_1 _33693_ (.Y(_10317_),
    .A(net1873),
    .B(net3987));
 sg13g2_nand2_1 _33694_ (.Y(_10318_),
    .A(net1873),
    .B(_12218_));
 sg13g2_nor2_1 _33695_ (.A(_10630_),
    .B(_10311_),
    .Y(_10319_));
 sg13g2_and2_1 _33696_ (.A(net1873),
    .B(_10319_),
    .X(_10320_));
 sg13g2_xor2_1 _33697_ (.B(_10319_),
    .A(net1873),
    .X(_10321_));
 sg13g2_a22oi_1 _33698_ (.Y(_10322_),
    .B1(_10321_),
    .B2(net3866),
    .A2(_10318_),
    .A1(_12220_));
 sg13g2_o21ai_1 _33699_ (.B1(_10317_),
    .Y(_01826_),
    .A1(net4239),
    .A2(_10322_));
 sg13g2_o21ai_1 _33700_ (.B1(net3866),
    .Y(_10323_),
    .A1(net3160),
    .A2(_10320_));
 sg13g2_a21oi_1 _33701_ (.A1(net3160),
    .A2(_10320_),
    .Y(_10324_),
    .B1(_10323_));
 sg13g2_o21ai_1 _33702_ (.B1(net3907),
    .Y(_10325_),
    .A1(_12220_),
    .A2(_10324_));
 sg13g2_o21ai_1 _33703_ (.B1(_10325_),
    .Y(_01827_),
    .A1(_10631_),
    .A2(net4039));
 sg13g2_dfrbpq_1 _33704_ (.RESET_B(net4815),
    .D(net1064),
    .Q(\u_inv.input_valid ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _33705_ (.RESET_B(net4815),
    .D(_00003_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _33706_ (.RESET_B(net4815),
    .D(_00004_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _33707_ (.RESET_B(net4824),
    .D(net1070),
    .Q(\byte_cnt[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33708_ (.RESET_B(net4824),
    .D(net1296),
    .Q(\byte_cnt[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33709_ (.RESET_B(net4824),
    .D(net2012),
    .Q(\byte_cnt[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _33710_ (.RESET_B(net4825),
    .D(net1104),
    .Q(\byte_cnt[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33711_ (.RESET_B(net4825),
    .D(_00009_),
    .Q(\byte_cnt[4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33712_ (.RESET_B(net4815),
    .D(net1217),
    .Q(inv_go),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _33713_ (.RESET_B(net4815),
    .D(net9),
    .Q(wr_prev),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33714_ (.RESET_B(net4815),
    .D(net10),
    .Q(rd_prev),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _33715_ (.RESET_B(net397),
    .D(_00010_),
    .Q(\u_inv.f_next[256] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _33716_ (.RESET_B(net4818),
    .D(_00011_),
    .Q(\shift_reg[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _33717_ (.RESET_B(net4820),
    .D(net1370),
    .Q(\shift_reg[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _33718_ (.RESET_B(net4820),
    .D(_00013_),
    .Q(\shift_reg[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _33719_ (.RESET_B(net4820),
    .D(net1830),
    .Q(\shift_reg[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _33720_ (.RESET_B(net4824),
    .D(net1170),
    .Q(\shift_reg[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _33721_ (.RESET_B(net4824),
    .D(net1348),
    .Q(\shift_reg[5] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _33722_ (.RESET_B(net4822),
    .D(_00017_),
    .Q(\shift_reg[6] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _33723_ (.RESET_B(net4822),
    .D(_00018_),
    .Q(\shift_reg[7] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _33724_ (.RESET_B(net4822),
    .D(net1447),
    .Q(\shift_reg[8] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _33725_ (.RESET_B(net4821),
    .D(net1250),
    .Q(\shift_reg[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _33726_ (.RESET_B(net4822),
    .D(net1594),
    .Q(\shift_reg[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _33727_ (.RESET_B(net4820),
    .D(net1242),
    .Q(\shift_reg[11] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _33728_ (.RESET_B(net4836),
    .D(net1213),
    .Q(\shift_reg[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _33729_ (.RESET_B(net4837),
    .D(net1144),
    .Q(\shift_reg[13] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _33730_ (.RESET_B(net4823),
    .D(_00025_),
    .Q(\shift_reg[14] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _33731_ (.RESET_B(net4836),
    .D(_00026_),
    .Q(\shift_reg[15] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _33732_ (.RESET_B(net4822),
    .D(_00027_),
    .Q(\shift_reg[16] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _33733_ (.RESET_B(net4822),
    .D(net2039),
    .Q(\shift_reg[17] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _33734_ (.RESET_B(net4836),
    .D(_00029_),
    .Q(\shift_reg[18] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _33735_ (.RESET_B(net4836),
    .D(_00030_),
    .Q(\shift_reg[19] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _33736_ (.RESET_B(net4838),
    .D(_00031_),
    .Q(\shift_reg[20] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _33737_ (.RESET_B(net4838),
    .D(net1252),
    .Q(\shift_reg[21] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _33738_ (.RESET_B(net4838),
    .D(net1360),
    .Q(\shift_reg[22] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _33739_ (.RESET_B(net4838),
    .D(net1488),
    .Q(\shift_reg[23] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _33740_ (.RESET_B(net4839),
    .D(net1634),
    .Q(\shift_reg[24] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _33741_ (.RESET_B(net4839),
    .D(net1231),
    .Q(\shift_reg[25] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _33742_ (.RESET_B(net4839),
    .D(net1211),
    .Q(\shift_reg[26] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _33743_ (.RESET_B(net4839),
    .D(net1585),
    .Q(\shift_reg[27] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33744_ (.RESET_B(net4839),
    .D(net1161),
    .Q(\shift_reg[28] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _33745_ (.RESET_B(net4841),
    .D(net1462),
    .Q(\shift_reg[29] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33746_ (.RESET_B(net4854),
    .D(net1156),
    .Q(\shift_reg[30] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33747_ (.RESET_B(net4854),
    .D(net1149),
    .Q(\shift_reg[31] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33748_ (.RESET_B(net4851),
    .D(net1385),
    .Q(\shift_reg[32] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33749_ (.RESET_B(net4854),
    .D(net1133),
    .Q(\shift_reg[33] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33750_ (.RESET_B(net4851),
    .D(net1389),
    .Q(\shift_reg[34] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _33751_ (.RESET_B(net4853),
    .D(net1163),
    .Q(\shift_reg[35] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _33752_ (.RESET_B(net4853),
    .D(net1430),
    .Q(\shift_reg[36] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _33753_ (.RESET_B(net4853),
    .D(net1356),
    .Q(\shift_reg[37] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _33754_ (.RESET_B(net4851),
    .D(net1262),
    .Q(\shift_reg[38] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _33755_ (.RESET_B(net4851),
    .D(net1480),
    .Q(\shift_reg[39] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _33756_ (.RESET_B(net4856),
    .D(net1337),
    .Q(\shift_reg[40] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _33757_ (.RESET_B(net4856),
    .D(net1311),
    .Q(\shift_reg[41] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _33758_ (.RESET_B(net4857),
    .D(net1275),
    .Q(\shift_reg[42] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _33759_ (.RESET_B(net4856),
    .D(_00054_),
    .Q(\shift_reg[43] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _33760_ (.RESET_B(net4857),
    .D(net1152),
    .Q(\shift_reg[44] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _33761_ (.RESET_B(net4856),
    .D(_00056_),
    .Q(\shift_reg[45] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _33762_ (.RESET_B(net4857),
    .D(_00057_),
    .Q(\shift_reg[46] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _33763_ (.RESET_B(net4857),
    .D(net1712),
    .Q(\shift_reg[47] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _33764_ (.RESET_B(net4862),
    .D(_00059_),
    .Q(\shift_reg[48] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _33765_ (.RESET_B(net4870),
    .D(net1421),
    .Q(\shift_reg[49] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _33766_ (.RESET_B(net4870),
    .D(net1199),
    .Q(\shift_reg[50] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _33767_ (.RESET_B(net4871),
    .D(net1124),
    .Q(\shift_reg[51] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _33768_ (.RESET_B(net4874),
    .D(_00063_),
    .Q(\shift_reg[52] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _33769_ (.RESET_B(net4870),
    .D(net1542),
    .Q(\shift_reg[53] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _33770_ (.RESET_B(net4872),
    .D(net1285),
    .Q(\shift_reg[54] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _33771_ (.RESET_B(net4876),
    .D(net1233),
    .Q(\shift_reg[55] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _33772_ (.RESET_B(net4872),
    .D(net1351),
    .Q(\shift_reg[56] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _33773_ (.RESET_B(net4873),
    .D(_00068_),
    .Q(\shift_reg[57] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _33774_ (.RESET_B(net4873),
    .D(net1573),
    .Q(\shift_reg[58] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _33775_ (.RESET_B(net4875),
    .D(_00070_),
    .Q(\shift_reg[59] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _33776_ (.RESET_B(net4873),
    .D(net1590),
    .Q(\shift_reg[60] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _33777_ (.RESET_B(net4873),
    .D(_00072_),
    .Q(\shift_reg[61] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _33778_ (.RESET_B(net4872),
    .D(_00073_),
    .Q(\shift_reg[62] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _33779_ (.RESET_B(net4872),
    .D(net1520),
    .Q(\shift_reg[63] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _33780_ (.RESET_B(net4884),
    .D(_00075_),
    .Q(\shift_reg[64] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _33781_ (.RESET_B(net4884),
    .D(net1474),
    .Q(\shift_reg[65] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _33782_ (.RESET_B(net4885),
    .D(net1486),
    .Q(\shift_reg[66] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _33783_ (.RESET_B(net4888),
    .D(net1387),
    .Q(\shift_reg[67] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _33784_ (.RESET_B(net4884),
    .D(net1287),
    .Q(\shift_reg[68] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _33785_ (.RESET_B(net4884),
    .D(net1158),
    .Q(\shift_reg[69] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33786_ (.RESET_B(net4886),
    .D(_00081_),
    .Q(\shift_reg[70] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _33787_ (.RESET_B(net4885),
    .D(net1258),
    .Q(\shift_reg[71] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _33788_ (.RESET_B(net4886),
    .D(net1209),
    .Q(\shift_reg[72] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _33789_ (.RESET_B(net4886),
    .D(net1571),
    .Q(\shift_reg[73] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _33790_ (.RESET_B(net4893),
    .D(net1239),
    .Q(\shift_reg[74] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _33791_ (.RESET_B(net4889),
    .D(net1403),
    .Q(\shift_reg[75] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _33792_ (.RESET_B(net4886),
    .D(net1460),
    .Q(\shift_reg[76] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33793_ (.RESET_B(net4889),
    .D(net1478),
    .Q(\shift_reg[77] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _33794_ (.RESET_B(net4886),
    .D(net1381),
    .Q(\shift_reg[78] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _33795_ (.RESET_B(net4889),
    .D(net1318),
    .Q(\shift_reg[79] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _33796_ (.RESET_B(net4889),
    .D(_00091_),
    .Q(\shift_reg[80] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _33797_ (.RESET_B(net4890),
    .D(net1283),
    .Q(\shift_reg[81] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _33798_ (.RESET_B(net4892),
    .D(net1466),
    .Q(\shift_reg[82] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _33799_ (.RESET_B(net4891),
    .D(net1344),
    .Q(\shift_reg[83] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _33800_ (.RESET_B(net4891),
    .D(net1472),
    .Q(\shift_reg[84] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33801_ (.RESET_B(net4890),
    .D(net1254),
    .Q(\shift_reg[85] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33802_ (.RESET_B(net4891),
    .D(_00097_),
    .Q(\shift_reg[86] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33803_ (.RESET_B(net4891),
    .D(net1248),
    .Q(\shift_reg[87] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _33804_ (.RESET_B(net4896),
    .D(net1292),
    .Q(\shift_reg[88] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _33805_ (.RESET_B(net4896),
    .D(net1329),
    .Q(\shift_reg[89] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _33806_ (.RESET_B(net4898),
    .D(net1379),
    .Q(\shift_reg[90] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _33807_ (.RESET_B(net4896),
    .D(_00102_),
    .Q(\shift_reg[91] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _33808_ (.RESET_B(net4891),
    .D(net1482),
    .Q(\shift_reg[92] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _33809_ (.RESET_B(net4896),
    .D(net1205),
    .Q(\shift_reg[93] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _33810_ (.RESET_B(net4896),
    .D(net1331),
    .Q(\shift_reg[94] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _33811_ (.RESET_B(net4897),
    .D(_00106_),
    .Q(\shift_reg[95] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _33812_ (.RESET_B(net4899),
    .D(_00107_),
    .Q(\shift_reg[96] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _33813_ (.RESET_B(net4900),
    .D(net1362),
    .Q(\shift_reg[97] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _33814_ (.RESET_B(net4899),
    .D(_00109_),
    .Q(\shift_reg[98] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _33815_ (.RESET_B(net4900),
    .D(net1470),
    .Q(\shift_reg[99] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33816_ (.RESET_B(net4900),
    .D(_00111_),
    .Q(\shift_reg[100] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33817_ (.RESET_B(net4899),
    .D(_00112_),
    .Q(\shift_reg[101] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _33818_ (.RESET_B(net4900),
    .D(_00113_),
    .Q(\shift_reg[102] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _33819_ (.RESET_B(net4899),
    .D(_00114_),
    .Q(\shift_reg[103] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _33820_ (.RESET_B(net4901),
    .D(_00115_),
    .Q(\shift_reg[104] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _33821_ (.RESET_B(net4914),
    .D(net1174),
    .Q(\shift_reg[105] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _33822_ (.RESET_B(net4910),
    .D(net1397),
    .Q(\shift_reg[106] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _33823_ (.RESET_B(net4914),
    .D(net1405),
    .Q(\shift_reg[107] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _33824_ (.RESET_B(net4917),
    .D(net1197),
    .Q(\shift_reg[108] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _33825_ (.RESET_B(net4915),
    .D(net1865),
    .Q(\shift_reg[109] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _33826_ (.RESET_B(net4910),
    .D(net1777),
    .Q(\shift_reg[110] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _33827_ (.RESET_B(net4904),
    .D(net2162),
    .Q(\shift_reg[111] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _33828_ (.RESET_B(net4919),
    .D(net1354),
    .Q(\shift_reg[112] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _33829_ (.RESET_B(net4942),
    .D(net1630),
    .Q(\shift_reg[113] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _33830_ (.RESET_B(net4916),
    .D(net1108),
    .Q(\shift_reg[114] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _33831_ (.RESET_B(net4915),
    .D(_00126_),
    .Q(\shift_reg[115] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _33832_ (.RESET_B(net4942),
    .D(_00127_),
    .Q(\shift_reg[116] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _33833_ (.RESET_B(net4945),
    .D(net1260),
    .Q(\shift_reg[117] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _33834_ (.RESET_B(net4916),
    .D(_00129_),
    .Q(\shift_reg[118] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33835_ (.RESET_B(net4939),
    .D(net1775),
    .Q(\shift_reg[119] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33836_ (.RESET_B(net4942),
    .D(net1890),
    .Q(\shift_reg[120] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _33837_ (.RESET_B(net4943),
    .D(net1501),
    .Q(\shift_reg[121] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _33838_ (.RESET_B(net4945),
    .D(net1418),
    .Q(\shift_reg[122] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _33839_ (.RESET_B(net4943),
    .D(net1699),
    .Q(\shift_reg[123] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _33840_ (.RESET_B(net4946),
    .D(net1181),
    .Q(\shift_reg[124] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _33841_ (.RESET_B(net4946),
    .D(_00136_),
    .Q(\shift_reg[125] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _33842_ (.RESET_B(net4941),
    .D(net1531),
    .Q(\shift_reg[126] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _33843_ (.RESET_B(net4946),
    .D(net1113),
    .Q(\shift_reg[127] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _33844_ (.RESET_B(net4925),
    .D(net1327),
    .Q(\shift_reg[128] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _33845_ (.RESET_B(net4933),
    .D(net1556),
    .Q(\shift_reg[129] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _33846_ (.RESET_B(net4933),
    .D(net1607),
    .Q(\shift_reg[130] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _33847_ (.RESET_B(net4933),
    .D(net1289),
    .Q(\shift_reg[131] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _33848_ (.RESET_B(net4928),
    .D(_00143_),
    .Q(\shift_reg[132] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _33849_ (.RESET_B(net4930),
    .D(net1266),
    .Q(\shift_reg[133] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _33850_ (.RESET_B(net4928),
    .D(net1415),
    .Q(\shift_reg[134] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _33851_ (.RESET_B(net4930),
    .D(net1395),
    .Q(\shift_reg[135] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _33852_ (.RESET_B(net4929),
    .D(net1222),
    .Q(\shift_reg[136] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _33853_ (.RESET_B(net4932),
    .D(_00148_),
    .Q(\shift_reg[137] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _33854_ (.RESET_B(net4930),
    .D(net1179),
    .Q(\shift_reg[138] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _33855_ (.RESET_B(net4929),
    .D(net1235),
    .Q(\shift_reg[139] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _33856_ (.RESET_B(net4928),
    .D(_00151_),
    .Q(\shift_reg[140] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _33857_ (.RESET_B(net4931),
    .D(_00152_),
    .Q(\shift_reg[141] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _33858_ (.RESET_B(net4929),
    .D(_00153_),
    .Q(\shift_reg[142] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _33859_ (.RESET_B(net4929),
    .D(net1649),
    .Q(\shift_reg[143] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _33860_ (.RESET_B(net4929),
    .D(net1537),
    .Q(\shift_reg[144] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _33861_ (.RESET_B(net4934),
    .D(net1490),
    .Q(\shift_reg[145] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _33862_ (.RESET_B(net4930),
    .D(_00157_),
    .Q(\shift_reg[146] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _33863_ (.RESET_B(net4933),
    .D(_00158_),
    .Q(\shift_reg[147] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _33864_ (.RESET_B(net4934),
    .D(_00159_),
    .Q(\shift_reg[148] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _33865_ (.RESET_B(net4933),
    .D(net1525),
    .Q(\shift_reg[149] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _33866_ (.RESET_B(net4924),
    .D(_00161_),
    .Q(\shift_reg[150] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _33867_ (.RESET_B(net4933),
    .D(net1601),
    .Q(\shift_reg[151] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _33868_ (.RESET_B(net4936),
    .D(_00163_),
    .Q(\shift_reg[152] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _33869_ (.RESET_B(net4934),
    .D(_00164_),
    .Q(\shift_reg[153] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _33870_ (.RESET_B(net4925),
    .D(net1658),
    .Q(\shift_reg[154] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _33871_ (.RESET_B(net4934),
    .D(net1645),
    .Q(\shift_reg[155] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _33872_ (.RESET_B(net4934),
    .D(_00167_),
    .Q(\shift_reg[156] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _33873_ (.RESET_B(net4946),
    .D(net1546),
    .Q(\shift_reg[157] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _33874_ (.RESET_B(net4940),
    .D(net1674),
    .Q(\shift_reg[158] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _33875_ (.RESET_B(net4946),
    .D(_00170_),
    .Q(\shift_reg[159] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _33876_ (.RESET_B(net4940),
    .D(net1277),
    .Q(\shift_reg[160] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _33877_ (.RESET_B(net4941),
    .D(net1366),
    .Q(\shift_reg[161] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _33878_ (.RESET_B(net4940),
    .D(net1313),
    .Q(\shift_reg[162] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33879_ (.RESET_B(net4941),
    .D(_00174_),
    .Q(\shift_reg[163] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _33880_ (.RESET_B(net4940),
    .D(net1244),
    .Q(\shift_reg[164] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _33881_ (.RESET_B(net4940),
    .D(net1652),
    .Q(\shift_reg[165] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33882_ (.RESET_B(net4940),
    .D(net1270),
    .Q(\shift_reg[166] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _33883_ (.RESET_B(net4938),
    .D(net1436),
    .Q(\shift_reg[167] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _33884_ (.RESET_B(net4938),
    .D(_00179_),
    .Q(\shift_reg[168] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _33885_ (.RESET_B(net4939),
    .D(net1442),
    .Q(\shift_reg[169] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _33886_ (.RESET_B(net4916),
    .D(_00181_),
    .Q(\shift_reg[170] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33887_ (.RESET_B(net4916),
    .D(net1407),
    .Q(\shift_reg[171] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _33888_ (.RESET_B(net4938),
    .D(_00183_),
    .Q(\shift_reg[172] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _33889_ (.RESET_B(net4917),
    .D(net1499),
    .Q(\shift_reg[173] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _33890_ (.RESET_B(net4916),
    .D(_00185_),
    .Q(\shift_reg[174] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _33891_ (.RESET_B(net4914),
    .D(net1305),
    .Q(\shift_reg[175] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _33892_ (.RESET_B(net4912),
    .D(net1504),
    .Q(\shift_reg[176] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _33893_ (.RESET_B(net4914),
    .D(net1273),
    .Q(\shift_reg[177] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _33894_ (.RESET_B(net4914),
    .D(_00189_),
    .Q(\shift_reg[178] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _33895_ (.RESET_B(net4912),
    .D(_00190_),
    .Q(\shift_reg[179] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _33896_ (.RESET_B(net4912),
    .D(net1617),
    .Q(\shift_reg[180] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _33897_ (.RESET_B(net4904),
    .D(net1423),
    .Q(\shift_reg[181] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _33898_ (.RESET_B(net4904),
    .D(net1597),
    .Q(\shift_reg[182] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _33899_ (.RESET_B(net4904),
    .D(net1168),
    .Q(\shift_reg[183] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _33900_ (.RESET_B(net4901),
    .D(_00195_),
    .Q(\shift_reg[184] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33901_ (.RESET_B(net4903),
    .D(_00196_),
    .Q(\shift_reg[185] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33902_ (.RESET_B(net4907),
    .D(net1688),
    .Q(\shift_reg[186] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33903_ (.RESET_B(net4901),
    .D(_00198_),
    .Q(\shift_reg[187] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _33904_ (.RESET_B(net4900),
    .D(net1514),
    .Q(\shift_reg[188] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _33905_ (.RESET_B(net4899),
    .D(_00200_),
    .Q(\shift_reg[189] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _33906_ (.RESET_B(net4898),
    .D(_00201_),
    .Q(\shift_reg[190] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _33907_ (.RESET_B(net4896),
    .D(net1346),
    .Q(\shift_reg[191] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _33908_ (.RESET_B(net4885),
    .D(net1660),
    .Q(\shift_reg[192] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _33909_ (.RESET_B(net4884),
    .D(net1281),
    .Q(\shift_reg[193] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _33910_ (.RESET_B(net4881),
    .D(net1399),
    .Q(\shift_reg[194] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _33911_ (.RESET_B(net4881),
    .D(_00206_),
    .Q(\shift_reg[195] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _33912_ (.RESET_B(net4879),
    .D(_00207_),
    .Q(\shift_reg[196] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _33913_ (.RESET_B(net4880),
    .D(net2058),
    .Q(\shift_reg[197] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _33914_ (.RESET_B(net4881),
    .D(_00209_),
    .Q(\shift_reg[198] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _33915_ (.RESET_B(net4887),
    .D(_00210_),
    .Q(\shift_reg[199] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _33916_ (.RESET_B(net4868),
    .D(_00211_),
    .Q(\shift_reg[200] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _33917_ (.RESET_B(net4867),
    .D(net1568),
    .Q(\shift_reg[201] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _33918_ (.RESET_B(net4866),
    .D(net1358),
    .Q(\shift_reg[202] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _33919_ (.RESET_B(net4867),
    .D(net1201),
    .Q(\shift_reg[203] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _33920_ (.RESET_B(net4864),
    .D(net1316),
    .Q(\shift_reg[204] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33921_ (.RESET_B(net4862),
    .D(net1425),
    .Q(\shift_reg[205] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _33922_ (.RESET_B(net4863),
    .D(net1806),
    .Q(\shift_reg[206] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33923_ (.RESET_B(net4861),
    .D(net1324),
    .Q(\shift_reg[207] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33924_ (.RESET_B(net4861),
    .D(net1372),
    .Q(\shift_reg[208] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _33925_ (.RESET_B(net4847),
    .D(net1165),
    .Q(\shift_reg[209] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _33926_ (.RESET_B(net4861),
    .D(_00221_),
    .Q(\shift_reg[210] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _33927_ (.RESET_B(net4864),
    .D(net1495),
    .Q(\shift_reg[211] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33928_ (.RESET_B(net4861),
    .D(_00223_),
    .Q(\shift_reg[212] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _33929_ (.RESET_B(net4861),
    .D(net1183),
    .Q(\shift_reg[213] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33930_ (.RESET_B(net4861),
    .D(net1307),
    .Q(\shift_reg[214] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _33931_ (.RESET_B(net4847),
    .D(net1137),
    .Q(\shift_reg[215] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _33932_ (.RESET_B(net4844),
    .D(net1126),
    .Q(\shift_reg[216] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _33933_ (.RESET_B(net4850),
    .D(_00228_),
    .Q(\shift_reg[217] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _33934_ (.RESET_B(net4850),
    .D(_00229_),
    .Q(\shift_reg[218] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _33935_ (.RESET_B(net4847),
    .D(net1588),
    .Q(\shift_reg[219] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _33936_ (.RESET_B(net4847),
    .D(_00231_),
    .Q(\shift_reg[220] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _33937_ (.RESET_B(net4847),
    .D(_00232_),
    .Q(\shift_reg[221] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _33938_ (.RESET_B(net4849),
    .D(_00233_),
    .Q(\shift_reg[222] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _33939_ (.RESET_B(net4832),
    .D(net1091),
    .Q(\shift_reg[223] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _33940_ (.RESET_B(net4846),
    .D(_00235_),
    .Q(\shift_reg[224] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _33941_ (.RESET_B(net4844),
    .D(_00236_),
    .Q(\shift_reg[225] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _33942_ (.RESET_B(net4845),
    .D(_00237_),
    .Q(\shift_reg[226] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _33943_ (.RESET_B(net4830),
    .D(net1147),
    .Q(\shift_reg[227] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _33944_ (.RESET_B(net4845),
    .D(net1686),
    .Q(\shift_reg[228] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _33945_ (.RESET_B(net4832),
    .D(net1193),
    .Q(\shift_reg[229] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _33946_ (.RESET_B(net4830),
    .D(net1203),
    .Q(\shift_reg[230] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _33947_ (.RESET_B(net4833),
    .D(_00242_),
    .Q(\shift_reg[231] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _33948_ (.RESET_B(net4830),
    .D(net1189),
    .Q(\shift_reg[232] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _33949_ (.RESET_B(net4830),
    .D(net1320),
    .Q(\shift_reg[233] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _33950_ (.RESET_B(net4830),
    .D(net1130),
    .Q(\shift_reg[234] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _33951_ (.RESET_B(net4830),
    .D(net1341),
    .Q(\shift_reg[235] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _33952_ (.RESET_B(net4829),
    .D(net1195),
    .Q(\shift_reg[236] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _33953_ (.RESET_B(net4831),
    .D(net1119),
    .Q(\shift_reg[237] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _33954_ (.RESET_B(net4829),
    .D(net1303),
    .Q(\shift_reg[238] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _33955_ (.RESET_B(net4809),
    .D(net1106),
    .Q(\shift_reg[239] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _33956_ (.RESET_B(net4827),
    .D(_00251_),
    .Q(\shift_reg[240] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _33957_ (.RESET_B(net4810),
    .D(net1139),
    .Q(\shift_reg[241] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _33958_ (.RESET_B(net4809),
    .D(net1550),
    .Q(\shift_reg[242] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _33959_ (.RESET_B(net4829),
    .D(_00254_),
    .Q(\shift_reg[243] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _33960_ (.RESET_B(net4827),
    .D(_00255_),
    .Q(\shift_reg[244] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _33961_ (.RESET_B(net4809),
    .D(net1640),
    .Q(\shift_reg[245] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _33962_ (.RESET_B(net4807),
    .D(net1565),
    .Q(\shift_reg[246] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _33963_ (.RESET_B(net4809),
    .D(net1707),
    .Q(\shift_reg[247] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _33964_ (.RESET_B(net4817),
    .D(net1128),
    .Q(\shift_reg[248] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _33965_ (.RESET_B(net4814),
    .D(net1098),
    .Q(\shift_reg[249] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _33966_ (.RESET_B(net4817),
    .D(net1087),
    .Q(\shift_reg[250] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _33967_ (.RESET_B(net4814),
    .D(net1116),
    .Q(\shift_reg[251] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _33968_ (.RESET_B(net4812),
    .D(net1154),
    .Q(\shift_reg[252] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _33969_ (.RESET_B(net4813),
    .D(net1122),
    .Q(\shift_reg[253] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _33970_ (.RESET_B(net4813),
    .D(net1100),
    .Q(\shift_reg[254] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _33971_ (.RESET_B(net4813),
    .D(net1110),
    .Q(\shift_reg[255] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _33972_ (.RESET_B(net4814),
    .D(net2222),
    .Q(inv_done),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _33973_ (.RESET_B(net4811),
    .D(_00267_),
    .Q(\u_inv.counter[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _33974_ (.RESET_B(net4812),
    .D(net1563),
    .Q(\u_inv.counter[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33975_ (.RESET_B(net4812),
    .D(net1632),
    .Q(\u_inv.counter[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33976_ (.RESET_B(net4812),
    .D(net1089),
    .Q(\u_inv.counter[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _33977_ (.RESET_B(net4811),
    .D(_00271_),
    .Q(\u_inv.counter[4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _33978_ (.RESET_B(net4811),
    .D(_00272_),
    .Q(\u_inv.counter[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _33979_ (.RESET_B(net4811),
    .D(_00273_),
    .Q(\u_inv.counter[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _33980_ (.RESET_B(net4811),
    .D(net1076),
    .Q(\u_inv.counter[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _33981_ (.RESET_B(net4811),
    .D(net1229),
    .Q(\u_inv.counter[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _33982_ (.RESET_B(net4811),
    .D(net1068),
    .Q(\u_inv.counter[9] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _33983_ (.RESET_B(net4814),
    .D(_17369_[0]),
    .Q(\u_inv.load_input ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _33984_ (.RESET_B(net396),
    .D(_00277_),
    .Q(\u_inv.d_next[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _33985_ (.RESET_B(net395),
    .D(_00278_),
    .Q(\u_inv.d_next[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _33986_ (.RESET_B(net394),
    .D(_00279_),
    .Q(\u_inv.d_next[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _33987_ (.RESET_B(net393),
    .D(_00280_),
    .Q(\u_inv.d_next[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _33988_ (.RESET_B(net392),
    .D(_00281_),
    .Q(\u_inv.d_next[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _33989_ (.RESET_B(net391),
    .D(_00282_),
    .Q(\u_inv.d_next[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _33990_ (.RESET_B(net390),
    .D(_00283_),
    .Q(\u_inv.d_next[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _33991_ (.RESET_B(net389),
    .D(_00284_),
    .Q(\u_inv.d_next[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _33992_ (.RESET_B(net388),
    .D(_00285_),
    .Q(\u_inv.d_next[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _33993_ (.RESET_B(net387),
    .D(_00286_),
    .Q(\u_inv.d_next[9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _33994_ (.RESET_B(net386),
    .D(_00287_),
    .Q(\u_inv.d_next[10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _33995_ (.RESET_B(net385),
    .D(_00288_),
    .Q(\u_inv.d_next[11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _33996_ (.RESET_B(net384),
    .D(_00289_),
    .Q(\u_inv.d_next[12] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _33997_ (.RESET_B(net383),
    .D(_00290_),
    .Q(\u_inv.d_next[13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _33998_ (.RESET_B(net382),
    .D(_00291_),
    .Q(\u_inv.d_next[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _33999_ (.RESET_B(net381),
    .D(_00292_),
    .Q(\u_inv.d_next[15] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _34000_ (.RESET_B(net380),
    .D(_00293_),
    .Q(\u_inv.d_next[16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _34001_ (.RESET_B(net379),
    .D(_00294_),
    .Q(\u_inv.d_next[17] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34002_ (.RESET_B(net378),
    .D(_00295_),
    .Q(\u_inv.d_next[18] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _34003_ (.RESET_B(net377),
    .D(_00296_),
    .Q(\u_inv.d_next[19] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _34004_ (.RESET_B(net376),
    .D(_00297_),
    .Q(\u_inv.d_next[20] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _34005_ (.RESET_B(net375),
    .D(_00298_),
    .Q(\u_inv.d_next[21] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _34006_ (.RESET_B(net374),
    .D(_00299_),
    .Q(\u_inv.d_next[22] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _34007_ (.RESET_B(net373),
    .D(_00300_),
    .Q(\u_inv.d_next[23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34008_ (.RESET_B(net372),
    .D(_00301_),
    .Q(\u_inv.d_next[24] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _34009_ (.RESET_B(net371),
    .D(_00302_),
    .Q(\u_inv.d_next[25] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34010_ (.RESET_B(net370),
    .D(_00303_),
    .Q(\u_inv.d_next[26] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34011_ (.RESET_B(net369),
    .D(_00304_),
    .Q(\u_inv.d_next[27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34012_ (.RESET_B(net368),
    .D(_00305_),
    .Q(\u_inv.d_next[28] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34013_ (.RESET_B(net367),
    .D(_00306_),
    .Q(\u_inv.d_next[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34014_ (.RESET_B(net366),
    .D(_00307_),
    .Q(\u_inv.d_next[30] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34015_ (.RESET_B(net365),
    .D(_00308_),
    .Q(\u_inv.d_next[31] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34016_ (.RESET_B(net364),
    .D(_00309_),
    .Q(\u_inv.d_next[32] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34017_ (.RESET_B(net363),
    .D(_00310_),
    .Q(\u_inv.d_next[33] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34018_ (.RESET_B(net362),
    .D(_00311_),
    .Q(\u_inv.d_next[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34019_ (.RESET_B(net361),
    .D(_00312_),
    .Q(\u_inv.d_next[35] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34020_ (.RESET_B(net360),
    .D(_00313_),
    .Q(\u_inv.d_next[36] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34021_ (.RESET_B(net359),
    .D(_00314_),
    .Q(\u_inv.d_next[37] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34022_ (.RESET_B(net358),
    .D(_00315_),
    .Q(\u_inv.d_next[38] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34023_ (.RESET_B(net357),
    .D(_00316_),
    .Q(\u_inv.d_next[39] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34024_ (.RESET_B(net356),
    .D(_00317_),
    .Q(\u_inv.d_next[40] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34025_ (.RESET_B(net355),
    .D(_00318_),
    .Q(\u_inv.d_next[41] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34026_ (.RESET_B(net354),
    .D(_00319_),
    .Q(\u_inv.d_next[42] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34027_ (.RESET_B(net353),
    .D(_00320_),
    .Q(\u_inv.d_next[43] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34028_ (.RESET_B(net352),
    .D(_00321_),
    .Q(\u_inv.d_next[44] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34029_ (.RESET_B(net351),
    .D(_00322_),
    .Q(\u_inv.d_next[45] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34030_ (.RESET_B(net350),
    .D(_00323_),
    .Q(\u_inv.d_next[46] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34031_ (.RESET_B(net349),
    .D(_00324_),
    .Q(\u_inv.d_next[47] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34032_ (.RESET_B(net348),
    .D(_00325_),
    .Q(\u_inv.d_next[48] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34033_ (.RESET_B(net347),
    .D(_00326_),
    .Q(\u_inv.d_next[49] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34034_ (.RESET_B(net346),
    .D(_00327_),
    .Q(\u_inv.d_next[50] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34035_ (.RESET_B(net345),
    .D(_00328_),
    .Q(\u_inv.d_next[51] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34036_ (.RESET_B(net344),
    .D(_00329_),
    .Q(\u_inv.d_next[52] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34037_ (.RESET_B(net343),
    .D(_00330_),
    .Q(\u_inv.d_next[53] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34038_ (.RESET_B(net342),
    .D(_00331_),
    .Q(\u_inv.d_next[54] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34039_ (.RESET_B(net341),
    .D(_00332_),
    .Q(\u_inv.d_next[55] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34040_ (.RESET_B(net340),
    .D(_00333_),
    .Q(\u_inv.d_next[56] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34041_ (.RESET_B(net339),
    .D(_00334_),
    .Q(\u_inv.d_next[57] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34042_ (.RESET_B(net338),
    .D(_00335_),
    .Q(\u_inv.d_next[58] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34043_ (.RESET_B(net337),
    .D(_00336_),
    .Q(\u_inv.d_next[59] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34044_ (.RESET_B(net336),
    .D(_00337_),
    .Q(\u_inv.d_next[60] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34045_ (.RESET_B(net335),
    .D(_00338_),
    .Q(\u_inv.d_next[61] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34046_ (.RESET_B(net334),
    .D(_00339_),
    .Q(\u_inv.d_next[62] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34047_ (.RESET_B(net333),
    .D(_00340_),
    .Q(\u_inv.d_next[63] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34048_ (.RESET_B(net332),
    .D(_00341_),
    .Q(\u_inv.d_next[64] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34049_ (.RESET_B(net331),
    .D(_00342_),
    .Q(\u_inv.d_next[65] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34050_ (.RESET_B(net330),
    .D(_00343_),
    .Q(\u_inv.d_next[66] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34051_ (.RESET_B(net329),
    .D(_00344_),
    .Q(\u_inv.d_next[67] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34052_ (.RESET_B(net328),
    .D(_00345_),
    .Q(\u_inv.d_next[68] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _34053_ (.RESET_B(net327),
    .D(_00346_),
    .Q(\u_inv.d_next[69] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34054_ (.RESET_B(net326),
    .D(_00347_),
    .Q(\u_inv.d_next[70] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34055_ (.RESET_B(net325),
    .D(_00348_),
    .Q(\u_inv.d_next[71] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34056_ (.RESET_B(net324),
    .D(_00349_),
    .Q(\u_inv.d_next[72] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34057_ (.RESET_B(net323),
    .D(_00350_),
    .Q(\u_inv.d_next[73] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34058_ (.RESET_B(net322),
    .D(_00351_),
    .Q(\u_inv.d_next[74] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34059_ (.RESET_B(net321),
    .D(_00352_),
    .Q(\u_inv.d_next[75] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34060_ (.RESET_B(net320),
    .D(_00353_),
    .Q(\u_inv.d_next[76] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34061_ (.RESET_B(net319),
    .D(_00354_),
    .Q(\u_inv.d_next[77] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34062_ (.RESET_B(net318),
    .D(_00355_),
    .Q(\u_inv.d_next[78] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34063_ (.RESET_B(net317),
    .D(_00356_),
    .Q(\u_inv.d_next[79] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34064_ (.RESET_B(net316),
    .D(_00357_),
    .Q(\u_inv.d_next[80] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34065_ (.RESET_B(net315),
    .D(_00358_),
    .Q(\u_inv.d_next[81] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34066_ (.RESET_B(net314),
    .D(_00359_),
    .Q(\u_inv.d_next[82] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34067_ (.RESET_B(net313),
    .D(_00360_),
    .Q(\u_inv.d_next[83] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34068_ (.RESET_B(net312),
    .D(_00361_),
    .Q(\u_inv.d_next[84] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34069_ (.RESET_B(net311),
    .D(_00362_),
    .Q(\u_inv.d_next[85] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34070_ (.RESET_B(net310),
    .D(_00363_),
    .Q(\u_inv.d_next[86] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34071_ (.RESET_B(net309),
    .D(_00364_),
    .Q(\u_inv.d_next[87] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34072_ (.RESET_B(net308),
    .D(_00365_),
    .Q(\u_inv.d_next[88] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34073_ (.RESET_B(net307),
    .D(_00366_),
    .Q(\u_inv.d_next[89] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34074_ (.RESET_B(net306),
    .D(_00367_),
    .Q(\u_inv.d_next[90] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34075_ (.RESET_B(net305),
    .D(_00368_),
    .Q(\u_inv.d_next[91] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34076_ (.RESET_B(net304),
    .D(_00369_),
    .Q(\u_inv.d_next[92] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34077_ (.RESET_B(net303),
    .D(_00370_),
    .Q(\u_inv.d_next[93] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34078_ (.RESET_B(net302),
    .D(_00371_),
    .Q(\u_inv.d_next[94] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34079_ (.RESET_B(net301),
    .D(_00372_),
    .Q(\u_inv.d_next[95] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34080_ (.RESET_B(net300),
    .D(_00373_),
    .Q(\u_inv.d_next[96] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34081_ (.RESET_B(net299),
    .D(_00374_),
    .Q(\u_inv.d_next[97] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34082_ (.RESET_B(net298),
    .D(_00375_),
    .Q(\u_inv.d_next[98] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34083_ (.RESET_B(net297),
    .D(_00376_),
    .Q(\u_inv.d_next[99] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34084_ (.RESET_B(net296),
    .D(_00377_),
    .Q(\u_inv.d_next[100] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34085_ (.RESET_B(net295),
    .D(_00378_),
    .Q(\u_inv.d_next[101] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _34086_ (.RESET_B(net294),
    .D(_00379_),
    .Q(\u_inv.d_next[102] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _34087_ (.RESET_B(net293),
    .D(_00380_),
    .Q(\u_inv.d_next[103] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _34088_ (.RESET_B(net292),
    .D(_00381_),
    .Q(\u_inv.d_next[104] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34089_ (.RESET_B(net291),
    .D(_00382_),
    .Q(\u_inv.d_next[105] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34090_ (.RESET_B(net290),
    .D(_00383_),
    .Q(\u_inv.d_next[106] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _34091_ (.RESET_B(net289),
    .D(_00384_),
    .Q(\u_inv.d_next[107] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34092_ (.RESET_B(net288),
    .D(_00385_),
    .Q(\u_inv.d_next[108] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34093_ (.RESET_B(net287),
    .D(_00386_),
    .Q(\u_inv.d_next[109] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34094_ (.RESET_B(net286),
    .D(_00387_),
    .Q(\u_inv.d_next[110] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34095_ (.RESET_B(net285),
    .D(_00388_),
    .Q(\u_inv.d_next[111] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34096_ (.RESET_B(net284),
    .D(_00389_),
    .Q(\u_inv.d_next[112] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34097_ (.RESET_B(net283),
    .D(_00390_),
    .Q(\u_inv.d_next[113] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34098_ (.RESET_B(net282),
    .D(_00391_),
    .Q(\u_inv.d_next[114] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34099_ (.RESET_B(net281),
    .D(_00392_),
    .Q(\u_inv.d_next[115] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34100_ (.RESET_B(net280),
    .D(_00393_),
    .Q(\u_inv.d_next[116] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34101_ (.RESET_B(net279),
    .D(_00394_),
    .Q(\u_inv.d_next[117] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34102_ (.RESET_B(net278),
    .D(_00395_),
    .Q(\u_inv.d_next[118] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34103_ (.RESET_B(net277),
    .D(_00396_),
    .Q(\u_inv.d_next[119] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34104_ (.RESET_B(net276),
    .D(_00397_),
    .Q(\u_inv.d_next[120] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34105_ (.RESET_B(net275),
    .D(_00398_),
    .Q(\u_inv.d_next[121] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34106_ (.RESET_B(net274),
    .D(_00399_),
    .Q(\u_inv.d_next[122] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34107_ (.RESET_B(net273),
    .D(_00400_),
    .Q(\u_inv.d_next[123] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34108_ (.RESET_B(net272),
    .D(_00401_),
    .Q(\u_inv.d_next[124] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34109_ (.RESET_B(net271),
    .D(_00402_),
    .Q(\u_inv.d_next[125] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34110_ (.RESET_B(net270),
    .D(_00403_),
    .Q(\u_inv.d_next[126] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34111_ (.RESET_B(net269),
    .D(_00404_),
    .Q(\u_inv.d_next[127] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34112_ (.RESET_B(net268),
    .D(_00405_),
    .Q(\u_inv.d_next[128] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34113_ (.RESET_B(net267),
    .D(_00406_),
    .Q(\u_inv.d_next[129] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34114_ (.RESET_B(net266),
    .D(_00407_),
    .Q(\u_inv.d_next[130] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34115_ (.RESET_B(net265),
    .D(_00408_),
    .Q(\u_inv.d_next[131] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34116_ (.RESET_B(net264),
    .D(_00409_),
    .Q(\u_inv.d_next[132] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34117_ (.RESET_B(net263),
    .D(_00410_),
    .Q(\u_inv.d_next[133] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34118_ (.RESET_B(net262),
    .D(_00411_),
    .Q(\u_inv.d_next[134] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34119_ (.RESET_B(net261),
    .D(_00412_),
    .Q(\u_inv.d_next[135] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34120_ (.RESET_B(net260),
    .D(_00413_),
    .Q(\u_inv.d_next[136] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34121_ (.RESET_B(net259),
    .D(_00414_),
    .Q(\u_inv.d_next[137] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34122_ (.RESET_B(net258),
    .D(_00415_),
    .Q(\u_inv.d_next[138] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34123_ (.RESET_B(net257),
    .D(_00416_),
    .Q(\u_inv.d_next[139] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34124_ (.RESET_B(net256),
    .D(_00417_),
    .Q(\u_inv.d_next[140] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34125_ (.RESET_B(net255),
    .D(_00418_),
    .Q(\u_inv.d_next[141] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34126_ (.RESET_B(net254),
    .D(_00419_),
    .Q(\u_inv.d_next[142] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34127_ (.RESET_B(net253),
    .D(_00420_),
    .Q(\u_inv.d_next[143] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34128_ (.RESET_B(net252),
    .D(_00421_),
    .Q(\u_inv.d_next[144] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34129_ (.RESET_B(net251),
    .D(_00422_),
    .Q(\u_inv.d_next[145] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34130_ (.RESET_B(net250),
    .D(_00423_),
    .Q(\u_inv.d_next[146] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34131_ (.RESET_B(net249),
    .D(_00424_),
    .Q(\u_inv.d_next[147] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34132_ (.RESET_B(net248),
    .D(_00425_),
    .Q(\u_inv.d_next[148] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _34133_ (.RESET_B(net247),
    .D(_00426_),
    .Q(\u_inv.d_next[149] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _34134_ (.RESET_B(net246),
    .D(_00427_),
    .Q(\u_inv.d_next[150] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34135_ (.RESET_B(net245),
    .D(_00428_),
    .Q(\u_inv.d_next[151] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34136_ (.RESET_B(net244),
    .D(_00429_),
    .Q(\u_inv.d_next[152] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34137_ (.RESET_B(net243),
    .D(_00430_),
    .Q(\u_inv.d_next[153] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34138_ (.RESET_B(net242),
    .D(_00431_),
    .Q(\u_inv.d_next[154] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34139_ (.RESET_B(net241),
    .D(_00432_),
    .Q(\u_inv.d_next[155] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34140_ (.RESET_B(net240),
    .D(_00433_),
    .Q(\u_inv.d_next[156] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34141_ (.RESET_B(net239),
    .D(_00434_),
    .Q(\u_inv.d_next[157] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34142_ (.RESET_B(net238),
    .D(_00435_),
    .Q(\u_inv.d_next[158] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34143_ (.RESET_B(net237),
    .D(_00436_),
    .Q(\u_inv.d_next[159] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34144_ (.RESET_B(net236),
    .D(_00437_),
    .Q(\u_inv.d_next[160] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34145_ (.RESET_B(net235),
    .D(_00438_),
    .Q(\u_inv.d_next[161] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _34146_ (.RESET_B(net234),
    .D(_00439_),
    .Q(\u_inv.d_next[162] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34147_ (.RESET_B(net233),
    .D(_00440_),
    .Q(\u_inv.d_next[163] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34148_ (.RESET_B(net232),
    .D(_00441_),
    .Q(\u_inv.d_next[164] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34149_ (.RESET_B(net231),
    .D(_00442_),
    .Q(\u_inv.d_next[165] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34150_ (.RESET_B(net230),
    .D(_00443_),
    .Q(\u_inv.d_next[166] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34151_ (.RESET_B(net229),
    .D(_00444_),
    .Q(\u_inv.d_next[167] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34152_ (.RESET_B(net228),
    .D(_00445_),
    .Q(\u_inv.d_next[168] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34153_ (.RESET_B(net227),
    .D(_00446_),
    .Q(\u_inv.d_next[169] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _34154_ (.RESET_B(net226),
    .D(_00447_),
    .Q(\u_inv.d_next[170] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _34155_ (.RESET_B(net225),
    .D(_00448_),
    .Q(\u_inv.d_next[171] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _34156_ (.RESET_B(net224),
    .D(_00449_),
    .Q(\u_inv.d_next[172] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _34157_ (.RESET_B(net223),
    .D(_00450_),
    .Q(\u_inv.d_next[173] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _34158_ (.RESET_B(net222),
    .D(_00451_),
    .Q(\u_inv.d_next[174] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _34159_ (.RESET_B(net221),
    .D(_00452_),
    .Q(\u_inv.d_next[175] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34160_ (.RESET_B(net220),
    .D(_00453_),
    .Q(\u_inv.d_next[176] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34161_ (.RESET_B(net219),
    .D(_00454_),
    .Q(\u_inv.d_next[177] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34162_ (.RESET_B(net218),
    .D(_00455_),
    .Q(\u_inv.d_next[178] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _34163_ (.RESET_B(net217),
    .D(_00456_),
    .Q(\u_inv.d_next[179] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34164_ (.RESET_B(net216),
    .D(_00457_),
    .Q(\u_inv.d_next[180] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _34165_ (.RESET_B(net215),
    .D(_00458_),
    .Q(\u_inv.d_next[181] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _34166_ (.RESET_B(net214),
    .D(_00459_),
    .Q(\u_inv.d_next[182] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34167_ (.RESET_B(net213),
    .D(_00460_),
    .Q(\u_inv.d_next[183] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34168_ (.RESET_B(net212),
    .D(_00461_),
    .Q(\u_inv.d_next[184] ),
    .CLK(clknet_6_54__leaf_clk));
 sg13g2_dfrbpq_2 _34169_ (.RESET_B(net211),
    .D(_00462_),
    .Q(\u_inv.d_next[185] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _34170_ (.RESET_B(net210),
    .D(_00463_),
    .Q(\u_inv.d_next[186] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _34171_ (.RESET_B(net209),
    .D(_00464_),
    .Q(\u_inv.d_next[187] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34172_ (.RESET_B(net208),
    .D(_00465_),
    .Q(\u_inv.d_next[188] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _34173_ (.RESET_B(net207),
    .D(_00466_),
    .Q(\u_inv.d_next[189] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34174_ (.RESET_B(net206),
    .D(_00467_),
    .Q(\u_inv.d_next[190] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34175_ (.RESET_B(net205),
    .D(_00468_),
    .Q(\u_inv.d_next[191] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34176_ (.RESET_B(net204),
    .D(_00469_),
    .Q(\u_inv.d_next[192] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _34177_ (.RESET_B(net203),
    .D(_00470_),
    .Q(\u_inv.d_next[193] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _34178_ (.RESET_B(net202),
    .D(_00471_),
    .Q(\u_inv.d_next[194] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34179_ (.RESET_B(net201),
    .D(_00472_),
    .Q(\u_inv.d_next[195] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34180_ (.RESET_B(net200),
    .D(_00473_),
    .Q(\u_inv.d_next[196] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34181_ (.RESET_B(net199),
    .D(_00474_),
    .Q(\u_inv.d_next[197] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34182_ (.RESET_B(net198),
    .D(_00475_),
    .Q(\u_inv.d_next[198] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34183_ (.RESET_B(net197),
    .D(_00476_),
    .Q(\u_inv.d_next[199] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34184_ (.RESET_B(net196),
    .D(_00477_),
    .Q(\u_inv.d_next[200] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _34185_ (.RESET_B(net195),
    .D(_00478_),
    .Q(\u_inv.d_next[201] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34186_ (.RESET_B(net194),
    .D(_00479_),
    .Q(\u_inv.d_next[202] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _34187_ (.RESET_B(net193),
    .D(_00480_),
    .Q(\u_inv.d_next[203] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _34188_ (.RESET_B(net192),
    .D(_00481_),
    .Q(\u_inv.d_next[204] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34189_ (.RESET_B(net191),
    .D(_00482_),
    .Q(\u_inv.d_next[205] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34190_ (.RESET_B(net190),
    .D(_00483_),
    .Q(\u_inv.d_next[206] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34191_ (.RESET_B(net189),
    .D(_00484_),
    .Q(\u_inv.d_next[207] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34192_ (.RESET_B(net188),
    .D(_00485_),
    .Q(\u_inv.d_next[208] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34193_ (.RESET_B(net187),
    .D(_00486_),
    .Q(\u_inv.d_next[209] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _34194_ (.RESET_B(net186),
    .D(_00487_),
    .Q(\u_inv.d_next[210] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34195_ (.RESET_B(net185),
    .D(_00488_),
    .Q(\u_inv.d_next[211] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34196_ (.RESET_B(net184),
    .D(_00489_),
    .Q(\u_inv.d_next[212] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34197_ (.RESET_B(net183),
    .D(_00490_),
    .Q(\u_inv.d_next[213] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34198_ (.RESET_B(net182),
    .D(_00491_),
    .Q(\u_inv.d_next[214] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34199_ (.RESET_B(net181),
    .D(_00492_),
    .Q(\u_inv.d_next[215] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34200_ (.RESET_B(net180),
    .D(_00493_),
    .Q(\u_inv.d_next[216] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34201_ (.RESET_B(net179),
    .D(_00494_),
    .Q(\u_inv.d_next[217] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34202_ (.RESET_B(net178),
    .D(_00495_),
    .Q(\u_inv.d_next[218] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34203_ (.RESET_B(net177),
    .D(_00496_),
    .Q(\u_inv.d_next[219] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34204_ (.RESET_B(net176),
    .D(_00497_),
    .Q(\u_inv.d_next[220] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _34205_ (.RESET_B(net175),
    .D(_00498_),
    .Q(\u_inv.d_next[221] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34206_ (.RESET_B(net174),
    .D(_00499_),
    .Q(\u_inv.d_next[222] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34207_ (.RESET_B(net173),
    .D(_00500_),
    .Q(\u_inv.d_next[223] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34208_ (.RESET_B(net172),
    .D(_00501_),
    .Q(\u_inv.d_next[224] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34209_ (.RESET_B(net171),
    .D(_00502_),
    .Q(\u_inv.d_next[225] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34210_ (.RESET_B(net170),
    .D(_00503_),
    .Q(\u_inv.d_next[226] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34211_ (.RESET_B(net169),
    .D(_00504_),
    .Q(\u_inv.d_next[227] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34212_ (.RESET_B(net168),
    .D(_00505_),
    .Q(\u_inv.d_next[228] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34213_ (.RESET_B(net167),
    .D(_00506_),
    .Q(\u_inv.d_next[229] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34214_ (.RESET_B(net166),
    .D(_00507_),
    .Q(\u_inv.d_next[230] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34215_ (.RESET_B(net165),
    .D(_00508_),
    .Q(\u_inv.d_next[231] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34216_ (.RESET_B(net164),
    .D(_00509_),
    .Q(\u_inv.d_next[232] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34217_ (.RESET_B(net163),
    .D(_00510_),
    .Q(\u_inv.d_next[233] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _34218_ (.RESET_B(net162),
    .D(_00511_),
    .Q(\u_inv.d_next[234] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34219_ (.RESET_B(net161),
    .D(_00512_),
    .Q(\u_inv.d_next[235] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34220_ (.RESET_B(net160),
    .D(_00513_),
    .Q(\u_inv.d_next[236] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34221_ (.RESET_B(net159),
    .D(_00514_),
    .Q(\u_inv.d_next[237] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34222_ (.RESET_B(net158),
    .D(_00515_),
    .Q(\u_inv.d_next[238] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34223_ (.RESET_B(net157),
    .D(_00516_),
    .Q(\u_inv.d_next[239] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34224_ (.RESET_B(net156),
    .D(_00517_),
    .Q(\u_inv.d_next[240] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34225_ (.RESET_B(net155),
    .D(_00518_),
    .Q(\u_inv.d_next[241] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34226_ (.RESET_B(net154),
    .D(_00519_),
    .Q(\u_inv.d_next[242] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34227_ (.RESET_B(net153),
    .D(_00520_),
    .Q(\u_inv.d_next[243] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34228_ (.RESET_B(net152),
    .D(_00521_),
    .Q(\u_inv.d_next[244] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34229_ (.RESET_B(net151),
    .D(_00522_),
    .Q(\u_inv.d_next[245] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34230_ (.RESET_B(net150),
    .D(_00523_),
    .Q(\u_inv.d_next[246] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34231_ (.RESET_B(net148),
    .D(_00524_),
    .Q(\u_inv.d_next[247] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34232_ (.RESET_B(net146),
    .D(_00525_),
    .Q(\u_inv.d_next[248] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34233_ (.RESET_B(net144),
    .D(_00526_),
    .Q(\u_inv.d_next[249] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34234_ (.RESET_B(net142),
    .D(_00527_),
    .Q(\u_inv.d_next[250] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34235_ (.RESET_B(net140),
    .D(_00528_),
    .Q(\u_inv.d_next[251] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _34236_ (.RESET_B(net138),
    .D(_00529_),
    .Q(\u_inv.d_next[252] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _34237_ (.RESET_B(net136),
    .D(_00530_),
    .Q(\u_inv.d_next[253] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _34238_ (.RESET_B(net134),
    .D(_00531_),
    .Q(\u_inv.d_next[254] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _34239_ (.RESET_B(net132),
    .D(_00532_),
    .Q(\u_inv.d_next[255] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34240_ (.RESET_B(net130),
    .D(_00533_),
    .Q(\u_inv.d_next[256] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _34241_ (.RESET_B(net128),
    .D(_00534_),
    .Q(\u_inv.d_reg[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _34242_ (.RESET_B(net126),
    .D(_00535_),
    .Q(\u_inv.d_reg[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _34243_ (.RESET_B(net124),
    .D(_00536_),
    .Q(\u_inv.d_reg[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _34244_ (.RESET_B(net122),
    .D(_00537_),
    .Q(\u_inv.d_reg[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _34245_ (.RESET_B(net120),
    .D(_00538_),
    .Q(\u_inv.d_reg[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _34246_ (.RESET_B(net118),
    .D(_00539_),
    .Q(\u_inv.d_reg[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _34247_ (.RESET_B(net116),
    .D(_00540_),
    .Q(\u_inv.d_reg[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _34248_ (.RESET_B(net114),
    .D(_00541_),
    .Q(\u_inv.d_reg[7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34249_ (.RESET_B(net112),
    .D(_00542_),
    .Q(\u_inv.d_reg[8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _34250_ (.RESET_B(net110),
    .D(_00543_),
    .Q(\u_inv.d_reg[9] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34251_ (.RESET_B(net108),
    .D(_00544_),
    .Q(\u_inv.d_reg[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _34252_ (.RESET_B(net106),
    .D(_00545_),
    .Q(\u_inv.d_reg[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _34253_ (.RESET_B(net104),
    .D(_00546_),
    .Q(\u_inv.d_reg[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _34254_ (.RESET_B(net102),
    .D(_00547_),
    .Q(\u_inv.d_reg[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34255_ (.RESET_B(net100),
    .D(_00548_),
    .Q(\u_inv.d_reg[14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34256_ (.RESET_B(net98),
    .D(_00549_),
    .Q(\u_inv.d_reg[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34257_ (.RESET_B(net96),
    .D(_00550_),
    .Q(\u_inv.d_reg[16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _34258_ (.RESET_B(net94),
    .D(_00551_),
    .Q(\u_inv.d_reg[17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _34259_ (.RESET_B(net92),
    .D(_00552_),
    .Q(\u_inv.d_reg[18] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _34260_ (.RESET_B(net90),
    .D(_00553_),
    .Q(\u_inv.d_reg[19] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _34261_ (.RESET_B(net88),
    .D(_00554_),
    .Q(\u_inv.d_reg[20] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _34262_ (.RESET_B(net86),
    .D(_00555_),
    .Q(\u_inv.d_reg[21] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _34263_ (.RESET_B(net84),
    .D(_00556_),
    .Q(\u_inv.d_reg[22] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _34264_ (.RESET_B(net82),
    .D(_00557_),
    .Q(\u_inv.d_reg[23] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _34265_ (.RESET_B(net80),
    .D(_00558_),
    .Q(\u_inv.d_reg[24] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _34266_ (.RESET_B(net78),
    .D(_00559_),
    .Q(\u_inv.d_reg[25] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _34267_ (.RESET_B(net76),
    .D(_00560_),
    .Q(\u_inv.d_reg[26] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34268_ (.RESET_B(net74),
    .D(_00561_),
    .Q(\u_inv.d_reg[27] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34269_ (.RESET_B(net72),
    .D(_00562_),
    .Q(\u_inv.d_reg[28] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _34270_ (.RESET_B(net70),
    .D(_00563_),
    .Q(\u_inv.d_reg[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34271_ (.RESET_B(net68),
    .D(_00564_),
    .Q(\u_inv.d_reg[30] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34272_ (.RESET_B(net66),
    .D(_00565_),
    .Q(\u_inv.d_reg[31] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34273_ (.RESET_B(net64),
    .D(_00566_),
    .Q(\u_inv.d_reg[32] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34274_ (.RESET_B(net62),
    .D(_00567_),
    .Q(\u_inv.d_reg[33] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34275_ (.RESET_B(net60),
    .D(_00568_),
    .Q(\u_inv.d_reg[34] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34276_ (.RESET_B(net58),
    .D(_00569_),
    .Q(\u_inv.d_reg[35] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34277_ (.RESET_B(net56),
    .D(_00570_),
    .Q(\u_inv.d_reg[36] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _34278_ (.RESET_B(net54),
    .D(_00571_),
    .Q(\u_inv.d_reg[37] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34279_ (.RESET_B(net52),
    .D(_00572_),
    .Q(\u_inv.d_reg[38] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34280_ (.RESET_B(net50),
    .D(_00573_),
    .Q(\u_inv.d_reg[39] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34281_ (.RESET_B(net48),
    .D(_00574_),
    .Q(\u_inv.d_reg[40] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34282_ (.RESET_B(net46),
    .D(_00575_),
    .Q(\u_inv.d_reg[41] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _34283_ (.RESET_B(net44),
    .D(_00576_),
    .Q(\u_inv.d_reg[42] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34284_ (.RESET_B(net42),
    .D(_00577_),
    .Q(\u_inv.d_reg[43] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34285_ (.RESET_B(net40),
    .D(_00578_),
    .Q(\u_inv.d_reg[44] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _34286_ (.RESET_B(net38),
    .D(_00579_),
    .Q(\u_inv.d_reg[45] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34287_ (.RESET_B(net36),
    .D(_00580_),
    .Q(\u_inv.d_reg[46] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34288_ (.RESET_B(net34),
    .D(_00581_),
    .Q(\u_inv.d_reg[47] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _34289_ (.RESET_B(net32),
    .D(_00582_),
    .Q(\u_inv.d_reg[48] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _34290_ (.RESET_B(net30),
    .D(_00583_),
    .Q(\u_inv.d_reg[49] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34291_ (.RESET_B(net28),
    .D(_00584_),
    .Q(\u_inv.d_reg[50] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34292_ (.RESET_B(net26),
    .D(_00585_),
    .Q(\u_inv.d_reg[51] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _34293_ (.RESET_B(net24),
    .D(_00586_),
    .Q(\u_inv.d_reg[52] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _34294_ (.RESET_B(net1060),
    .D(_00587_),
    .Q(\u_inv.d_reg[53] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _34295_ (.RESET_B(net1058),
    .D(_00588_),
    .Q(\u_inv.d_reg[54] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34296_ (.RESET_B(net1056),
    .D(_00589_),
    .Q(\u_inv.d_reg[55] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34297_ (.RESET_B(net1054),
    .D(_00590_),
    .Q(\u_inv.d_reg[56] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34298_ (.RESET_B(net1052),
    .D(_00591_),
    .Q(\u_inv.d_reg[57] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34299_ (.RESET_B(net1050),
    .D(_00592_),
    .Q(\u_inv.d_reg[58] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34300_ (.RESET_B(net1048),
    .D(_00593_),
    .Q(\u_inv.d_reg[59] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34301_ (.RESET_B(net1046),
    .D(_00594_),
    .Q(\u_inv.d_reg[60] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34302_ (.RESET_B(net1044),
    .D(_00595_),
    .Q(\u_inv.d_reg[61] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34303_ (.RESET_B(net1042),
    .D(_00596_),
    .Q(\u_inv.d_reg[62] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _34304_ (.RESET_B(net1040),
    .D(_00597_),
    .Q(\u_inv.d_reg[63] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _34305_ (.RESET_B(net1038),
    .D(_00598_),
    .Q(\u_inv.d_reg[64] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _34306_ (.RESET_B(net1036),
    .D(_00599_),
    .Q(\u_inv.d_reg[65] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34307_ (.RESET_B(net1034),
    .D(_00600_),
    .Q(\u_inv.d_reg[66] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _34308_ (.RESET_B(net1032),
    .D(_00601_),
    .Q(\u_inv.d_reg[67] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34309_ (.RESET_B(net1030),
    .D(_00602_),
    .Q(\u_inv.d_reg[68] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34310_ (.RESET_B(net1028),
    .D(_00603_),
    .Q(\u_inv.d_reg[69] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34311_ (.RESET_B(net1026),
    .D(_00604_),
    .Q(\u_inv.d_reg[70] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34312_ (.RESET_B(net1024),
    .D(_00605_),
    .Q(\u_inv.d_reg[71] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34313_ (.RESET_B(net1022),
    .D(_00606_),
    .Q(\u_inv.d_reg[72] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34314_ (.RESET_B(net1020),
    .D(_00607_),
    .Q(\u_inv.d_reg[73] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34315_ (.RESET_B(net1018),
    .D(_00608_),
    .Q(\u_inv.d_reg[74] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _34316_ (.RESET_B(net1016),
    .D(_00609_),
    .Q(\u_inv.d_reg[75] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _34317_ (.RESET_B(net1014),
    .D(_00610_),
    .Q(\u_inv.d_reg[76] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _34318_ (.RESET_B(net1012),
    .D(_00611_),
    .Q(\u_inv.d_reg[77] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _34319_ (.RESET_B(net1010),
    .D(_00612_),
    .Q(\u_inv.d_reg[78] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34320_ (.RESET_B(net1008),
    .D(_00613_),
    .Q(\u_inv.d_reg[79] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34321_ (.RESET_B(net1006),
    .D(_00614_),
    .Q(\u_inv.d_reg[80] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34322_ (.RESET_B(net1004),
    .D(_00615_),
    .Q(\u_inv.d_reg[81] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34323_ (.RESET_B(net1002),
    .D(_00616_),
    .Q(\u_inv.d_reg[82] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34324_ (.RESET_B(net1000),
    .D(_00617_),
    .Q(\u_inv.d_reg[83] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34325_ (.RESET_B(net998),
    .D(_00618_),
    .Q(\u_inv.d_reg[84] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34326_ (.RESET_B(net996),
    .D(_00619_),
    .Q(\u_inv.d_reg[85] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _34327_ (.RESET_B(net994),
    .D(_00620_),
    .Q(\u_inv.d_reg[86] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34328_ (.RESET_B(net992),
    .D(_00621_),
    .Q(\u_inv.d_reg[87] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34329_ (.RESET_B(net990),
    .D(_00622_),
    .Q(\u_inv.d_reg[88] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34330_ (.RESET_B(net988),
    .D(_00623_),
    .Q(\u_inv.d_reg[89] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _34331_ (.RESET_B(net986),
    .D(_00624_),
    .Q(\u_inv.d_reg[90] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34332_ (.RESET_B(net984),
    .D(_00625_),
    .Q(\u_inv.d_reg[91] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34333_ (.RESET_B(net982),
    .D(_00626_),
    .Q(\u_inv.d_reg[92] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _34334_ (.RESET_B(net980),
    .D(_00627_),
    .Q(\u_inv.d_reg[93] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34335_ (.RESET_B(net978),
    .D(_00628_),
    .Q(\u_inv.d_reg[94] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34336_ (.RESET_B(net976),
    .D(_00629_),
    .Q(\u_inv.d_reg[95] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34337_ (.RESET_B(net974),
    .D(_00630_),
    .Q(\u_inv.d_reg[96] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34338_ (.RESET_B(net972),
    .D(_00631_),
    .Q(\u_inv.d_reg[97] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _34339_ (.RESET_B(net970),
    .D(_00632_),
    .Q(\u_inv.d_reg[98] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34340_ (.RESET_B(net968),
    .D(_00633_),
    .Q(\u_inv.d_reg[99] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _34341_ (.RESET_B(net966),
    .D(_00634_),
    .Q(\u_inv.d_reg[100] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34342_ (.RESET_B(net964),
    .D(_00635_),
    .Q(\u_inv.d_reg[101] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34343_ (.RESET_B(net962),
    .D(_00636_),
    .Q(\u_inv.d_reg[102] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _34344_ (.RESET_B(net960),
    .D(_00637_),
    .Q(\u_inv.d_reg[103] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _34345_ (.RESET_B(net958),
    .D(_00638_),
    .Q(\u_inv.d_reg[104] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34346_ (.RESET_B(net956),
    .D(_00639_),
    .Q(\u_inv.d_reg[105] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34347_ (.RESET_B(net954),
    .D(_00640_),
    .Q(\u_inv.d_reg[106] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _34348_ (.RESET_B(net952),
    .D(_00641_),
    .Q(\u_inv.d_reg[107] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34349_ (.RESET_B(net950),
    .D(_00642_),
    .Q(\u_inv.d_reg[108] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34350_ (.RESET_B(net948),
    .D(_00643_),
    .Q(\u_inv.d_reg[109] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34351_ (.RESET_B(net946),
    .D(_00644_),
    .Q(\u_inv.d_reg[110] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34352_ (.RESET_B(net944),
    .D(_00645_),
    .Q(\u_inv.d_reg[111] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _34353_ (.RESET_B(net942),
    .D(_00646_),
    .Q(\u_inv.d_reg[112] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34354_ (.RESET_B(net940),
    .D(_00647_),
    .Q(\u_inv.d_reg[113] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34355_ (.RESET_B(net938),
    .D(_00648_),
    .Q(\u_inv.d_reg[114] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34356_ (.RESET_B(net936),
    .D(_00649_),
    .Q(\u_inv.d_reg[115] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34357_ (.RESET_B(net934),
    .D(_00650_),
    .Q(\u_inv.d_reg[116] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _34358_ (.RESET_B(net932),
    .D(_00651_),
    .Q(\u_inv.d_reg[117] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34359_ (.RESET_B(net930),
    .D(_00652_),
    .Q(\u_inv.d_reg[118] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34360_ (.RESET_B(net928),
    .D(_00653_),
    .Q(\u_inv.d_reg[119] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _34361_ (.RESET_B(net926),
    .D(_00654_),
    .Q(\u_inv.d_reg[120] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34362_ (.RESET_B(net924),
    .D(_00655_),
    .Q(\u_inv.d_reg[121] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34363_ (.RESET_B(net922),
    .D(_00656_),
    .Q(\u_inv.d_reg[122] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34364_ (.RESET_B(net920),
    .D(_00657_),
    .Q(\u_inv.d_reg[123] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34365_ (.RESET_B(net918),
    .D(_00658_),
    .Q(\u_inv.d_reg[124] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34366_ (.RESET_B(net916),
    .D(_00659_),
    .Q(\u_inv.d_reg[125] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34367_ (.RESET_B(net914),
    .D(_00660_),
    .Q(\u_inv.d_reg[126] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34368_ (.RESET_B(net912),
    .D(_00661_),
    .Q(\u_inv.d_reg[127] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34369_ (.RESET_B(net910),
    .D(_00662_),
    .Q(\u_inv.d_reg[128] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34370_ (.RESET_B(net908),
    .D(_00663_),
    .Q(\u_inv.d_reg[129] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _34371_ (.RESET_B(net906),
    .D(_00664_),
    .Q(\u_inv.d_reg[130] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _34372_ (.RESET_B(net904),
    .D(_00665_),
    .Q(\u_inv.d_reg[131] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34373_ (.RESET_B(net902),
    .D(_00666_),
    .Q(\u_inv.d_reg[132] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34374_ (.RESET_B(net900),
    .D(_00667_),
    .Q(\u_inv.d_reg[133] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34375_ (.RESET_B(net898),
    .D(_00668_),
    .Q(\u_inv.d_reg[134] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34376_ (.RESET_B(net896),
    .D(_00669_),
    .Q(\u_inv.d_reg[135] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34377_ (.RESET_B(net894),
    .D(_00670_),
    .Q(\u_inv.d_reg[136] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _34378_ (.RESET_B(net892),
    .D(_00671_),
    .Q(\u_inv.d_reg[137] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _34379_ (.RESET_B(net890),
    .D(_00672_),
    .Q(\u_inv.d_reg[138] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34380_ (.RESET_B(net888),
    .D(_00673_),
    .Q(\u_inv.d_reg[139] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34381_ (.RESET_B(net886),
    .D(_00674_),
    .Q(\u_inv.d_reg[140] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34382_ (.RESET_B(net884),
    .D(_00675_),
    .Q(\u_inv.d_reg[141] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34383_ (.RESET_B(net882),
    .D(_00676_),
    .Q(\u_inv.d_reg[142] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34384_ (.RESET_B(net880),
    .D(_00677_),
    .Q(\u_inv.d_reg[143] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34385_ (.RESET_B(net878),
    .D(_00678_),
    .Q(\u_inv.d_reg[144] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34386_ (.RESET_B(net876),
    .D(_00679_),
    .Q(\u_inv.d_reg[145] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _34387_ (.RESET_B(net874),
    .D(_00680_),
    .Q(\u_inv.d_reg[146] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _34388_ (.RESET_B(net872),
    .D(_00681_),
    .Q(\u_inv.d_reg[147] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _34389_ (.RESET_B(net870),
    .D(_00682_),
    .Q(\u_inv.d_reg[148] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _34390_ (.RESET_B(net868),
    .D(_00683_),
    .Q(\u_inv.d_reg[149] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _34391_ (.RESET_B(net866),
    .D(_00684_),
    .Q(\u_inv.d_reg[150] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _34392_ (.RESET_B(net864),
    .D(_00685_),
    .Q(\u_inv.d_reg[151] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _34393_ (.RESET_B(net862),
    .D(_00686_),
    .Q(\u_inv.d_reg[152] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34394_ (.RESET_B(net860),
    .D(_00687_),
    .Q(\u_inv.d_reg[153] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34395_ (.RESET_B(net858),
    .D(_00688_),
    .Q(\u_inv.d_reg[154] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34396_ (.RESET_B(net856),
    .D(_00689_),
    .Q(\u_inv.d_reg[155] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _34397_ (.RESET_B(net854),
    .D(_00690_),
    .Q(\u_inv.d_reg[156] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34398_ (.RESET_B(net852),
    .D(_00691_),
    .Q(\u_inv.d_reg[157] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34399_ (.RESET_B(net850),
    .D(_00692_),
    .Q(\u_inv.d_reg[158] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34400_ (.RESET_B(net848),
    .D(_00693_),
    .Q(\u_inv.d_reg[159] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _34401_ (.RESET_B(net846),
    .D(_00694_),
    .Q(\u_inv.d_reg[160] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _34402_ (.RESET_B(net844),
    .D(_00695_),
    .Q(\u_inv.d_reg[161] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34403_ (.RESET_B(net842),
    .D(_00696_),
    .Q(\u_inv.d_reg[162] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34404_ (.RESET_B(net840),
    .D(_00697_),
    .Q(\u_inv.d_reg[163] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _34405_ (.RESET_B(net838),
    .D(_00698_),
    .Q(\u_inv.d_reg[164] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34406_ (.RESET_B(net836),
    .D(_00699_),
    .Q(\u_inv.d_reg[165] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34407_ (.RESET_B(net834),
    .D(_00700_),
    .Q(\u_inv.d_reg[166] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34408_ (.RESET_B(net832),
    .D(_00701_),
    .Q(\u_inv.d_reg[167] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34409_ (.RESET_B(net830),
    .D(_00702_),
    .Q(\u_inv.d_reg[168] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _34410_ (.RESET_B(net828),
    .D(_00703_),
    .Q(\u_inv.d_reg[169] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _34411_ (.RESET_B(net826),
    .D(_00704_),
    .Q(\u_inv.d_reg[170] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _34412_ (.RESET_B(net824),
    .D(_00705_),
    .Q(\u_inv.d_reg[171] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _34413_ (.RESET_B(net822),
    .D(_00706_),
    .Q(\u_inv.d_reg[172] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _34414_ (.RESET_B(net820),
    .D(_00707_),
    .Q(\u_inv.d_reg[173] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _34415_ (.RESET_B(net818),
    .D(_00708_),
    .Q(\u_inv.d_reg[174] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _34416_ (.RESET_B(net816),
    .D(_00709_),
    .Q(\u_inv.d_reg[175] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34417_ (.RESET_B(net814),
    .D(_00710_),
    .Q(\u_inv.d_reg[176] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34418_ (.RESET_B(net812),
    .D(_00711_),
    .Q(\u_inv.d_reg[177] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34419_ (.RESET_B(net810),
    .D(_00712_),
    .Q(\u_inv.d_reg[178] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _34420_ (.RESET_B(net808),
    .D(_00713_),
    .Q(\u_inv.d_reg[179] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _34421_ (.RESET_B(net806),
    .D(_00714_),
    .Q(\u_inv.d_reg[180] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _34422_ (.RESET_B(net804),
    .D(_00715_),
    .Q(\u_inv.d_reg[181] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _34423_ (.RESET_B(net802),
    .D(_00716_),
    .Q(\u_inv.d_reg[182] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _34424_ (.RESET_B(net800),
    .D(_00717_),
    .Q(\u_inv.d_reg[183] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34425_ (.RESET_B(net798),
    .D(_00718_),
    .Q(\u_inv.d_reg[184] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _34426_ (.RESET_B(net796),
    .D(_00719_),
    .Q(\u_inv.d_reg[185] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34427_ (.RESET_B(net794),
    .D(_00720_),
    .Q(\u_inv.d_reg[186] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _34428_ (.RESET_B(net792),
    .D(_00721_),
    .Q(\u_inv.d_reg[187] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _34429_ (.RESET_B(net790),
    .D(_00722_),
    .Q(\u_inv.d_reg[188] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _34430_ (.RESET_B(net788),
    .D(_00723_),
    .Q(\u_inv.d_reg[189] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _34431_ (.RESET_B(net786),
    .D(_00724_),
    .Q(\u_inv.d_reg[190] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34432_ (.RESET_B(net784),
    .D(_00725_),
    .Q(\u_inv.d_reg[191] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _34433_ (.RESET_B(net782),
    .D(_00726_),
    .Q(\u_inv.d_reg[192] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34434_ (.RESET_B(net780),
    .D(_00727_),
    .Q(\u_inv.d_reg[193] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _34435_ (.RESET_B(net778),
    .D(_00728_),
    .Q(\u_inv.d_reg[194] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _34436_ (.RESET_B(net776),
    .D(_00729_),
    .Q(\u_inv.d_reg[195] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _34437_ (.RESET_B(net774),
    .D(_00730_),
    .Q(\u_inv.d_reg[196] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34438_ (.RESET_B(net772),
    .D(_00731_),
    .Q(\u_inv.d_reg[197] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34439_ (.RESET_B(net770),
    .D(_00732_),
    .Q(\u_inv.d_reg[198] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34440_ (.RESET_B(net768),
    .D(_00733_),
    .Q(\u_inv.d_reg[199] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _34441_ (.RESET_B(net766),
    .D(_00734_),
    .Q(\u_inv.d_reg[200] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34442_ (.RESET_B(net764),
    .D(_00735_),
    .Q(\u_inv.d_reg[201] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _34443_ (.RESET_B(net762),
    .D(_00736_),
    .Q(\u_inv.d_reg[202] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34444_ (.RESET_B(net760),
    .D(_00737_),
    .Q(\u_inv.d_reg[203] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34445_ (.RESET_B(net758),
    .D(_00738_),
    .Q(\u_inv.d_reg[204] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34446_ (.RESET_B(net756),
    .D(_00739_),
    .Q(\u_inv.d_reg[205] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34447_ (.RESET_B(net754),
    .D(_00740_),
    .Q(\u_inv.d_reg[206] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34448_ (.RESET_B(net752),
    .D(_00741_),
    .Q(\u_inv.d_reg[207] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34449_ (.RESET_B(net750),
    .D(_00742_),
    .Q(\u_inv.d_reg[208] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34450_ (.RESET_B(net748),
    .D(_00743_),
    .Q(\u_inv.d_reg[209] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34451_ (.RESET_B(net746),
    .D(_00744_),
    .Q(\u_inv.d_reg[210] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _34452_ (.RESET_B(net744),
    .D(_00745_),
    .Q(\u_inv.d_reg[211] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34453_ (.RESET_B(net742),
    .D(_00746_),
    .Q(\u_inv.d_reg[212] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _34454_ (.RESET_B(net740),
    .D(_00747_),
    .Q(\u_inv.d_reg[213] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34455_ (.RESET_B(net738),
    .D(_00748_),
    .Q(\u_inv.d_reg[214] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _34456_ (.RESET_B(net736),
    .D(_00749_),
    .Q(\u_inv.d_reg[215] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34457_ (.RESET_B(net734),
    .D(_00750_),
    .Q(\u_inv.d_reg[216] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34458_ (.RESET_B(net732),
    .D(_00751_),
    .Q(\u_inv.d_reg[217] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _34459_ (.RESET_B(net730),
    .D(_00752_),
    .Q(\u_inv.d_reg[218] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _34460_ (.RESET_B(net728),
    .D(_00753_),
    .Q(\u_inv.d_reg[219] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34461_ (.RESET_B(net726),
    .D(_00754_),
    .Q(\u_inv.d_reg[220] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34462_ (.RESET_B(net724),
    .D(_00755_),
    .Q(\u_inv.d_reg[221] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _34463_ (.RESET_B(net722),
    .D(_00756_),
    .Q(\u_inv.d_reg[222] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34464_ (.RESET_B(net720),
    .D(_00757_),
    .Q(\u_inv.d_reg[223] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34465_ (.RESET_B(net718),
    .D(_00758_),
    .Q(\u_inv.d_reg[224] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34466_ (.RESET_B(net716),
    .D(_00759_),
    .Q(\u_inv.d_reg[225] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _34467_ (.RESET_B(net714),
    .D(_00760_),
    .Q(\u_inv.d_reg[226] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _34468_ (.RESET_B(net712),
    .D(_00761_),
    .Q(\u_inv.d_reg[227] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _34469_ (.RESET_B(net710),
    .D(_00762_),
    .Q(\u_inv.d_reg[228] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _34470_ (.RESET_B(net708),
    .D(_00763_),
    .Q(\u_inv.d_reg[229] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34471_ (.RESET_B(net706),
    .D(_00764_),
    .Q(\u_inv.d_reg[230] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34472_ (.RESET_B(net704),
    .D(_00765_),
    .Q(\u_inv.d_reg[231] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34473_ (.RESET_B(net702),
    .D(_00766_),
    .Q(\u_inv.d_reg[232] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34474_ (.RESET_B(net700),
    .D(_00767_),
    .Q(\u_inv.d_reg[233] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _34475_ (.RESET_B(net698),
    .D(_00768_),
    .Q(\u_inv.d_reg[234] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34476_ (.RESET_B(net696),
    .D(_00769_),
    .Q(\u_inv.d_reg[235] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34477_ (.RESET_B(net694),
    .D(_00770_),
    .Q(\u_inv.d_reg[236] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _34478_ (.RESET_B(net692),
    .D(_00771_),
    .Q(\u_inv.d_reg[237] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34479_ (.RESET_B(net690),
    .D(_00772_),
    .Q(\u_inv.d_reg[238] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34480_ (.RESET_B(net688),
    .D(_00773_),
    .Q(\u_inv.d_reg[239] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _34481_ (.RESET_B(net686),
    .D(_00774_),
    .Q(\u_inv.d_reg[240] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _34482_ (.RESET_B(net684),
    .D(_00775_),
    .Q(\u_inv.d_reg[241] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34483_ (.RESET_B(net682),
    .D(_00776_),
    .Q(\u_inv.d_reg[242] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34484_ (.RESET_B(net680),
    .D(_00777_),
    .Q(\u_inv.d_reg[243] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34485_ (.RESET_B(net678),
    .D(_00778_),
    .Q(\u_inv.d_reg[244] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34486_ (.RESET_B(net676),
    .D(_00779_),
    .Q(\u_inv.d_reg[245] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34487_ (.RESET_B(net675),
    .D(_00780_),
    .Q(\u_inv.d_reg[246] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34488_ (.RESET_B(net674),
    .D(_00781_),
    .Q(\u_inv.d_reg[247] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34489_ (.RESET_B(net673),
    .D(_00782_),
    .Q(\u_inv.d_reg[248] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _34490_ (.RESET_B(net672),
    .D(_00783_),
    .Q(\u_inv.d_reg[249] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _34491_ (.RESET_B(net671),
    .D(_00784_),
    .Q(\u_inv.d_reg[250] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _34492_ (.RESET_B(net670),
    .D(_00785_),
    .Q(\u_inv.d_reg[251] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _34493_ (.RESET_B(net669),
    .D(_00786_),
    .Q(\u_inv.d_reg[252] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _34494_ (.RESET_B(net668),
    .D(_00787_),
    .Q(\u_inv.d_reg[253] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _34495_ (.RESET_B(net667),
    .D(_00788_),
    .Q(\u_inv.d_reg[254] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _34496_ (.RESET_B(net666),
    .D(_00789_),
    .Q(\u_inv.d_reg[255] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _34497_ (.RESET_B(net665),
    .D(_00790_),
    .Q(\u_inv.d_reg[256] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _34498_ (.RESET_B(net664),
    .D(_00791_),
    .Q(\u_inv.f_reg[0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _34499_ (.RESET_B(net663),
    .D(net2584),
    .Q(\u_inv.f_reg[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _34500_ (.RESET_B(net662),
    .D(net1985),
    .Q(\u_inv.f_reg[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _34501_ (.RESET_B(net661),
    .D(net2187),
    .Q(\u_inv.f_reg[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _34502_ (.RESET_B(net660),
    .D(_00795_),
    .Q(\u_inv.f_reg[4] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _34503_ (.RESET_B(net659),
    .D(net2123),
    .Q(\u_inv.f_reg[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _34504_ (.RESET_B(net658),
    .D(_00797_),
    .Q(\u_inv.f_reg[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _34505_ (.RESET_B(net657),
    .D(_00798_),
    .Q(\u_inv.f_reg[7] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _34506_ (.RESET_B(net656),
    .D(_00799_),
    .Q(\u_inv.f_reg[8] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _34507_ (.RESET_B(net655),
    .D(_00800_),
    .Q(\u_inv.f_reg[9] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _34508_ (.RESET_B(net654),
    .D(net2602),
    .Q(\u_inv.f_reg[10] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _34509_ (.RESET_B(net653),
    .D(_00802_),
    .Q(\u_inv.f_reg[11] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _34510_ (.RESET_B(net652),
    .D(_00803_),
    .Q(\u_inv.f_reg[12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _34511_ (.RESET_B(net651),
    .D(net2574),
    .Q(\u_inv.f_reg[13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _34512_ (.RESET_B(net650),
    .D(net3089),
    .Q(\u_inv.f_reg[14] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _34513_ (.RESET_B(net649),
    .D(net2296),
    .Q(\u_inv.f_reg[15] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _34514_ (.RESET_B(net648),
    .D(net2719),
    .Q(\u_inv.f_reg[16] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _34515_ (.RESET_B(net647),
    .D(_00808_),
    .Q(\u_inv.f_reg[17] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _34516_ (.RESET_B(net646),
    .D(net2291),
    .Q(\u_inv.f_reg[18] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _34517_ (.RESET_B(net645),
    .D(net2048),
    .Q(\u_inv.f_reg[19] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _34518_ (.RESET_B(net644),
    .D(net2588),
    .Q(\u_inv.f_reg[20] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _34519_ (.RESET_B(net643),
    .D(net2251),
    .Q(\u_inv.f_reg[21] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _34520_ (.RESET_B(net642),
    .D(net2228),
    .Q(\u_inv.f_reg[22] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _34521_ (.RESET_B(net641),
    .D(net2431),
    .Q(\u_inv.f_reg[23] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _34522_ (.RESET_B(net640),
    .D(_00815_),
    .Q(\u_inv.f_reg[24] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _34523_ (.RESET_B(net639),
    .D(_00816_),
    .Q(\u_inv.f_reg[25] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _34524_ (.RESET_B(net638),
    .D(net2680),
    .Q(\u_inv.f_reg[26] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _34525_ (.RESET_B(net637),
    .D(net3134),
    .Q(\u_inv.f_reg[27] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _34526_ (.RESET_B(net636),
    .D(net2518),
    .Q(\u_inv.f_reg[28] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _34527_ (.RESET_B(net635),
    .D(_00820_),
    .Q(\u_inv.f_reg[29] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _34528_ (.RESET_B(net634),
    .D(net2579),
    .Q(\u_inv.f_reg[30] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _34529_ (.RESET_B(net633),
    .D(net2713),
    .Q(\u_inv.f_reg[31] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _34530_ (.RESET_B(net632),
    .D(_00823_),
    .Q(\u_inv.f_reg[32] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _34531_ (.RESET_B(net631),
    .D(net2092),
    .Q(\u_inv.f_reg[33] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _34532_ (.RESET_B(net630),
    .D(net2711),
    .Q(\u_inv.f_reg[34] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _34533_ (.RESET_B(net629),
    .D(net2802),
    .Q(\u_inv.f_reg[35] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _34534_ (.RESET_B(net628),
    .D(_00827_),
    .Q(\u_inv.f_reg[36] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _34535_ (.RESET_B(net627),
    .D(net2503),
    .Q(\u_inv.f_reg[37] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _34536_ (.RESET_B(net626),
    .D(net2154),
    .Q(\u_inv.f_reg[38] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _34537_ (.RESET_B(net625),
    .D(net2514),
    .Q(\u_inv.f_reg[39] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _34538_ (.RESET_B(net624),
    .D(_00831_),
    .Q(\u_inv.f_reg[40] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _34539_ (.RESET_B(net623),
    .D(_00832_),
    .Q(\u_inv.f_reg[41] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _34540_ (.RESET_B(net622),
    .D(_00833_),
    .Q(\u_inv.f_reg[42] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _34541_ (.RESET_B(net621),
    .D(net3254),
    .Q(\u_inv.f_reg[43] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _34542_ (.RESET_B(net620),
    .D(net2260),
    .Q(\u_inv.f_reg[44] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _34543_ (.RESET_B(net619),
    .D(net2594),
    .Q(\u_inv.f_reg[45] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _34544_ (.RESET_B(net618),
    .D(net2457),
    .Q(\u_inv.f_reg[46] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _34545_ (.RESET_B(net617),
    .D(net2921),
    .Q(\u_inv.f_reg[47] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _34546_ (.RESET_B(net616),
    .D(net2486),
    .Q(\u_inv.f_reg[48] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _34547_ (.RESET_B(net615),
    .D(net2262),
    .Q(\u_inv.f_reg[49] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _34548_ (.RESET_B(net614),
    .D(_00841_),
    .Q(\u_inv.f_reg[50] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _34549_ (.RESET_B(net613),
    .D(_00842_),
    .Q(\u_inv.f_reg[51] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _34550_ (.RESET_B(net612),
    .D(_00843_),
    .Q(\u_inv.f_reg[52] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _34551_ (.RESET_B(net611),
    .D(_00844_),
    .Q(\u_inv.f_reg[53] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _34552_ (.RESET_B(net610),
    .D(net2552),
    .Q(\u_inv.f_reg[54] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _34553_ (.RESET_B(net609),
    .D(net2314),
    .Q(\u_inv.f_reg[55] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _34554_ (.RESET_B(net608),
    .D(_00847_),
    .Q(\u_inv.f_reg[56] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _34555_ (.RESET_B(net607),
    .D(net3179),
    .Q(\u_inv.f_reg[57] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _34556_ (.RESET_B(net606),
    .D(net2200),
    .Q(\u_inv.f_reg[58] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _34557_ (.RESET_B(net605),
    .D(net2640),
    .Q(\u_inv.f_reg[59] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _34558_ (.RESET_B(net604),
    .D(net2356),
    .Q(\u_inv.f_reg[60] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _34559_ (.RESET_B(net603),
    .D(net2474),
    .Q(\u_inv.f_reg[61] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _34560_ (.RESET_B(net602),
    .D(_00853_),
    .Q(\u_inv.f_reg[62] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _34561_ (.RESET_B(net601),
    .D(net3130),
    .Q(\u_inv.f_reg[63] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _34562_ (.RESET_B(net600),
    .D(_00855_),
    .Q(\u_inv.f_reg[64] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _34563_ (.RESET_B(net599),
    .D(_00856_),
    .Q(\u_inv.f_reg[65] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _34564_ (.RESET_B(net598),
    .D(net2218),
    .Q(\u_inv.f_reg[66] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _34565_ (.RESET_B(net597),
    .D(net2350),
    .Q(\u_inv.f_reg[67] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _34566_ (.RESET_B(net596),
    .D(_00859_),
    .Q(\u_inv.f_reg[68] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _34567_ (.RESET_B(net595),
    .D(net2555),
    .Q(\u_inv.f_reg[69] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _34568_ (.RESET_B(net594),
    .D(_00861_),
    .Q(\u_inv.f_reg[70] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _34569_ (.RESET_B(net593),
    .D(net2318),
    .Q(\u_inv.f_reg[71] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _34570_ (.RESET_B(net592),
    .D(_00863_),
    .Q(\u_inv.f_reg[72] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _34571_ (.RESET_B(net591),
    .D(_00864_),
    .Q(\u_inv.f_reg[73] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _34572_ (.RESET_B(net590),
    .D(net2572),
    .Q(\u_inv.f_reg[74] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _34573_ (.RESET_B(net589),
    .D(net2980),
    .Q(\u_inv.f_reg[75] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _34574_ (.RESET_B(net588),
    .D(net2303),
    .Q(\u_inv.f_reg[76] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _34575_ (.RESET_B(net587),
    .D(net2770),
    .Q(\u_inv.f_reg[77] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _34576_ (.RESET_B(net586),
    .D(net2272),
    .Q(\u_inv.f_reg[78] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _34577_ (.RESET_B(net585),
    .D(net2569),
    .Q(\u_inv.f_reg[79] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _34578_ (.RESET_B(net584),
    .D(net3072),
    .Q(\u_inv.f_reg[80] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _34579_ (.RESET_B(net583),
    .D(net2142),
    .Q(\u_inv.f_reg[81] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _34580_ (.RESET_B(net582),
    .D(net2383),
    .Q(\u_inv.f_reg[82] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _34581_ (.RESET_B(net581),
    .D(_00874_),
    .Q(\u_inv.f_reg[83] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _34582_ (.RESET_B(net580),
    .D(net2533),
    .Q(\u_inv.f_reg[84] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _34583_ (.RESET_B(net579),
    .D(net3157),
    .Q(\u_inv.f_reg[85] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _34584_ (.RESET_B(net578),
    .D(net1901),
    .Q(\u_inv.f_reg[86] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _34585_ (.RESET_B(net577),
    .D(net2742),
    .Q(\u_inv.f_reg[87] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _34586_ (.RESET_B(net576),
    .D(net2378),
    .Q(\u_inv.f_reg[88] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _34587_ (.RESET_B(net575),
    .D(net2866),
    .Q(\u_inv.f_reg[89] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _34588_ (.RESET_B(net574),
    .D(net2522),
    .Q(\u_inv.f_reg[90] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _34589_ (.RESET_B(net573),
    .D(_00882_),
    .Q(\u_inv.f_reg[91] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _34590_ (.RESET_B(net572),
    .D(_00883_),
    .Q(\u_inv.f_reg[92] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _34591_ (.RESET_B(net571),
    .D(net2843),
    .Q(\u_inv.f_reg[93] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _34592_ (.RESET_B(net570),
    .D(_00885_),
    .Q(\u_inv.f_reg[94] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _34593_ (.RESET_B(net569),
    .D(net2381),
    .Q(\u_inv.f_reg[95] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _34594_ (.RESET_B(net568),
    .D(net2500),
    .Q(\u_inv.f_reg[96] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _34595_ (.RESET_B(net567),
    .D(net2687),
    .Q(\u_inv.f_reg[97] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _34596_ (.RESET_B(net566),
    .D(_00889_),
    .Q(\u_inv.f_reg[98] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _34597_ (.RESET_B(net565),
    .D(_00890_),
    .Q(\u_inv.f_reg[99] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _34598_ (.RESET_B(net564),
    .D(net2888),
    .Q(\u_inv.f_reg[100] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _34599_ (.RESET_B(net563),
    .D(_00892_),
    .Q(\u_inv.f_reg[101] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _34600_ (.RESET_B(net562),
    .D(net1977),
    .Q(\u_inv.f_reg[102] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _34601_ (.RESET_B(net561),
    .D(_00894_),
    .Q(\u_inv.f_reg[103] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _34602_ (.RESET_B(net560),
    .D(net2596),
    .Q(\u_inv.f_reg[104] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _34603_ (.RESET_B(net559),
    .D(net2986),
    .Q(\u_inv.f_reg[105] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _34604_ (.RESET_B(net558),
    .D(net2373),
    .Q(\u_inv.f_reg[106] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _34605_ (.RESET_B(net557),
    .D(net2586),
    .Q(\u_inv.f_reg[107] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _34606_ (.RESET_B(net556),
    .D(net2415),
    .Q(\u_inv.f_reg[108] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _34607_ (.RESET_B(net555),
    .D(net2527),
    .Q(\u_inv.f_reg[109] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _34608_ (.RESET_B(net554),
    .D(_00901_),
    .Q(\u_inv.f_reg[110] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _34609_ (.RESET_B(net553),
    .D(net2149),
    .Q(\u_inv.f_reg[111] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _34610_ (.RESET_B(net552),
    .D(_00903_),
    .Q(\u_inv.f_reg[112] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _34611_ (.RESET_B(net551),
    .D(_00904_),
    .Q(\u_inv.f_reg[113] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _34612_ (.RESET_B(net550),
    .D(net2405),
    .Q(\u_inv.f_reg[114] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _34613_ (.RESET_B(net549),
    .D(_00906_),
    .Q(\u_inv.f_reg[115] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34614_ (.RESET_B(net548),
    .D(net2224),
    .Q(\u_inv.f_reg[116] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _34615_ (.RESET_B(net547),
    .D(_00908_),
    .Q(\u_inv.f_reg[117] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34616_ (.RESET_B(net546),
    .D(net2035),
    .Q(\u_inv.f_reg[118] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _34617_ (.RESET_B(net545),
    .D(net2470),
    .Q(\u_inv.f_reg[119] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _34618_ (.RESET_B(net544),
    .D(net2387),
    .Q(\u_inv.f_reg[120] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _34619_ (.RESET_B(net543),
    .D(net2421),
    .Q(\u_inv.f_reg[121] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _34620_ (.RESET_B(net542),
    .D(_00913_),
    .Q(\u_inv.f_reg[122] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _34621_ (.RESET_B(net541),
    .D(net2885),
    .Q(\u_inv.f_reg[123] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _34622_ (.RESET_B(net540),
    .D(_00915_),
    .Q(\u_inv.f_reg[124] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _34623_ (.RESET_B(net539),
    .D(net2172),
    .Q(\u_inv.f_reg[125] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _34624_ (.RESET_B(net538),
    .D(net2103),
    .Q(\u_inv.f_reg[126] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _34625_ (.RESET_B(net537),
    .D(net2546),
    .Q(\u_inv.f_reg[127] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _34626_ (.RESET_B(net536),
    .D(_00919_),
    .Q(\u_inv.f_reg[128] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _34627_ (.RESET_B(net535),
    .D(_00920_),
    .Q(\u_inv.f_reg[129] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _34628_ (.RESET_B(net534),
    .D(net2814),
    .Q(\u_inv.f_reg[130] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _34629_ (.RESET_B(net533),
    .D(_00922_),
    .Q(\u_inv.f_reg[131] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _34630_ (.RESET_B(net532),
    .D(_00923_),
    .Q(\u_inv.f_reg[132] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _34631_ (.RESET_B(net531),
    .D(_00924_),
    .Q(\u_inv.f_reg[133] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _34632_ (.RESET_B(net530),
    .D(_00925_),
    .Q(\u_inv.f_reg[134] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _34633_ (.RESET_B(net529),
    .D(_00926_),
    .Q(\u_inv.f_reg[135] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _34634_ (.RESET_B(net528),
    .D(net2159),
    .Q(\u_inv.f_reg[136] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _34635_ (.RESET_B(net527),
    .D(_00928_),
    .Q(\u_inv.f_reg[137] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _34636_ (.RESET_B(net526),
    .D(net2168),
    .Q(\u_inv.f_reg[138] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _34637_ (.RESET_B(net525),
    .D(net3142),
    .Q(\u_inv.f_reg[139] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _34638_ (.RESET_B(net524),
    .D(_00931_),
    .Q(\u_inv.f_reg[140] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _34639_ (.RESET_B(net523),
    .D(net2407),
    .Q(\u_inv.f_reg[141] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _34640_ (.RESET_B(net522),
    .D(_00933_),
    .Q(\u_inv.f_reg[142] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _34641_ (.RESET_B(net521),
    .D(_00934_),
    .Q(\u_inv.f_reg[143] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _34642_ (.RESET_B(net520),
    .D(_00935_),
    .Q(\u_inv.f_reg[144] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _34643_ (.RESET_B(net519),
    .D(net2684),
    .Q(\u_inv.f_reg[145] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _34644_ (.RESET_B(net518),
    .D(net3101),
    .Q(\u_inv.f_reg[146] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _34645_ (.RESET_B(net517),
    .D(net3019),
    .Q(\u_inv.f_reg[147] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _34646_ (.RESET_B(net516),
    .D(_00939_),
    .Q(\u_inv.f_reg[148] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _34647_ (.RESET_B(net515),
    .D(net2793),
    .Q(\u_inv.f_reg[149] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _34648_ (.RESET_B(net514),
    .D(net3078),
    .Q(\u_inv.f_reg[150] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _34649_ (.RESET_B(net513),
    .D(net3043),
    .Q(\u_inv.f_reg[151] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _34650_ (.RESET_B(net512),
    .D(net2335),
    .Q(\u_inv.f_reg[152] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _34651_ (.RESET_B(net511),
    .D(_00944_),
    .Q(\u_inv.f_reg[153] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _34652_ (.RESET_B(net510),
    .D(net2412),
    .Q(\u_inv.f_reg[154] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _34653_ (.RESET_B(net509),
    .D(net2828),
    .Q(\u_inv.f_reg[155] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _34654_ (.RESET_B(net508),
    .D(_00947_),
    .Q(\u_inv.f_reg[156] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _34655_ (.RESET_B(net507),
    .D(net3029),
    .Q(\u_inv.f_reg[157] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _34656_ (.RESET_B(net506),
    .D(_00949_),
    .Q(\u_inv.f_reg[158] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _34657_ (.RESET_B(net505),
    .D(net1957),
    .Q(\u_inv.f_reg[159] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _34658_ (.RESET_B(net504),
    .D(net2435),
    .Q(\u_inv.f_reg[160] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _34659_ (.RESET_B(net503),
    .D(_00952_),
    .Q(\u_inv.f_reg[161] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _34660_ (.RESET_B(net502),
    .D(_00953_),
    .Q(\u_inv.f_reg[162] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _34661_ (.RESET_B(net501),
    .D(_00954_),
    .Q(\u_inv.f_reg[163] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _34662_ (.RESET_B(net500),
    .D(_00955_),
    .Q(\u_inv.f_reg[164] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34663_ (.RESET_B(net499),
    .D(_00956_),
    .Q(\u_inv.f_reg[165] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34664_ (.RESET_B(net498),
    .D(net2003),
    .Q(\u_inv.f_reg[166] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _34665_ (.RESET_B(net497),
    .D(net2505),
    .Q(\u_inv.f_reg[167] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _34666_ (.RESET_B(net496),
    .D(_00959_),
    .Q(\u_inv.f_reg[168] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _34667_ (.RESET_B(net495),
    .D(_00960_),
    .Q(\u_inv.f_reg[169] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34668_ (.RESET_B(net494),
    .D(net2751),
    .Q(\u_inv.f_reg[170] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _34669_ (.RESET_B(net493),
    .D(net2785),
    .Q(\u_inv.f_reg[171] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _34670_ (.RESET_B(net492),
    .D(net2288),
    .Q(\u_inv.f_reg[172] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _34671_ (.RESET_B(net491),
    .D(net2203),
    .Q(\u_inv.f_reg[173] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _34672_ (.RESET_B(net490),
    .D(net2604),
    .Q(\u_inv.f_reg[174] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _34673_ (.RESET_B(net489),
    .D(_00966_),
    .Q(\u_inv.f_reg[175] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _34674_ (.RESET_B(net488),
    .D(_00967_),
    .Q(\u_inv.f_reg[176] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _34675_ (.RESET_B(net487),
    .D(_00968_),
    .Q(\u_inv.f_reg[177] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _34676_ (.RESET_B(net486),
    .D(net2248),
    .Q(\u_inv.f_reg[178] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _34677_ (.RESET_B(net485),
    .D(net2472),
    .Q(\u_inv.f_reg[179] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _34678_ (.RESET_B(net484),
    .D(net2498),
    .Q(\u_inv.f_reg[180] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _34679_ (.RESET_B(net483),
    .D(net2617),
    .Q(\u_inv.f_reg[181] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _34680_ (.RESET_B(net482),
    .D(_00973_),
    .Q(\u_inv.f_reg[182] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _34681_ (.RESET_B(net481),
    .D(_00974_),
    .Q(\u_inv.f_reg[183] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _34682_ (.RESET_B(net480),
    .D(_00975_),
    .Q(\u_inv.f_reg[184] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _34683_ (.RESET_B(net479),
    .D(_00976_),
    .Q(\u_inv.f_reg[185] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _34684_ (.RESET_B(net478),
    .D(net1942),
    .Q(\u_inv.f_reg[186] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _34685_ (.RESET_B(net477),
    .D(_00978_),
    .Q(\u_inv.f_reg[187] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _34686_ (.RESET_B(net476),
    .D(_00979_),
    .Q(\u_inv.f_reg[188] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _34687_ (.RESET_B(net475),
    .D(_00980_),
    .Q(\u_inv.f_reg[189] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _34688_ (.RESET_B(net474),
    .D(_00981_),
    .Q(\u_inv.f_reg[190] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _34689_ (.RESET_B(net473),
    .D(net2576),
    .Q(\u_inv.f_reg[191] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _34690_ (.RESET_B(net472),
    .D(_00983_),
    .Q(\u_inv.f_reg[192] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _34691_ (.RESET_B(net471),
    .D(net2772),
    .Q(\u_inv.f_reg[193] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _34692_ (.RESET_B(net470),
    .D(net2359),
    .Q(\u_inv.f_reg[194] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _34693_ (.RESET_B(net469),
    .D(net2441),
    .Q(\u_inv.f_reg[195] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _34694_ (.RESET_B(net468),
    .D(_00987_),
    .Q(\u_inv.f_reg[196] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _34695_ (.RESET_B(net467),
    .D(_00988_),
    .Q(\u_inv.f_reg[197] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _34696_ (.RESET_B(net466),
    .D(_00989_),
    .Q(\u_inv.f_reg[198] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _34697_ (.RESET_B(net465),
    .D(net2678),
    .Q(\u_inv.f_reg[199] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _34698_ (.RESET_B(net464),
    .D(_00991_),
    .Q(\u_inv.f_reg[200] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _34699_ (.RESET_B(net463),
    .D(_00992_),
    .Q(\u_inv.f_reg[201] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _34700_ (.RESET_B(net462),
    .D(_00993_),
    .Q(\u_inv.f_reg[202] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _34701_ (.RESET_B(net461),
    .D(net3260),
    .Q(\u_inv.f_reg[203] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _34702_ (.RESET_B(net460),
    .D(net2255),
    .Q(\u_inv.f_reg[204] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _34703_ (.RESET_B(net459),
    .D(net2944),
    .Q(\u_inv.f_reg[205] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _34704_ (.RESET_B(net458),
    .D(_00997_),
    .Q(\u_inv.f_reg[206] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _34705_ (.RESET_B(net457),
    .D(_00998_),
    .Q(\u_inv.f_reg[207] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _34706_ (.RESET_B(net456),
    .D(net2483),
    .Q(\u_inv.f_reg[208] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _34707_ (.RESET_B(net455),
    .D(_01000_),
    .Q(\u_inv.f_reg[209] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _34708_ (.RESET_B(net454),
    .D(_01001_),
    .Q(\u_inv.f_reg[210] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _34709_ (.RESET_B(net453),
    .D(net2833),
    .Q(\u_inv.f_reg[211] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _34710_ (.RESET_B(net452),
    .D(net2321),
    .Q(\u_inv.f_reg[212] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _34711_ (.RESET_B(net451),
    .D(net2478),
    .Q(\u_inv.f_reg[213] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _34712_ (.RESET_B(net450),
    .D(_01005_),
    .Q(\u_inv.f_reg[214] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _34713_ (.RESET_B(net449),
    .D(_01006_),
    .Q(\u_inv.f_reg[215] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _34714_ (.RESET_B(net448),
    .D(_01007_),
    .Q(\u_inv.f_reg[216] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _34715_ (.RESET_B(net447),
    .D(_01008_),
    .Q(\u_inv.f_reg[217] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _34716_ (.RESET_B(net446),
    .D(_01009_),
    .Q(\u_inv.f_reg[218] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _34717_ (.RESET_B(net445),
    .D(_01010_),
    .Q(\u_inv.f_reg[219] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _34718_ (.RESET_B(net444),
    .D(_01011_),
    .Q(\u_inv.f_reg[220] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _34719_ (.RESET_B(net443),
    .D(_01012_),
    .Q(\u_inv.f_reg[221] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _34720_ (.RESET_B(net442),
    .D(_01013_),
    .Q(\u_inv.f_reg[222] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _34721_ (.RESET_B(net441),
    .D(net2339),
    .Q(\u_inv.f_reg[223] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _34722_ (.RESET_B(net440),
    .D(_01015_),
    .Q(\u_inv.f_reg[224] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _34723_ (.RESET_B(net439),
    .D(_01016_),
    .Q(\u_inv.f_reg[225] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _34724_ (.RESET_B(net438),
    .D(net2362),
    .Q(\u_inv.f_reg[226] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _34725_ (.RESET_B(net437),
    .D(net3194),
    .Q(\u_inv.f_reg[227] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _34726_ (.RESET_B(net436),
    .D(net3278),
    .Q(\u_inv.f_reg[228] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _34727_ (.RESET_B(net435),
    .D(_01020_),
    .Q(\u_inv.f_reg[229] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _34728_ (.RESET_B(net434),
    .D(net2965),
    .Q(\u_inv.f_reg[230] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _34729_ (.RESET_B(net433),
    .D(net3250),
    .Q(\u_inv.f_reg[231] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _34730_ (.RESET_B(net432),
    .D(net2682),
    .Q(\u_inv.f_reg[232] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _34731_ (.RESET_B(net431),
    .D(_01024_),
    .Q(\u_inv.f_reg[233] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _34732_ (.RESET_B(net430),
    .D(_01025_),
    .Q(\u_inv.f_reg[234] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _34733_ (.RESET_B(net429),
    .D(net2348),
    .Q(\u_inv.f_reg[235] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _34734_ (.RESET_B(net428),
    .D(_01027_),
    .Q(\u_inv.f_reg[236] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _34735_ (.RESET_B(net427),
    .D(_01028_),
    .Q(\u_inv.f_reg[237] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _34736_ (.RESET_B(net426),
    .D(net2146),
    .Q(\u_inv.f_reg[238] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _34737_ (.RESET_B(net425),
    .D(net2765),
    .Q(\u_inv.f_reg[239] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _34738_ (.RESET_B(net424),
    .D(_01031_),
    .Q(\u_inv.f_reg[240] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _34739_ (.RESET_B(net423),
    .D(net3185),
    .Q(\u_inv.f_reg[241] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _34740_ (.RESET_B(net422),
    .D(_01033_),
    .Q(\u_inv.f_reg[242] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _34741_ (.RESET_B(net421),
    .D(_01034_),
    .Q(\u_inv.f_reg[243] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _34742_ (.RESET_B(net420),
    .D(_01035_),
    .Q(\u_inv.f_reg[244] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _34743_ (.RESET_B(net419),
    .D(_01036_),
    .Q(\u_inv.f_reg[245] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _34744_ (.RESET_B(net418),
    .D(_01037_),
    .Q(\u_inv.f_reg[246] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _34745_ (.RESET_B(net416),
    .D(_01038_),
    .Q(\u_inv.f_reg[247] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _34746_ (.RESET_B(net414),
    .D(_01039_),
    .Q(\u_inv.f_reg[248] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _34747_ (.RESET_B(net412),
    .D(net3092),
    .Q(\u_inv.f_reg[249] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _34748_ (.RESET_B(net410),
    .D(net2428),
    .Q(\u_inv.f_reg[250] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _34749_ (.RESET_B(net408),
    .D(net3076),
    .Q(\u_inv.f_reg[251] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _34750_ (.RESET_B(net407),
    .D(_01043_),
    .Q(\u_inv.f_reg[252] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _34751_ (.RESET_B(net405),
    .D(net2341),
    .Q(\u_inv.f_reg[253] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _34752_ (.RESET_B(net403),
    .D(net2536),
    .Q(\u_inv.f_reg[254] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _34753_ (.RESET_B(net401),
    .D(_01046_),
    .Q(\u_inv.f_reg[255] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _34754_ (.RESET_B(net399),
    .D(_01047_),
    .Q(\u_inv.f_reg[256] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34755_ (.RESET_B(net4818),
    .D(net1428),
    .Q(\inv_result[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _34756_ (.RESET_B(net4817),
    .D(_01049_),
    .Q(\inv_result[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _34757_ (.RESET_B(net4818),
    .D(_01050_),
    .Q(\inv_result[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _34758_ (.RESET_B(net4818),
    .D(_01051_),
    .Q(\inv_result[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _34759_ (.RESET_B(net4809),
    .D(net1691),
    .Q(\inv_result[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _34760_ (.RESET_B(net4818),
    .D(_01053_),
    .Q(\inv_result[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _34761_ (.RESET_B(net4818),
    .D(_01054_),
    .Q(\inv_result[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34762_ (.RESET_B(net4819),
    .D(_01055_),
    .Q(\inv_result[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _34763_ (.RESET_B(net4819),
    .D(_01056_),
    .Q(\inv_result[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34764_ (.RESET_B(net4819),
    .D(net1207),
    .Q(\inv_result[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34765_ (.RESET_B(net4819),
    .D(_01058_),
    .Q(\inv_result[10] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _34766_ (.RESET_B(net4818),
    .D(_01059_),
    .Q(\inv_result[11] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34767_ (.RESET_B(net4821),
    .D(_01060_),
    .Q(\inv_result[12] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34768_ (.RESET_B(net4821),
    .D(_01061_),
    .Q(\inv_result[13] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _34769_ (.RESET_B(net4821),
    .D(_01062_),
    .Q(\inv_result[14] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _34770_ (.RESET_B(net4823),
    .D(_01063_),
    .Q(\inv_result[15] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _34771_ (.RESET_B(net4821),
    .D(_01064_),
    .Q(\inv_result[16] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _34772_ (.RESET_B(net4821),
    .D(_01065_),
    .Q(\inv_result[17] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _34773_ (.RESET_B(net4821),
    .D(_01066_),
    .Q(\inv_result[18] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _34774_ (.RESET_B(net4821),
    .D(net1669),
    .Q(\inv_result[19] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _34775_ (.RESET_B(net4841),
    .D(_01068_),
    .Q(\inv_result[20] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _34776_ (.RESET_B(net4838),
    .D(_01069_),
    .Q(\inv_result[21] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _34777_ (.RESET_B(net4840),
    .D(_01070_),
    .Q(\inv_result[22] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _34778_ (.RESET_B(net4838),
    .D(_01071_),
    .Q(\inv_result[23] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _34779_ (.RESET_B(net4840),
    .D(_01072_),
    .Q(\inv_result[24] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _34780_ (.RESET_B(net4833),
    .D(_01073_),
    .Q(\inv_result[25] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _34781_ (.RESET_B(net4840),
    .D(_01074_),
    .Q(\inv_result[26] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _34782_ (.RESET_B(net4840),
    .D(_01075_),
    .Q(\inv_result[27] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _34783_ (.RESET_B(net4840),
    .D(_01076_),
    .Q(\inv_result[28] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _34784_ (.RESET_B(net4840),
    .D(_01077_),
    .Q(\inv_result[29] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _34785_ (.RESET_B(net4840),
    .D(_01078_),
    .Q(\inv_result[30] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _34786_ (.RESET_B(net4832),
    .D(_01079_),
    .Q(\inv_result[31] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _34787_ (.RESET_B(net4852),
    .D(_01080_),
    .Q(\inv_result[32] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34788_ (.RESET_B(net4852),
    .D(_01081_),
    .Q(\inv_result[33] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34789_ (.RESET_B(net4852),
    .D(_01082_),
    .Q(\inv_result[34] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34790_ (.RESET_B(net4852),
    .D(_01083_),
    .Q(\inv_result[35] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34791_ (.RESET_B(net4852),
    .D(_01084_),
    .Q(\inv_result[36] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _34792_ (.RESET_B(net4852),
    .D(_01085_),
    .Q(\inv_result[37] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34793_ (.RESET_B(net4852),
    .D(_01086_),
    .Q(\inv_result[38] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _34794_ (.RESET_B(net4845),
    .D(_01087_),
    .Q(\inv_result[39] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _34795_ (.RESET_B(net4849),
    .D(_01088_),
    .Q(\inv_result[40] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _34796_ (.RESET_B(net4849),
    .D(_01089_),
    .Q(\inv_result[41] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34797_ (.RESET_B(net4852),
    .D(_01090_),
    .Q(\inv_result[42] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _34798_ (.RESET_B(net4856),
    .D(_01091_),
    .Q(\inv_result[43] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _34799_ (.RESET_B(net4857),
    .D(_01092_),
    .Q(\inv_result[44] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _34800_ (.RESET_B(net4849),
    .D(_01093_),
    .Q(\inv_result[45] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34801_ (.RESET_B(net4847),
    .D(_01094_),
    .Q(\inv_result[46] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _34802_ (.RESET_B(net4848),
    .D(_01095_),
    .Q(\inv_result[47] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _34803_ (.RESET_B(net4862),
    .D(_01096_),
    .Q(\inv_result[48] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _34804_ (.RESET_B(net4862),
    .D(_01097_),
    .Q(\inv_result[49] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34805_ (.RESET_B(net4863),
    .D(_01098_),
    .Q(\inv_result[50] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34806_ (.RESET_B(net4863),
    .D(_01099_),
    .Q(\inv_result[51] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _34807_ (.RESET_B(net4867),
    .D(_01100_),
    .Q(\inv_result[52] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34808_ (.RESET_B(net4867),
    .D(_01101_),
    .Q(\inv_result[53] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34809_ (.RESET_B(net4869),
    .D(_01102_),
    .Q(\inv_result[54] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _34810_ (.RESET_B(net4867),
    .D(_01103_),
    .Q(\inv_result[55] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _34811_ (.RESET_B(net4868),
    .D(_01104_),
    .Q(\inv_result[56] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34812_ (.RESET_B(net4868),
    .D(_01105_),
    .Q(\inv_result[57] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34813_ (.RESET_B(net4868),
    .D(_01106_),
    .Q(\inv_result[58] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _34814_ (.RESET_B(net4868),
    .D(_01107_),
    .Q(\inv_result[59] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _34815_ (.RESET_B(net4868),
    .D(_01108_),
    .Q(\inv_result[60] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34816_ (.RESET_B(net4872),
    .D(_01109_),
    .Q(\inv_result[61] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34817_ (.RESET_B(net4881),
    .D(_01110_),
    .Q(\inv_result[62] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _34818_ (.RESET_B(net4872),
    .D(_01111_),
    .Q(\inv_result[63] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _34819_ (.RESET_B(net4868),
    .D(_01112_),
    .Q(\inv_result[64] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _34820_ (.RESET_B(net4881),
    .D(_01113_),
    .Q(\inv_result[65] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _34821_ (.RESET_B(net4881),
    .D(_01114_),
    .Q(\inv_result[66] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34822_ (.RESET_B(net4884),
    .D(_01115_),
    .Q(\inv_result[67] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _34823_ (.RESET_B(net4884),
    .D(_01116_),
    .Q(\inv_result[68] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34824_ (.RESET_B(net4884),
    .D(_01117_),
    .Q(\inv_result[69] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34825_ (.RESET_B(net4886),
    .D(_01118_),
    .Q(\inv_result[70] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _34826_ (.RESET_B(net4886),
    .D(net1433),
    .Q(\inv_result[71] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34827_ (.RESET_B(net4879),
    .D(_01120_),
    .Q(\inv_result[72] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34828_ (.RESET_B(net4879),
    .D(_01121_),
    .Q(\inv_result[73] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34829_ (.RESET_B(net4889),
    .D(_01122_),
    .Q(\inv_result[74] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34830_ (.RESET_B(net4882),
    .D(_01123_),
    .Q(\inv_result[75] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34831_ (.RESET_B(net4889),
    .D(_01124_),
    .Q(\inv_result[76] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _34832_ (.RESET_B(net4879),
    .D(_01125_),
    .Q(\inv_result[77] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _34833_ (.RESET_B(net4894),
    .D(_01126_),
    .Q(\inv_result[78] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _34834_ (.RESET_B(net4894),
    .D(net1822),
    .Q(\inv_result[79] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34835_ (.RESET_B(net4882),
    .D(_01128_),
    .Q(\inv_result[80] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34836_ (.RESET_B(net4882),
    .D(_01129_),
    .Q(\inv_result[81] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34837_ (.RESET_B(net4892),
    .D(_01130_),
    .Q(\inv_result[82] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34838_ (.RESET_B(net4882),
    .D(_01131_),
    .Q(\inv_result[83] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34839_ (.RESET_B(net4882),
    .D(_01132_),
    .Q(\inv_result[84] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34840_ (.RESET_B(net4882),
    .D(_01133_),
    .Q(\inv_result[85] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34841_ (.RESET_B(net4882),
    .D(_01134_),
    .Q(\inv_result[86] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34842_ (.RESET_B(net4891),
    .D(_01135_),
    .Q(\inv_result[87] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34843_ (.RESET_B(net4894),
    .D(_01136_),
    .Q(\inv_result[88] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34844_ (.RESET_B(net4894),
    .D(net1769),
    .Q(\inv_result[89] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34845_ (.RESET_B(net4896),
    .D(_01138_),
    .Q(\inv_result[90] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _34846_ (.RESET_B(net4892),
    .D(_01139_),
    .Q(\inv_result[91] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _34847_ (.RESET_B(net4883),
    .D(_01140_),
    .Q(\inv_result[92] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34848_ (.RESET_B(net4883),
    .D(_01141_),
    .Q(\inv_result[93] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34849_ (.RESET_B(net4894),
    .D(_01142_),
    .Q(\inv_result[94] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34850_ (.RESET_B(net4891),
    .D(_01143_),
    .Q(\inv_result[95] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _34851_ (.RESET_B(net4894),
    .D(_01144_),
    .Q(\inv_result[96] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34852_ (.RESET_B(net4895),
    .D(_01145_),
    .Q(\inv_result[97] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _34853_ (.RESET_B(net4895),
    .D(_01146_),
    .Q(\inv_result[98] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34854_ (.RESET_B(net4895),
    .D(_01147_),
    .Q(\inv_result[99] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _34855_ (.RESET_B(net4900),
    .D(_01148_),
    .Q(\inv_result[100] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34856_ (.RESET_B(net4895),
    .D(_01149_),
    .Q(\inv_result[101] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _34857_ (.RESET_B(net4894),
    .D(_01150_),
    .Q(\inv_result[102] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _34858_ (.RESET_B(net4894),
    .D(_01151_),
    .Q(\inv_result[103] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34859_ (.RESET_B(net4901),
    .D(_01152_),
    .Q(\inv_result[104] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _34860_ (.RESET_B(net4902),
    .D(_01153_),
    .Q(\inv_result[105] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34861_ (.RESET_B(net4902),
    .D(_01154_),
    .Q(\inv_result[106] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _34862_ (.RESET_B(net4908),
    .D(_01155_),
    .Q(\inv_result[107] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _34863_ (.RESET_B(net4902),
    .D(_01156_),
    .Q(\inv_result[108] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34864_ (.RESET_B(net4905),
    .D(_01157_),
    .Q(\inv_result[109] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34865_ (.RESET_B(net4902),
    .D(_01158_),
    .Q(\inv_result[110] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _34866_ (.RESET_B(net4903),
    .D(_01159_),
    .Q(\inv_result[111] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34867_ (.RESET_B(net4913),
    .D(_01160_),
    .Q(\inv_result[112] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _34868_ (.RESET_B(net4915),
    .D(_01161_),
    .Q(\inv_result[113] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34869_ (.RESET_B(net4912),
    .D(_01162_),
    .Q(\inv_result[114] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34870_ (.RESET_B(net4920),
    .D(_01163_),
    .Q(\inv_result[115] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _34871_ (.RESET_B(net4927),
    .D(_01164_),
    .Q(\inv_result[116] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _34872_ (.RESET_B(net4925),
    .D(_01165_),
    .Q(\inv_result[117] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34873_ (.RESET_B(net4920),
    .D(_01166_),
    .Q(\inv_result[118] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _34874_ (.RESET_B(net4920),
    .D(_01167_),
    .Q(\inv_result[119] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _34875_ (.RESET_B(net4920),
    .D(_01168_),
    .Q(\inv_result[120] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34876_ (.RESET_B(net4920),
    .D(_01169_),
    .Q(\inv_result[121] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _34877_ (.RESET_B(net4917),
    .D(_01170_),
    .Q(\inv_result[122] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _34878_ (.RESET_B(net4915),
    .D(_01171_),
    .Q(\inv_result[123] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34879_ (.RESET_B(net4926),
    .D(_01172_),
    .Q(\inv_result[124] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34880_ (.RESET_B(net4941),
    .D(_01173_),
    .Q(\inv_result[125] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34881_ (.RESET_B(net4925),
    .D(_01174_),
    .Q(\inv_result[126] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34882_ (.RESET_B(net4925),
    .D(_01175_),
    .Q(\inv_result[127] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34883_ (.RESET_B(net4927),
    .D(_01176_),
    .Q(\inv_result[128] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34884_ (.RESET_B(net4924),
    .D(_01177_),
    .Q(\inv_result[129] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34885_ (.RESET_B(net4924),
    .D(_01178_),
    .Q(\inv_result[130] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34886_ (.RESET_B(net4927),
    .D(_01179_),
    .Q(\inv_result[131] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34887_ (.RESET_B(net4929),
    .D(_01180_),
    .Q(\inv_result[132] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34888_ (.RESET_B(net4921),
    .D(_01181_),
    .Q(\inv_result[133] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34889_ (.RESET_B(net4921),
    .D(_01182_),
    .Q(\inv_result[134] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34890_ (.RESET_B(net4928),
    .D(_01183_),
    .Q(\inv_result[135] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _34891_ (.RESET_B(net4923),
    .D(_01184_),
    .Q(\inv_result[136] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _34892_ (.RESET_B(net4923),
    .D(_01185_),
    .Q(\inv_result[137] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _34893_ (.RESET_B(net4921),
    .D(_01186_),
    .Q(\inv_result[138] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _34894_ (.RESET_B(net4929),
    .D(_01187_),
    .Q(\inv_result[139] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _34895_ (.RESET_B(net4928),
    .D(_01188_),
    .Q(\inv_result[140] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _34896_ (.RESET_B(net4921),
    .D(_01189_),
    .Q(\inv_result[141] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34897_ (.RESET_B(net4921),
    .D(_01190_),
    .Q(\inv_result[142] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _34898_ (.RESET_B(net4923),
    .D(_01191_),
    .Q(\inv_result[143] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34899_ (.RESET_B(net4921),
    .D(_01192_),
    .Q(\inv_result[144] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _34900_ (.RESET_B(net4922),
    .D(_01193_),
    .Q(\inv_result[145] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34901_ (.RESET_B(net4929),
    .D(_01194_),
    .Q(\inv_result[146] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _34902_ (.RESET_B(net4922),
    .D(_01195_),
    .Q(\inv_result[147] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34903_ (.RESET_B(net4928),
    .D(_01196_),
    .Q(\inv_result[148] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _34904_ (.RESET_B(net4922),
    .D(_01197_),
    .Q(\inv_result[149] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _34905_ (.RESET_B(net4922),
    .D(_01198_),
    .Q(\inv_result[150] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34906_ (.RESET_B(net4921),
    .D(_01199_),
    .Q(\inv_result[151] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _34907_ (.RESET_B(net4921),
    .D(_01200_),
    .Q(\inv_result[152] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _34908_ (.RESET_B(net4924),
    .D(_01201_),
    .Q(\inv_result[153] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _34909_ (.RESET_B(net4924),
    .D(net1614),
    .Q(\inv_result[154] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34910_ (.RESET_B(net4924),
    .D(_01203_),
    .Q(\inv_result[155] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _34911_ (.RESET_B(net4926),
    .D(_01204_),
    .Q(\inv_result[156] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34912_ (.RESET_B(net4925),
    .D(_01205_),
    .Q(\inv_result[157] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _34913_ (.RESET_B(net4924),
    .D(_01206_),
    .Q(\inv_result[158] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34914_ (.RESET_B(net4924),
    .D(_01207_),
    .Q(\inv_result[159] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34915_ (.RESET_B(net4926),
    .D(_01208_),
    .Q(\inv_result[160] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34916_ (.RESET_B(net4926),
    .D(_01209_),
    .Q(\inv_result[161] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _34917_ (.RESET_B(net4925),
    .D(net1449),
    .Q(\inv_result[162] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34918_ (.RESET_B(net4925),
    .D(_01211_),
    .Q(\inv_result[163] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _34919_ (.RESET_B(net4927),
    .D(_01212_),
    .Q(\inv_result[164] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _34920_ (.RESET_B(net4927),
    .D(_01213_),
    .Q(\inv_result[165] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34921_ (.RESET_B(net4940),
    .D(_01214_),
    .Q(\inv_result[166] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _34922_ (.RESET_B(net4938),
    .D(_01215_),
    .Q(\inv_result[167] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _34923_ (.RESET_B(net4939),
    .D(_01216_),
    .Q(\inv_result[168] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _34924_ (.RESET_B(net4938),
    .D(_01217_),
    .Q(\inv_result[169] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _34925_ (.RESET_B(net4938),
    .D(_01218_),
    .Q(\inv_result[170] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34926_ (.RESET_B(net4917),
    .D(_01219_),
    .Q(\inv_result[171] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _34927_ (.RESET_B(net4938),
    .D(_01220_),
    .Q(\inv_result[172] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34928_ (.RESET_B(net4938),
    .D(_01221_),
    .Q(\inv_result[173] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _34929_ (.RESET_B(net4917),
    .D(_01222_),
    .Q(\inv_result[174] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _34930_ (.RESET_B(net4917),
    .D(_01223_),
    .Q(\inv_result[175] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _34931_ (.RESET_B(net4915),
    .D(_01224_),
    .Q(\inv_result[176] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34932_ (.RESET_B(net4911),
    .D(_01225_),
    .Q(\inv_result[177] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34933_ (.RESET_B(net4911),
    .D(_01226_),
    .Q(\inv_result[178] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _34934_ (.RESET_B(net4911),
    .D(_01227_),
    .Q(\inv_result[179] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _34935_ (.RESET_B(net4911),
    .D(_01228_),
    .Q(\inv_result[180] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _34936_ (.RESET_B(net4911),
    .D(net2209),
    .Q(\inv_result[181] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _34937_ (.RESET_B(net4912),
    .D(_01230_),
    .Q(\inv_result[182] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _34938_ (.RESET_B(net4911),
    .D(_01231_),
    .Q(\inv_result[183] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _34939_ (.RESET_B(net4905),
    .D(_01232_),
    .Q(\inv_result[184] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34940_ (.RESET_B(net4902),
    .D(_01233_),
    .Q(\inv_result[185] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34941_ (.RESET_B(net4902),
    .D(_01234_),
    .Q(\inv_result[186] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _34942_ (.RESET_B(net4902),
    .D(_01235_),
    .Q(\inv_result[187] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _34943_ (.RESET_B(net4900),
    .D(_01236_),
    .Q(\inv_result[188] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _34944_ (.RESET_B(net4902),
    .D(_01237_),
    .Q(\inv_result[189] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _34945_ (.RESET_B(net4905),
    .D(_01238_),
    .Q(\inv_result[190] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _34946_ (.RESET_B(net4905),
    .D(_01239_),
    .Q(\inv_result[191] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _34947_ (.RESET_B(net4879),
    .D(_01240_),
    .Q(\inv_result[192] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34948_ (.RESET_B(net4879),
    .D(_01241_),
    .Q(\inv_result[193] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34949_ (.RESET_B(net4881),
    .D(_01242_),
    .Q(\inv_result[194] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34950_ (.RESET_B(net4880),
    .D(_01243_),
    .Q(\inv_result[195] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34951_ (.RESET_B(net4879),
    .D(_01244_),
    .Q(\inv_result[196] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34952_ (.RESET_B(net4880),
    .D(_01245_),
    .Q(\inv_result[197] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _34953_ (.RESET_B(net4879),
    .D(_01246_),
    .Q(\inv_result[198] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _34954_ (.RESET_B(net4882),
    .D(_01247_),
    .Q(\inv_result[199] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _34955_ (.RESET_B(net4868),
    .D(_01248_),
    .Q(\inv_result[200] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _34956_ (.RESET_B(net4866),
    .D(_01249_),
    .Q(\inv_result[201] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34957_ (.RESET_B(net4866),
    .D(_01250_),
    .Q(\inv_result[202] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34958_ (.RESET_B(net4866),
    .D(_01251_),
    .Q(\inv_result[203] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34959_ (.RESET_B(net4866),
    .D(_01252_),
    .Q(\inv_result[204] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34960_ (.RESET_B(net4864),
    .D(_01253_),
    .Q(\inv_result[205] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34961_ (.RESET_B(net4864),
    .D(_01254_),
    .Q(\inv_result[206] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34962_ (.RESET_B(net4864),
    .D(_01255_),
    .Q(\inv_result[207] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34963_ (.RESET_B(net4861),
    .D(net1456),
    .Q(\inv_result[208] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _34964_ (.RESET_B(net4865),
    .D(_01257_),
    .Q(\inv_result[209] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34965_ (.RESET_B(net4864),
    .D(_01258_),
    .Q(\inv_result[210] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _34966_ (.RESET_B(net4864),
    .D(_01259_),
    .Q(\inv_result[211] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34967_ (.RESET_B(net4865),
    .D(_01260_),
    .Q(\inv_result[212] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34968_ (.RESET_B(net4860),
    .D(_01261_),
    .Q(\inv_result[213] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34969_ (.RESET_B(net4861),
    .D(_01262_),
    .Q(\inv_result[214] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _34970_ (.RESET_B(net4860),
    .D(_01263_),
    .Q(\inv_result[215] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34971_ (.RESET_B(net4860),
    .D(_01264_),
    .Q(\inv_result[216] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34972_ (.RESET_B(net4860),
    .D(_01265_),
    .Q(\inv_result[217] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34973_ (.RESET_B(net4850),
    .D(_01266_),
    .Q(\inv_result[218] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34974_ (.RESET_B(net4860),
    .D(_01267_),
    .Q(\inv_result[219] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34975_ (.RESET_B(net4860),
    .D(_01268_),
    .Q(\inv_result[220] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34976_ (.RESET_B(net4860),
    .D(_01269_),
    .Q(\inv_result[221] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34977_ (.RESET_B(net4860),
    .D(_01270_),
    .Q(\inv_result[222] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _34978_ (.RESET_B(net4850),
    .D(_01271_),
    .Q(\inv_result[223] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34979_ (.RESET_B(net4844),
    .D(_01272_),
    .Q(\inv_result[224] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _34980_ (.RESET_B(net4844),
    .D(_01273_),
    .Q(\inv_result[225] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34981_ (.RESET_B(net4844),
    .D(_01274_),
    .Q(\inv_result[226] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34982_ (.RESET_B(net4844),
    .D(_01275_),
    .Q(\inv_result[227] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _34983_ (.RESET_B(net4844),
    .D(_01276_),
    .Q(\inv_result[228] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _34984_ (.RESET_B(net4844),
    .D(_01277_),
    .Q(\inv_result[229] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _34985_ (.RESET_B(net4833),
    .D(_01278_),
    .Q(\inv_result[230] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _34986_ (.RESET_B(net4833),
    .D(_01279_),
    .Q(\inv_result[231] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _34987_ (.RESET_B(net4834),
    .D(_01280_),
    .Q(\inv_result[232] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _34988_ (.RESET_B(net4834),
    .D(_01281_),
    .Q(\inv_result[233] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _34989_ (.RESET_B(net4828),
    .D(_01282_),
    .Q(\inv_result[234] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _34990_ (.RESET_B(net4828),
    .D(_01283_),
    .Q(\inv_result[235] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _34991_ (.RESET_B(net4834),
    .D(_01284_),
    .Q(\inv_result[236] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _34992_ (.RESET_B(net4828),
    .D(_01285_),
    .Q(\inv_result[237] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _34993_ (.RESET_B(net4828),
    .D(_01286_),
    .Q(\inv_result[238] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _34994_ (.RESET_B(net4828),
    .D(_01287_),
    .Q(\inv_result[239] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _34995_ (.RESET_B(net4827),
    .D(net2033),
    .Q(\inv_result[240] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _34996_ (.RESET_B(net4828),
    .D(net1226),
    .Q(\inv_result[241] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _34997_ (.RESET_B(net4827),
    .D(_01290_),
    .Q(\inv_result[242] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _34998_ (.RESET_B(net4827),
    .D(_01291_),
    .Q(\inv_result[243] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _34999_ (.RESET_B(net4827),
    .D(net1376),
    .Q(\inv_result[244] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _35000_ (.RESET_B(net4827),
    .D(net2346),
    .Q(\inv_result[245] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _35001_ (.RESET_B(net4827),
    .D(net2107),
    .Q(\inv_result[246] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _35002_ (.RESET_B(net4808),
    .D(_01295_),
    .Q(\inv_result[247] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _35003_ (.RESET_B(net4808),
    .D(_01296_),
    .Q(\inv_result[248] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _35004_ (.RESET_B(net4808),
    .D(_01297_),
    .Q(\inv_result[249] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _35005_ (.RESET_B(net4808),
    .D(_01298_),
    .Q(\inv_result[250] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _35006_ (.RESET_B(net4808),
    .D(_01299_),
    .Q(\inv_result[251] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _35007_ (.RESET_B(net4808),
    .D(_01300_),
    .Q(\inv_result[252] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _35008_ (.RESET_B(net4808),
    .D(_01301_),
    .Q(\inv_result[253] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _35009_ (.RESET_B(net4808),
    .D(_01302_),
    .Q(\inv_result[254] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _35010_ (.RESET_B(net4809),
    .D(_01303_),
    .Q(\inv_result[255] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _35011_ (.RESET_B(net149),
    .D(_01304_),
    .Q(\u_inv.f_next[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _35012_ (.RESET_B(net147),
    .D(_01305_),
    .Q(\u_inv.f_next[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _35013_ (.RESET_B(net145),
    .D(_01306_),
    .Q(\u_inv.f_next[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _35014_ (.RESET_B(net143),
    .D(_01307_),
    .Q(\u_inv.f_next[3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _35015_ (.RESET_B(net141),
    .D(_01308_),
    .Q(\u_inv.f_next[4] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _35016_ (.RESET_B(net139),
    .D(_01309_),
    .Q(\u_inv.f_next[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _35017_ (.RESET_B(net137),
    .D(_01310_),
    .Q(\u_inv.f_next[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _35018_ (.RESET_B(net135),
    .D(net2706),
    .Q(\u_inv.f_next[7] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _35019_ (.RESET_B(net133),
    .D(_01312_),
    .Q(\u_inv.f_next[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _35020_ (.RESET_B(net131),
    .D(net2395),
    .Q(\u_inv.f_next[9] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _35021_ (.RESET_B(net129),
    .D(_01314_),
    .Q(\u_inv.f_next[10] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _35022_ (.RESET_B(net127),
    .D(_01315_),
    .Q(\u_inv.f_next[11] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _35023_ (.RESET_B(net125),
    .D(net2529),
    .Q(\u_inv.f_next[12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _35024_ (.RESET_B(net123),
    .D(_01317_),
    .Q(\u_inv.f_next[13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _35025_ (.RESET_B(net121),
    .D(_01318_),
    .Q(\u_inv.f_next[14] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _35026_ (.RESET_B(net119),
    .D(net3065),
    .Q(\u_inv.f_next[15] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _35027_ (.RESET_B(net117),
    .D(_01320_),
    .Q(\u_inv.f_next[16] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _35028_ (.RESET_B(net115),
    .D(net1745),
    .Q(\u_inv.f_next[17] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _35029_ (.RESET_B(net113),
    .D(_01322_),
    .Q(\u_inv.f_next[18] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _35030_ (.RESET_B(net111),
    .D(_01323_),
    .Q(\u_inv.f_next[19] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _35031_ (.RESET_B(net109),
    .D(_01324_),
    .Q(\u_inv.f_next[20] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _35032_ (.RESET_B(net107),
    .D(_01325_),
    .Q(\u_inv.f_next[21] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _35033_ (.RESET_B(net105),
    .D(_01326_),
    .Q(\u_inv.f_next[22] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _35034_ (.RESET_B(net103),
    .D(_01327_),
    .Q(\u_inv.f_next[23] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _35035_ (.RESET_B(net101),
    .D(net1755),
    .Q(\u_inv.f_next[24] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _35036_ (.RESET_B(net99),
    .D(net2723),
    .Q(\u_inv.f_next[25] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _35037_ (.RESET_B(net97),
    .D(_01330_),
    .Q(\u_inv.f_next[26] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _35038_ (.RESET_B(net95),
    .D(_01331_),
    .Q(\u_inv.f_next[27] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _35039_ (.RESET_B(net93),
    .D(_01332_),
    .Q(\u_inv.f_next[28] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _35040_ (.RESET_B(net91),
    .D(net3120),
    .Q(\u_inv.f_next[29] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _35041_ (.RESET_B(net89),
    .D(_01334_),
    .Q(\u_inv.f_next[30] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _35042_ (.RESET_B(net87),
    .D(_01335_),
    .Q(\u_inv.f_next[31] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _35043_ (.RESET_B(net85),
    .D(net2281),
    .Q(\u_inv.f_next[32] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _35044_ (.RESET_B(net83),
    .D(_01337_),
    .Q(\u_inv.f_next[33] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _35045_ (.RESET_B(net81),
    .D(_01338_),
    .Q(\u_inv.f_next[34] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _35046_ (.RESET_B(net79),
    .D(_01339_),
    .Q(\u_inv.f_next[35] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _35047_ (.RESET_B(net77),
    .D(net2078),
    .Q(\u_inv.f_next[36] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _35048_ (.RESET_B(net75),
    .D(_01341_),
    .Q(\u_inv.f_next[37] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _35049_ (.RESET_B(net73),
    .D(net2611),
    .Q(\u_inv.f_next[38] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35050_ (.RESET_B(net71),
    .D(_01343_),
    .Q(\u_inv.f_next[39] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _35051_ (.RESET_B(net69),
    .D(_01344_),
    .Q(\u_inv.f_next[40] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _35052_ (.RESET_B(net67),
    .D(net1906),
    .Q(\u_inv.f_next[41] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _35053_ (.RESET_B(net65),
    .D(net2307),
    .Q(\u_inv.f_next[42] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35054_ (.RESET_B(net63),
    .D(_01347_),
    .Q(\u_inv.f_next[43] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35055_ (.RESET_B(net61),
    .D(net3014),
    .Q(\u_inv.f_next[44] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35056_ (.RESET_B(net59),
    .D(_01349_),
    .Q(\u_inv.f_next[45] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _35057_ (.RESET_B(net57),
    .D(_01350_),
    .Q(\u_inv.f_next[46] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _35058_ (.RESET_B(net55),
    .D(_01351_),
    .Q(\u_inv.f_next[47] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35059_ (.RESET_B(net53),
    .D(_01352_),
    .Q(\u_inv.f_next[48] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _35060_ (.RESET_B(net51),
    .D(_01353_),
    .Q(\u_inv.f_next[49] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _35061_ (.RESET_B(net49),
    .D(net2235),
    .Q(\u_inv.f_next[50] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _35062_ (.RESET_B(net47),
    .D(_01355_),
    .Q(\u_inv.f_next[51] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _35063_ (.RESET_B(net45),
    .D(net2403),
    .Q(\u_inv.f_next[52] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _35064_ (.RESET_B(net43),
    .D(net2858),
    .Q(\u_inv.f_next[53] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _35065_ (.RESET_B(net41),
    .D(_01358_),
    .Q(\u_inv.f_next[54] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _35066_ (.RESET_B(net39),
    .D(_01359_),
    .Q(\u_inv.f_next[55] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _35067_ (.RESET_B(net37),
    .D(net2690),
    .Q(\u_inv.f_next[56] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _35068_ (.RESET_B(net35),
    .D(_01361_),
    .Q(\u_inv.f_next[57] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _35069_ (.RESET_B(net33),
    .D(_01362_),
    .Q(\u_inv.f_next[58] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _35070_ (.RESET_B(net31),
    .D(net2656),
    .Q(\u_inv.f_next[59] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _35071_ (.RESET_B(net29),
    .D(net3125),
    .Q(\u_inv.f_next[60] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _35072_ (.RESET_B(net27),
    .D(_01365_),
    .Q(\u_inv.f_next[61] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _35073_ (.RESET_B(net25),
    .D(net1970),
    .Q(\u_inv.f_next[62] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _35074_ (.RESET_B(net23),
    .D(_01367_),
    .Q(\u_inv.f_next[63] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _35075_ (.RESET_B(net1059),
    .D(_01368_),
    .Q(\u_inv.f_next[64] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _35076_ (.RESET_B(net1057),
    .D(net2052),
    .Q(\u_inv.f_next[65] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _35077_ (.RESET_B(net1055),
    .D(_01370_),
    .Q(\u_inv.f_next[66] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _35078_ (.RESET_B(net1053),
    .D(_01371_),
    .Q(\u_inv.f_next[67] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _35079_ (.RESET_B(net1051),
    .D(net2061),
    .Q(\u_inv.f_next[68] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _35080_ (.RESET_B(net1049),
    .D(_01373_),
    .Q(\u_inv.f_next[69] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _35081_ (.RESET_B(net1047),
    .D(net1540),
    .Q(\u_inv.f_next[70] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _35082_ (.RESET_B(net1045),
    .D(_01375_),
    .Q(\u_inv.f_next[71] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _35083_ (.RESET_B(net1043),
    .D(net2068),
    .Q(\u_inv.f_next[72] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _35084_ (.RESET_B(net1041),
    .D(net2309),
    .Q(\u_inv.f_next[73] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _35085_ (.RESET_B(net1039),
    .D(_01378_),
    .Q(\u_inv.f_next[74] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _35086_ (.RESET_B(net1037),
    .D(_01379_),
    .Q(\u_inv.f_next[75] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _35087_ (.RESET_B(net1035),
    .D(_01380_),
    .Q(\u_inv.f_next[76] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _35088_ (.RESET_B(net1033),
    .D(_01381_),
    .Q(\u_inv.f_next[77] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _35089_ (.RESET_B(net1031),
    .D(_01382_),
    .Q(\u_inv.f_next[78] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _35090_ (.RESET_B(net1029),
    .D(_01383_),
    .Q(\u_inv.f_next[79] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _35091_ (.RESET_B(net1027),
    .D(_01384_),
    .Q(\u_inv.f_next[80] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _35092_ (.RESET_B(net1025),
    .D(net2376),
    .Q(\u_inv.f_next[81] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _35093_ (.RESET_B(net1023),
    .D(_01386_),
    .Q(\u_inv.f_next[82] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _35094_ (.RESET_B(net1021),
    .D(_01387_),
    .Q(\u_inv.f_next[83] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _35095_ (.RESET_B(net1019),
    .D(net3154),
    .Q(\u_inv.f_next[84] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _35096_ (.RESET_B(net1017),
    .D(_01389_),
    .Q(\u_inv.f_next[85] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _35097_ (.RESET_B(net1015),
    .D(_01390_),
    .Q(\u_inv.f_next[86] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _35098_ (.RESET_B(net1013),
    .D(net2820),
    .Q(\u_inv.f_next[87] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _35099_ (.RESET_B(net1011),
    .D(_01392_),
    .Q(\u_inv.f_next[88] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _35100_ (.RESET_B(net1009),
    .D(_01393_),
    .Q(\u_inv.f_next[89] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _35101_ (.RESET_B(net1007),
    .D(_01394_),
    .Q(\u_inv.f_next[90] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _35102_ (.RESET_B(net1005),
    .D(_01395_),
    .Q(\u_inv.f_next[91] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _35103_ (.RESET_B(net1003),
    .D(net2354),
    .Q(\u_inv.f_next[92] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _35104_ (.RESET_B(net1001),
    .D(_01397_),
    .Q(\u_inv.f_next[93] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _35105_ (.RESET_B(net999),
    .D(net1800),
    .Q(\u_inv.f_next[94] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _35106_ (.RESET_B(net997),
    .D(_01399_),
    .Q(\u_inv.f_next[95] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _35107_ (.RESET_B(net995),
    .D(_01400_),
    .Q(\u_inv.f_next[96] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _35108_ (.RESET_B(net993),
    .D(_01401_),
    .Q(\u_inv.f_next[97] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _35109_ (.RESET_B(net991),
    .D(_01402_),
    .Q(\u_inv.f_next[98] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35110_ (.RESET_B(net989),
    .D(net1762),
    .Q(\u_inv.f_next[99] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _35111_ (.RESET_B(net987),
    .D(_01404_),
    .Q(\u_inv.f_next[100] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _35112_ (.RESET_B(net985),
    .D(net2019),
    .Q(\u_inv.f_next[101] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _35113_ (.RESET_B(net983),
    .D(_01406_),
    .Q(\u_inv.f_next[102] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _35114_ (.RESET_B(net981),
    .D(net2329),
    .Q(\u_inv.f_next[103] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _35115_ (.RESET_B(net979),
    .D(net3163),
    .Q(\u_inv.f_next[104] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _35116_ (.RESET_B(net977),
    .D(_01409_),
    .Q(\u_inv.f_next[105] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _35117_ (.RESET_B(net975),
    .D(net3285),
    .Q(\u_inv.f_next[106] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _35118_ (.RESET_B(net973),
    .D(_01411_),
    .Q(\u_inv.f_next[107] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _35119_ (.RESET_B(net971),
    .D(_01412_),
    .Q(\u_inv.f_next[108] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _35120_ (.RESET_B(net969),
    .D(_01413_),
    .Q(\u_inv.f_next[109] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _35121_ (.RESET_B(net967),
    .D(net2101),
    .Q(\u_inv.f_next[110] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _35122_ (.RESET_B(net965),
    .D(_01415_),
    .Q(\u_inv.f_next[111] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _35123_ (.RESET_B(net963),
    .D(net1528),
    .Q(\u_inv.f_next[112] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _35124_ (.RESET_B(net961),
    .D(_01417_),
    .Q(\u_inv.f_next[113] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _35125_ (.RESET_B(net959),
    .D(_01418_),
    .Q(\u_inv.f_next[114] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _35126_ (.RESET_B(net957),
    .D(_01419_),
    .Q(\u_inv.f_next[115] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _35127_ (.RESET_B(net955),
    .D(_01420_),
    .Q(\u_inv.f_next[116] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _35128_ (.RESET_B(net953),
    .D(net2990),
    .Q(\u_inv.f_next[117] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _35129_ (.RESET_B(net951),
    .D(_01422_),
    .Q(\u_inv.f_next[118] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _35130_ (.RESET_B(net949),
    .D(net2768),
    .Q(\u_inv.f_next[119] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _35131_ (.RESET_B(net947),
    .D(_01424_),
    .Q(\u_inv.f_next[120] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _35132_ (.RESET_B(net945),
    .D(_01425_),
    .Q(\u_inv.f_next[121] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _35133_ (.RESET_B(net943),
    .D(net2165),
    .Q(\u_inv.f_next[122] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _35134_ (.RESET_B(net941),
    .D(_01427_),
    .Q(\u_inv.f_next[123] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _35135_ (.RESET_B(net939),
    .D(net1559),
    .Q(\u_inv.f_next[124] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _35136_ (.RESET_B(net937),
    .D(_01429_),
    .Q(\u_inv.f_next[125] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _35137_ (.RESET_B(net935),
    .D(_01430_),
    .Q(\u_inv.f_next[126] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _35138_ (.RESET_B(net933),
    .D(_01431_),
    .Q(\u_inv.f_next[127] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _35139_ (.RESET_B(net931),
    .D(_01432_),
    .Q(\u_inv.f_next[128] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _35140_ (.RESET_B(net929),
    .D(net1879),
    .Q(\u_inv.f_next[129] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _35141_ (.RESET_B(net927),
    .D(_01434_),
    .Q(\u_inv.f_next[130] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _35142_ (.RESET_B(net925),
    .D(_01435_),
    .Q(\u_inv.f_next[131] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _35143_ (.RESET_B(net923),
    .D(net2098),
    .Q(\u_inv.f_next[132] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _35144_ (.RESET_B(net921),
    .D(net2401),
    .Q(\u_inv.f_next[133] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _35145_ (.RESET_B(net919),
    .D(net2619),
    .Q(\u_inv.f_next[134] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _35146_ (.RESET_B(net917),
    .D(net2869),
    .Q(\u_inv.f_next[135] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _35147_ (.RESET_B(net915),
    .D(_01440_),
    .Q(\u_inv.f_next[136] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _35148_ (.RESET_B(net913),
    .D(net2333),
    .Q(\u_inv.f_next[137] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _35149_ (.RESET_B(net911),
    .D(net2543),
    .Q(\u_inv.f_next[138] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _35150_ (.RESET_B(net909),
    .D(_01443_),
    .Q(\u_inv.f_next[139] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _35151_ (.RESET_B(net907),
    .D(net1729),
    .Q(\u_inv.f_next[140] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _35152_ (.RESET_B(net905),
    .D(_01445_),
    .Q(\u_inv.f_next[141] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _35153_ (.RESET_B(net903),
    .D(_01446_),
    .Q(\u_inv.f_next[142] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _35154_ (.RESET_B(net901),
    .D(_01447_),
    .Q(\u_inv.f_next[143] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _35155_ (.RESET_B(net899),
    .D(net2074),
    .Q(\u_inv.f_next[144] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _35156_ (.RESET_B(net897),
    .D(net2739),
    .Q(\u_inv.f_next[145] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _35157_ (.RESET_B(net895),
    .D(_01450_),
    .Q(\u_inv.f_next[146] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _35158_ (.RESET_B(net893),
    .D(_01451_),
    .Q(\u_inv.f_next[147] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _35159_ (.RESET_B(net891),
    .D(_01452_),
    .Q(\u_inv.f_next[148] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _35160_ (.RESET_B(net889),
    .D(_01453_),
    .Q(\u_inv.f_next[149] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _35161_ (.RESET_B(net887),
    .D(_01454_),
    .Q(\u_inv.f_next[150] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _35162_ (.RESET_B(net885),
    .D(_01455_),
    .Q(\u_inv.f_next[151] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _35163_ (.RESET_B(net883),
    .D(_01456_),
    .Q(\u_inv.f_next[152] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _35164_ (.RESET_B(net881),
    .D(_01457_),
    .Q(\u_inv.f_next[153] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _35165_ (.RESET_B(net879),
    .D(_01458_),
    .Q(\u_inv.f_next[154] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _35166_ (.RESET_B(net877),
    .D(_01459_),
    .Q(\u_inv.f_next[155] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _35167_ (.RESET_B(net875),
    .D(net1749),
    .Q(\u_inv.f_next[156] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _35168_ (.RESET_B(net873),
    .D(_01461_),
    .Q(\u_inv.f_next[157] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _35169_ (.RESET_B(net871),
    .D(net1476),
    .Q(\u_inv.f_next[158] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _35170_ (.RESET_B(net869),
    .D(net1220),
    .Q(\u_inv.f_next[159] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _35171_ (.RESET_B(net867),
    .D(net3272),
    .Q(\u_inv.f_next[160] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _35172_ (.RESET_B(net865),
    .D(_01465_),
    .Q(\u_inv.f_next[161] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _35173_ (.RESET_B(net863),
    .D(net1773),
    .Q(\u_inv.f_next[162] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _35174_ (.RESET_B(net861),
    .D(net1909),
    .Q(\u_inv.f_next[163] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _35175_ (.RESET_B(net859),
    .D(net2257),
    .Q(\u_inv.f_next[164] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _35176_ (.RESET_B(net857),
    .D(_01469_),
    .Q(\u_inv.f_next[165] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _35177_ (.RESET_B(net855),
    .D(net2022),
    .Q(\u_inv.f_next[166] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _35178_ (.RESET_B(net853),
    .D(_01471_),
    .Q(\u_inv.f_next[167] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _35179_ (.RESET_B(net851),
    .D(_01472_),
    .Q(\u_inv.f_next[168] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _35180_ (.RESET_B(net849),
    .D(net2084),
    .Q(\u_inv.f_next[169] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _35181_ (.RESET_B(net847),
    .D(_01474_),
    .Q(\u_inv.f_next[170] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _35182_ (.RESET_B(net845),
    .D(_01475_),
    .Q(\u_inv.f_next[171] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _35183_ (.RESET_B(net843),
    .D(_01476_),
    .Q(\u_inv.f_next[172] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _35184_ (.RESET_B(net841),
    .D(_01477_),
    .Q(\u_inv.f_next[173] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _35185_ (.RESET_B(net839),
    .D(_01478_),
    .Q(\u_inv.f_next[174] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _35186_ (.RESET_B(net837),
    .D(net2192),
    .Q(\u_inv.f_next[175] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _35187_ (.RESET_B(net835),
    .D(net2045),
    .Q(\u_inv.f_next[176] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _35188_ (.RESET_B(net833),
    .D(net2232),
    .Q(\u_inv.f_next[177] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35189_ (.RESET_B(net831),
    .D(_01482_),
    .Q(\u_inv.f_next[178] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _35190_ (.RESET_B(net829),
    .D(_01483_),
    .Q(\u_inv.f_next[179] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _35191_ (.RESET_B(net827),
    .D(_01484_),
    .Q(\u_inv.f_next[180] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _35192_ (.RESET_B(net825),
    .D(_01485_),
    .Q(\u_inv.f_next[181] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _35193_ (.RESET_B(net823),
    .D(_01486_),
    .Q(\u_inv.f_next[182] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _35194_ (.RESET_B(net821),
    .D(_01487_),
    .Q(\u_inv.f_next[183] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _35195_ (.RESET_B(net819),
    .D(net2152),
    .Q(\u_inv.f_next[184] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35196_ (.RESET_B(net817),
    .D(net2176),
    .Q(\u_inv.f_next[185] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35197_ (.RESET_B(net815),
    .D(_01490_),
    .Q(\u_inv.f_next[186] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _35198_ (.RESET_B(net813),
    .D(_01491_),
    .Q(\u_inv.f_next[187] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _35199_ (.RESET_B(net811),
    .D(_01492_),
    .Q(\u_inv.f_next[188] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _35200_ (.RESET_B(net809),
    .D(net2130),
    .Q(\u_inv.f_next[189] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _35201_ (.RESET_B(net807),
    .D(_01494_),
    .Q(\u_inv.f_next[190] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35202_ (.RESET_B(net805),
    .D(_01495_),
    .Q(\u_inv.f_next[191] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _35203_ (.RESET_B(net803),
    .D(net2243),
    .Q(\u_inv.f_next[192] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _35204_ (.RESET_B(net801),
    .D(_01497_),
    .Q(\u_inv.f_next[193] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _35205_ (.RESET_B(net799),
    .D(_01498_),
    .Q(\u_inv.f_next[194] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _35206_ (.RESET_B(net797),
    .D(_01499_),
    .Q(\u_inv.f_next[195] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _35207_ (.RESET_B(net795),
    .D(net1771),
    .Q(\u_inv.f_next[196] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _35208_ (.RESET_B(net793),
    .D(net1705),
    .Q(\u_inv.f_next[197] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _35209_ (.RESET_B(net791),
    .D(net1628),
    .Q(\u_inv.f_next[198] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _35210_ (.RESET_B(net789),
    .D(_01503_),
    .Q(\u_inv.f_next[199] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _35211_ (.RESET_B(net787),
    .D(_01504_),
    .Q(\u_inv.f_next[200] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _35212_ (.RESET_B(net785),
    .D(_01505_),
    .Q(\u_inv.f_next[201] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _35213_ (.RESET_B(net783),
    .D(net1960),
    .Q(\u_inv.f_next[202] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _35214_ (.RESET_B(net781),
    .D(_01507_),
    .Q(\u_inv.f_next[203] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _35215_ (.RESET_B(net779),
    .D(_01508_),
    .Q(\u_inv.f_next[204] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _35216_ (.RESET_B(net777),
    .D(_01509_),
    .Q(\u_inv.f_next[205] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _35217_ (.RESET_B(net775),
    .D(_01510_),
    .Q(\u_inv.f_next[206] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _35218_ (.RESET_B(net773),
    .D(net2178),
    .Q(\u_inv.f_next[207] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _35219_ (.RESET_B(net771),
    .D(_01512_),
    .Q(\u_inv.f_next[208] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _35220_ (.RESET_B(net769),
    .D(_01513_),
    .Q(\u_inv.f_next[209] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _35221_ (.RESET_B(net767),
    .D(net2207),
    .Q(\u_inv.f_next[210] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _35222_ (.RESET_B(net765),
    .D(_01515_),
    .Q(\u_inv.f_next[211] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _35223_ (.RESET_B(net763),
    .D(_01516_),
    .Q(\u_inv.f_next[212] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _35224_ (.RESET_B(net761),
    .D(_01517_),
    .Q(\u_inv.f_next[213] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _35225_ (.RESET_B(net759),
    .D(net1697),
    .Q(\u_inv.f_next[214] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _35226_ (.RESET_B(net757),
    .D(net2125),
    .Q(\u_inv.f_next[215] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _35227_ (.RESET_B(net755),
    .D(net2196),
    .Q(\u_inv.f_next[216] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _35228_ (.RESET_B(net753),
    .D(_01521_),
    .Q(\u_inv.f_next[217] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _35229_ (.RESET_B(net751),
    .D(net2110),
    .Q(\u_inv.f_next[218] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _35230_ (.RESET_B(net749),
    .D(_01523_),
    .Q(\u_inv.f_next[219] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _35231_ (.RESET_B(net747),
    .D(net1710),
    .Q(\u_inv.f_next[220] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _35232_ (.RESET_B(net745),
    .D(_01525_),
    .Q(\u_inv.f_next[221] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _35233_ (.RESET_B(net743),
    .D(net1464),
    .Q(\u_inv.f_next[222] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _35234_ (.RESET_B(net741),
    .D(_01527_),
    .Q(\u_inv.f_next[223] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _35235_ (.RESET_B(net739),
    .D(_01528_),
    .Q(\u_inv.f_next[224] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _35236_ (.RESET_B(net737),
    .D(net2267),
    .Q(\u_inv.f_next[225] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _35237_ (.RESET_B(net735),
    .D(net2701),
    .Q(\u_inv.f_next[226] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _35238_ (.RESET_B(net733),
    .D(_01531_),
    .Q(\u_inv.f_next[227] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _35239_ (.RESET_B(net731),
    .D(_01532_),
    .Q(\u_inv.f_next[228] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _35240_ (.RESET_B(net729),
    .D(net2213),
    .Q(\u_inv.f_next[229] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _35241_ (.RESET_B(net727),
    .D(net3264),
    .Q(\u_inv.f_next[230] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _35242_ (.RESET_B(net725),
    .D(_01535_),
    .Q(\u_inv.f_next[231] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _35243_ (.RESET_B(net723),
    .D(_01536_),
    .Q(\u_inv.f_next[232] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _35244_ (.RESET_B(net721),
    .D(_01537_),
    .Q(\u_inv.f_next[233] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _35245_ (.RESET_B(net719),
    .D(net1413),
    .Q(\u_inv.f_next[234] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _35246_ (.RESET_B(net717),
    .D(_01539_),
    .Q(\u_inv.f_next[235] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _35247_ (.RESET_B(net715),
    .D(net1626),
    .Q(\u_inv.f_next[236] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _35248_ (.RESET_B(net713),
    .D(net1968),
    .Q(\u_inv.f_next[237] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _35249_ (.RESET_B(net711),
    .D(_01542_),
    .Q(\u_inv.f_next[238] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _35250_ (.RESET_B(net709),
    .D(_01543_),
    .Q(\u_inv.f_next[239] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _35251_ (.RESET_B(net707),
    .D(net2697),
    .Q(\u_inv.f_next[240] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _35252_ (.RESET_B(net705),
    .D(_01545_),
    .Q(\u_inv.f_next[241] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _35253_ (.RESET_B(net703),
    .D(net1827),
    .Q(\u_inv.f_next[242] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _35254_ (.RESET_B(net701),
    .D(_01547_),
    .Q(\u_inv.f_next[243] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _35255_ (.RESET_B(net699),
    .D(net1440),
    .Q(\u_inv.f_next[244] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _35256_ (.RESET_B(net697),
    .D(_01549_),
    .Q(\u_inv.f_next[245] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _35257_ (.RESET_B(net695),
    .D(net1662),
    .Q(\u_inv.f_next[246] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _35258_ (.RESET_B(net693),
    .D(net2337),
    .Q(\u_inv.f_next[247] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _35259_ (.RESET_B(net691),
    .D(net2891),
    .Q(\u_inv.f_next[248] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _35260_ (.RESET_B(net689),
    .D(net3172),
    .Q(\u_inv.f_next[249] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _35261_ (.RESET_B(net687),
    .D(net3181),
    .Q(\u_inv.f_next[250] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _35262_ (.RESET_B(net685),
    .D(_01555_),
    .Q(\u_inv.f_next[251] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _35263_ (.RESET_B(net683),
    .D(net2245),
    .Q(\u_inv.f_next[252] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _35264_ (.RESET_B(net681),
    .D(_01557_),
    .Q(\u_inv.f_next[253] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _35265_ (.RESET_B(net679),
    .D(_01558_),
    .Q(\u_inv.f_next[254] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _35266_ (.RESET_B(net677),
    .D(net2531),
    .Q(\u_inv.f_next[255] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _35267_ (.RESET_B(net4814),
    .D(_01560_),
    .Q(\u_inv.state[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _35268_ (.RESET_B(net4814),
    .D(_01561_),
    .Q(\u_inv.state[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _35269_ (.RESET_B(net4818),
    .D(net1492),
    .Q(\u_inv.input_reg[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _35270_ (.RESET_B(net4820),
    .D(_01563_),
    .Q(\u_inv.input_reg[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _35271_ (.RESET_B(net4820),
    .D(net1622),
    .Q(\u_inv.input_reg[2] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _35272_ (.RESET_B(net4824),
    .D(net1268),
    .Q(\u_inv.input_reg[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35273_ (.RESET_B(net4824),
    .D(_01566_),
    .Q(\u_inv.input_reg[4] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35274_ (.RESET_B(net4824),
    .D(net1301),
    .Q(\u_inv.input_reg[5] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _35275_ (.RESET_B(net4825),
    .D(net1191),
    .Q(\u_inv.input_reg[6] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35276_ (.RESET_B(net4825),
    .D(_01569_),
    .Q(\u_inv.input_reg[7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35277_ (.RESET_B(net4822),
    .D(_01570_),
    .Q(\u_inv.input_reg[8] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35278_ (.RESET_B(net4822),
    .D(_01571_),
    .Q(\u_inv.input_reg[9] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35279_ (.RESET_B(net4823),
    .D(_01572_),
    .Q(\u_inv.input_reg[10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35280_ (.RESET_B(net4825),
    .D(_01573_),
    .Q(\u_inv.input_reg[11] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _35281_ (.RESET_B(net4837),
    .D(_01574_),
    .Q(\u_inv.input_reg[12] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _35282_ (.RESET_B(net4837),
    .D(_01575_),
    .Q(\u_inv.input_reg[13] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _35283_ (.RESET_B(net4836),
    .D(net1812),
    .Q(\u_inv.input_reg[14] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _35284_ (.RESET_B(net4837),
    .D(net1786),
    .Q(\u_inv.input_reg[15] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _35285_ (.RESET_B(net4836),
    .D(net1684),
    .Q(\u_inv.input_reg[16] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _35286_ (.RESET_B(net4836),
    .D(net1846),
    .Q(\u_inv.input_reg[17] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _35287_ (.RESET_B(net4836),
    .D(net1620),
    .Q(\u_inv.input_reg[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _35288_ (.RESET_B(net4837),
    .D(net1856),
    .Q(\u_inv.input_reg[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _35289_ (.RESET_B(net4842),
    .D(_01582_),
    .Q(\u_inv.input_reg[20] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _35290_ (.RESET_B(net4842),
    .D(_01583_),
    .Q(\u_inv.input_reg[21] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _35291_ (.RESET_B(net4838),
    .D(_01584_),
    .Q(\u_inv.input_reg[22] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35292_ (.RESET_B(net4842),
    .D(_01585_),
    .Q(\u_inv.input_reg[23] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35293_ (.RESET_B(net4839),
    .D(_01586_),
    .Q(\u_inv.input_reg[24] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35294_ (.RESET_B(net4842),
    .D(_01587_),
    .Q(\u_inv.input_reg[25] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35295_ (.RESET_B(net4839),
    .D(_01588_),
    .Q(\u_inv.input_reg[26] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35296_ (.RESET_B(net4842),
    .D(_01589_),
    .Q(\u_inv.input_reg[27] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35297_ (.RESET_B(net4842),
    .D(_01590_),
    .Q(\u_inv.input_reg[28] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _35298_ (.RESET_B(net4839),
    .D(_01591_),
    .Q(\u_inv.input_reg[29] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35299_ (.RESET_B(net4854),
    .D(_01592_),
    .Q(\u_inv.input_reg[30] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35300_ (.RESET_B(net4855),
    .D(_01593_),
    .Q(\u_inv.input_reg[31] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35301_ (.RESET_B(net4854),
    .D(_01594_),
    .Q(\u_inv.input_reg[32] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35302_ (.RESET_B(net4854),
    .D(_01595_),
    .Q(\u_inv.input_reg[33] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _35303_ (.RESET_B(net4851),
    .D(_01596_),
    .Q(\u_inv.input_reg[34] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _35304_ (.RESET_B(net4851),
    .D(_01597_),
    .Q(\u_inv.input_reg[35] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _35305_ (.RESET_B(net4851),
    .D(_01598_),
    .Q(\u_inv.input_reg[36] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _35306_ (.RESET_B(net4855),
    .D(_01599_),
    .Q(\u_inv.input_reg[37] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _35307_ (.RESET_B(net4851),
    .D(_01600_),
    .Q(\u_inv.input_reg[38] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _35308_ (.RESET_B(net4855),
    .D(_01601_),
    .Q(\u_inv.input_reg[39] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _35309_ (.RESET_B(net4856),
    .D(_01602_),
    .Q(\u_inv.input_reg[40] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _35310_ (.RESET_B(net4856),
    .D(_01603_),
    .Q(\u_inv.input_reg[41] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _35311_ (.RESET_B(net4855),
    .D(_01604_),
    .Q(\u_inv.input_reg[42] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _35312_ (.RESET_B(net4856),
    .D(_01605_),
    .Q(\u_inv.input_reg[43] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _35313_ (.RESET_B(net4858),
    .D(_01606_),
    .Q(\u_inv.input_reg[44] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _35314_ (.RESET_B(net4858),
    .D(net1979),
    .Q(\u_inv.input_reg[45] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _35315_ (.RESET_B(net4857),
    .D(net1721),
    .Q(\u_inv.input_reg[46] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _35316_ (.RESET_B(net4858),
    .D(_01609_),
    .Q(\u_inv.input_reg[47] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _35317_ (.RESET_B(net4870),
    .D(net1719),
    .Q(\u_inv.input_reg[48] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _35318_ (.RESET_B(net4870),
    .D(_01611_),
    .Q(\u_inv.input_reg[49] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _35319_ (.RESET_B(net4870),
    .D(_01612_),
    .Q(\u_inv.input_reg[50] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _35320_ (.RESET_B(net4871),
    .D(_01613_),
    .Q(\u_inv.input_reg[51] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _35321_ (.RESET_B(net4870),
    .D(_01614_),
    .Q(\u_inv.input_reg[52] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35322_ (.RESET_B(net4870),
    .D(_01615_),
    .Q(\u_inv.input_reg[53] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _35323_ (.RESET_B(net4873),
    .D(_01616_),
    .Q(\u_inv.input_reg[54] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _35324_ (.RESET_B(net4871),
    .D(_01617_),
    .Q(\u_inv.input_reg[55] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35325_ (.RESET_B(net4874),
    .D(_01618_),
    .Q(\u_inv.input_reg[56] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35326_ (.RESET_B(net4874),
    .D(_01619_),
    .Q(\u_inv.input_reg[57] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35327_ (.RESET_B(net4875),
    .D(_01620_),
    .Q(\u_inv.input_reg[58] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _35328_ (.RESET_B(net4875),
    .D(_01621_),
    .Q(\u_inv.input_reg[59] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35329_ (.RESET_B(net4875),
    .D(_01622_),
    .Q(\u_inv.input_reg[60] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _35330_ (.RESET_B(net4875),
    .D(net1765),
    .Q(\u_inv.input_reg[61] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35331_ (.RESET_B(net4873),
    .D(_01624_),
    .Q(\u_inv.input_reg[62] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _35332_ (.RESET_B(net4875),
    .D(_01625_),
    .Q(\u_inv.input_reg[63] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _35333_ (.RESET_B(net4875),
    .D(_01626_),
    .Q(\u_inv.input_reg[64] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _35334_ (.RESET_B(net4875),
    .D(_01627_),
    .Q(\u_inv.input_reg[65] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _35335_ (.RESET_B(net4885),
    .D(_01628_),
    .Q(\u_inv.input_reg[66] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _35336_ (.RESET_B(net4888),
    .D(_01629_),
    .Q(\u_inv.input_reg[67] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _35337_ (.RESET_B(net4885),
    .D(_01630_),
    .Q(\u_inv.input_reg[68] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _35338_ (.RESET_B(net4885),
    .D(_01631_),
    .Q(\u_inv.input_reg[69] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _35339_ (.RESET_B(net4887),
    .D(_01632_),
    .Q(\u_inv.input_reg[70] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _35340_ (.RESET_B(net4885),
    .D(_01633_),
    .Q(\u_inv.input_reg[71] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _35341_ (.RESET_B(net4886),
    .D(_01634_),
    .Q(\u_inv.input_reg[72] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _35342_ (.RESET_B(net4887),
    .D(_01635_),
    .Q(\u_inv.input_reg[73] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _35343_ (.RESET_B(net4892),
    .D(_01636_),
    .Q(\u_inv.input_reg[74] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35344_ (.RESET_B(net4887),
    .D(_01637_),
    .Q(\u_inv.input_reg[75] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _35345_ (.RESET_B(net4887),
    .D(_01638_),
    .Q(\u_inv.input_reg[76] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _35346_ (.RESET_B(net4889),
    .D(_01639_),
    .Q(\u_inv.input_reg[77] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35347_ (.RESET_B(net4887),
    .D(_01640_),
    .Q(\u_inv.input_reg[78] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35348_ (.RESET_B(net4890),
    .D(_01641_),
    .Q(\u_inv.input_reg[79] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35349_ (.RESET_B(net4890),
    .D(_01642_),
    .Q(\u_inv.input_reg[80] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35350_ (.RESET_B(net4889),
    .D(_01643_),
    .Q(\u_inv.input_reg[81] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35351_ (.RESET_B(net4892),
    .D(_01644_),
    .Q(\u_inv.input_reg[82] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35352_ (.RESET_B(net4890),
    .D(_01645_),
    .Q(\u_inv.input_reg[83] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35353_ (.RESET_B(net4890),
    .D(_01646_),
    .Q(\u_inv.input_reg[84] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _35354_ (.RESET_B(net4891),
    .D(_01647_),
    .Q(\u_inv.input_reg[85] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35355_ (.RESET_B(net4892),
    .D(_01648_),
    .Q(\u_inv.input_reg[86] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35356_ (.RESET_B(net4892),
    .D(_01649_),
    .Q(\u_inv.input_reg[87] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35357_ (.RESET_B(net4897),
    .D(_01650_),
    .Q(\u_inv.input_reg[88] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35358_ (.RESET_B(net4897),
    .D(_01651_),
    .Q(\u_inv.input_reg[89] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _35359_ (.RESET_B(net4898),
    .D(_01652_),
    .Q(\u_inv.input_reg[90] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35360_ (.RESET_B(net4897),
    .D(_01653_),
    .Q(\u_inv.input_reg[91] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35361_ (.RESET_B(net4897),
    .D(_01654_),
    .Q(\u_inv.input_reg[92] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _35362_ (.RESET_B(net4897),
    .D(_01655_),
    .Q(\u_inv.input_reg[93] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35363_ (.RESET_B(net4896),
    .D(_01656_),
    .Q(\u_inv.input_reg[94] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35364_ (.RESET_B(net4897),
    .D(net1638),
    .Q(\u_inv.input_reg[95] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35365_ (.RESET_B(net4910),
    .D(_01658_),
    .Q(\u_inv.input_reg[96] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _35366_ (.RESET_B(net4901),
    .D(_01659_),
    .Q(\u_inv.input_reg[97] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35367_ (.RESET_B(net4910),
    .D(_01660_),
    .Q(\u_inv.input_reg[98] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _35368_ (.RESET_B(net4904),
    .D(_01661_),
    .Q(\u_inv.input_reg[99] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35369_ (.RESET_B(net4910),
    .D(_01662_),
    .Q(\u_inv.input_reg[100] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35370_ (.RESET_B(net4911),
    .D(net1877),
    .Q(\u_inv.input_reg[101] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _35371_ (.RESET_B(net4910),
    .D(_01664_),
    .Q(\u_inv.input_reg[102] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _35372_ (.RESET_B(net4910),
    .D(_01665_),
    .Q(\u_inv.input_reg[103] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35373_ (.RESET_B(net4918),
    .D(_01666_),
    .Q(\u_inv.input_reg[104] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35374_ (.RESET_B(net4918),
    .D(_01667_),
    .Q(\u_inv.input_reg[105] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35375_ (.RESET_B(net4918),
    .D(_01668_),
    .Q(\u_inv.input_reg[106] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _35376_ (.RESET_B(net4916),
    .D(_01669_),
    .Q(\u_inv.input_reg[107] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _35377_ (.RESET_B(net4939),
    .D(_01670_),
    .Q(\u_inv.input_reg[108] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _35378_ (.RESET_B(net4942),
    .D(_01671_),
    .Q(\u_inv.input_reg[109] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _35379_ (.RESET_B(net4916),
    .D(_01672_),
    .Q(\u_inv.input_reg[110] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _35380_ (.RESET_B(net4918),
    .D(_01673_),
    .Q(\u_inv.input_reg[111] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _35381_ (.RESET_B(net4918),
    .D(_01674_),
    .Q(\u_inv.input_reg[112] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _35382_ (.RESET_B(net4945),
    .D(_01675_),
    .Q(\u_inv.input_reg[113] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _35383_ (.RESET_B(net4917),
    .D(_01676_),
    .Q(\u_inv.input_reg[114] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _35384_ (.RESET_B(net4948),
    .D(_01677_),
    .Q(\u_inv.input_reg[115] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35385_ (.RESET_B(net4948),
    .D(_01678_),
    .Q(\u_inv.input_reg[116] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35386_ (.RESET_B(net4947),
    .D(_01679_),
    .Q(\u_inv.input_reg[117] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35387_ (.RESET_B(net4948),
    .D(_01680_),
    .Q(\u_inv.input_reg[118] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35388_ (.RESET_B(net4948),
    .D(_01681_),
    .Q(\u_inv.input_reg[119] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _35389_ (.RESET_B(net4945),
    .D(_01682_),
    .Q(\u_inv.input_reg[120] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _35390_ (.RESET_B(net4945),
    .D(_01683_),
    .Q(\u_inv.input_reg[121] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35391_ (.RESET_B(net4945),
    .D(_01684_),
    .Q(\u_inv.input_reg[122] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _35392_ (.RESET_B(net4945),
    .D(_01685_),
    .Q(\u_inv.input_reg[123] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _35393_ (.RESET_B(net4947),
    .D(_01686_),
    .Q(\u_inv.input_reg[124] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _35394_ (.RESET_B(net4945),
    .D(_01687_),
    .Q(\u_inv.input_reg[125] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _35395_ (.RESET_B(net4947),
    .D(_01688_),
    .Q(\u_inv.input_reg[126] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35396_ (.RESET_B(net4946),
    .D(_01689_),
    .Q(\u_inv.input_reg[127] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _35397_ (.RESET_B(net4934),
    .D(_01690_),
    .Q(\u_inv.input_reg[128] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _35398_ (.RESET_B(net4934),
    .D(_01691_),
    .Q(\u_inv.input_reg[129] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _35399_ (.RESET_B(net4933),
    .D(_01692_),
    .Q(\u_inv.input_reg[130] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _35400_ (.RESET_B(net4933),
    .D(_01693_),
    .Q(\u_inv.input_reg[131] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _35401_ (.RESET_B(net4928),
    .D(_01694_),
    .Q(\u_inv.input_reg[132] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _35402_ (.RESET_B(net4931),
    .D(_01695_),
    .Q(\u_inv.input_reg[133] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _35403_ (.RESET_B(net4928),
    .D(_01696_),
    .Q(\u_inv.input_reg[134] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _35404_ (.RESET_B(net4931),
    .D(_01697_),
    .Q(\u_inv.input_reg[135] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _35405_ (.RESET_B(net4931),
    .D(_01698_),
    .Q(\u_inv.input_reg[136] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _35406_ (.RESET_B(net4932),
    .D(net1752),
    .Q(\u_inv.input_reg[137] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _35407_ (.RESET_B(net4931),
    .D(_01700_),
    .Q(\u_inv.input_reg[138] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _35408_ (.RESET_B(net4932),
    .D(_01701_),
    .Q(\u_inv.input_reg[139] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _35409_ (.RESET_B(net4931),
    .D(_01702_),
    .Q(\u_inv.input_reg[140] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _35410_ (.RESET_B(net4932),
    .D(_01703_),
    .Q(\u_inv.input_reg[141] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _35411_ (.RESET_B(net4932),
    .D(_01704_),
    .Q(\u_inv.input_reg[142] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _35412_ (.RESET_B(net4931),
    .D(_01705_),
    .Q(\u_inv.input_reg[143] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _35413_ (.RESET_B(net4931),
    .D(_01706_),
    .Q(\u_inv.input_reg[144] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _35414_ (.RESET_B(net4935),
    .D(_01707_),
    .Q(\u_inv.input_reg[145] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _35415_ (.RESET_B(net4935),
    .D(_01708_),
    .Q(\u_inv.input_reg[146] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _35416_ (.RESET_B(net4935),
    .D(_01709_),
    .Q(\u_inv.input_reg[147] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _35417_ (.RESET_B(net4935),
    .D(_01710_),
    .Q(\u_inv.input_reg[148] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _35418_ (.RESET_B(net4936),
    .D(_01711_),
    .Q(\u_inv.input_reg[149] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _35419_ (.RESET_B(net4935),
    .D(_01712_),
    .Q(\u_inv.input_reg[150] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _35420_ (.RESET_B(net4935),
    .D(_01713_),
    .Q(\u_inv.input_reg[151] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _35421_ (.RESET_B(net4936),
    .D(_01714_),
    .Q(\u_inv.input_reg[152] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _35422_ (.RESET_B(net4935),
    .D(net1820),
    .Q(\u_inv.input_reg[153] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _35423_ (.RESET_B(net4947),
    .D(_01716_),
    .Q(\u_inv.input_reg[154] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _35424_ (.RESET_B(net4947),
    .D(_01717_),
    .Q(\u_inv.input_reg[155] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _35425_ (.RESET_B(net4935),
    .D(net1832),
    .Q(\u_inv.input_reg[156] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _35426_ (.RESET_B(net4946),
    .D(_01719_),
    .Q(\u_inv.input_reg[157] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _35427_ (.RESET_B(net4947),
    .D(_01720_),
    .Q(\u_inv.input_reg[158] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _35428_ (.RESET_B(net4946),
    .D(_01721_),
    .Q(\u_inv.input_reg[159] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _35429_ (.RESET_B(net4943),
    .D(_01722_),
    .Q(\u_inv.input_reg[160] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _35430_ (.RESET_B(net4943),
    .D(_01723_),
    .Q(\u_inv.input_reg[161] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _35431_ (.RESET_B(net4942),
    .D(_01724_),
    .Q(\u_inv.input_reg[162] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _35432_ (.RESET_B(net4942),
    .D(_01725_),
    .Q(\u_inv.input_reg[163] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _35433_ (.RESET_B(net4940),
    .D(_01726_),
    .Q(\u_inv.input_reg[164] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _35434_ (.RESET_B(net4942),
    .D(_01727_),
    .Q(\u_inv.input_reg[165] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _35435_ (.RESET_B(net4942),
    .D(_01728_),
    .Q(\u_inv.input_reg[166] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _35436_ (.RESET_B(net4939),
    .D(_01729_),
    .Q(\u_inv.input_reg[167] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _35437_ (.RESET_B(net4939),
    .D(_01730_),
    .Q(\u_inv.input_reg[168] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _35438_ (.RESET_B(net4916),
    .D(_01731_),
    .Q(\u_inv.input_reg[169] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _35439_ (.RESET_B(net4918),
    .D(_01732_),
    .Q(\u_inv.input_reg[170] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _35440_ (.RESET_B(net4914),
    .D(_01733_),
    .Q(\u_inv.input_reg[171] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35441_ (.RESET_B(net4915),
    .D(_01734_),
    .Q(\u_inv.input_reg[172] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _35442_ (.RESET_B(net4914),
    .D(_01735_),
    .Q(\u_inv.input_reg[173] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35443_ (.RESET_B(net4914),
    .D(_01736_),
    .Q(\u_inv.input_reg[174] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35444_ (.RESET_B(net4911),
    .D(_01737_),
    .Q(\u_inv.input_reg[175] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _35445_ (.RESET_B(net4904),
    .D(_01738_),
    .Q(\u_inv.input_reg[176] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _35446_ (.RESET_B(net4919),
    .D(_01739_),
    .Q(\u_inv.input_reg[177] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _35447_ (.RESET_B(net4910),
    .D(_01740_),
    .Q(\u_inv.input_reg[178] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _35448_ (.RESET_B(net4904),
    .D(_01741_),
    .Q(\u_inv.input_reg[179] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35449_ (.RESET_B(net4904),
    .D(_01742_),
    .Q(\u_inv.input_reg[180] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35450_ (.RESET_B(net4901),
    .D(_01743_),
    .Q(\u_inv.input_reg[181] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35451_ (.RESET_B(net4906),
    .D(_01744_),
    .Q(\u_inv.input_reg[182] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _35452_ (.RESET_B(net4903),
    .D(_01745_),
    .Q(\u_inv.input_reg[183] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _35453_ (.RESET_B(net4901),
    .D(net1892),
    .Q(\u_inv.input_reg[184] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _35454_ (.RESET_B(net4901),
    .D(net1791),
    .Q(\u_inv.input_reg[185] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35455_ (.RESET_B(net4899),
    .D(_01748_),
    .Q(\u_inv.input_reg[186] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _35456_ (.RESET_B(net4899),
    .D(_01749_),
    .Q(\u_inv.input_reg[187] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _35457_ (.RESET_B(net4898),
    .D(_01750_),
    .Q(\u_inv.input_reg[188] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35458_ (.RESET_B(net4897),
    .D(_01751_),
    .Q(\u_inv.input_reg[189] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _35459_ (.RESET_B(net4899),
    .D(_01752_),
    .Q(\u_inv.input_reg[190] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35460_ (.RESET_B(net4893),
    .D(_01753_),
    .Q(\u_inv.input_reg[191] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _35461_ (.RESET_B(net4872),
    .D(_01754_),
    .Q(\u_inv.input_reg[192] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _35462_ (.RESET_B(net4872),
    .D(_01755_),
    .Q(\u_inv.input_reg[193] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _35463_ (.RESET_B(net4866),
    .D(_01756_),
    .Q(\u_inv.input_reg[194] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _35464_ (.RESET_B(net4866),
    .D(_01757_),
    .Q(\u_inv.input_reg[195] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _35465_ (.RESET_B(net4866),
    .D(_01758_),
    .Q(\u_inv.input_reg[196] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _35466_ (.RESET_B(net4863),
    .D(net1834),
    .Q(\u_inv.input_reg[197] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _35467_ (.RESET_B(net4863),
    .D(net1840),
    .Q(\u_inv.input_reg[198] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _35468_ (.RESET_B(net4871),
    .D(net1916),
    .Q(\u_inv.input_reg[199] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _35469_ (.RESET_B(net4863),
    .D(_01762_),
    .Q(\u_inv.input_reg[200] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _35470_ (.RESET_B(net4862),
    .D(_01763_),
    .Q(\u_inv.input_reg[201] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _35471_ (.RESET_B(net4862),
    .D(_01764_),
    .Q(\u_inv.input_reg[202] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _35472_ (.RESET_B(net4863),
    .D(_01765_),
    .Q(\u_inv.input_reg[203] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _35473_ (.RESET_B(net4863),
    .D(_01766_),
    .Q(\u_inv.input_reg[204] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _35474_ (.RESET_B(net4862),
    .D(_01767_),
    .Q(\u_inv.input_reg[205] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _35475_ (.RESET_B(net4862),
    .D(net1782),
    .Q(\u_inv.input_reg[206] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _35476_ (.RESET_B(net4848),
    .D(_01769_),
    .Q(\u_inv.input_reg[207] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _35477_ (.RESET_B(net4847),
    .D(_01770_),
    .Q(\u_inv.input_reg[208] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _35478_ (.RESET_B(net4847),
    .D(_01771_),
    .Q(\u_inv.input_reg[209] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _35479_ (.RESET_B(net4849),
    .D(_01772_),
    .Q(\u_inv.input_reg[210] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _35480_ (.RESET_B(net4848),
    .D(_01773_),
    .Q(\u_inv.input_reg[211] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _35481_ (.RESET_B(net4848),
    .D(_01774_),
    .Q(\u_inv.input_reg[212] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _35482_ (.RESET_B(net4848),
    .D(_01775_),
    .Q(\u_inv.input_reg[213] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _35483_ (.RESET_B(net4848),
    .D(_01776_),
    .Q(\u_inv.input_reg[214] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _35484_ (.RESET_B(net4846),
    .D(_01777_),
    .Q(\u_inv.input_reg[215] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _35485_ (.RESET_B(net4846),
    .D(_01778_),
    .Q(\u_inv.input_reg[216] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _35486_ (.RESET_B(net4845),
    .D(_01779_),
    .Q(\u_inv.input_reg[217] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _35487_ (.RESET_B(net4845),
    .D(_01780_),
    .Q(\u_inv.input_reg[218] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _35488_ (.RESET_B(net4845),
    .D(_01781_),
    .Q(\u_inv.input_reg[219] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _35489_ (.RESET_B(net4845),
    .D(_01782_),
    .Q(\u_inv.input_reg[220] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _35490_ (.RESET_B(net4845),
    .D(net2082),
    .Q(\u_inv.input_reg[221] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _35491_ (.RESET_B(net4833),
    .D(_01784_),
    .Q(\u_inv.input_reg[222] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35492_ (.RESET_B(net4833),
    .D(_01785_),
    .Q(\u_inv.input_reg[223] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35493_ (.RESET_B(net4832),
    .D(net1836),
    .Q(\u_inv.input_reg[224] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _35494_ (.RESET_B(net4832),
    .D(_01787_),
    .Q(\u_inv.input_reg[225] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35495_ (.RESET_B(net4832),
    .D(_01788_),
    .Q(\u_inv.input_reg[226] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35496_ (.RESET_B(net4832),
    .D(_01789_),
    .Q(\u_inv.input_reg[227] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35497_ (.RESET_B(net4832),
    .D(_01790_),
    .Q(\u_inv.input_reg[228] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35498_ (.RESET_B(net4831),
    .D(_01791_),
    .Q(\u_inv.input_reg[229] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35499_ (.RESET_B(net4830),
    .D(_01792_),
    .Q(\u_inv.input_reg[230] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _35500_ (.RESET_B(net4831),
    .D(_01793_),
    .Q(\u_inv.input_reg[231] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35501_ (.RESET_B(net4830),
    .D(_01794_),
    .Q(\u_inv.input_reg[232] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35502_ (.RESET_B(net4829),
    .D(_01795_),
    .Q(\u_inv.input_reg[233] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35503_ (.RESET_B(net4829),
    .D(_01796_),
    .Q(\u_inv.input_reg[234] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _35504_ (.RESET_B(net4829),
    .D(_01797_),
    .Q(\u_inv.input_reg[235] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35505_ (.RESET_B(net4829),
    .D(_01798_),
    .Q(\u_inv.input_reg[236] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _35506_ (.RESET_B(net4831),
    .D(_01799_),
    .Q(\u_inv.input_reg[237] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _35507_ (.RESET_B(net4829),
    .D(_01800_),
    .Q(\u_inv.input_reg[238] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _35508_ (.RESET_B(net4809),
    .D(_01801_),
    .Q(\u_inv.input_reg[239] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _35509_ (.RESET_B(net4810),
    .D(net2005),
    .Q(\u_inv.input_reg[240] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _35510_ (.RESET_B(net4807),
    .D(_01803_),
    .Q(\u_inv.input_reg[241] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _35511_ (.RESET_B(net4807),
    .D(_01804_),
    .Q(\u_inv.input_reg[242] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _35512_ (.RESET_B(net4807),
    .D(net1933),
    .Q(\u_inv.input_reg[243] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _35513_ (.RESET_B(net4807),
    .D(net1789),
    .Q(\u_inv.input_reg[244] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _35514_ (.RESET_B(net4807),
    .D(_01807_),
    .Q(\u_inv.input_reg[245] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _35515_ (.RESET_B(net4807),
    .D(_01808_),
    .Q(\u_inv.input_reg[246] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _35516_ (.RESET_B(net4807),
    .D(_01809_),
    .Q(\u_inv.input_reg[247] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _35517_ (.RESET_B(net4817),
    .D(_01810_),
    .Q(\u_inv.input_reg[248] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _35518_ (.RESET_B(net4814),
    .D(_01811_),
    .Q(\u_inv.input_reg[249] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _35519_ (.RESET_B(net4817),
    .D(_01812_),
    .Q(\u_inv.input_reg[250] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _35520_ (.RESET_B(net4814),
    .D(_01813_),
    .Q(\u_inv.input_reg[251] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _35521_ (.RESET_B(net4813),
    .D(_01814_),
    .Q(\u_inv.input_reg[252] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _35522_ (.RESET_B(net4813),
    .D(_01815_),
    .Q(\u_inv.input_reg[253] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _35523_ (.RESET_B(net4813),
    .D(_01816_),
    .Q(\u_inv.input_reg[254] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _35524_ (.RESET_B(net4813),
    .D(_01817_),
    .Q(\u_inv.input_reg[255] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _35525_ (.RESET_B(net417),
    .D(_01818_),
    .Q(\u_inv.delta_reg[0] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _35526_ (.RESET_B(net413),
    .D(net1604),
    .Q(\u_inv.delta_reg[1] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _35527_ (.RESET_B(net409),
    .D(_01820_),
    .Q(\u_inv.delta_reg[2] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _35528_ (.RESET_B(net406),
    .D(_01821_),
    .Q(\u_inv.delta_reg[3] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _35529_ (.RESET_B(net402),
    .D(_01822_),
    .Q(\u_inv.delta_reg[4] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _35530_ (.RESET_B(net398),
    .D(_01823_),
    .Q(\u_inv.delta_reg[5] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _35531_ (.RESET_B(net411),
    .D(net1522),
    .Q(\u_inv.delta_reg[6] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _35532_ (.RESET_B(net404),
    .D(_01825_),
    .Q(\u_inv.delta_reg[7] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _35533_ (.RESET_B(net415),
    .D(net1874),
    .Q(\u_inv.delta_reg[8] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _35534_ (.RESET_B(net400),
    .D(_01827_),
    .Q(\u_inv.delta_reg[9] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_tiehi _34293__24 (.L_HI(net24));
 sg13g2_tiehi _35073__25 (.L_HI(net25));
 sg13g2_tiehi _34292__26 (.L_HI(net26));
 sg13g2_tiehi _35072__27 (.L_HI(net27));
 sg13g2_tiehi _34291__28 (.L_HI(net28));
 sg13g2_tiehi _35071__29 (.L_HI(net29));
 sg13g2_tiehi _34290__30 (.L_HI(net30));
 sg13g2_tiehi _35070__31 (.L_HI(net31));
 sg13g2_tiehi _34289__32 (.L_HI(net32));
 sg13g2_tiehi _35069__33 (.L_HI(net33));
 sg13g2_tiehi _34288__34 (.L_HI(net34));
 sg13g2_tiehi _35068__35 (.L_HI(net35));
 sg13g2_tiehi _34287__36 (.L_HI(net36));
 sg13g2_tiehi _35067__37 (.L_HI(net37));
 sg13g2_tiehi _34286__38 (.L_HI(net38));
 sg13g2_tiehi _35066__39 (.L_HI(net39));
 sg13g2_tiehi _34285__40 (.L_HI(net40));
 sg13g2_tiehi _35065__41 (.L_HI(net41));
 sg13g2_tiehi _34284__42 (.L_HI(net42));
 sg13g2_tiehi _35064__43 (.L_HI(net43));
 sg13g2_tiehi _34283__44 (.L_HI(net44));
 sg13g2_tiehi _35063__45 (.L_HI(net45));
 sg13g2_tiehi _34282__46 (.L_HI(net46));
 sg13g2_tiehi _35062__47 (.L_HI(net47));
 sg13g2_tiehi _34281__48 (.L_HI(net48));
 sg13g2_tiehi _35061__49 (.L_HI(net49));
 sg13g2_tiehi _34280__50 (.L_HI(net50));
 sg13g2_tiehi _35060__51 (.L_HI(net51));
 sg13g2_tiehi _34279__52 (.L_HI(net52));
 sg13g2_tiehi _35059__53 (.L_HI(net53));
 sg13g2_tiehi _34278__54 (.L_HI(net54));
 sg13g2_tiehi _35058__55 (.L_HI(net55));
 sg13g2_tiehi _34277__56 (.L_HI(net56));
 sg13g2_tiehi _35057__57 (.L_HI(net57));
 sg13g2_tiehi _34276__58 (.L_HI(net58));
 sg13g2_tiehi _35056__59 (.L_HI(net59));
 sg13g2_tiehi _34275__60 (.L_HI(net60));
 sg13g2_tiehi _35055__61 (.L_HI(net61));
 sg13g2_tiehi _34274__62 (.L_HI(net62));
 sg13g2_tiehi _35054__63 (.L_HI(net63));
 sg13g2_tiehi _34273__64 (.L_HI(net64));
 sg13g2_tiehi _35053__65 (.L_HI(net65));
 sg13g2_tiehi _34272__66 (.L_HI(net66));
 sg13g2_tiehi _35052__67 (.L_HI(net67));
 sg13g2_tiehi _34271__68 (.L_HI(net68));
 sg13g2_tiehi _35051__69 (.L_HI(net69));
 sg13g2_tiehi _34270__70 (.L_HI(net70));
 sg13g2_tiehi _35050__71 (.L_HI(net71));
 sg13g2_tiehi _34269__72 (.L_HI(net72));
 sg13g2_tiehi _35049__73 (.L_HI(net73));
 sg13g2_tiehi _34268__74 (.L_HI(net74));
 sg13g2_tiehi _35048__75 (.L_HI(net75));
 sg13g2_tiehi _34267__76 (.L_HI(net76));
 sg13g2_tiehi _35047__77 (.L_HI(net77));
 sg13g2_tiehi _34266__78 (.L_HI(net78));
 sg13g2_tiehi _35046__79 (.L_HI(net79));
 sg13g2_tiehi _34265__80 (.L_HI(net80));
 sg13g2_tiehi _35045__81 (.L_HI(net81));
 sg13g2_tiehi _34264__82 (.L_HI(net82));
 sg13g2_tiehi _35044__83 (.L_HI(net83));
 sg13g2_tiehi _34263__84 (.L_HI(net84));
 sg13g2_tiehi _35043__85 (.L_HI(net85));
 sg13g2_tiehi _34262__86 (.L_HI(net86));
 sg13g2_tiehi _35042__87 (.L_HI(net87));
 sg13g2_tiehi _34261__88 (.L_HI(net88));
 sg13g2_tiehi _35041__89 (.L_HI(net89));
 sg13g2_tiehi _34260__90 (.L_HI(net90));
 sg13g2_tiehi _35040__91 (.L_HI(net91));
 sg13g2_tiehi _34259__92 (.L_HI(net92));
 sg13g2_tiehi _35039__93 (.L_HI(net93));
 sg13g2_tiehi _34258__94 (.L_HI(net94));
 sg13g2_tiehi _35038__95 (.L_HI(net95));
 sg13g2_tiehi _34257__96 (.L_HI(net96));
 sg13g2_tiehi _35037__97 (.L_HI(net97));
 sg13g2_tiehi _34256__98 (.L_HI(net98));
 sg13g2_tiehi _35036__99 (.L_HI(net99));
 sg13g2_tiehi _34255__100 (.L_HI(net100));
 sg13g2_tiehi _35035__101 (.L_HI(net101));
 sg13g2_tiehi _34254__102 (.L_HI(net102));
 sg13g2_tiehi _35034__103 (.L_HI(net103));
 sg13g2_tiehi _34253__104 (.L_HI(net104));
 sg13g2_tiehi _35033__105 (.L_HI(net105));
 sg13g2_tiehi _34252__106 (.L_HI(net106));
 sg13g2_tiehi _35032__107 (.L_HI(net107));
 sg13g2_tiehi _34251__108 (.L_HI(net108));
 sg13g2_tiehi _35031__109 (.L_HI(net109));
 sg13g2_tiehi _34250__110 (.L_HI(net110));
 sg13g2_tiehi _35030__111 (.L_HI(net111));
 sg13g2_tiehi _34249__112 (.L_HI(net112));
 sg13g2_tiehi _35029__113 (.L_HI(net113));
 sg13g2_tiehi _34248__114 (.L_HI(net114));
 sg13g2_tiehi _35028__115 (.L_HI(net115));
 sg13g2_tiehi _34247__116 (.L_HI(net116));
 sg13g2_tiehi _35027__117 (.L_HI(net117));
 sg13g2_tiehi _34246__118 (.L_HI(net118));
 sg13g2_tiehi _35026__119 (.L_HI(net119));
 sg13g2_tiehi _34245__120 (.L_HI(net120));
 sg13g2_tiehi _35025__121 (.L_HI(net121));
 sg13g2_tiehi _34244__122 (.L_HI(net122));
 sg13g2_tiehi _35024__123 (.L_HI(net123));
 sg13g2_tiehi _34243__124 (.L_HI(net124));
 sg13g2_tiehi _35023__125 (.L_HI(net125));
 sg13g2_tiehi _34242__126 (.L_HI(net126));
 sg13g2_tiehi _35022__127 (.L_HI(net127));
 sg13g2_tiehi _34241__128 (.L_HI(net128));
 sg13g2_tiehi _35021__129 (.L_HI(net129));
 sg13g2_tiehi _34240__130 (.L_HI(net130));
 sg13g2_tiehi _35020__131 (.L_HI(net131));
 sg13g2_tiehi _34239__132 (.L_HI(net132));
 sg13g2_tiehi _35019__133 (.L_HI(net133));
 sg13g2_tiehi _34238__134 (.L_HI(net134));
 sg13g2_tiehi _35018__135 (.L_HI(net135));
 sg13g2_tiehi _34237__136 (.L_HI(net136));
 sg13g2_tiehi _35017__137 (.L_HI(net137));
 sg13g2_tiehi _34236__138 (.L_HI(net138));
 sg13g2_tiehi _35016__139 (.L_HI(net139));
 sg13g2_tiehi _34235__140 (.L_HI(net140));
 sg13g2_tiehi _35015__141 (.L_HI(net141));
 sg13g2_tiehi _34234__142 (.L_HI(net142));
 sg13g2_tiehi _35014__143 (.L_HI(net143));
 sg13g2_tiehi _34233__144 (.L_HI(net144));
 sg13g2_tiehi _35013__145 (.L_HI(net145));
 sg13g2_tiehi _34232__146 (.L_HI(net146));
 sg13g2_tiehi _35012__147 (.L_HI(net147));
 sg13g2_tiehi _34231__148 (.L_HI(net148));
 sg13g2_tiehi _35011__149 (.L_HI(net149));
 sg13g2_tiehi _34230__150 (.L_HI(net150));
 sg13g2_tiehi _34229__151 (.L_HI(net151));
 sg13g2_tiehi _34228__152 (.L_HI(net152));
 sg13g2_tiehi _34227__153 (.L_HI(net153));
 sg13g2_tiehi _34226__154 (.L_HI(net154));
 sg13g2_tiehi _34225__155 (.L_HI(net155));
 sg13g2_tiehi _34224__156 (.L_HI(net156));
 sg13g2_tiehi _34223__157 (.L_HI(net157));
 sg13g2_tiehi _34222__158 (.L_HI(net158));
 sg13g2_tiehi _34221__159 (.L_HI(net159));
 sg13g2_tiehi _34220__160 (.L_HI(net160));
 sg13g2_tiehi _34219__161 (.L_HI(net161));
 sg13g2_tiehi _34218__162 (.L_HI(net162));
 sg13g2_tiehi _34217__163 (.L_HI(net163));
 sg13g2_tiehi _34216__164 (.L_HI(net164));
 sg13g2_tiehi _34215__165 (.L_HI(net165));
 sg13g2_tiehi _34214__166 (.L_HI(net166));
 sg13g2_tiehi _34213__167 (.L_HI(net167));
 sg13g2_tiehi _34212__168 (.L_HI(net168));
 sg13g2_tiehi _34211__169 (.L_HI(net169));
 sg13g2_tiehi _34210__170 (.L_HI(net170));
 sg13g2_tiehi _34209__171 (.L_HI(net171));
 sg13g2_tiehi _34208__172 (.L_HI(net172));
 sg13g2_tiehi _34207__173 (.L_HI(net173));
 sg13g2_tiehi _34206__174 (.L_HI(net174));
 sg13g2_tiehi _34205__175 (.L_HI(net175));
 sg13g2_tiehi _34204__176 (.L_HI(net176));
 sg13g2_tiehi _34203__177 (.L_HI(net177));
 sg13g2_tiehi _34202__178 (.L_HI(net178));
 sg13g2_tiehi _34201__179 (.L_HI(net179));
 sg13g2_tiehi _34200__180 (.L_HI(net180));
 sg13g2_tiehi _34199__181 (.L_HI(net181));
 sg13g2_tiehi _34198__182 (.L_HI(net182));
 sg13g2_tiehi _34197__183 (.L_HI(net183));
 sg13g2_tiehi _34196__184 (.L_HI(net184));
 sg13g2_tiehi _34195__185 (.L_HI(net185));
 sg13g2_tiehi _34194__186 (.L_HI(net186));
 sg13g2_tiehi _34193__187 (.L_HI(net187));
 sg13g2_tiehi _34192__188 (.L_HI(net188));
 sg13g2_tiehi _34191__189 (.L_HI(net189));
 sg13g2_tiehi _34190__190 (.L_HI(net190));
 sg13g2_tiehi _34189__191 (.L_HI(net191));
 sg13g2_tiehi _34188__192 (.L_HI(net192));
 sg13g2_tiehi _34187__193 (.L_HI(net193));
 sg13g2_tiehi _34186__194 (.L_HI(net194));
 sg13g2_tiehi _34185__195 (.L_HI(net195));
 sg13g2_tiehi _34184__196 (.L_HI(net196));
 sg13g2_tiehi _34183__197 (.L_HI(net197));
 sg13g2_tiehi _34182__198 (.L_HI(net198));
 sg13g2_tiehi _34181__199 (.L_HI(net199));
 sg13g2_tiehi _34180__200 (.L_HI(net200));
 sg13g2_tiehi _34179__201 (.L_HI(net201));
 sg13g2_tiehi _34178__202 (.L_HI(net202));
 sg13g2_tiehi _34177__203 (.L_HI(net203));
 sg13g2_tiehi _34176__204 (.L_HI(net204));
 sg13g2_tiehi _34175__205 (.L_HI(net205));
 sg13g2_tiehi _34174__206 (.L_HI(net206));
 sg13g2_tiehi _34173__207 (.L_HI(net207));
 sg13g2_tiehi _34172__208 (.L_HI(net208));
 sg13g2_tiehi _34171__209 (.L_HI(net209));
 sg13g2_tiehi _34170__210 (.L_HI(net210));
 sg13g2_tiehi _34169__211 (.L_HI(net211));
 sg13g2_tiehi _34168__212 (.L_HI(net212));
 sg13g2_tiehi _34167__213 (.L_HI(net213));
 sg13g2_tiehi _34166__214 (.L_HI(net214));
 sg13g2_tiehi _34165__215 (.L_HI(net215));
 sg13g2_tiehi _34164__216 (.L_HI(net216));
 sg13g2_tiehi _34163__217 (.L_HI(net217));
 sg13g2_tiehi _34162__218 (.L_HI(net218));
 sg13g2_tiehi _34161__219 (.L_HI(net219));
 sg13g2_tiehi _34160__220 (.L_HI(net220));
 sg13g2_tiehi _34159__221 (.L_HI(net221));
 sg13g2_tiehi _34158__222 (.L_HI(net222));
 sg13g2_tiehi _34157__223 (.L_HI(net223));
 sg13g2_tiehi _34156__224 (.L_HI(net224));
 sg13g2_tiehi _34155__225 (.L_HI(net225));
 sg13g2_tiehi _34154__226 (.L_HI(net226));
 sg13g2_tiehi _34153__227 (.L_HI(net227));
 sg13g2_tiehi _34152__228 (.L_HI(net228));
 sg13g2_tiehi _34151__229 (.L_HI(net229));
 sg13g2_tiehi _34150__230 (.L_HI(net230));
 sg13g2_tiehi _34149__231 (.L_HI(net231));
 sg13g2_tiehi _34148__232 (.L_HI(net232));
 sg13g2_tiehi _34147__233 (.L_HI(net233));
 sg13g2_tiehi _34146__234 (.L_HI(net234));
 sg13g2_tiehi _34145__235 (.L_HI(net235));
 sg13g2_tiehi _34144__236 (.L_HI(net236));
 sg13g2_tiehi _34143__237 (.L_HI(net237));
 sg13g2_tiehi _34142__238 (.L_HI(net238));
 sg13g2_tiehi _34141__239 (.L_HI(net239));
 sg13g2_tiehi _34140__240 (.L_HI(net240));
 sg13g2_tiehi _34139__241 (.L_HI(net241));
 sg13g2_tiehi _34138__242 (.L_HI(net242));
 sg13g2_tiehi _34137__243 (.L_HI(net243));
 sg13g2_tiehi _34136__244 (.L_HI(net244));
 sg13g2_tiehi _34135__245 (.L_HI(net245));
 sg13g2_tiehi _34134__246 (.L_HI(net246));
 sg13g2_tiehi _34133__247 (.L_HI(net247));
 sg13g2_tiehi _34132__248 (.L_HI(net248));
 sg13g2_tiehi _34131__249 (.L_HI(net249));
 sg13g2_tiehi _34130__250 (.L_HI(net250));
 sg13g2_tiehi _34129__251 (.L_HI(net251));
 sg13g2_tiehi _34128__252 (.L_HI(net252));
 sg13g2_tiehi _34127__253 (.L_HI(net253));
 sg13g2_tiehi _34126__254 (.L_HI(net254));
 sg13g2_tiehi _34125__255 (.L_HI(net255));
 sg13g2_tiehi _34124__256 (.L_HI(net256));
 sg13g2_tiehi _34123__257 (.L_HI(net257));
 sg13g2_tiehi _34122__258 (.L_HI(net258));
 sg13g2_tiehi _34121__259 (.L_HI(net259));
 sg13g2_tiehi _34120__260 (.L_HI(net260));
 sg13g2_tiehi _34119__261 (.L_HI(net261));
 sg13g2_tiehi _34118__262 (.L_HI(net262));
 sg13g2_tiehi _34117__263 (.L_HI(net263));
 sg13g2_tiehi _34116__264 (.L_HI(net264));
 sg13g2_tiehi _34115__265 (.L_HI(net265));
 sg13g2_tiehi _34114__266 (.L_HI(net266));
 sg13g2_tiehi _34113__267 (.L_HI(net267));
 sg13g2_tiehi _34112__268 (.L_HI(net268));
 sg13g2_tiehi _34111__269 (.L_HI(net269));
 sg13g2_tiehi _34110__270 (.L_HI(net270));
 sg13g2_tiehi _34109__271 (.L_HI(net271));
 sg13g2_tiehi _34108__272 (.L_HI(net272));
 sg13g2_tiehi _34107__273 (.L_HI(net273));
 sg13g2_tiehi _34106__274 (.L_HI(net274));
 sg13g2_tiehi _34105__275 (.L_HI(net275));
 sg13g2_tiehi _34104__276 (.L_HI(net276));
 sg13g2_tiehi _34103__277 (.L_HI(net277));
 sg13g2_tiehi _34102__278 (.L_HI(net278));
 sg13g2_tiehi _34101__279 (.L_HI(net279));
 sg13g2_tiehi _34100__280 (.L_HI(net280));
 sg13g2_tiehi _34099__281 (.L_HI(net281));
 sg13g2_tiehi _34098__282 (.L_HI(net282));
 sg13g2_tiehi _34097__283 (.L_HI(net283));
 sg13g2_tiehi _34096__284 (.L_HI(net284));
 sg13g2_tiehi _34095__285 (.L_HI(net285));
 sg13g2_tiehi _34094__286 (.L_HI(net286));
 sg13g2_tiehi _34093__287 (.L_HI(net287));
 sg13g2_tiehi _34092__288 (.L_HI(net288));
 sg13g2_tiehi _34091__289 (.L_HI(net289));
 sg13g2_tiehi _34090__290 (.L_HI(net290));
 sg13g2_tiehi _34089__291 (.L_HI(net291));
 sg13g2_tiehi _34088__292 (.L_HI(net292));
 sg13g2_tiehi _34087__293 (.L_HI(net293));
 sg13g2_tiehi _34086__294 (.L_HI(net294));
 sg13g2_tiehi _34085__295 (.L_HI(net295));
 sg13g2_tiehi _34084__296 (.L_HI(net296));
 sg13g2_tiehi _34083__297 (.L_HI(net297));
 sg13g2_tiehi _34082__298 (.L_HI(net298));
 sg13g2_tiehi _34081__299 (.L_HI(net299));
 sg13g2_tiehi _34080__300 (.L_HI(net300));
 sg13g2_tiehi _34079__301 (.L_HI(net301));
 sg13g2_tiehi _34078__302 (.L_HI(net302));
 sg13g2_tiehi _34077__303 (.L_HI(net303));
 sg13g2_tiehi _34076__304 (.L_HI(net304));
 sg13g2_tiehi _34075__305 (.L_HI(net305));
 sg13g2_tiehi _34074__306 (.L_HI(net306));
 sg13g2_tiehi _34073__307 (.L_HI(net307));
 sg13g2_tiehi _34072__308 (.L_HI(net308));
 sg13g2_tiehi _34071__309 (.L_HI(net309));
 sg13g2_tiehi _34070__310 (.L_HI(net310));
 sg13g2_tiehi _34069__311 (.L_HI(net311));
 sg13g2_tiehi _34068__312 (.L_HI(net312));
 sg13g2_tiehi _34067__313 (.L_HI(net313));
 sg13g2_tiehi _34066__314 (.L_HI(net314));
 sg13g2_tiehi _34065__315 (.L_HI(net315));
 sg13g2_tiehi _34064__316 (.L_HI(net316));
 sg13g2_tiehi _34063__317 (.L_HI(net317));
 sg13g2_tiehi _34062__318 (.L_HI(net318));
 sg13g2_tiehi _34061__319 (.L_HI(net319));
 sg13g2_tiehi _34060__320 (.L_HI(net320));
 sg13g2_tiehi _34059__321 (.L_HI(net321));
 sg13g2_tiehi _34058__322 (.L_HI(net322));
 sg13g2_tiehi _34057__323 (.L_HI(net323));
 sg13g2_tiehi _34056__324 (.L_HI(net324));
 sg13g2_tiehi _34055__325 (.L_HI(net325));
 sg13g2_tiehi _34054__326 (.L_HI(net326));
 sg13g2_tiehi _34053__327 (.L_HI(net327));
 sg13g2_tiehi _34052__328 (.L_HI(net328));
 sg13g2_tiehi _34051__329 (.L_HI(net329));
 sg13g2_tiehi _34050__330 (.L_HI(net330));
 sg13g2_tiehi _34049__331 (.L_HI(net331));
 sg13g2_tiehi _34048__332 (.L_HI(net332));
 sg13g2_tiehi _34047__333 (.L_HI(net333));
 sg13g2_tiehi _34046__334 (.L_HI(net334));
 sg13g2_tiehi _34045__335 (.L_HI(net335));
 sg13g2_tiehi _34044__336 (.L_HI(net336));
 sg13g2_tiehi _34043__337 (.L_HI(net337));
 sg13g2_tiehi _34042__338 (.L_HI(net338));
 sg13g2_tiehi _34041__339 (.L_HI(net339));
 sg13g2_tiehi _34040__340 (.L_HI(net340));
 sg13g2_tiehi _34039__341 (.L_HI(net341));
 sg13g2_tiehi _34038__342 (.L_HI(net342));
 sg13g2_tiehi _34037__343 (.L_HI(net343));
 sg13g2_tiehi _34036__344 (.L_HI(net344));
 sg13g2_tiehi _34035__345 (.L_HI(net345));
 sg13g2_tiehi _34034__346 (.L_HI(net346));
 sg13g2_tiehi _34033__347 (.L_HI(net347));
 sg13g2_tiehi _34032__348 (.L_HI(net348));
 sg13g2_tiehi _34031__349 (.L_HI(net349));
 sg13g2_tiehi _34030__350 (.L_HI(net350));
 sg13g2_tiehi _34029__351 (.L_HI(net351));
 sg13g2_tiehi _34028__352 (.L_HI(net352));
 sg13g2_tiehi _34027__353 (.L_HI(net353));
 sg13g2_tiehi _34026__354 (.L_HI(net354));
 sg13g2_tiehi _34025__355 (.L_HI(net355));
 sg13g2_tiehi _34024__356 (.L_HI(net356));
 sg13g2_tiehi _34023__357 (.L_HI(net357));
 sg13g2_tiehi _34022__358 (.L_HI(net358));
 sg13g2_tiehi _34021__359 (.L_HI(net359));
 sg13g2_tiehi _34020__360 (.L_HI(net360));
 sg13g2_tiehi _34019__361 (.L_HI(net361));
 sg13g2_tiehi _34018__362 (.L_HI(net362));
 sg13g2_tiehi _34017__363 (.L_HI(net363));
 sg13g2_tiehi _34016__364 (.L_HI(net364));
 sg13g2_tiehi _34015__365 (.L_HI(net365));
 sg13g2_tiehi _34014__366 (.L_HI(net366));
 sg13g2_tiehi _34013__367 (.L_HI(net367));
 sg13g2_tiehi _34012__368 (.L_HI(net368));
 sg13g2_tiehi _34011__369 (.L_HI(net369));
 sg13g2_tiehi _34010__370 (.L_HI(net370));
 sg13g2_tiehi _34009__371 (.L_HI(net371));
 sg13g2_tiehi _34008__372 (.L_HI(net372));
 sg13g2_tiehi _34007__373 (.L_HI(net373));
 sg13g2_tiehi _34006__374 (.L_HI(net374));
 sg13g2_tiehi _34005__375 (.L_HI(net375));
 sg13g2_tiehi _34004__376 (.L_HI(net376));
 sg13g2_tiehi _34003__377 (.L_HI(net377));
 sg13g2_tiehi _34002__378 (.L_HI(net378));
 sg13g2_tiehi _34001__379 (.L_HI(net379));
 sg13g2_tiehi _34000__380 (.L_HI(net380));
 sg13g2_tiehi _33999__381 (.L_HI(net381));
 sg13g2_tiehi _33998__382 (.L_HI(net382));
 sg13g2_tiehi _33997__383 (.L_HI(net383));
 sg13g2_tiehi _33996__384 (.L_HI(net384));
 sg13g2_tiehi _33995__385 (.L_HI(net385));
 sg13g2_tiehi _33994__386 (.L_HI(net386));
 sg13g2_tiehi _33993__387 (.L_HI(net387));
 sg13g2_tiehi _33992__388 (.L_HI(net388));
 sg13g2_tiehi _33991__389 (.L_HI(net389));
 sg13g2_tiehi _33990__390 (.L_HI(net390));
 sg13g2_tiehi _33989__391 (.L_HI(net391));
 sg13g2_tiehi _33988__392 (.L_HI(net392));
 sg13g2_tiehi _33987__393 (.L_HI(net393));
 sg13g2_tiehi _33986__394 (.L_HI(net394));
 sg13g2_tiehi _33985__395 (.L_HI(net395));
 sg13g2_tiehi _33984__396 (.L_HI(net396));
 sg13g2_tiehi _33715__397 (.L_HI(net397));
 sg13g2_tiehi _35530__398 (.L_HI(net398));
 sg13g2_tiehi _34754__399 (.L_HI(net399));
 sg13g2_tiehi _35534__400 (.L_HI(net400));
 sg13g2_tiehi _34753__401 (.L_HI(net401));
 sg13g2_tiehi _35529__402 (.L_HI(net402));
 sg13g2_tiehi _34752__403 (.L_HI(net403));
 sg13g2_tiehi _35532__404 (.L_HI(net404));
 sg13g2_tiehi _34751__405 (.L_HI(net405));
 sg13g2_tiehi _35528__406 (.L_HI(net406));
 sg13g2_tiehi _34750__407 (.L_HI(net407));
 sg13g2_tiehi _34749__408 (.L_HI(net408));
 sg13g2_tiehi _35527__409 (.L_HI(net409));
 sg13g2_tiehi _34748__410 (.L_HI(net410));
 sg13g2_tiehi _35531__411 (.L_HI(net411));
 sg13g2_tiehi _34747__412 (.L_HI(net412));
 sg13g2_tiehi _35526__413 (.L_HI(net413));
 sg13g2_tiehi _34746__414 (.L_HI(net414));
 sg13g2_tiehi _35533__415 (.L_HI(net415));
 sg13g2_tiehi _34745__416 (.L_HI(net416));
 sg13g2_tiehi _35525__417 (.L_HI(net417));
 sg13g2_tiehi _34744__418 (.L_HI(net418));
 sg13g2_tiehi _34743__419 (.L_HI(net419));
 sg13g2_tiehi _34742__420 (.L_HI(net420));
 sg13g2_tiehi _34741__421 (.L_HI(net421));
 sg13g2_tiehi _34740__422 (.L_HI(net422));
 sg13g2_tiehi _34739__423 (.L_HI(net423));
 sg13g2_tiehi _34738__424 (.L_HI(net424));
 sg13g2_tiehi _34737__425 (.L_HI(net425));
 sg13g2_tiehi _34736__426 (.L_HI(net426));
 sg13g2_tiehi _34735__427 (.L_HI(net427));
 sg13g2_tiehi _34734__428 (.L_HI(net428));
 sg13g2_tiehi _34733__429 (.L_HI(net429));
 sg13g2_tiehi _34732__430 (.L_HI(net430));
 sg13g2_tiehi _34731__431 (.L_HI(net431));
 sg13g2_tiehi _34730__432 (.L_HI(net432));
 sg13g2_tiehi _34729__433 (.L_HI(net433));
 sg13g2_tiehi _34728__434 (.L_HI(net434));
 sg13g2_tiehi _34727__435 (.L_HI(net435));
 sg13g2_tiehi _34726__436 (.L_HI(net436));
 sg13g2_tiehi _34725__437 (.L_HI(net437));
 sg13g2_tiehi _34724__438 (.L_HI(net438));
 sg13g2_tiehi _34723__439 (.L_HI(net439));
 sg13g2_tiehi _34722__440 (.L_HI(net440));
 sg13g2_tiehi _34721__441 (.L_HI(net441));
 sg13g2_tiehi _34720__442 (.L_HI(net442));
 sg13g2_tiehi _34719__443 (.L_HI(net443));
 sg13g2_tiehi _34718__444 (.L_HI(net444));
 sg13g2_tiehi _34717__445 (.L_HI(net445));
 sg13g2_tiehi _34716__446 (.L_HI(net446));
 sg13g2_tiehi _34715__447 (.L_HI(net447));
 sg13g2_tiehi _34714__448 (.L_HI(net448));
 sg13g2_tiehi _34713__449 (.L_HI(net449));
 sg13g2_tiehi _34712__450 (.L_HI(net450));
 sg13g2_tiehi _34711__451 (.L_HI(net451));
 sg13g2_tiehi _34710__452 (.L_HI(net452));
 sg13g2_tiehi _34709__453 (.L_HI(net453));
 sg13g2_tiehi _34708__454 (.L_HI(net454));
 sg13g2_tiehi _34707__455 (.L_HI(net455));
 sg13g2_tiehi _34706__456 (.L_HI(net456));
 sg13g2_tiehi _34705__457 (.L_HI(net457));
 sg13g2_tiehi _34704__458 (.L_HI(net458));
 sg13g2_tiehi _34703__459 (.L_HI(net459));
 sg13g2_tiehi _34702__460 (.L_HI(net460));
 sg13g2_tiehi _34701__461 (.L_HI(net461));
 sg13g2_tiehi _34700__462 (.L_HI(net462));
 sg13g2_tiehi _34699__463 (.L_HI(net463));
 sg13g2_tiehi _34698__464 (.L_HI(net464));
 sg13g2_tiehi _34697__465 (.L_HI(net465));
 sg13g2_tiehi _34696__466 (.L_HI(net466));
 sg13g2_tiehi _34695__467 (.L_HI(net467));
 sg13g2_tiehi _34694__468 (.L_HI(net468));
 sg13g2_tiehi _34693__469 (.L_HI(net469));
 sg13g2_tiehi _34692__470 (.L_HI(net470));
 sg13g2_tiehi _34691__471 (.L_HI(net471));
 sg13g2_tiehi _34690__472 (.L_HI(net472));
 sg13g2_tiehi _34689__473 (.L_HI(net473));
 sg13g2_tiehi _34688__474 (.L_HI(net474));
 sg13g2_tiehi _34687__475 (.L_HI(net475));
 sg13g2_tiehi _34686__476 (.L_HI(net476));
 sg13g2_tiehi _34685__477 (.L_HI(net477));
 sg13g2_tiehi _34684__478 (.L_HI(net478));
 sg13g2_tiehi _34683__479 (.L_HI(net479));
 sg13g2_tiehi _34682__480 (.L_HI(net480));
 sg13g2_tiehi _34681__481 (.L_HI(net481));
 sg13g2_tiehi _34680__482 (.L_HI(net482));
 sg13g2_tiehi _34679__483 (.L_HI(net483));
 sg13g2_tiehi _34678__484 (.L_HI(net484));
 sg13g2_tiehi _34677__485 (.L_HI(net485));
 sg13g2_tiehi _34676__486 (.L_HI(net486));
 sg13g2_tiehi _34675__487 (.L_HI(net487));
 sg13g2_tiehi _34674__488 (.L_HI(net488));
 sg13g2_tiehi _34673__489 (.L_HI(net489));
 sg13g2_tiehi _34672__490 (.L_HI(net490));
 sg13g2_tiehi _34671__491 (.L_HI(net491));
 sg13g2_tiehi _34670__492 (.L_HI(net492));
 sg13g2_tiehi _34669__493 (.L_HI(net493));
 sg13g2_tiehi _34668__494 (.L_HI(net494));
 sg13g2_tiehi _34667__495 (.L_HI(net495));
 sg13g2_tiehi _34666__496 (.L_HI(net496));
 sg13g2_tiehi _34665__497 (.L_HI(net497));
 sg13g2_tiehi _34664__498 (.L_HI(net498));
 sg13g2_tiehi _34663__499 (.L_HI(net499));
 sg13g2_tiehi _34662__500 (.L_HI(net500));
 sg13g2_tiehi _34661__501 (.L_HI(net501));
 sg13g2_tiehi _34660__502 (.L_HI(net502));
 sg13g2_tiehi _34659__503 (.L_HI(net503));
 sg13g2_tiehi _34658__504 (.L_HI(net504));
 sg13g2_tiehi _34657__505 (.L_HI(net505));
 sg13g2_tiehi _34656__506 (.L_HI(net506));
 sg13g2_tiehi _34655__507 (.L_HI(net507));
 sg13g2_tiehi _34654__508 (.L_HI(net508));
 sg13g2_tiehi _34653__509 (.L_HI(net509));
 sg13g2_tiehi _34652__510 (.L_HI(net510));
 sg13g2_tiehi _34651__511 (.L_HI(net511));
 sg13g2_tiehi _34650__512 (.L_HI(net512));
 sg13g2_tiehi _34649__513 (.L_HI(net513));
 sg13g2_tiehi _34648__514 (.L_HI(net514));
 sg13g2_tiehi _34647__515 (.L_HI(net515));
 sg13g2_tiehi _34646__516 (.L_HI(net516));
 sg13g2_tiehi _34645__517 (.L_HI(net517));
 sg13g2_tiehi _34644__518 (.L_HI(net518));
 sg13g2_tiehi _34643__519 (.L_HI(net519));
 sg13g2_tiehi _34642__520 (.L_HI(net520));
 sg13g2_tiehi _34641__521 (.L_HI(net521));
 sg13g2_tiehi _34640__522 (.L_HI(net522));
 sg13g2_tiehi _34639__523 (.L_HI(net523));
 sg13g2_tiehi _34638__524 (.L_HI(net524));
 sg13g2_tiehi _34637__525 (.L_HI(net525));
 sg13g2_tiehi _34636__526 (.L_HI(net526));
 sg13g2_tiehi _34635__527 (.L_HI(net527));
 sg13g2_tiehi _34634__528 (.L_HI(net528));
 sg13g2_tiehi _34633__529 (.L_HI(net529));
 sg13g2_tiehi _34632__530 (.L_HI(net530));
 sg13g2_tiehi _34631__531 (.L_HI(net531));
 sg13g2_tiehi _34630__532 (.L_HI(net532));
 sg13g2_tiehi _34629__533 (.L_HI(net533));
 sg13g2_tiehi _34628__534 (.L_HI(net534));
 sg13g2_tiehi _34627__535 (.L_HI(net535));
 sg13g2_tiehi _34626__536 (.L_HI(net536));
 sg13g2_tiehi _34625__537 (.L_HI(net537));
 sg13g2_tiehi _34624__538 (.L_HI(net538));
 sg13g2_tiehi _34623__539 (.L_HI(net539));
 sg13g2_tiehi _34622__540 (.L_HI(net540));
 sg13g2_tiehi _34621__541 (.L_HI(net541));
 sg13g2_tiehi _34620__542 (.L_HI(net542));
 sg13g2_tiehi _34619__543 (.L_HI(net543));
 sg13g2_tiehi _34618__544 (.L_HI(net544));
 sg13g2_tiehi _34617__545 (.L_HI(net545));
 sg13g2_tiehi _34616__546 (.L_HI(net546));
 sg13g2_tiehi _34615__547 (.L_HI(net547));
 sg13g2_tiehi _34614__548 (.L_HI(net548));
 sg13g2_tiehi _34613__549 (.L_HI(net549));
 sg13g2_tiehi _34612__550 (.L_HI(net550));
 sg13g2_tiehi _34611__551 (.L_HI(net551));
 sg13g2_tiehi _34610__552 (.L_HI(net552));
 sg13g2_tiehi _34609__553 (.L_HI(net553));
 sg13g2_tiehi _34608__554 (.L_HI(net554));
 sg13g2_tiehi _34607__555 (.L_HI(net555));
 sg13g2_tiehi _34606__556 (.L_HI(net556));
 sg13g2_tiehi _34605__557 (.L_HI(net557));
 sg13g2_tiehi _34604__558 (.L_HI(net558));
 sg13g2_tiehi _34603__559 (.L_HI(net559));
 sg13g2_tiehi _34602__560 (.L_HI(net560));
 sg13g2_tiehi _34601__561 (.L_HI(net561));
 sg13g2_tiehi _34600__562 (.L_HI(net562));
 sg13g2_tiehi _34599__563 (.L_HI(net563));
 sg13g2_tiehi _34598__564 (.L_HI(net564));
 sg13g2_tiehi _34597__565 (.L_HI(net565));
 sg13g2_tiehi _34596__566 (.L_HI(net566));
 sg13g2_tiehi _34595__567 (.L_HI(net567));
 sg13g2_tiehi _34594__568 (.L_HI(net568));
 sg13g2_tiehi _34593__569 (.L_HI(net569));
 sg13g2_tiehi _34592__570 (.L_HI(net570));
 sg13g2_tiehi _34591__571 (.L_HI(net571));
 sg13g2_tiehi _34590__572 (.L_HI(net572));
 sg13g2_tiehi _34589__573 (.L_HI(net573));
 sg13g2_tiehi _34588__574 (.L_HI(net574));
 sg13g2_tiehi _34587__575 (.L_HI(net575));
 sg13g2_tiehi _34586__576 (.L_HI(net576));
 sg13g2_tiehi _34585__577 (.L_HI(net577));
 sg13g2_tiehi _34584__578 (.L_HI(net578));
 sg13g2_tiehi _34583__579 (.L_HI(net579));
 sg13g2_tiehi _34582__580 (.L_HI(net580));
 sg13g2_tiehi _34581__581 (.L_HI(net581));
 sg13g2_tiehi _34580__582 (.L_HI(net582));
 sg13g2_tiehi _34579__583 (.L_HI(net583));
 sg13g2_tiehi _34578__584 (.L_HI(net584));
 sg13g2_tiehi _34577__585 (.L_HI(net585));
 sg13g2_tiehi _34576__586 (.L_HI(net586));
 sg13g2_tiehi _34575__587 (.L_HI(net587));
 sg13g2_tiehi _34574__588 (.L_HI(net588));
 sg13g2_tiehi _34573__589 (.L_HI(net589));
 sg13g2_tiehi _34572__590 (.L_HI(net590));
 sg13g2_tiehi _34571__591 (.L_HI(net591));
 sg13g2_tiehi _34570__592 (.L_HI(net592));
 sg13g2_tiehi _34569__593 (.L_HI(net593));
 sg13g2_tiehi _34568__594 (.L_HI(net594));
 sg13g2_tiehi _34567__595 (.L_HI(net595));
 sg13g2_tiehi _34566__596 (.L_HI(net596));
 sg13g2_tiehi _34565__597 (.L_HI(net597));
 sg13g2_tiehi _34564__598 (.L_HI(net598));
 sg13g2_tiehi _34563__599 (.L_HI(net599));
 sg13g2_tiehi _34562__600 (.L_HI(net600));
 sg13g2_tiehi _34561__601 (.L_HI(net601));
 sg13g2_tiehi _34560__602 (.L_HI(net602));
 sg13g2_tiehi _34559__603 (.L_HI(net603));
 sg13g2_tiehi _34558__604 (.L_HI(net604));
 sg13g2_tiehi _34557__605 (.L_HI(net605));
 sg13g2_tiehi _34556__606 (.L_HI(net606));
 sg13g2_tiehi _34555__607 (.L_HI(net607));
 sg13g2_tiehi _34554__608 (.L_HI(net608));
 sg13g2_tiehi _34553__609 (.L_HI(net609));
 sg13g2_tiehi _34552__610 (.L_HI(net610));
 sg13g2_tiehi _34551__611 (.L_HI(net611));
 sg13g2_tiehi _34550__612 (.L_HI(net612));
 sg13g2_tiehi _34549__613 (.L_HI(net613));
 sg13g2_tiehi _34548__614 (.L_HI(net614));
 sg13g2_tiehi _34547__615 (.L_HI(net615));
 sg13g2_tiehi _34546__616 (.L_HI(net616));
 sg13g2_tiehi _34545__617 (.L_HI(net617));
 sg13g2_tiehi _34544__618 (.L_HI(net618));
 sg13g2_tiehi _34543__619 (.L_HI(net619));
 sg13g2_tiehi _34542__620 (.L_HI(net620));
 sg13g2_tiehi _34541__621 (.L_HI(net621));
 sg13g2_tiehi _34540__622 (.L_HI(net622));
 sg13g2_tiehi _34539__623 (.L_HI(net623));
 sg13g2_tiehi _34538__624 (.L_HI(net624));
 sg13g2_tiehi _34537__625 (.L_HI(net625));
 sg13g2_tiehi _34536__626 (.L_HI(net626));
 sg13g2_tiehi _34535__627 (.L_HI(net627));
 sg13g2_tiehi _34534__628 (.L_HI(net628));
 sg13g2_tiehi _34533__629 (.L_HI(net629));
 sg13g2_tiehi _34532__630 (.L_HI(net630));
 sg13g2_tiehi _34531__631 (.L_HI(net631));
 sg13g2_tiehi _34530__632 (.L_HI(net632));
 sg13g2_tiehi _34529__633 (.L_HI(net633));
 sg13g2_tiehi _34528__634 (.L_HI(net634));
 sg13g2_tiehi _34527__635 (.L_HI(net635));
 sg13g2_tiehi _34526__636 (.L_HI(net636));
 sg13g2_tiehi _34525__637 (.L_HI(net637));
 sg13g2_tiehi _34524__638 (.L_HI(net638));
 sg13g2_tiehi _34523__639 (.L_HI(net639));
 sg13g2_tiehi _34522__640 (.L_HI(net640));
 sg13g2_tiehi _34521__641 (.L_HI(net641));
 sg13g2_tiehi _34520__642 (.L_HI(net642));
 sg13g2_tiehi _34519__643 (.L_HI(net643));
 sg13g2_tiehi _34518__644 (.L_HI(net644));
 sg13g2_tiehi _34517__645 (.L_HI(net645));
 sg13g2_tiehi _34516__646 (.L_HI(net646));
 sg13g2_tiehi _34515__647 (.L_HI(net647));
 sg13g2_tiehi _34514__648 (.L_HI(net648));
 sg13g2_tiehi _34513__649 (.L_HI(net649));
 sg13g2_tiehi _34512__650 (.L_HI(net650));
 sg13g2_tiehi _34511__651 (.L_HI(net651));
 sg13g2_tiehi _34510__652 (.L_HI(net652));
 sg13g2_tiehi _34509__653 (.L_HI(net653));
 sg13g2_tiehi _34508__654 (.L_HI(net654));
 sg13g2_tiehi _34507__655 (.L_HI(net655));
 sg13g2_tiehi _34506__656 (.L_HI(net656));
 sg13g2_tiehi _34505__657 (.L_HI(net657));
 sg13g2_tiehi _34504__658 (.L_HI(net658));
 sg13g2_tiehi _34503__659 (.L_HI(net659));
 sg13g2_tiehi _34502__660 (.L_HI(net660));
 sg13g2_tiehi _34501__661 (.L_HI(net661));
 sg13g2_tiehi _34500__662 (.L_HI(net662));
 sg13g2_tiehi _34499__663 (.L_HI(net663));
 sg13g2_tiehi _34498__664 (.L_HI(net664));
 sg13g2_tiehi _34497__665 (.L_HI(net665));
 sg13g2_tiehi _34496__666 (.L_HI(net666));
 sg13g2_tiehi _34495__667 (.L_HI(net667));
 sg13g2_tiehi _34494__668 (.L_HI(net668));
 sg13g2_tiehi _34493__669 (.L_HI(net669));
 sg13g2_tiehi _34492__670 (.L_HI(net670));
 sg13g2_tiehi _34491__671 (.L_HI(net671));
 sg13g2_tiehi _34490__672 (.L_HI(net672));
 sg13g2_tiehi _34489__673 (.L_HI(net673));
 sg13g2_tiehi _34488__674 (.L_HI(net674));
 sg13g2_tiehi _34487__675 (.L_HI(net675));
 sg13g2_tiehi _34486__676 (.L_HI(net676));
 sg13g2_tiehi _35266__677 (.L_HI(net677));
 sg13g2_tiehi _34485__678 (.L_HI(net678));
 sg13g2_tiehi _35265__679 (.L_HI(net679));
 sg13g2_tiehi _34484__680 (.L_HI(net680));
 sg13g2_tiehi _35264__681 (.L_HI(net681));
 sg13g2_tiehi _34483__682 (.L_HI(net682));
 sg13g2_tiehi _35263__683 (.L_HI(net683));
 sg13g2_tiehi _34482__684 (.L_HI(net684));
 sg13g2_tiehi _35262__685 (.L_HI(net685));
 sg13g2_tiehi _34481__686 (.L_HI(net686));
 sg13g2_tiehi _35261__687 (.L_HI(net687));
 sg13g2_tiehi _34480__688 (.L_HI(net688));
 sg13g2_tiehi _35260__689 (.L_HI(net689));
 sg13g2_tiehi _34479__690 (.L_HI(net690));
 sg13g2_tiehi _35259__691 (.L_HI(net691));
 sg13g2_tiehi _34478__692 (.L_HI(net692));
 sg13g2_tiehi _35258__693 (.L_HI(net693));
 sg13g2_tiehi _34477__694 (.L_HI(net694));
 sg13g2_tiehi _35257__695 (.L_HI(net695));
 sg13g2_tiehi _34476__696 (.L_HI(net696));
 sg13g2_tiehi _35256__697 (.L_HI(net697));
 sg13g2_tiehi _34475__698 (.L_HI(net698));
 sg13g2_tiehi _35255__699 (.L_HI(net699));
 sg13g2_tiehi _34474__700 (.L_HI(net700));
 sg13g2_tiehi _35254__701 (.L_HI(net701));
 sg13g2_tiehi _34473__702 (.L_HI(net702));
 sg13g2_tiehi _35253__703 (.L_HI(net703));
 sg13g2_tiehi _34472__704 (.L_HI(net704));
 sg13g2_tiehi _35252__705 (.L_HI(net705));
 sg13g2_tiehi _34471__706 (.L_HI(net706));
 sg13g2_tiehi _35251__707 (.L_HI(net707));
 sg13g2_tiehi _34470__708 (.L_HI(net708));
 sg13g2_tiehi _35250__709 (.L_HI(net709));
 sg13g2_tiehi _34469__710 (.L_HI(net710));
 sg13g2_tiehi _35249__711 (.L_HI(net711));
 sg13g2_tiehi _34468__712 (.L_HI(net712));
 sg13g2_tiehi _35248__713 (.L_HI(net713));
 sg13g2_tiehi _34467__714 (.L_HI(net714));
 sg13g2_tiehi _35247__715 (.L_HI(net715));
 sg13g2_tiehi _34466__716 (.L_HI(net716));
 sg13g2_tiehi _35246__717 (.L_HI(net717));
 sg13g2_tiehi _34465__718 (.L_HI(net718));
 sg13g2_tiehi _35245__719 (.L_HI(net719));
 sg13g2_tiehi _34464__720 (.L_HI(net720));
 sg13g2_tiehi _35244__721 (.L_HI(net721));
 sg13g2_tiehi _34463__722 (.L_HI(net722));
 sg13g2_tiehi _35243__723 (.L_HI(net723));
 sg13g2_tiehi _34462__724 (.L_HI(net724));
 sg13g2_tiehi _35242__725 (.L_HI(net725));
 sg13g2_tiehi _34461__726 (.L_HI(net726));
 sg13g2_tiehi _35241__727 (.L_HI(net727));
 sg13g2_tiehi _34460__728 (.L_HI(net728));
 sg13g2_tiehi _35240__729 (.L_HI(net729));
 sg13g2_tiehi _34459__730 (.L_HI(net730));
 sg13g2_tiehi _35239__731 (.L_HI(net731));
 sg13g2_tiehi _34458__732 (.L_HI(net732));
 sg13g2_tiehi _35238__733 (.L_HI(net733));
 sg13g2_tiehi _34457__734 (.L_HI(net734));
 sg13g2_tiehi _35237__735 (.L_HI(net735));
 sg13g2_tiehi _34456__736 (.L_HI(net736));
 sg13g2_tiehi _35236__737 (.L_HI(net737));
 sg13g2_tiehi _34455__738 (.L_HI(net738));
 sg13g2_tiehi _35235__739 (.L_HI(net739));
 sg13g2_tiehi _34454__740 (.L_HI(net740));
 sg13g2_tiehi _35234__741 (.L_HI(net741));
 sg13g2_tiehi _34453__742 (.L_HI(net742));
 sg13g2_tiehi _35233__743 (.L_HI(net743));
 sg13g2_tiehi _34452__744 (.L_HI(net744));
 sg13g2_tiehi _35232__745 (.L_HI(net745));
 sg13g2_tiehi _34451__746 (.L_HI(net746));
 sg13g2_tiehi _35231__747 (.L_HI(net747));
 sg13g2_tiehi _34450__748 (.L_HI(net748));
 sg13g2_tiehi _35230__749 (.L_HI(net749));
 sg13g2_tiehi _34449__750 (.L_HI(net750));
 sg13g2_tiehi _35229__751 (.L_HI(net751));
 sg13g2_tiehi _34448__752 (.L_HI(net752));
 sg13g2_tiehi _35228__753 (.L_HI(net753));
 sg13g2_tiehi _34447__754 (.L_HI(net754));
 sg13g2_tiehi _35227__755 (.L_HI(net755));
 sg13g2_tiehi _34446__756 (.L_HI(net756));
 sg13g2_tiehi _35226__757 (.L_HI(net757));
 sg13g2_tiehi _34445__758 (.L_HI(net758));
 sg13g2_tiehi _35225__759 (.L_HI(net759));
 sg13g2_tiehi _34444__760 (.L_HI(net760));
 sg13g2_tiehi _35224__761 (.L_HI(net761));
 sg13g2_tiehi _34443__762 (.L_HI(net762));
 sg13g2_tiehi _35223__763 (.L_HI(net763));
 sg13g2_tiehi _34442__764 (.L_HI(net764));
 sg13g2_tiehi _35222__765 (.L_HI(net765));
 sg13g2_tiehi _34441__766 (.L_HI(net766));
 sg13g2_tiehi _35221__767 (.L_HI(net767));
 sg13g2_tiehi _34440__768 (.L_HI(net768));
 sg13g2_tiehi _35220__769 (.L_HI(net769));
 sg13g2_tiehi _34439__770 (.L_HI(net770));
 sg13g2_tiehi _35219__771 (.L_HI(net771));
 sg13g2_tiehi _34438__772 (.L_HI(net772));
 sg13g2_tiehi _35218__773 (.L_HI(net773));
 sg13g2_tiehi _34437__774 (.L_HI(net774));
 sg13g2_tiehi _35217__775 (.L_HI(net775));
 sg13g2_tiehi _34436__776 (.L_HI(net776));
 sg13g2_tiehi _35216__777 (.L_HI(net777));
 sg13g2_tiehi _34435__778 (.L_HI(net778));
 sg13g2_tiehi _35215__779 (.L_HI(net779));
 sg13g2_tiehi _34434__780 (.L_HI(net780));
 sg13g2_tiehi _35214__781 (.L_HI(net781));
 sg13g2_tiehi _34433__782 (.L_HI(net782));
 sg13g2_tiehi _35213__783 (.L_HI(net783));
 sg13g2_tiehi _34432__784 (.L_HI(net784));
 sg13g2_tiehi _35212__785 (.L_HI(net785));
 sg13g2_tiehi _34431__786 (.L_HI(net786));
 sg13g2_tiehi _35211__787 (.L_HI(net787));
 sg13g2_tiehi _34430__788 (.L_HI(net788));
 sg13g2_tiehi _35210__789 (.L_HI(net789));
 sg13g2_tiehi _34429__790 (.L_HI(net790));
 sg13g2_tiehi _35209__791 (.L_HI(net791));
 sg13g2_tiehi _34428__792 (.L_HI(net792));
 sg13g2_tiehi _35208__793 (.L_HI(net793));
 sg13g2_tiehi _34427__794 (.L_HI(net794));
 sg13g2_tiehi _35207__795 (.L_HI(net795));
 sg13g2_tiehi _34426__796 (.L_HI(net796));
 sg13g2_tiehi _35206__797 (.L_HI(net797));
 sg13g2_tiehi _34425__798 (.L_HI(net798));
 sg13g2_tiehi _35205__799 (.L_HI(net799));
 sg13g2_tiehi _34424__800 (.L_HI(net800));
 sg13g2_tiehi _35204__801 (.L_HI(net801));
 sg13g2_tiehi _34423__802 (.L_HI(net802));
 sg13g2_tiehi _35203__803 (.L_HI(net803));
 sg13g2_tiehi _34422__804 (.L_HI(net804));
 sg13g2_tiehi _35202__805 (.L_HI(net805));
 sg13g2_tiehi _34421__806 (.L_HI(net806));
 sg13g2_tiehi _35201__807 (.L_HI(net807));
 sg13g2_tiehi _34420__808 (.L_HI(net808));
 sg13g2_tiehi _35200__809 (.L_HI(net809));
 sg13g2_tiehi _34419__810 (.L_HI(net810));
 sg13g2_tiehi _35199__811 (.L_HI(net811));
 sg13g2_tiehi _34418__812 (.L_HI(net812));
 sg13g2_tiehi _35198__813 (.L_HI(net813));
 sg13g2_tiehi _34417__814 (.L_HI(net814));
 sg13g2_tiehi _35197__815 (.L_HI(net815));
 sg13g2_tiehi _34416__816 (.L_HI(net816));
 sg13g2_tiehi _35196__817 (.L_HI(net817));
 sg13g2_tiehi _34415__818 (.L_HI(net818));
 sg13g2_tiehi _35195__819 (.L_HI(net819));
 sg13g2_tiehi _34414__820 (.L_HI(net820));
 sg13g2_tiehi _35194__821 (.L_HI(net821));
 sg13g2_tiehi _34413__822 (.L_HI(net822));
 sg13g2_tiehi _35193__823 (.L_HI(net823));
 sg13g2_tiehi _34412__824 (.L_HI(net824));
 sg13g2_tiehi _35192__825 (.L_HI(net825));
 sg13g2_tiehi _34411__826 (.L_HI(net826));
 sg13g2_tiehi _35191__827 (.L_HI(net827));
 sg13g2_tiehi _34410__828 (.L_HI(net828));
 sg13g2_tiehi _35190__829 (.L_HI(net829));
 sg13g2_tiehi _34409__830 (.L_HI(net830));
 sg13g2_tiehi _35189__831 (.L_HI(net831));
 sg13g2_tiehi _34408__832 (.L_HI(net832));
 sg13g2_tiehi _35188__833 (.L_HI(net833));
 sg13g2_tiehi _34407__834 (.L_HI(net834));
 sg13g2_tiehi _35187__835 (.L_HI(net835));
 sg13g2_tiehi _34406__836 (.L_HI(net836));
 sg13g2_tiehi _35186__837 (.L_HI(net837));
 sg13g2_tiehi _34405__838 (.L_HI(net838));
 sg13g2_tiehi _35185__839 (.L_HI(net839));
 sg13g2_tiehi _34404__840 (.L_HI(net840));
 sg13g2_tiehi _35184__841 (.L_HI(net841));
 sg13g2_tiehi _34403__842 (.L_HI(net842));
 sg13g2_tiehi _35183__843 (.L_HI(net843));
 sg13g2_tiehi _34402__844 (.L_HI(net844));
 sg13g2_tiehi _35182__845 (.L_HI(net845));
 sg13g2_tiehi _34401__846 (.L_HI(net846));
 sg13g2_tiehi _35181__847 (.L_HI(net847));
 sg13g2_tiehi _34400__848 (.L_HI(net848));
 sg13g2_tiehi _35180__849 (.L_HI(net849));
 sg13g2_tiehi _34399__850 (.L_HI(net850));
 sg13g2_tiehi _35179__851 (.L_HI(net851));
 sg13g2_tiehi _34398__852 (.L_HI(net852));
 sg13g2_tiehi _35178__853 (.L_HI(net853));
 sg13g2_tiehi _34397__854 (.L_HI(net854));
 sg13g2_tiehi _35177__855 (.L_HI(net855));
 sg13g2_tiehi _34396__856 (.L_HI(net856));
 sg13g2_tiehi _35176__857 (.L_HI(net857));
 sg13g2_tiehi _34395__858 (.L_HI(net858));
 sg13g2_tiehi _35175__859 (.L_HI(net859));
 sg13g2_tiehi _34394__860 (.L_HI(net860));
 sg13g2_tiehi _35174__861 (.L_HI(net861));
 sg13g2_tiehi _34393__862 (.L_HI(net862));
 sg13g2_tiehi _35173__863 (.L_HI(net863));
 sg13g2_tiehi _34392__864 (.L_HI(net864));
 sg13g2_tiehi _35172__865 (.L_HI(net865));
 sg13g2_tiehi _34391__866 (.L_HI(net866));
 sg13g2_tiehi _35171__867 (.L_HI(net867));
 sg13g2_tiehi _34390__868 (.L_HI(net868));
 sg13g2_tiehi _35170__869 (.L_HI(net869));
 sg13g2_tiehi _34389__870 (.L_HI(net870));
 sg13g2_tiehi _35169__871 (.L_HI(net871));
 sg13g2_tiehi _34388__872 (.L_HI(net872));
 sg13g2_tiehi _35168__873 (.L_HI(net873));
 sg13g2_tiehi _34387__874 (.L_HI(net874));
 sg13g2_tiehi _35167__875 (.L_HI(net875));
 sg13g2_tiehi _34386__876 (.L_HI(net876));
 sg13g2_tiehi _35166__877 (.L_HI(net877));
 sg13g2_tiehi _34385__878 (.L_HI(net878));
 sg13g2_tiehi _35165__879 (.L_HI(net879));
 sg13g2_tiehi _34384__880 (.L_HI(net880));
 sg13g2_tiehi _35164__881 (.L_HI(net881));
 sg13g2_tiehi _34383__882 (.L_HI(net882));
 sg13g2_tiehi _35163__883 (.L_HI(net883));
 sg13g2_tiehi _34382__884 (.L_HI(net884));
 sg13g2_tiehi _35162__885 (.L_HI(net885));
 sg13g2_tiehi _34381__886 (.L_HI(net886));
 sg13g2_tiehi _35161__887 (.L_HI(net887));
 sg13g2_tiehi _34380__888 (.L_HI(net888));
 sg13g2_tiehi _35160__889 (.L_HI(net889));
 sg13g2_tiehi _34379__890 (.L_HI(net890));
 sg13g2_tiehi _35159__891 (.L_HI(net891));
 sg13g2_tiehi _34378__892 (.L_HI(net892));
 sg13g2_tiehi _35158__893 (.L_HI(net893));
 sg13g2_tiehi _34377__894 (.L_HI(net894));
 sg13g2_tiehi _35157__895 (.L_HI(net895));
 sg13g2_tiehi _34376__896 (.L_HI(net896));
 sg13g2_tiehi _35156__897 (.L_HI(net897));
 sg13g2_tiehi _34375__898 (.L_HI(net898));
 sg13g2_tiehi _35155__899 (.L_HI(net899));
 sg13g2_tiehi _34374__900 (.L_HI(net900));
 sg13g2_tiehi _35154__901 (.L_HI(net901));
 sg13g2_tiehi _34373__902 (.L_HI(net902));
 sg13g2_tiehi _35153__903 (.L_HI(net903));
 sg13g2_tiehi _34372__904 (.L_HI(net904));
 sg13g2_tiehi _35152__905 (.L_HI(net905));
 sg13g2_tiehi _34371__906 (.L_HI(net906));
 sg13g2_tiehi _35151__907 (.L_HI(net907));
 sg13g2_tiehi _34370__908 (.L_HI(net908));
 sg13g2_tiehi _35150__909 (.L_HI(net909));
 sg13g2_tiehi _34369__910 (.L_HI(net910));
 sg13g2_tiehi _35149__911 (.L_HI(net911));
 sg13g2_tiehi _34368__912 (.L_HI(net912));
 sg13g2_tiehi _35148__913 (.L_HI(net913));
 sg13g2_tiehi _34367__914 (.L_HI(net914));
 sg13g2_tiehi _35147__915 (.L_HI(net915));
 sg13g2_tiehi _34366__916 (.L_HI(net916));
 sg13g2_tiehi _35146__917 (.L_HI(net917));
 sg13g2_tiehi _34365__918 (.L_HI(net918));
 sg13g2_tiehi _35145__919 (.L_HI(net919));
 sg13g2_tiehi _34364__920 (.L_HI(net920));
 sg13g2_tiehi _35144__921 (.L_HI(net921));
 sg13g2_tiehi _34363__922 (.L_HI(net922));
 sg13g2_tiehi _35143__923 (.L_HI(net923));
 sg13g2_tiehi _34362__924 (.L_HI(net924));
 sg13g2_tiehi _35142__925 (.L_HI(net925));
 sg13g2_tiehi _34361__926 (.L_HI(net926));
 sg13g2_tiehi _35141__927 (.L_HI(net927));
 sg13g2_tiehi _34360__928 (.L_HI(net928));
 sg13g2_tiehi _35140__929 (.L_HI(net929));
 sg13g2_tiehi _34359__930 (.L_HI(net930));
 sg13g2_tiehi _35139__931 (.L_HI(net931));
 sg13g2_tiehi _34358__932 (.L_HI(net932));
 sg13g2_tiehi _35138__933 (.L_HI(net933));
 sg13g2_tiehi _34357__934 (.L_HI(net934));
 sg13g2_tiehi _35137__935 (.L_HI(net935));
 sg13g2_tiehi _34356__936 (.L_HI(net936));
 sg13g2_tiehi _35136__937 (.L_HI(net937));
 sg13g2_tiehi _34355__938 (.L_HI(net938));
 sg13g2_tiehi _35135__939 (.L_HI(net939));
 sg13g2_tiehi _34354__940 (.L_HI(net940));
 sg13g2_tiehi _35134__941 (.L_HI(net941));
 sg13g2_tiehi _34353__942 (.L_HI(net942));
 sg13g2_tiehi _35133__943 (.L_HI(net943));
 sg13g2_tiehi _34352__944 (.L_HI(net944));
 sg13g2_tiehi _35132__945 (.L_HI(net945));
 sg13g2_tiehi _34351__946 (.L_HI(net946));
 sg13g2_tiehi _35131__947 (.L_HI(net947));
 sg13g2_tiehi _34350__948 (.L_HI(net948));
 sg13g2_tiehi _35130__949 (.L_HI(net949));
 sg13g2_tiehi _34349__950 (.L_HI(net950));
 sg13g2_tiehi _35129__951 (.L_HI(net951));
 sg13g2_tiehi _34348__952 (.L_HI(net952));
 sg13g2_tiehi _35128__953 (.L_HI(net953));
 sg13g2_tiehi _34347__954 (.L_HI(net954));
 sg13g2_tiehi _35127__955 (.L_HI(net955));
 sg13g2_tiehi _34346__956 (.L_HI(net956));
 sg13g2_tiehi _35126__957 (.L_HI(net957));
 sg13g2_tiehi _34345__958 (.L_HI(net958));
 sg13g2_tiehi _35125__959 (.L_HI(net959));
 sg13g2_tiehi _34344__960 (.L_HI(net960));
 sg13g2_tiehi _35124__961 (.L_HI(net961));
 sg13g2_tiehi _34343__962 (.L_HI(net962));
 sg13g2_tiehi _35123__963 (.L_HI(net963));
 sg13g2_tiehi _34342__964 (.L_HI(net964));
 sg13g2_tiehi _35122__965 (.L_HI(net965));
 sg13g2_tiehi _34341__966 (.L_HI(net966));
 sg13g2_tiehi _35121__967 (.L_HI(net967));
 sg13g2_tiehi _34340__968 (.L_HI(net968));
 sg13g2_tiehi _35120__969 (.L_HI(net969));
 sg13g2_tiehi _34339__970 (.L_HI(net970));
 sg13g2_tiehi _35119__971 (.L_HI(net971));
 sg13g2_tiehi _34338__972 (.L_HI(net972));
 sg13g2_tiehi _35118__973 (.L_HI(net973));
 sg13g2_tiehi _34337__974 (.L_HI(net974));
 sg13g2_tiehi _35117__975 (.L_HI(net975));
 sg13g2_tiehi _34336__976 (.L_HI(net976));
 sg13g2_tiehi _35116__977 (.L_HI(net977));
 sg13g2_tiehi _34335__978 (.L_HI(net978));
 sg13g2_tiehi _35115__979 (.L_HI(net979));
 sg13g2_tiehi _34334__980 (.L_HI(net980));
 sg13g2_tiehi _35114__981 (.L_HI(net981));
 sg13g2_tiehi _34333__982 (.L_HI(net982));
 sg13g2_tiehi _35113__983 (.L_HI(net983));
 sg13g2_tiehi _34332__984 (.L_HI(net984));
 sg13g2_tiehi _35112__985 (.L_HI(net985));
 sg13g2_tiehi _34331__986 (.L_HI(net986));
 sg13g2_tiehi _35111__987 (.L_HI(net987));
 sg13g2_tiehi _34330__988 (.L_HI(net988));
 sg13g2_tiehi _35110__989 (.L_HI(net989));
 sg13g2_tiehi _34329__990 (.L_HI(net990));
 sg13g2_tiehi _35109__991 (.L_HI(net991));
 sg13g2_tiehi _34328__992 (.L_HI(net992));
 sg13g2_tiehi _35108__993 (.L_HI(net993));
 sg13g2_tiehi _34327__994 (.L_HI(net994));
 sg13g2_tiehi _35107__995 (.L_HI(net995));
 sg13g2_tiehi _34326__996 (.L_HI(net996));
 sg13g2_tiehi _35106__997 (.L_HI(net997));
 sg13g2_tiehi _34325__998 (.L_HI(net998));
 sg13g2_tiehi _35105__999 (.L_HI(net999));
 sg13g2_tiehi _34324__1000 (.L_HI(net1000));
 sg13g2_tiehi _35104__1001 (.L_HI(net1001));
 sg13g2_tiehi _34323__1002 (.L_HI(net1002));
 sg13g2_tiehi _35103__1003 (.L_HI(net1003));
 sg13g2_tiehi _34322__1004 (.L_HI(net1004));
 sg13g2_tiehi _35102__1005 (.L_HI(net1005));
 sg13g2_tiehi _34321__1006 (.L_HI(net1006));
 sg13g2_tiehi _35101__1007 (.L_HI(net1007));
 sg13g2_tiehi _34320__1008 (.L_HI(net1008));
 sg13g2_tiehi _35100__1009 (.L_HI(net1009));
 sg13g2_tiehi _34319__1010 (.L_HI(net1010));
 sg13g2_tiehi _35099__1011 (.L_HI(net1011));
 sg13g2_tiehi _34318__1012 (.L_HI(net1012));
 sg13g2_tiehi _35098__1013 (.L_HI(net1013));
 sg13g2_tiehi _34317__1014 (.L_HI(net1014));
 sg13g2_tiehi _35097__1015 (.L_HI(net1015));
 sg13g2_tiehi _34316__1016 (.L_HI(net1016));
 sg13g2_tiehi _35096__1017 (.L_HI(net1017));
 sg13g2_tiehi _34315__1018 (.L_HI(net1018));
 sg13g2_tiehi _35095__1019 (.L_HI(net1019));
 sg13g2_tiehi _34314__1020 (.L_HI(net1020));
 sg13g2_tiehi _35094__1021 (.L_HI(net1021));
 sg13g2_tiehi _34313__1022 (.L_HI(net1022));
 sg13g2_tiehi _35093__1023 (.L_HI(net1023));
 sg13g2_tiehi _34312__1024 (.L_HI(net1024));
 sg13g2_tiehi _35092__1025 (.L_HI(net1025));
 sg13g2_tiehi _34311__1026 (.L_HI(net1026));
 sg13g2_tiehi _35091__1027 (.L_HI(net1027));
 sg13g2_tiehi _34310__1028 (.L_HI(net1028));
 sg13g2_tiehi _35090__1029 (.L_HI(net1029));
 sg13g2_tiehi _34309__1030 (.L_HI(net1030));
 sg13g2_tiehi _35089__1031 (.L_HI(net1031));
 sg13g2_tiehi _34308__1032 (.L_HI(net1032));
 sg13g2_tiehi _35088__1033 (.L_HI(net1033));
 sg13g2_tiehi _34307__1034 (.L_HI(net1034));
 sg13g2_tiehi _35087__1035 (.L_HI(net1035));
 sg13g2_tiehi _34306__1036 (.L_HI(net1036));
 sg13g2_tiehi _35086__1037 (.L_HI(net1037));
 sg13g2_tiehi _34305__1038 (.L_HI(net1038));
 sg13g2_tiehi _35085__1039 (.L_HI(net1039));
 sg13g2_tiehi _34304__1040 (.L_HI(net1040));
 sg13g2_tiehi _35084__1041 (.L_HI(net1041));
 sg13g2_tiehi _34303__1042 (.L_HI(net1042));
 sg13g2_tiehi _35083__1043 (.L_HI(net1043));
 sg13g2_tiehi _34302__1044 (.L_HI(net1044));
 sg13g2_tiehi _35082__1045 (.L_HI(net1045));
 sg13g2_tiehi _34301__1046 (.L_HI(net1046));
 sg13g2_tiehi _35081__1047 (.L_HI(net1047));
 sg13g2_tiehi _34300__1048 (.L_HI(net1048));
 sg13g2_tiehi _35080__1049 (.L_HI(net1049));
 sg13g2_tiehi _34299__1050 (.L_HI(net1050));
 sg13g2_tiehi _35079__1051 (.L_HI(net1051));
 sg13g2_tiehi _34298__1052 (.L_HI(net1052));
 sg13g2_tiehi _35078__1053 (.L_HI(net1053));
 sg13g2_tiehi _34297__1054 (.L_HI(net1054));
 sg13g2_tiehi _35077__1055 (.L_HI(net1055));
 sg13g2_tiehi _34296__1056 (.L_HI(net1056));
 sg13g2_tiehi _35076__1057 (.L_HI(net1057));
 sg13g2_tiehi _34295__1058 (.L_HI(net1058));
 sg13g2_tiehi _35075__1059 (.L_HI(net1059));
 sg13g2_tiehi _34294__1060 (.L_HI(net1060));
 sg13g2_tiehi tt_um_corey_1061 (.L_HI(net1061));
 sg13g2_tiehi tt_um_corey_1062 (.L_HI(net1062));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_corey_12 (.L_LO(net12));
 sg13g2_tielo tt_um_corey_13 (.L_LO(net13));
 sg13g2_tielo tt_um_corey_14 (.L_LO(net14));
 sg13g2_tielo tt_um_corey_15 (.L_LO(net15));
 sg13g2_tielo tt_um_corey_16 (.L_LO(net16));
 sg13g2_tielo tt_um_corey_17 (.L_LO(net17));
 sg13g2_tielo tt_um_corey_18 (.L_LO(net18));
 sg13g2_tielo tt_um_corey_19 (.L_LO(net19));
 sg13g2_tielo tt_um_corey_20 (.L_LO(net20));
 sg13g2_tielo tt_um_corey_21 (.L_LO(net21));
 sg13g2_tielo tt_um_corey_22 (.L_LO(net22));
 sg13g2_tiehi _35074__23 (.L_HI(net23));
 sg13g2_buf_1 _36587_ (.A(\shift_reg[248] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _36588_ (.A(\shift_reg[249] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _36589_ (.A(\shift_reg[250] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _36590_ (.A(\shift_reg[251] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _36591_ (.A(\shift_reg[252] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _36592_ (.A(\shift_reg[253] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _36593_ (.A(\shift_reg[254] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _36594_ (.A(\shift_reg[255] ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout3310 (.A(net3312),
    .X(net3310));
 sg13g2_buf_8 fanout3311 (.A(net3312),
    .X(net3311));
 sg13g2_buf_8 fanout3312 (.A(_06643_),
    .X(net3312));
 sg13g2_buf_8 fanout3313 (.A(net3317),
    .X(net3313));
 sg13g2_buf_8 fanout3314 (.A(net3315),
    .X(net3314));
 sg13g2_buf_8 fanout3315 (.A(net3316),
    .X(net3315));
 sg13g2_buf_8 fanout3316 (.A(net3317),
    .X(net3316));
 sg13g2_buf_8 fanout3317 (.A(_06643_),
    .X(net3317));
 sg13g2_buf_8 fanout3318 (.A(net3319),
    .X(net3318));
 sg13g2_buf_8 fanout3319 (.A(net3322),
    .X(net3319));
 sg13g2_buf_8 fanout3320 (.A(net3321),
    .X(net3320));
 sg13g2_buf_8 fanout3321 (.A(net3322),
    .X(net3321));
 sg13g2_buf_8 fanout3322 (.A(net3329),
    .X(net3322));
 sg13g2_buf_8 fanout3323 (.A(net3324),
    .X(net3323));
 sg13g2_buf_8 fanout3324 (.A(net3329),
    .X(net3324));
 sg13g2_buf_8 fanout3325 (.A(net3328),
    .X(net3325));
 sg13g2_buf_8 fanout3326 (.A(net3328),
    .X(net3326));
 sg13g2_buf_1 fanout3327 (.A(net3328),
    .X(net3327));
 sg13g2_buf_8 fanout3328 (.A(net3329),
    .X(net3328));
 sg13g2_buf_8 fanout3329 (.A(_06642_),
    .X(net3329));
 sg13g2_buf_8 fanout3330 (.A(net3331),
    .X(net3330));
 sg13g2_buf_8 fanout3331 (.A(_06641_),
    .X(net3331));
 sg13g2_buf_8 fanout3332 (.A(net3333),
    .X(net3332));
 sg13g2_buf_8 fanout3333 (.A(net3335),
    .X(net3333));
 sg13g2_buf_8 fanout3334 (.A(net3335),
    .X(net3334));
 sg13g2_buf_8 fanout3335 (.A(net3339),
    .X(net3335));
 sg13g2_buf_8 fanout3336 (.A(net3339),
    .X(net3336));
 sg13g2_buf_1 fanout3337 (.A(net3339),
    .X(net3337));
 sg13g2_buf_8 fanout3338 (.A(net3339),
    .X(net3338));
 sg13g2_buf_8 fanout3339 (.A(_06640_),
    .X(net3339));
 sg13g2_buf_8 fanout3340 (.A(net3341),
    .X(net3340));
 sg13g2_buf_8 fanout3341 (.A(net3344),
    .X(net3341));
 sg13g2_buf_8 fanout3342 (.A(net3343),
    .X(net3342));
 sg13g2_buf_8 fanout3343 (.A(net3344),
    .X(net3343));
 sg13g2_buf_8 fanout3344 (.A(_06640_),
    .X(net3344));
 sg13g2_buf_8 fanout3345 (.A(net3346),
    .X(net3345));
 sg13g2_buf_8 fanout3346 (.A(net3351),
    .X(net3346));
 sg13g2_buf_8 fanout3347 (.A(net3351),
    .X(net3347));
 sg13g2_buf_8 fanout3348 (.A(net3350),
    .X(net3348));
 sg13g2_buf_1 fanout3349 (.A(net3350),
    .X(net3349));
 sg13g2_buf_8 fanout3350 (.A(net3351),
    .X(net3350));
 sg13g2_buf_8 fanout3351 (.A(net3375),
    .X(net3351));
 sg13g2_buf_8 fanout3352 (.A(net3353),
    .X(net3352));
 sg13g2_buf_8 fanout3353 (.A(net3375),
    .X(net3353));
 sg13g2_buf_8 fanout3354 (.A(net3355),
    .X(net3354));
 sg13g2_buf_1 fanout3355 (.A(net3356),
    .X(net3355));
 sg13g2_buf_1 fanout3356 (.A(net3357),
    .X(net3356));
 sg13g2_buf_1 fanout3357 (.A(net3358),
    .X(net3357));
 sg13g2_buf_8 fanout3358 (.A(net3375),
    .X(net3358));
 sg13g2_buf_8 fanout3359 (.A(net3360),
    .X(net3359));
 sg13g2_buf_8 fanout3360 (.A(net3364),
    .X(net3360));
 sg13g2_buf_8 fanout3361 (.A(net3363),
    .X(net3361));
 sg13g2_buf_8 fanout3362 (.A(net3363),
    .X(net3362));
 sg13g2_buf_8 fanout3363 (.A(net3364),
    .X(net3363));
 sg13g2_buf_8 fanout3364 (.A(net3374),
    .X(net3364));
 sg13g2_buf_8 fanout3365 (.A(net3374),
    .X(net3365));
 sg13g2_buf_8 fanout3366 (.A(net3374),
    .X(net3366));
 sg13g2_buf_8 fanout3367 (.A(net3373),
    .X(net3367));
 sg13g2_buf_8 fanout3368 (.A(net3373),
    .X(net3368));
 sg13g2_buf_8 fanout3369 (.A(net3373),
    .X(net3369));
 sg13g2_buf_8 fanout3370 (.A(net3371),
    .X(net3370));
 sg13g2_buf_8 fanout3371 (.A(net3372),
    .X(net3371));
 sg13g2_buf_8 fanout3372 (.A(net3373),
    .X(net3372));
 sg13g2_buf_8 fanout3373 (.A(net3374),
    .X(net3373));
 sg13g2_buf_8 fanout3374 (.A(net3375),
    .X(net3374));
 sg13g2_buf_8 fanout3375 (.A(_05890_),
    .X(net3375));
 sg13g2_buf_8 fanout3376 (.A(net3378),
    .X(net3376));
 sg13g2_buf_1 fanout3377 (.A(net3378),
    .X(net3377));
 sg13g2_buf_8 fanout3378 (.A(net3380),
    .X(net3378));
 sg13g2_buf_8 fanout3379 (.A(net3380),
    .X(net3379));
 sg13g2_buf_8 fanout3380 (.A(net3383),
    .X(net3380));
 sg13g2_buf_8 fanout3381 (.A(net3383),
    .X(net3381));
 sg13g2_buf_8 fanout3382 (.A(net3383),
    .X(net3382));
 sg13g2_buf_8 fanout3383 (.A(net3392),
    .X(net3383));
 sg13g2_buf_8 fanout3384 (.A(net3388),
    .X(net3384));
 sg13g2_buf_2 fanout3385 (.A(net3388),
    .X(net3385));
 sg13g2_buf_8 fanout3386 (.A(net3388),
    .X(net3386));
 sg13g2_buf_8 fanout3387 (.A(net3388),
    .X(net3387));
 sg13g2_buf_8 fanout3388 (.A(net3392),
    .X(net3388));
 sg13g2_buf_8 fanout3389 (.A(net3390),
    .X(net3389));
 sg13g2_buf_8 fanout3390 (.A(net3391),
    .X(net3390));
 sg13g2_buf_8 fanout3391 (.A(net3392),
    .X(net3391));
 sg13g2_buf_8 fanout3392 (.A(_05889_),
    .X(net3392));
 sg13g2_buf_8 fanout3393 (.A(net3397),
    .X(net3393));
 sg13g2_buf_1 fanout3394 (.A(net3397),
    .X(net3394));
 sg13g2_buf_8 fanout3395 (.A(net3397),
    .X(net3395));
 sg13g2_buf_1 fanout3396 (.A(net3397),
    .X(net3396));
 sg13g2_buf_8 fanout3397 (.A(net3409),
    .X(net3397));
 sg13g2_buf_8 fanout3398 (.A(net3399),
    .X(net3398));
 sg13g2_buf_8 fanout3399 (.A(net3409),
    .X(net3399));
 sg13g2_buf_8 fanout3400 (.A(net3401),
    .X(net3400));
 sg13g2_buf_8 fanout3401 (.A(net3404),
    .X(net3401));
 sg13g2_buf_8 fanout3402 (.A(net3403),
    .X(net3402));
 sg13g2_buf_8 fanout3403 (.A(net3404),
    .X(net3403));
 sg13g2_buf_8 fanout3404 (.A(net3409),
    .X(net3404));
 sg13g2_buf_8 fanout3405 (.A(net3406),
    .X(net3405));
 sg13g2_buf_8 fanout3406 (.A(net3408),
    .X(net3406));
 sg13g2_buf_8 fanout3407 (.A(net3408),
    .X(net3407));
 sg13g2_buf_2 fanout3408 (.A(net3409),
    .X(net3408));
 sg13g2_buf_8 fanout3409 (.A(_15649_),
    .X(net3409));
 sg13g2_buf_8 fanout3410 (.A(net3411),
    .X(net3410));
 sg13g2_buf_8 fanout3411 (.A(net3422),
    .X(net3411));
 sg13g2_buf_8 fanout3412 (.A(net3414),
    .X(net3412));
 sg13g2_buf_1 fanout3413 (.A(net3414),
    .X(net3413));
 sg13g2_buf_1 fanout3414 (.A(net3415),
    .X(net3414));
 sg13g2_buf_8 fanout3415 (.A(net3422),
    .X(net3415));
 sg13g2_buf_8 fanout3416 (.A(net3417),
    .X(net3416));
 sg13g2_buf_8 fanout3417 (.A(net3418),
    .X(net3417));
 sg13g2_buf_8 fanout3418 (.A(net3421),
    .X(net3418));
 sg13g2_buf_8 fanout3419 (.A(net3421),
    .X(net3419));
 sg13g2_buf_1 fanout3420 (.A(net3421),
    .X(net3420));
 sg13g2_buf_8 fanout3421 (.A(net3422),
    .X(net3421));
 sg13g2_buf_8 fanout3422 (.A(_15649_),
    .X(net3422));
 sg13g2_buf_8 fanout3423 (.A(net3425),
    .X(net3423));
 sg13g2_buf_8 fanout3424 (.A(net3425),
    .X(net3424));
 sg13g2_buf_8 fanout3425 (.A(net3426),
    .X(net3425));
 sg13g2_buf_8 fanout3426 (.A(net3432),
    .X(net3426));
 sg13g2_buf_8 fanout3427 (.A(net3432),
    .X(net3427));
 sg13g2_buf_8 fanout3428 (.A(net3432),
    .X(net3428));
 sg13g2_buf_8 fanout3429 (.A(net3431),
    .X(net3429));
 sg13g2_buf_8 fanout3430 (.A(net3431),
    .X(net3430));
 sg13g2_buf_8 fanout3431 (.A(net3432),
    .X(net3431));
 sg13g2_buf_8 fanout3432 (.A(net3447),
    .X(net3432));
 sg13g2_buf_8 fanout3433 (.A(net3434),
    .X(net3433));
 sg13g2_buf_8 fanout3434 (.A(net3447),
    .X(net3434));
 sg13g2_buf_8 fanout3435 (.A(net3441),
    .X(net3435));
 sg13g2_buf_8 fanout3436 (.A(net3441),
    .X(net3436));
 sg13g2_buf_1 fanout3437 (.A(net3438),
    .X(net3437));
 sg13g2_buf_8 fanout3438 (.A(net3441),
    .X(net3438));
 sg13g2_buf_8 fanout3439 (.A(net3440),
    .X(net3439));
 sg13g2_buf_8 fanout3440 (.A(net3441),
    .X(net3440));
 sg13g2_buf_8 fanout3441 (.A(net3447),
    .X(net3441));
 sg13g2_buf_8 fanout3442 (.A(net3446),
    .X(net3442));
 sg13g2_buf_8 fanout3443 (.A(net3446),
    .X(net3443));
 sg13g2_buf_1 fanout3444 (.A(net3445),
    .X(net3444));
 sg13g2_buf_8 fanout3445 (.A(net3446),
    .X(net3445));
 sg13g2_buf_8 fanout3446 (.A(net3447),
    .X(net3446));
 sg13g2_buf_8 fanout3447 (.A(net3466),
    .X(net3447));
 sg13g2_buf_8 fanout3448 (.A(net3459),
    .X(net3448));
 sg13g2_buf_8 fanout3449 (.A(net3459),
    .X(net3449));
 sg13g2_buf_8 fanout3450 (.A(net3451),
    .X(net3450));
 sg13g2_buf_8 fanout3451 (.A(net3453),
    .X(net3451));
 sg13g2_buf_8 fanout3452 (.A(net3453),
    .X(net3452));
 sg13g2_buf_8 fanout3453 (.A(net3459),
    .X(net3453));
 sg13g2_buf_8 fanout3454 (.A(net3455),
    .X(net3454));
 sg13g2_buf_8 fanout3455 (.A(net3459),
    .X(net3455));
 sg13g2_buf_8 fanout3456 (.A(net3458),
    .X(net3456));
 sg13g2_buf_8 fanout3457 (.A(net3458),
    .X(net3457));
 sg13g2_buf_8 fanout3458 (.A(net3459),
    .X(net3458));
 sg13g2_buf_8 fanout3459 (.A(net3466),
    .X(net3459));
 sg13g2_buf_8 fanout3460 (.A(net3461),
    .X(net3460));
 sg13g2_buf_8 fanout3461 (.A(net3466),
    .X(net3461));
 sg13g2_buf_8 fanout3462 (.A(net3465),
    .X(net3462));
 sg13g2_buf_1 fanout3463 (.A(net3465),
    .X(net3463));
 sg13g2_buf_8 fanout3464 (.A(net3465),
    .X(net3464));
 sg13g2_buf_8 fanout3465 (.A(net3466),
    .X(net3465));
 sg13g2_buf_8 fanout3466 (.A(_15649_),
    .X(net3466));
 sg13g2_buf_8 fanout3467 (.A(net3468),
    .X(net3467));
 sg13g2_buf_8 fanout3468 (.A(net3469),
    .X(net3468));
 sg13g2_buf_8 fanout3469 (.A(net3470),
    .X(net3469));
 sg13g2_buf_8 fanout3470 (.A(net3476),
    .X(net3470));
 sg13g2_buf_8 fanout3471 (.A(net3476),
    .X(net3471));
 sg13g2_buf_8 fanout3472 (.A(net3476),
    .X(net3472));
 sg13g2_buf_8 fanout3473 (.A(net3476),
    .X(net3473));
 sg13g2_buf_8 fanout3474 (.A(net3475),
    .X(net3474));
 sg13g2_buf_8 fanout3475 (.A(net3476),
    .X(net3475));
 sg13g2_buf_8 fanout3476 (.A(_15648_),
    .X(net3476));
 sg13g2_buf_8 fanout3477 (.A(net3478),
    .X(net3477));
 sg13g2_buf_8 fanout3478 (.A(net3479),
    .X(net3478));
 sg13g2_buf_8 fanout3479 (.A(net3488),
    .X(net3479));
 sg13g2_buf_8 fanout3480 (.A(net3481),
    .X(net3480));
 sg13g2_buf_8 fanout3481 (.A(net3483),
    .X(net3481));
 sg13g2_buf_8 fanout3482 (.A(net3483),
    .X(net3482));
 sg13g2_buf_8 fanout3483 (.A(net3488),
    .X(net3483));
 sg13g2_buf_8 fanout3484 (.A(net3486),
    .X(net3484));
 sg13g2_buf_8 fanout3485 (.A(net3486),
    .X(net3485));
 sg13g2_buf_8 fanout3486 (.A(net3487),
    .X(net3486));
 sg13g2_buf_8 fanout3487 (.A(net3488),
    .X(net3487));
 sg13g2_buf_8 fanout3488 (.A(_15648_),
    .X(net3488));
 sg13g2_buf_8 fanout3489 (.A(_05814_),
    .X(net3489));
 sg13g2_buf_8 fanout3490 (.A(_15647_),
    .X(net3490));
 sg13g2_buf_8 fanout3491 (.A(_15034_),
    .X(net3491));
 sg13g2_buf_8 fanout3492 (.A(_05794_),
    .X(net3492));
 sg13g2_buf_8 fanout3493 (.A(_05763_),
    .X(net3493));
 sg13g2_buf_8 fanout3494 (.A(net3502),
    .X(net3494));
 sg13g2_buf_8 fanout3495 (.A(net3496),
    .X(net3495));
 sg13g2_buf_8 fanout3496 (.A(net3502),
    .X(net3496));
 sg13g2_buf_8 fanout3497 (.A(net3498),
    .X(net3497));
 sg13g2_buf_8 fanout3498 (.A(net3499),
    .X(net3498));
 sg13g2_buf_8 fanout3499 (.A(net3501),
    .X(net3499));
 sg13g2_buf_8 fanout3500 (.A(net3501),
    .X(net3500));
 sg13g2_buf_8 fanout3501 (.A(net3502),
    .X(net3501));
 sg13g2_buf_8 fanout3502 (.A(net3585),
    .X(net3502));
 sg13g2_buf_8 fanout3503 (.A(net3514),
    .X(net3503));
 sg13g2_buf_1 fanout3504 (.A(net3514),
    .X(net3504));
 sg13g2_buf_8 fanout3505 (.A(net3507),
    .X(net3505));
 sg13g2_buf_8 fanout3506 (.A(net3507),
    .X(net3506));
 sg13g2_buf_8 fanout3507 (.A(net3514),
    .X(net3507));
 sg13g2_buf_8 fanout3508 (.A(net3511),
    .X(net3508));
 sg13g2_buf_1 fanout3509 (.A(net3511),
    .X(net3509));
 sg13g2_buf_8 fanout3510 (.A(net3511),
    .X(net3510));
 sg13g2_buf_8 fanout3511 (.A(net3514),
    .X(net3511));
 sg13g2_buf_8 fanout3512 (.A(net3513),
    .X(net3512));
 sg13g2_buf_8 fanout3513 (.A(net3514),
    .X(net3513));
 sg13g2_buf_8 fanout3514 (.A(net3585),
    .X(net3514));
 sg13g2_buf_8 fanout3515 (.A(net3516),
    .X(net3515));
 sg13g2_buf_8 fanout3516 (.A(net3519),
    .X(net3516));
 sg13g2_buf_8 fanout3517 (.A(net3518),
    .X(net3517));
 sg13g2_buf_8 fanout3518 (.A(net3519),
    .X(net3518));
 sg13g2_buf_8 fanout3519 (.A(net3537),
    .X(net3519));
 sg13g2_buf_8 fanout3520 (.A(net3523),
    .X(net3520));
 sg13g2_buf_8 fanout3521 (.A(net3523),
    .X(net3521));
 sg13g2_buf_1 fanout3522 (.A(net3523),
    .X(net3522));
 sg13g2_buf_8 fanout3523 (.A(net3537),
    .X(net3523));
 sg13g2_buf_8 fanout3524 (.A(net3527),
    .X(net3524));
 sg13g2_buf_8 fanout3525 (.A(net3527),
    .X(net3525));
 sg13g2_buf_1 fanout3526 (.A(net3527),
    .X(net3526));
 sg13g2_buf_8 fanout3527 (.A(net3537),
    .X(net3527));
 sg13g2_buf_8 fanout3528 (.A(net3532),
    .X(net3528));
 sg13g2_buf_8 fanout3529 (.A(net3531),
    .X(net3529));
 sg13g2_buf_8 fanout3530 (.A(net3531),
    .X(net3530));
 sg13g2_buf_8 fanout3531 (.A(net3532),
    .X(net3531));
 sg13g2_buf_8 fanout3532 (.A(net3537),
    .X(net3532));
 sg13g2_buf_8 fanout3533 (.A(net3534),
    .X(net3533));
 sg13g2_buf_8 fanout3534 (.A(net3537),
    .X(net3534));
 sg13g2_buf_8 fanout3535 (.A(net3536),
    .X(net3535));
 sg13g2_buf_8 fanout3536 (.A(net3537),
    .X(net3536));
 sg13g2_buf_8 fanout3537 (.A(net3585),
    .X(net3537));
 sg13g2_buf_8 fanout3538 (.A(net3543),
    .X(net3538));
 sg13g2_buf_8 fanout3539 (.A(net3543),
    .X(net3539));
 sg13g2_buf_8 fanout3540 (.A(net3542),
    .X(net3540));
 sg13g2_buf_8 fanout3541 (.A(net3542),
    .X(net3541));
 sg13g2_buf_8 fanout3542 (.A(net3543),
    .X(net3542));
 sg13g2_buf_8 fanout3543 (.A(net3548),
    .X(net3543));
 sg13g2_buf_8 fanout3544 (.A(net3548),
    .X(net3544));
 sg13g2_buf_1 fanout3545 (.A(net3548),
    .X(net3545));
 sg13g2_buf_8 fanout3546 (.A(net3547),
    .X(net3546));
 sg13g2_buf_1 fanout3547 (.A(net3548),
    .X(net3547));
 sg13g2_buf_8 fanout3548 (.A(net3584),
    .X(net3548));
 sg13g2_buf_8 fanout3549 (.A(net3551),
    .X(net3549));
 sg13g2_buf_1 fanout3550 (.A(net3551),
    .X(net3550));
 sg13g2_buf_8 fanout3551 (.A(net3555),
    .X(net3551));
 sg13g2_buf_8 fanout3552 (.A(net3553),
    .X(net3552));
 sg13g2_buf_8 fanout3553 (.A(net3555),
    .X(net3553));
 sg13g2_buf_8 fanout3554 (.A(net3555),
    .X(net3554));
 sg13g2_buf_8 fanout3555 (.A(net3584),
    .X(net3555));
 sg13g2_buf_8 fanout3556 (.A(net3560),
    .X(net3556));
 sg13g2_buf_8 fanout3557 (.A(net3560),
    .X(net3557));
 sg13g2_buf_1 fanout3558 (.A(net3559),
    .X(net3558));
 sg13g2_buf_8 fanout3559 (.A(net3560),
    .X(net3559));
 sg13g2_buf_8 fanout3560 (.A(net3584),
    .X(net3560));
 sg13g2_buf_8 fanout3561 (.A(net3562),
    .X(net3561));
 sg13g2_buf_8 fanout3562 (.A(net3571),
    .X(net3562));
 sg13g2_buf_8 fanout3563 (.A(net3564),
    .X(net3563));
 sg13g2_buf_8 fanout3564 (.A(net3565),
    .X(net3564));
 sg13g2_buf_8 fanout3565 (.A(net3571),
    .X(net3565));
 sg13g2_buf_8 fanout3566 (.A(net3567),
    .X(net3566));
 sg13g2_buf_8 fanout3567 (.A(net3571),
    .X(net3567));
 sg13g2_buf_8 fanout3568 (.A(net3570),
    .X(net3568));
 sg13g2_buf_1 fanout3569 (.A(net3570),
    .X(net3569));
 sg13g2_buf_8 fanout3570 (.A(net3571),
    .X(net3570));
 sg13g2_buf_8 fanout3571 (.A(net3584),
    .X(net3571));
 sg13g2_buf_8 fanout3572 (.A(net3583),
    .X(net3572));
 sg13g2_buf_1 fanout3573 (.A(net3574),
    .X(net3573));
 sg13g2_buf_8 fanout3574 (.A(net3575),
    .X(net3574));
 sg13g2_buf_8 fanout3575 (.A(net3583),
    .X(net3575));
 sg13g2_buf_8 fanout3576 (.A(net3578),
    .X(net3576));
 sg13g2_buf_1 fanout3577 (.A(net3578),
    .X(net3577));
 sg13g2_buf_8 fanout3578 (.A(net3583),
    .X(net3578));
 sg13g2_buf_8 fanout3579 (.A(net3582),
    .X(net3579));
 sg13g2_buf_1 fanout3580 (.A(net3582),
    .X(net3580));
 sg13g2_buf_8 fanout3581 (.A(net3582),
    .X(net3581));
 sg13g2_buf_8 fanout3582 (.A(net3583),
    .X(net3582));
 sg13g2_buf_8 fanout3583 (.A(net3584),
    .X(net3583));
 sg13g2_buf_8 fanout3584 (.A(net3585),
    .X(net3584));
 sg13g2_buf_8 fanout3585 (.A(_05431_),
    .X(net3585));
 sg13g2_buf_8 fanout3586 (.A(_15630_),
    .X(net3586));
 sg13g2_buf_8 fanout3587 (.A(net3595),
    .X(net3587));
 sg13g2_buf_8 fanout3588 (.A(net3589),
    .X(net3588));
 sg13g2_buf_8 fanout3589 (.A(net3595),
    .X(net3589));
 sg13g2_buf_8 fanout3590 (.A(net3591),
    .X(net3590));
 sg13g2_buf_8 fanout3591 (.A(net3592),
    .X(net3591));
 sg13g2_buf_8 fanout3592 (.A(net3594),
    .X(net3592));
 sg13g2_buf_8 fanout3593 (.A(net3594),
    .X(net3593));
 sg13g2_buf_8 fanout3594 (.A(net3595),
    .X(net3594));
 sg13g2_buf_8 fanout3595 (.A(net3678),
    .X(net3595));
 sg13g2_buf_8 fanout3596 (.A(net3607),
    .X(net3596));
 sg13g2_buf_1 fanout3597 (.A(net3607),
    .X(net3597));
 sg13g2_buf_8 fanout3598 (.A(net3600),
    .X(net3598));
 sg13g2_buf_8 fanout3599 (.A(net3600),
    .X(net3599));
 sg13g2_buf_8 fanout3600 (.A(net3607),
    .X(net3600));
 sg13g2_buf_8 fanout3601 (.A(net3604),
    .X(net3601));
 sg13g2_buf_2 fanout3602 (.A(net3604),
    .X(net3602));
 sg13g2_buf_8 fanout3603 (.A(net3604),
    .X(net3603));
 sg13g2_buf_8 fanout3604 (.A(net3607),
    .X(net3604));
 sg13g2_buf_8 fanout3605 (.A(net3606),
    .X(net3605));
 sg13g2_buf_8 fanout3606 (.A(net3607),
    .X(net3606));
 sg13g2_buf_8 fanout3607 (.A(net3678),
    .X(net3607));
 sg13g2_buf_8 fanout3608 (.A(net3609),
    .X(net3608));
 sg13g2_buf_8 fanout3609 (.A(net3612),
    .X(net3609));
 sg13g2_buf_8 fanout3610 (.A(net3611),
    .X(net3610));
 sg13g2_buf_8 fanout3611 (.A(net3612),
    .X(net3611));
 sg13g2_buf_8 fanout3612 (.A(net3630),
    .X(net3612));
 sg13g2_buf_8 fanout3613 (.A(net3616),
    .X(net3613));
 sg13g2_buf_8 fanout3614 (.A(net3616),
    .X(net3614));
 sg13g2_buf_1 fanout3615 (.A(net3616),
    .X(net3615));
 sg13g2_buf_8 fanout3616 (.A(net3630),
    .X(net3616));
 sg13g2_buf_8 fanout3617 (.A(net3620),
    .X(net3617));
 sg13g2_buf_8 fanout3618 (.A(net3620),
    .X(net3618));
 sg13g2_buf_1 fanout3619 (.A(net3620),
    .X(net3619));
 sg13g2_buf_8 fanout3620 (.A(net3630),
    .X(net3620));
 sg13g2_buf_8 fanout3621 (.A(net3625),
    .X(net3621));
 sg13g2_buf_8 fanout3622 (.A(net3624),
    .X(net3622));
 sg13g2_buf_8 fanout3623 (.A(net3624),
    .X(net3623));
 sg13g2_buf_8 fanout3624 (.A(net3625),
    .X(net3624));
 sg13g2_buf_8 fanout3625 (.A(net3630),
    .X(net3625));
 sg13g2_buf_8 fanout3626 (.A(net3627),
    .X(net3626));
 sg13g2_buf_8 fanout3627 (.A(net3630),
    .X(net3627));
 sg13g2_buf_8 fanout3628 (.A(net3629),
    .X(net3628));
 sg13g2_buf_8 fanout3629 (.A(net3630),
    .X(net3629));
 sg13g2_buf_8 fanout3630 (.A(net3678),
    .X(net3630));
 sg13g2_buf_8 fanout3631 (.A(net3636),
    .X(net3631));
 sg13g2_buf_8 fanout3632 (.A(net3636),
    .X(net3632));
 sg13g2_buf_8 fanout3633 (.A(net3635),
    .X(net3633));
 sg13g2_buf_8 fanout3634 (.A(net3635),
    .X(net3634));
 sg13g2_buf_8 fanout3635 (.A(net3636),
    .X(net3635));
 sg13g2_buf_8 fanout3636 (.A(net3641),
    .X(net3636));
 sg13g2_buf_8 fanout3637 (.A(net3641),
    .X(net3637));
 sg13g2_buf_1 fanout3638 (.A(net3641),
    .X(net3638));
 sg13g2_buf_8 fanout3639 (.A(net3640),
    .X(net3639));
 sg13g2_buf_2 fanout3640 (.A(net3641),
    .X(net3640));
 sg13g2_buf_8 fanout3641 (.A(net3677),
    .X(net3641));
 sg13g2_buf_8 fanout3642 (.A(net3644),
    .X(net3642));
 sg13g2_buf_1 fanout3643 (.A(net3644),
    .X(net3643));
 sg13g2_buf_8 fanout3644 (.A(net3648),
    .X(net3644));
 sg13g2_buf_8 fanout3645 (.A(net3646),
    .X(net3645));
 sg13g2_buf_8 fanout3646 (.A(net3648),
    .X(net3646));
 sg13g2_buf_8 fanout3647 (.A(net3648),
    .X(net3647));
 sg13g2_buf_8 fanout3648 (.A(net3677),
    .X(net3648));
 sg13g2_buf_8 fanout3649 (.A(net3653),
    .X(net3649));
 sg13g2_buf_8 fanout3650 (.A(net3653),
    .X(net3650));
 sg13g2_buf_1 fanout3651 (.A(net3652),
    .X(net3651));
 sg13g2_buf_8 fanout3652 (.A(net3653),
    .X(net3652));
 sg13g2_buf_8 fanout3653 (.A(net3677),
    .X(net3653));
 sg13g2_buf_8 fanout3654 (.A(net3655),
    .X(net3654));
 sg13g2_buf_8 fanout3655 (.A(net3664),
    .X(net3655));
 sg13g2_buf_8 fanout3656 (.A(net3657),
    .X(net3656));
 sg13g2_buf_8 fanout3657 (.A(net3658),
    .X(net3657));
 sg13g2_buf_8 fanout3658 (.A(net3664),
    .X(net3658));
 sg13g2_buf_8 fanout3659 (.A(net3660),
    .X(net3659));
 sg13g2_buf_8 fanout3660 (.A(net3664),
    .X(net3660));
 sg13g2_buf_8 fanout3661 (.A(net3663),
    .X(net3661));
 sg13g2_buf_2 fanout3662 (.A(net3663),
    .X(net3662));
 sg13g2_buf_8 fanout3663 (.A(net3664),
    .X(net3663));
 sg13g2_buf_8 fanout3664 (.A(net3677),
    .X(net3664));
 sg13g2_buf_8 fanout3665 (.A(net3676),
    .X(net3665));
 sg13g2_buf_1 fanout3666 (.A(net3667),
    .X(net3666));
 sg13g2_buf_8 fanout3667 (.A(net3668),
    .X(net3667));
 sg13g2_buf_8 fanout3668 (.A(net3676),
    .X(net3668));
 sg13g2_buf_8 fanout3669 (.A(net3671),
    .X(net3669));
 sg13g2_buf_1 fanout3670 (.A(net3671),
    .X(net3670));
 sg13g2_buf_8 fanout3671 (.A(net3676),
    .X(net3671));
 sg13g2_buf_8 fanout3672 (.A(net3675),
    .X(net3672));
 sg13g2_buf_1 fanout3673 (.A(net3675),
    .X(net3673));
 sg13g2_buf_8 fanout3674 (.A(net3675),
    .X(net3674));
 sg13g2_buf_8 fanout3675 (.A(net3676),
    .X(net3675));
 sg13g2_buf_8 fanout3676 (.A(net3677),
    .X(net3676));
 sg13g2_buf_8 fanout3677 (.A(net3678),
    .X(net3677));
 sg13g2_buf_8 fanout3678 (.A(_05434_),
    .X(net3678));
 sg13g2_buf_8 fanout3679 (.A(net3682),
    .X(net3679));
 sg13g2_buf_8 fanout3680 (.A(net3682),
    .X(net3680));
 sg13g2_buf_8 fanout3681 (.A(net3682),
    .X(net3681));
 sg13g2_buf_8 fanout3682 (.A(net3688),
    .X(net3682));
 sg13g2_buf_8 fanout3683 (.A(net3688),
    .X(net3683));
 sg13g2_buf_1 fanout3684 (.A(net3688),
    .X(net3684));
 sg13g2_buf_8 fanout3685 (.A(net3687),
    .X(net3685));
 sg13g2_buf_8 fanout3686 (.A(net3687),
    .X(net3686));
 sg13g2_buf_8 fanout3687 (.A(net3688),
    .X(net3687));
 sg13g2_buf_8 fanout3688 (.A(_05433_),
    .X(net3688));
 sg13g2_buf_8 fanout3689 (.A(net3690),
    .X(net3689));
 sg13g2_buf_8 fanout3690 (.A(net3692),
    .X(net3690));
 sg13g2_buf_8 fanout3691 (.A(net3692),
    .X(net3691));
 sg13g2_buf_8 fanout3692 (.A(net3700),
    .X(net3692));
 sg13g2_buf_8 fanout3693 (.A(net3694),
    .X(net3693));
 sg13g2_buf_8 fanout3694 (.A(net3700),
    .X(net3694));
 sg13g2_buf_8 fanout3695 (.A(net3696),
    .X(net3695));
 sg13g2_buf_8 fanout3696 (.A(net3700),
    .X(net3696));
 sg13g2_buf_8 fanout3697 (.A(net3699),
    .X(net3697));
 sg13g2_buf_8 fanout3698 (.A(net3699),
    .X(net3698));
 sg13g2_buf_8 fanout3699 (.A(net3700),
    .X(net3699));
 sg13g2_buf_8 fanout3700 (.A(_05432_),
    .X(net3700));
 sg13g2_buf_8 fanout3701 (.A(net3702),
    .X(net3701));
 sg13g2_buf_8 fanout3702 (.A(net3710),
    .X(net3702));
 sg13g2_buf_8 fanout3703 (.A(net3710),
    .X(net3703));
 sg13g2_buf_8 fanout3704 (.A(net3710),
    .X(net3704));
 sg13g2_buf_8 fanout3705 (.A(net3706),
    .X(net3705));
 sg13g2_buf_8 fanout3706 (.A(net3710),
    .X(net3706));
 sg13g2_buf_8 fanout3707 (.A(net3708),
    .X(net3707));
 sg13g2_buf_8 fanout3708 (.A(net3709),
    .X(net3708));
 sg13g2_buf_8 fanout3709 (.A(net3710),
    .X(net3709));
 sg13g2_buf_8 fanout3710 (.A(_05430_),
    .X(net3710));
 sg13g2_buf_8 fanout3711 (.A(net3713),
    .X(net3711));
 sg13g2_buf_8 fanout3712 (.A(net3713),
    .X(net3712));
 sg13g2_buf_8 fanout3713 (.A(_05429_),
    .X(net3713));
 sg13g2_buf_8 fanout3714 (.A(net3715),
    .X(net3714));
 sg13g2_buf_8 fanout3715 (.A(net3716),
    .X(net3715));
 sg13g2_buf_8 fanout3716 (.A(_05429_),
    .X(net3716));
 sg13g2_buf_8 fanout3717 (.A(net3721),
    .X(net3717));
 sg13g2_buf_8 fanout3718 (.A(net3719),
    .X(net3718));
 sg13g2_buf_8 fanout3719 (.A(net3720),
    .X(net3719));
 sg13g2_buf_8 fanout3720 (.A(net3721),
    .X(net3720));
 sg13g2_buf_8 fanout3721 (.A(_05429_),
    .X(net3721));
 sg13g2_buf_8 fanout3722 (.A(net3723),
    .X(net3722));
 sg13g2_buf_8 fanout3723 (.A(net3724),
    .X(net3723));
 sg13g2_buf_8 fanout3724 (.A(net3729),
    .X(net3724));
 sg13g2_buf_8 fanout3725 (.A(net3726),
    .X(net3725));
 sg13g2_buf_8 fanout3726 (.A(net3729),
    .X(net3726));
 sg13g2_buf_8 fanout3727 (.A(net3728),
    .X(net3727));
 sg13g2_buf_8 fanout3728 (.A(net3729),
    .X(net3728));
 sg13g2_buf_8 fanout3729 (.A(net3736),
    .X(net3729));
 sg13g2_buf_8 fanout3730 (.A(net3736),
    .X(net3730));
 sg13g2_buf_8 fanout3731 (.A(net3736),
    .X(net3731));
 sg13g2_buf_8 fanout3732 (.A(net3733),
    .X(net3732));
 sg13g2_buf_8 fanout3733 (.A(net3734),
    .X(net3733));
 sg13g2_buf_8 fanout3734 (.A(net3735),
    .X(net3734));
 sg13g2_buf_8 fanout3735 (.A(net3736),
    .X(net3735));
 sg13g2_buf_8 fanout3736 (.A(_12225_),
    .X(net3736));
 sg13g2_buf_8 fanout3737 (.A(net3738),
    .X(net3737));
 sg13g2_buf_8 fanout3738 (.A(net3743),
    .X(net3738));
 sg13g2_buf_8 fanout3739 (.A(net3740),
    .X(net3739));
 sg13g2_buf_2 fanout3740 (.A(net3741),
    .X(net3740));
 sg13g2_buf_8 fanout3741 (.A(net3743),
    .X(net3741));
 sg13g2_buf_8 fanout3742 (.A(net3743),
    .X(net3742));
 sg13g2_buf_8 fanout3743 (.A(net3776),
    .X(net3743));
 sg13g2_buf_8 fanout3744 (.A(net3745),
    .X(net3744));
 sg13g2_buf_8 fanout3745 (.A(net3751),
    .X(net3745));
 sg13g2_buf_8 fanout3746 (.A(net3751),
    .X(net3746));
 sg13g2_buf_8 fanout3747 (.A(net3748),
    .X(net3747));
 sg13g2_buf_2 fanout3748 (.A(net3751),
    .X(net3748));
 sg13g2_buf_8 fanout3749 (.A(net3751),
    .X(net3749));
 sg13g2_buf_2 fanout3750 (.A(net3751),
    .X(net3750));
 sg13g2_buf_8 fanout3751 (.A(net3776),
    .X(net3751));
 sg13g2_buf_8 fanout3752 (.A(net3754),
    .X(net3752));
 sg13g2_buf_1 fanout3753 (.A(net3754),
    .X(net3753));
 sg13g2_buf_8 fanout3754 (.A(net3776),
    .X(net3754));
 sg13g2_buf_8 fanout3755 (.A(net3756),
    .X(net3755));
 sg13g2_buf_8 fanout3756 (.A(net3758),
    .X(net3756));
 sg13g2_buf_8 fanout3757 (.A(net3758),
    .X(net3757));
 sg13g2_buf_8 fanout3758 (.A(net3761),
    .X(net3758));
 sg13g2_buf_8 fanout3759 (.A(net3760),
    .X(net3759));
 sg13g2_buf_8 fanout3760 (.A(net3761),
    .X(net3760));
 sg13g2_buf_2 fanout3761 (.A(net3775),
    .X(net3761));
 sg13g2_buf_8 fanout3762 (.A(net3764),
    .X(net3762));
 sg13g2_buf_8 fanout3763 (.A(net3764),
    .X(net3763));
 sg13g2_buf_8 fanout3764 (.A(net3775),
    .X(net3764));
 sg13g2_buf_8 fanout3765 (.A(net3767),
    .X(net3765));
 sg13g2_buf_2 fanout3766 (.A(net3767),
    .X(net3766));
 sg13g2_buf_8 fanout3767 (.A(net3773),
    .X(net3767));
 sg13g2_buf_8 fanout3768 (.A(net3770),
    .X(net3768));
 sg13g2_buf_1 fanout3769 (.A(net3770),
    .X(net3769));
 sg13g2_buf_8 fanout3770 (.A(net3773),
    .X(net3770));
 sg13g2_buf_8 fanout3771 (.A(net3773),
    .X(net3771));
 sg13g2_buf_2 fanout3772 (.A(net3773),
    .X(net3772));
 sg13g2_buf_8 fanout3773 (.A(net3775),
    .X(net3773));
 sg13g2_buf_8 fanout3774 (.A(net3775),
    .X(net3774));
 sg13g2_buf_8 fanout3775 (.A(net3776),
    .X(net3775));
 sg13g2_buf_8 fanout3776 (.A(_12222_),
    .X(net3776));
 sg13g2_buf_8 fanout3777 (.A(net3779),
    .X(net3777));
 sg13g2_buf_1 fanout3778 (.A(net3779),
    .X(net3778));
 sg13g2_buf_8 fanout3779 (.A(net3787),
    .X(net3779));
 sg13g2_buf_8 fanout3780 (.A(net3787),
    .X(net3780));
 sg13g2_buf_1 fanout3781 (.A(net3787),
    .X(net3781));
 sg13g2_buf_8 fanout3782 (.A(net3783),
    .X(net3782));
 sg13g2_buf_8 fanout3783 (.A(net3784),
    .X(net3783));
 sg13g2_buf_8 fanout3784 (.A(net3787),
    .X(net3784));
 sg13g2_buf_8 fanout3785 (.A(net3787),
    .X(net3785));
 sg13g2_buf_1 fanout3786 (.A(net3787),
    .X(net3786));
 sg13g2_buf_8 fanout3787 (.A(net3822),
    .X(net3787));
 sg13g2_buf_8 fanout3788 (.A(net3789),
    .X(net3788));
 sg13g2_buf_8 fanout3789 (.A(net3798),
    .X(net3789));
 sg13g2_buf_8 fanout3790 (.A(net3798),
    .X(net3790));
 sg13g2_buf_1 fanout3791 (.A(net3798),
    .X(net3791));
 sg13g2_buf_8 fanout3792 (.A(net3794),
    .X(net3792));
 sg13g2_buf_1 fanout3793 (.A(net3794),
    .X(net3793));
 sg13g2_buf_8 fanout3794 (.A(net3797),
    .X(net3794));
 sg13g2_buf_8 fanout3795 (.A(net3797),
    .X(net3795));
 sg13g2_buf_8 fanout3796 (.A(net3797),
    .X(net3796));
 sg13g2_buf_8 fanout3797 (.A(net3798),
    .X(net3797));
 sg13g2_buf_8 fanout3798 (.A(net3803),
    .X(net3798));
 sg13g2_buf_8 fanout3799 (.A(net3803),
    .X(net3799));
 sg13g2_buf_8 fanout3800 (.A(net3802),
    .X(net3800));
 sg13g2_buf_1 fanout3801 (.A(net3802),
    .X(net3801));
 sg13g2_buf_8 fanout3802 (.A(net3803),
    .X(net3802));
 sg13g2_buf_8 fanout3803 (.A(net3822),
    .X(net3803));
 sg13g2_buf_8 fanout3804 (.A(net3805),
    .X(net3804));
 sg13g2_buf_8 fanout3805 (.A(net3806),
    .X(net3805));
 sg13g2_buf_8 fanout3806 (.A(net3811),
    .X(net3806));
 sg13g2_buf_8 fanout3807 (.A(net3809),
    .X(net3807));
 sg13g2_buf_1 fanout3808 (.A(net3809),
    .X(net3808));
 sg13g2_buf_8 fanout3809 (.A(net3811),
    .X(net3809));
 sg13g2_buf_8 fanout3810 (.A(net3811),
    .X(net3810));
 sg13g2_buf_8 fanout3811 (.A(net3822),
    .X(net3811));
 sg13g2_buf_8 fanout3812 (.A(net3813),
    .X(net3812));
 sg13g2_buf_8 fanout3813 (.A(net3815),
    .X(net3813));
 sg13g2_buf_8 fanout3814 (.A(net3815),
    .X(net3814));
 sg13g2_buf_8 fanout3815 (.A(net3822),
    .X(net3815));
 sg13g2_buf_8 fanout3816 (.A(net3817),
    .X(net3816));
 sg13g2_buf_8 fanout3817 (.A(net3819),
    .X(net3817));
 sg13g2_buf_8 fanout3818 (.A(net3819),
    .X(net3818));
 sg13g2_buf_8 fanout3819 (.A(net3821),
    .X(net3819));
 sg13g2_buf_8 fanout3820 (.A(net3821),
    .X(net3820));
 sg13g2_buf_8 fanout3821 (.A(net3822),
    .X(net3821));
 sg13g2_buf_8 fanout3822 (.A(_12222_),
    .X(net3822));
 sg13g2_buf_8 fanout3823 (.A(net3834),
    .X(net3823));
 sg13g2_buf_1 fanout3824 (.A(net3834),
    .X(net3824));
 sg13g2_buf_8 fanout3825 (.A(net3826),
    .X(net3825));
 sg13g2_buf_8 fanout3826 (.A(net3827),
    .X(net3826));
 sg13g2_buf_8 fanout3827 (.A(net3828),
    .X(net3827));
 sg13g2_buf_8 fanout3828 (.A(net3834),
    .X(net3828));
 sg13g2_buf_8 fanout3829 (.A(net3834),
    .X(net3829));
 sg13g2_buf_2 fanout3830 (.A(net3834),
    .X(net3830));
 sg13g2_buf_8 fanout3831 (.A(net3832),
    .X(net3831));
 sg13g2_buf_8 fanout3832 (.A(net3833),
    .X(net3832));
 sg13g2_buf_8 fanout3833 (.A(net3834),
    .X(net3833));
 sg13g2_buf_8 fanout3834 (.A(_12221_),
    .X(net3834));
 sg13g2_buf_8 fanout3835 (.A(net3848),
    .X(net3835));
 sg13g2_buf_8 fanout3836 (.A(net3848),
    .X(net3836));
 sg13g2_buf_8 fanout3837 (.A(net3838),
    .X(net3837));
 sg13g2_buf_8 fanout3838 (.A(net3840),
    .X(net3838));
 sg13g2_buf_8 fanout3839 (.A(net3840),
    .X(net3839));
 sg13g2_buf_8 fanout3840 (.A(net3848),
    .X(net3840));
 sg13g2_buf_8 fanout3841 (.A(net3842),
    .X(net3841));
 sg13g2_buf_8 fanout3842 (.A(net3847),
    .X(net3842));
 sg13g2_buf_8 fanout3843 (.A(net3846),
    .X(net3843));
 sg13g2_buf_2 fanout3844 (.A(net3846),
    .X(net3844));
 sg13g2_buf_8 fanout3845 (.A(net3846),
    .X(net3845));
 sg13g2_buf_8 fanout3846 (.A(net3847),
    .X(net3846));
 sg13g2_buf_8 fanout3847 (.A(net3848),
    .X(net3847));
 sg13g2_buf_8 fanout3848 (.A(_12221_),
    .X(net3848));
 sg13g2_buf_8 fanout3849 (.A(net3850),
    .X(net3849));
 sg13g2_buf_8 fanout3850 (.A(net3858),
    .X(net3850));
 sg13g2_buf_8 fanout3851 (.A(net3852),
    .X(net3851));
 sg13g2_buf_8 fanout3852 (.A(net3858),
    .X(net3852));
 sg13g2_buf_8 fanout3853 (.A(net3854),
    .X(net3853));
 sg13g2_buf_8 fanout3854 (.A(net3857),
    .X(net3854));
 sg13g2_buf_8 fanout3855 (.A(net3857),
    .X(net3855));
 sg13g2_buf_8 fanout3856 (.A(net3857),
    .X(net3856));
 sg13g2_buf_8 fanout3857 (.A(net3858),
    .X(net3857));
 sg13g2_buf_8 fanout3858 (.A(net3873),
    .X(net3858));
 sg13g2_buf_8 fanout3859 (.A(net3864),
    .X(net3859));
 sg13g2_buf_8 fanout3860 (.A(net3863),
    .X(net3860));
 sg13g2_buf_8 fanout3861 (.A(net3862),
    .X(net3861));
 sg13g2_buf_8 fanout3862 (.A(net3863),
    .X(net3862));
 sg13g2_buf_8 fanout3863 (.A(net3864),
    .X(net3863));
 sg13g2_buf_8 fanout3864 (.A(net3873),
    .X(net3864));
 sg13g2_buf_8 fanout3865 (.A(net3866),
    .X(net3865));
 sg13g2_buf_8 fanout3866 (.A(net3868),
    .X(net3866));
 sg13g2_buf_1 fanout3867 (.A(net3868),
    .X(net3867));
 sg13g2_buf_8 fanout3868 (.A(net3873),
    .X(net3868));
 sg13g2_buf_8 fanout3869 (.A(net3872),
    .X(net3869));
 sg13g2_buf_8 fanout3870 (.A(net3872),
    .X(net3870));
 sg13g2_buf_8 fanout3871 (.A(net3872),
    .X(net3871));
 sg13g2_buf_8 fanout3872 (.A(net3873),
    .X(net3872));
 sg13g2_buf_8 fanout3873 (.A(_12221_),
    .X(net3873));
 sg13g2_buf_8 fanout3874 (.A(net3875),
    .X(net3874));
 sg13g2_buf_8 fanout3875 (.A(net3877),
    .X(net3875));
 sg13g2_buf_8 fanout3876 (.A(net3877),
    .X(net3876));
 sg13g2_buf_8 fanout3877 (.A(net3889),
    .X(net3877));
 sg13g2_buf_8 fanout3878 (.A(net3879),
    .X(net3878));
 sg13g2_buf_8 fanout3879 (.A(net3880),
    .X(net3879));
 sg13g2_buf_8 fanout3880 (.A(net3889),
    .X(net3880));
 sg13g2_buf_1 fanout3881 (.A(net3889),
    .X(net3881));
 sg13g2_buf_8 fanout3882 (.A(net3884),
    .X(net3882));
 sg13g2_buf_8 fanout3883 (.A(net3884),
    .X(net3883));
 sg13g2_buf_8 fanout3884 (.A(net3888),
    .X(net3884));
 sg13g2_buf_8 fanout3885 (.A(net3886),
    .X(net3885));
 sg13g2_buf_8 fanout3886 (.A(net3887),
    .X(net3886));
 sg13g2_buf_8 fanout3887 (.A(net3888),
    .X(net3887));
 sg13g2_buf_8 fanout3888 (.A(net3889),
    .X(net3888));
 sg13g2_buf_8 fanout3889 (.A(_12817_),
    .X(net3889));
 sg13g2_buf_8 fanout3890 (.A(net3895),
    .X(net3890));
 sg13g2_buf_2 fanout3891 (.A(net3895),
    .X(net3891));
 sg13g2_buf_8 fanout3892 (.A(net3893),
    .X(net3892));
 sg13g2_buf_8 fanout3893 (.A(net3895),
    .X(net3893));
 sg13g2_buf_8 fanout3894 (.A(net3895),
    .X(net3894));
 sg13g2_buf_8 fanout3895 (.A(net3911),
    .X(net3895));
 sg13g2_buf_8 fanout3896 (.A(net3899),
    .X(net3896));
 sg13g2_buf_8 fanout3897 (.A(net3899),
    .X(net3897));
 sg13g2_buf_1 fanout3898 (.A(net3899),
    .X(net3898));
 sg13g2_buf_8 fanout3899 (.A(net3911),
    .X(net3899));
 sg13g2_buf_8 fanout3900 (.A(net3902),
    .X(net3900));
 sg13g2_buf_1 fanout3901 (.A(net3902),
    .X(net3901));
 sg13g2_buf_8 fanout3902 (.A(net3911),
    .X(net3902));
 sg13g2_buf_8 fanout3903 (.A(net3904),
    .X(net3903));
 sg13g2_buf_8 fanout3904 (.A(net3905),
    .X(net3904));
 sg13g2_buf_8 fanout3905 (.A(net3910),
    .X(net3905));
 sg13g2_buf_8 fanout3906 (.A(net3910),
    .X(net3906));
 sg13g2_buf_8 fanout3907 (.A(net3908),
    .X(net3907));
 sg13g2_buf_2 fanout3908 (.A(net3910),
    .X(net3908));
 sg13g2_buf_8 fanout3909 (.A(net3910),
    .X(net3909));
 sg13g2_buf_8 fanout3910 (.A(net3911),
    .X(net3910));
 sg13g2_buf_8 fanout3911 (.A(_12817_),
    .X(net3911));
 sg13g2_buf_8 fanout3912 (.A(net3913),
    .X(net3912));
 sg13g2_buf_8 fanout3913 (.A(net3914),
    .X(net3913));
 sg13g2_buf_8 fanout3914 (.A(net3920),
    .X(net3914));
 sg13g2_buf_8 fanout3915 (.A(net3916),
    .X(net3915));
 sg13g2_buf_8 fanout3916 (.A(net3920),
    .X(net3916));
 sg13g2_buf_8 fanout3917 (.A(net3920),
    .X(net3917));
 sg13g2_buf_8 fanout3918 (.A(net3919),
    .X(net3918));
 sg13g2_buf_8 fanout3919 (.A(net3920),
    .X(net3919));
 sg13g2_buf_8 fanout3920 (.A(net3999),
    .X(net3920));
 sg13g2_buf_8 fanout3921 (.A(net3925),
    .X(net3921));
 sg13g2_buf_1 fanout3922 (.A(net3925),
    .X(net3922));
 sg13g2_buf_8 fanout3923 (.A(net3924),
    .X(net3923));
 sg13g2_buf_8 fanout3924 (.A(net3925),
    .X(net3924));
 sg13g2_buf_8 fanout3925 (.A(net3931),
    .X(net3925));
 sg13g2_buf_8 fanout3926 (.A(net3928),
    .X(net3926));
 sg13g2_buf_8 fanout3927 (.A(net3928),
    .X(net3927));
 sg13g2_buf_8 fanout3928 (.A(net3931),
    .X(net3928));
 sg13g2_buf_8 fanout3929 (.A(net3931),
    .X(net3929));
 sg13g2_buf_1 fanout3930 (.A(net3931),
    .X(net3930));
 sg13g2_buf_8 fanout3931 (.A(net3999),
    .X(net3931));
 sg13g2_buf_8 fanout3932 (.A(net3933),
    .X(net3932));
 sg13g2_buf_8 fanout3933 (.A(net3935),
    .X(net3933));
 sg13g2_buf_8 fanout3934 (.A(net3935),
    .X(net3934));
 sg13g2_buf_8 fanout3935 (.A(net3952),
    .X(net3935));
 sg13g2_buf_8 fanout3936 (.A(net3942),
    .X(net3936));
 sg13g2_buf_1 fanout3937 (.A(net3938),
    .X(net3937));
 sg13g2_buf_8 fanout3938 (.A(net3942),
    .X(net3938));
 sg13g2_buf_8 fanout3939 (.A(net3940),
    .X(net3939));
 sg13g2_buf_8 fanout3940 (.A(net3942),
    .X(net3940));
 sg13g2_buf_8 fanout3941 (.A(net3942),
    .X(net3941));
 sg13g2_buf_8 fanout3942 (.A(net3952),
    .X(net3942));
 sg13g2_buf_8 fanout3943 (.A(net3946),
    .X(net3943));
 sg13g2_buf_8 fanout3944 (.A(net3946),
    .X(net3944));
 sg13g2_buf_8 fanout3945 (.A(net3946),
    .X(net3945));
 sg13g2_buf_8 fanout3946 (.A(net3952),
    .X(net3946));
 sg13g2_buf_8 fanout3947 (.A(net3951),
    .X(net3947));
 sg13g2_buf_8 fanout3948 (.A(net3949),
    .X(net3948));
 sg13g2_buf_8 fanout3949 (.A(net3951),
    .X(net3949));
 sg13g2_buf_8 fanout3950 (.A(net3951),
    .X(net3950));
 sg13g2_buf_8 fanout3951 (.A(net3952),
    .X(net3951));
 sg13g2_buf_8 fanout3952 (.A(net3999),
    .X(net3952));
 sg13g2_buf_8 fanout3953 (.A(net3964),
    .X(net3953));
 sg13g2_buf_8 fanout3954 (.A(net3964),
    .X(net3954));
 sg13g2_buf_8 fanout3955 (.A(net3957),
    .X(net3955));
 sg13g2_buf_8 fanout3956 (.A(net3957),
    .X(net3956));
 sg13g2_buf_8 fanout3957 (.A(net3964),
    .X(net3957));
 sg13g2_buf_8 fanout3958 (.A(net3959),
    .X(net3958));
 sg13g2_buf_8 fanout3959 (.A(net3963),
    .X(net3959));
 sg13g2_buf_8 fanout3960 (.A(net3963),
    .X(net3960));
 sg13g2_buf_1 fanout3961 (.A(net3963),
    .X(net3961));
 sg13g2_buf_8 fanout3962 (.A(net3963),
    .X(net3962));
 sg13g2_buf_8 fanout3963 (.A(net3964),
    .X(net3963));
 sg13g2_buf_8 fanout3964 (.A(net3998),
    .X(net3964));
 sg13g2_buf_8 fanout3965 (.A(net3970),
    .X(net3965));
 sg13g2_buf_2 fanout3966 (.A(net3970),
    .X(net3966));
 sg13g2_buf_8 fanout3967 (.A(net3968),
    .X(net3967));
 sg13g2_buf_8 fanout3968 (.A(net3970),
    .X(net3968));
 sg13g2_buf_1 fanout3969 (.A(net3970),
    .X(net3969));
 sg13g2_buf_8 fanout3970 (.A(net3998),
    .X(net3970));
 sg13g2_buf_8 fanout3971 (.A(net3975),
    .X(net3971));
 sg13g2_buf_8 fanout3972 (.A(net3974),
    .X(net3972));
 sg13g2_buf_1 fanout3973 (.A(net3974),
    .X(net3973));
 sg13g2_buf_8 fanout3974 (.A(net3975),
    .X(net3974));
 sg13g2_buf_8 fanout3975 (.A(net3998),
    .X(net3975));
 sg13g2_buf_8 fanout3976 (.A(net3977),
    .X(net3976));
 sg13g2_buf_8 fanout3977 (.A(net3979),
    .X(net3977));
 sg13g2_buf_8 fanout3978 (.A(net3979),
    .X(net3978));
 sg13g2_buf_8 fanout3979 (.A(net3997),
    .X(net3979));
 sg13g2_buf_8 fanout3980 (.A(net3981),
    .X(net3980));
 sg13g2_buf_8 fanout3981 (.A(net3997),
    .X(net3981));
 sg13g2_buf_8 fanout3982 (.A(net3984),
    .X(net3982));
 sg13g2_buf_2 fanout3983 (.A(net3984),
    .X(net3983));
 sg13g2_buf_8 fanout3984 (.A(net3997),
    .X(net3984));
 sg13g2_buf_8 fanout3985 (.A(net3996),
    .X(net3985));
 sg13g2_buf_8 fanout3986 (.A(net3990),
    .X(net3986));
 sg13g2_buf_1 fanout3987 (.A(net3990),
    .X(net3987));
 sg13g2_buf_8 fanout3988 (.A(net3990),
    .X(net3988));
 sg13g2_buf_8 fanout3989 (.A(net3990),
    .X(net3989));
 sg13g2_buf_8 fanout3990 (.A(net3996),
    .X(net3990));
 sg13g2_buf_8 fanout3991 (.A(net3992),
    .X(net3991));
 sg13g2_buf_8 fanout3992 (.A(net3996),
    .X(net3992));
 sg13g2_buf_8 fanout3993 (.A(net3995),
    .X(net3993));
 sg13g2_buf_2 fanout3994 (.A(net3995),
    .X(net3994));
 sg13g2_buf_8 fanout3995 (.A(net3996),
    .X(net3995));
 sg13g2_buf_8 fanout3996 (.A(net3997),
    .X(net3996));
 sg13g2_buf_8 fanout3997 (.A(net3998),
    .X(net3997));
 sg13g2_buf_8 fanout3998 (.A(net3999),
    .X(net3998));
 sg13g2_buf_8 fanout3999 (.A(_11067_),
    .X(net3999));
 sg13g2_buf_8 fanout4000 (.A(net4004),
    .X(net4000));
 sg13g2_buf_1 fanout4001 (.A(net4004),
    .X(net4001));
 sg13g2_buf_8 fanout4002 (.A(net4004),
    .X(net4002));
 sg13g2_buf_1 fanout4003 (.A(net4004),
    .X(net4003));
 sg13g2_buf_8 fanout4004 (.A(net4005),
    .X(net4004));
 sg13g2_buf_8 fanout4005 (.A(net4026),
    .X(net4005));
 sg13g2_buf_8 fanout4006 (.A(net4010),
    .X(net4006));
 sg13g2_buf_1 fanout4007 (.A(net4010),
    .X(net4007));
 sg13g2_buf_8 fanout4008 (.A(net4010),
    .X(net4008));
 sg13g2_buf_1 fanout4009 (.A(net4010),
    .X(net4009));
 sg13g2_buf_8 fanout4010 (.A(net4013),
    .X(net4010));
 sg13g2_buf_8 fanout4011 (.A(net4012),
    .X(net4011));
 sg13g2_buf_8 fanout4012 (.A(net4013),
    .X(net4012));
 sg13g2_buf_8 fanout4013 (.A(net4026),
    .X(net4013));
 sg13g2_buf_8 fanout4014 (.A(net4019),
    .X(net4014));
 sg13g2_buf_8 fanout4015 (.A(net4016),
    .X(net4015));
 sg13g2_buf_8 fanout4016 (.A(net4019),
    .X(net4016));
 sg13g2_buf_8 fanout4017 (.A(net4019),
    .X(net4017));
 sg13g2_buf_1 fanout4018 (.A(net4019),
    .X(net4018));
 sg13g2_buf_8 fanout4019 (.A(net4026),
    .X(net4019));
 sg13g2_buf_8 fanout4020 (.A(net4022),
    .X(net4020));
 sg13g2_buf_8 fanout4021 (.A(net4022),
    .X(net4021));
 sg13g2_buf_8 fanout4022 (.A(net4024),
    .X(net4022));
 sg13g2_buf_8 fanout4023 (.A(net4024),
    .X(net4023));
 sg13g2_buf_8 fanout4024 (.A(net4025),
    .X(net4024));
 sg13g2_buf_8 fanout4025 (.A(net4026),
    .X(net4025));
 sg13g2_buf_8 fanout4026 (.A(net4052),
    .X(net4026));
 sg13g2_buf_8 fanout4027 (.A(net4028),
    .X(net4027));
 sg13g2_buf_8 fanout4028 (.A(net4029),
    .X(net4028));
 sg13g2_buf_8 fanout4029 (.A(net4052),
    .X(net4029));
 sg13g2_buf_8 fanout4030 (.A(net4033),
    .X(net4030));
 sg13g2_buf_8 fanout4031 (.A(net4032),
    .X(net4031));
 sg13g2_buf_8 fanout4032 (.A(net4033),
    .X(net4032));
 sg13g2_buf_2 fanout4033 (.A(net4034),
    .X(net4033));
 sg13g2_buf_8 fanout4034 (.A(net4052),
    .X(net4034));
 sg13g2_buf_8 fanout4035 (.A(net4038),
    .X(net4035));
 sg13g2_buf_8 fanout4036 (.A(net4037),
    .X(net4036));
 sg13g2_buf_8 fanout4037 (.A(net4038),
    .X(net4037));
 sg13g2_buf_8 fanout4038 (.A(net4051),
    .X(net4038));
 sg13g2_buf_8 fanout4039 (.A(net4042),
    .X(net4039));
 sg13g2_buf_8 fanout4040 (.A(net4042),
    .X(net4040));
 sg13g2_buf_8 fanout4041 (.A(net4042),
    .X(net4041));
 sg13g2_buf_8 fanout4042 (.A(net4043),
    .X(net4042));
 sg13g2_buf_8 fanout4043 (.A(net4051),
    .X(net4043));
 sg13g2_buf_8 fanout4044 (.A(net4045),
    .X(net4044));
 sg13g2_buf_2 fanout4045 (.A(net4046),
    .X(net4045));
 sg13g2_buf_2 fanout4046 (.A(net4051),
    .X(net4046));
 sg13g2_buf_8 fanout4047 (.A(net4048),
    .X(net4047));
 sg13g2_buf_8 fanout4048 (.A(net4050),
    .X(net4048));
 sg13g2_buf_8 fanout4049 (.A(net4050),
    .X(net4049));
 sg13g2_buf_8 fanout4050 (.A(net4051),
    .X(net4050));
 sg13g2_buf_8 fanout4051 (.A(net4052),
    .X(net4051));
 sg13g2_buf_8 fanout4052 (.A(_11066_),
    .X(net4052));
 sg13g2_buf_8 fanout4053 (.A(net4063),
    .X(net4053));
 sg13g2_buf_1 fanout4054 (.A(net4063),
    .X(net4054));
 sg13g2_buf_8 fanout4055 (.A(net4056),
    .X(net4055));
 sg13g2_buf_8 fanout4056 (.A(net4057),
    .X(net4056));
 sg13g2_buf_1 fanout4057 (.A(net4063),
    .X(net4057));
 sg13g2_buf_8 fanout4058 (.A(net4059),
    .X(net4058));
 sg13g2_buf_8 fanout4059 (.A(net4063),
    .X(net4059));
 sg13g2_buf_8 fanout4060 (.A(net4061),
    .X(net4060));
 sg13g2_buf_1 fanout4061 (.A(net4062),
    .X(net4061));
 sg13g2_buf_1 fanout4062 (.A(net4063),
    .X(net4062));
 sg13g2_buf_8 fanout4063 (.A(net4072),
    .X(net4063));
 sg13g2_buf_8 fanout4064 (.A(net4066),
    .X(net4064));
 sg13g2_buf_8 fanout4065 (.A(net4066),
    .X(net4065));
 sg13g2_buf_8 fanout4066 (.A(net4067),
    .X(net4066));
 sg13g2_buf_8 fanout4067 (.A(net4072),
    .X(net4067));
 sg13g2_buf_8 fanout4068 (.A(net4069),
    .X(net4068));
 sg13g2_buf_8 fanout4069 (.A(net4070),
    .X(net4069));
 sg13g2_buf_8 fanout4070 (.A(net4071),
    .X(net4070));
 sg13g2_buf_8 fanout4071 (.A(net4072),
    .X(net4071));
 sg13g2_buf_8 fanout4072 (.A(_12822_),
    .X(net4072));
 sg13g2_buf_8 fanout4073 (.A(net4076),
    .X(net4073));
 sg13g2_buf_8 fanout4074 (.A(net4076),
    .X(net4074));
 sg13g2_buf_1 fanout4075 (.A(net4076),
    .X(net4075));
 sg13g2_buf_8 fanout4076 (.A(net4093),
    .X(net4076));
 sg13g2_buf_8 fanout4077 (.A(net4081),
    .X(net4077));
 sg13g2_buf_8 fanout4078 (.A(net4081),
    .X(net4078));
 sg13g2_buf_8 fanout4079 (.A(net4080),
    .X(net4079));
 sg13g2_buf_8 fanout4080 (.A(net4081),
    .X(net4080));
 sg13g2_buf_8 fanout4081 (.A(net4093),
    .X(net4081));
 sg13g2_buf_8 fanout4082 (.A(net4084),
    .X(net4082));
 sg13g2_buf_1 fanout4083 (.A(net4084),
    .X(net4083));
 sg13g2_buf_8 fanout4084 (.A(net4085),
    .X(net4084));
 sg13g2_buf_8 fanout4085 (.A(net4087),
    .X(net4085));
 sg13g2_buf_8 fanout4086 (.A(net4087),
    .X(net4086));
 sg13g2_buf_8 fanout4087 (.A(net4093),
    .X(net4087));
 sg13g2_buf_8 fanout4088 (.A(net4092),
    .X(net4088));
 sg13g2_buf_8 fanout4089 (.A(net4090),
    .X(net4089));
 sg13g2_buf_2 fanout4090 (.A(net4091),
    .X(net4090));
 sg13g2_buf_8 fanout4091 (.A(net4092),
    .X(net4091));
 sg13g2_buf_2 fanout4092 (.A(net4093),
    .X(net4092));
 sg13g2_buf_8 fanout4093 (.A(_12822_),
    .X(net4093));
 sg13g2_buf_8 fanout4094 (.A(net4104),
    .X(net4094));
 sg13g2_buf_8 fanout4095 (.A(net4096),
    .X(net4095));
 sg13g2_buf_8 fanout4096 (.A(net4098),
    .X(net4096));
 sg13g2_buf_8 fanout4097 (.A(net4098),
    .X(net4097));
 sg13g2_buf_8 fanout4098 (.A(net4099),
    .X(net4098));
 sg13g2_buf_2 fanout4099 (.A(net4104),
    .X(net4099));
 sg13g2_buf_8 fanout4100 (.A(net4103),
    .X(net4100));
 sg13g2_buf_8 fanout4101 (.A(net4103),
    .X(net4101));
 sg13g2_buf_8 fanout4102 (.A(net4103),
    .X(net4102));
 sg13g2_buf_8 fanout4103 (.A(net4104),
    .X(net4103));
 sg13g2_buf_8 fanout4104 (.A(net4143),
    .X(net4104));
 sg13g2_buf_8 fanout4105 (.A(net4106),
    .X(net4105));
 sg13g2_buf_8 fanout4106 (.A(net4109),
    .X(net4106));
 sg13g2_buf_8 fanout4107 (.A(net4109),
    .X(net4107));
 sg13g2_buf_1 fanout4108 (.A(net4109),
    .X(net4108));
 sg13g2_buf_2 fanout4109 (.A(net4114),
    .X(net4109));
 sg13g2_buf_8 fanout4110 (.A(net4111),
    .X(net4110));
 sg13g2_buf_2 fanout4111 (.A(net4112),
    .X(net4111));
 sg13g2_buf_1 fanout4112 (.A(net4114),
    .X(net4112));
 sg13g2_buf_8 fanout4113 (.A(net4114),
    .X(net4113));
 sg13g2_buf_1 fanout4114 (.A(net4143),
    .X(net4114));
 sg13g2_buf_8 fanout4115 (.A(net4120),
    .X(net4115));
 sg13g2_buf_1 fanout4116 (.A(net4120),
    .X(net4116));
 sg13g2_buf_8 fanout4117 (.A(net4119),
    .X(net4117));
 sg13g2_buf_2 fanout4118 (.A(net4119),
    .X(net4118));
 sg13g2_buf_8 fanout4119 (.A(net4120),
    .X(net4119));
 sg13g2_buf_2 fanout4120 (.A(net4143),
    .X(net4120));
 sg13g2_buf_8 fanout4121 (.A(net4122),
    .X(net4121));
 sg13g2_buf_8 fanout4122 (.A(net4125),
    .X(net4122));
 sg13g2_buf_8 fanout4123 (.A(net4124),
    .X(net4123));
 sg13g2_buf_8 fanout4124 (.A(net4125),
    .X(net4124));
 sg13g2_buf_8 fanout4125 (.A(net4142),
    .X(net4125));
 sg13g2_buf_8 fanout4126 (.A(net4128),
    .X(net4126));
 sg13g2_buf_1 fanout4127 (.A(net4128),
    .X(net4127));
 sg13g2_buf_8 fanout4128 (.A(net4129),
    .X(net4128));
 sg13g2_buf_8 fanout4129 (.A(net4142),
    .X(net4129));
 sg13g2_buf_8 fanout4130 (.A(net4131),
    .X(net4130));
 sg13g2_buf_1 fanout4131 (.A(net4134),
    .X(net4131));
 sg13g2_buf_8 fanout4132 (.A(net4134),
    .X(net4132));
 sg13g2_buf_1 fanout4133 (.A(net4134),
    .X(net4133));
 sg13g2_buf_8 fanout4134 (.A(net4142),
    .X(net4134));
 sg13g2_buf_8 fanout4135 (.A(net4138),
    .X(net4135));
 sg13g2_buf_1 fanout4136 (.A(net4138),
    .X(net4136));
 sg13g2_buf_8 fanout4137 (.A(net4138),
    .X(net4137));
 sg13g2_buf_2 fanout4138 (.A(net4141),
    .X(net4138));
 sg13g2_buf_8 fanout4139 (.A(net4141),
    .X(net4139));
 sg13g2_buf_1 fanout4140 (.A(net4141),
    .X(net4140));
 sg13g2_buf_8 fanout4141 (.A(net4142),
    .X(net4141));
 sg13g2_buf_8 fanout4142 (.A(net4143),
    .X(net4142));
 sg13g2_buf_8 fanout4143 (.A(_12822_),
    .X(net4143));
 sg13g2_buf_8 fanout4144 (.A(net4147),
    .X(net4144));
 sg13g2_buf_8 fanout4145 (.A(net4146),
    .X(net4145));
 sg13g2_buf_8 fanout4146 (.A(net4147),
    .X(net4146));
 sg13g2_buf_8 fanout4147 (.A(net4150),
    .X(net4147));
 sg13g2_buf_8 fanout4148 (.A(net4149),
    .X(net4148));
 sg13g2_buf_8 fanout4149 (.A(net4150),
    .X(net4149));
 sg13g2_buf_8 fanout4150 (.A(_05700_),
    .X(net4150));
 sg13g2_buf_8 fanout4151 (.A(net4153),
    .X(net4151));
 sg13g2_buf_8 fanout4152 (.A(net4153),
    .X(net4152));
 sg13g2_buf_8 fanout4153 (.A(net4157),
    .X(net4153));
 sg13g2_buf_8 fanout4154 (.A(net4157),
    .X(net4154));
 sg13g2_buf_8 fanout4155 (.A(net4156),
    .X(net4155));
 sg13g2_buf_8 fanout4156 (.A(net4157),
    .X(net4156));
 sg13g2_buf_8 fanout4157 (.A(_05700_),
    .X(net4157));
 sg13g2_buf_8 fanout4158 (.A(net4160),
    .X(net4158));
 sg13g2_buf_8 fanout4159 (.A(net4160),
    .X(net4159));
 sg13g2_buf_8 fanout4160 (.A(net4173),
    .X(net4160));
 sg13g2_buf_8 fanout4161 (.A(net4173),
    .X(net4161));
 sg13g2_buf_8 fanout4162 (.A(net4173),
    .X(net4162));
 sg13g2_buf_8 fanout4163 (.A(net4164),
    .X(net4163));
 sg13g2_buf_8 fanout4164 (.A(net4165),
    .X(net4164));
 sg13g2_buf_8 fanout4165 (.A(net4173),
    .X(net4165));
 sg13g2_buf_8 fanout4166 (.A(net4171),
    .X(net4166));
 sg13g2_buf_1 fanout4167 (.A(net4168),
    .X(net4167));
 sg13g2_buf_8 fanout4168 (.A(net4171),
    .X(net4168));
 sg13g2_buf_8 fanout4169 (.A(net4170),
    .X(net4169));
 sg13g2_buf_8 fanout4170 (.A(net4171),
    .X(net4170));
 sg13g2_buf_8 fanout4171 (.A(net4172),
    .X(net4171));
 sg13g2_buf_2 fanout4172 (.A(net4173),
    .X(net4172));
 sg13g2_buf_8 fanout4173 (.A(_05700_),
    .X(net4173));
 sg13g2_buf_8 fanout4174 (.A(net4175),
    .X(net4174));
 sg13g2_buf_1 fanout4175 (.A(net4180),
    .X(net4175));
 sg13g2_buf_8 fanout4176 (.A(net4180),
    .X(net4176));
 sg13g2_buf_2 fanout4177 (.A(net4180),
    .X(net4177));
 sg13g2_buf_8 fanout4178 (.A(net4180),
    .X(net4178));
 sg13g2_buf_8 fanout4179 (.A(net4180),
    .X(net4179));
 sg13g2_buf_8 fanout4180 (.A(net4201),
    .X(net4180));
 sg13g2_buf_8 fanout4181 (.A(net4183),
    .X(net4181));
 sg13g2_buf_8 fanout4182 (.A(net4183),
    .X(net4182));
 sg13g2_buf_8 fanout4183 (.A(net4201),
    .X(net4183));
 sg13g2_buf_8 fanout4184 (.A(net4186),
    .X(net4184));
 sg13g2_buf_1 fanout4185 (.A(net4186),
    .X(net4185));
 sg13g2_buf_2 fanout4186 (.A(net4187),
    .X(net4186));
 sg13g2_buf_1 fanout4187 (.A(net4201),
    .X(net4187));
 sg13g2_buf_8 fanout4188 (.A(net4189),
    .X(net4188));
 sg13g2_buf_1 fanout4189 (.A(net4200),
    .X(net4189));
 sg13g2_buf_8 fanout4190 (.A(net4191),
    .X(net4190));
 sg13g2_buf_8 fanout4191 (.A(net4192),
    .X(net4191));
 sg13g2_buf_8 fanout4192 (.A(net4200),
    .X(net4192));
 sg13g2_buf_8 fanout4193 (.A(net4195),
    .X(net4193));
 sg13g2_buf_1 fanout4194 (.A(net4195),
    .X(net4194));
 sg13g2_buf_8 fanout4195 (.A(net4196),
    .X(net4195));
 sg13g2_buf_8 fanout4196 (.A(net4200),
    .X(net4196));
 sg13g2_buf_8 fanout4197 (.A(net4198),
    .X(net4197));
 sg13g2_buf_1 fanout4198 (.A(net4199),
    .X(net4198));
 sg13g2_buf_1 fanout4199 (.A(net4200),
    .X(net4199));
 sg13g2_buf_8 fanout4200 (.A(net4201),
    .X(net4200));
 sg13g2_buf_8 fanout4201 (.A(_05699_),
    .X(net4201));
 sg13g2_buf_8 fanout4202 (.A(net4204),
    .X(net4202));
 sg13g2_buf_1 fanout4203 (.A(net4204),
    .X(net4203));
 sg13g2_buf_8 fanout4204 (.A(net4205),
    .X(net4204));
 sg13g2_buf_8 fanout4205 (.A(net4215),
    .X(net4205));
 sg13g2_buf_8 fanout4206 (.A(net4208),
    .X(net4206));
 sg13g2_buf_1 fanout4207 (.A(net4208),
    .X(net4207));
 sg13g2_buf_8 fanout4208 (.A(net4215),
    .X(net4208));
 sg13g2_buf_8 fanout4209 (.A(net4210),
    .X(net4209));
 sg13g2_buf_2 fanout4210 (.A(net4211),
    .X(net4210));
 sg13g2_buf_8 fanout4211 (.A(net4215),
    .X(net4211));
 sg13g2_buf_8 fanout4212 (.A(net4213),
    .X(net4212));
 sg13g2_buf_8 fanout4213 (.A(net4214),
    .X(net4213));
 sg13g2_buf_8 fanout4214 (.A(net4215),
    .X(net4214));
 sg13g2_buf_8 fanout4215 (.A(_05699_),
    .X(net4215));
 sg13g2_buf_8 fanout4216 (.A(net4217),
    .X(net4216));
 sg13g2_buf_8 fanout4217 (.A(net4231),
    .X(net4217));
 sg13g2_buf_8 fanout4218 (.A(net4231),
    .X(net4218));
 sg13g2_buf_8 fanout4219 (.A(net4225),
    .X(net4219));
 sg13g2_buf_8 fanout4220 (.A(net4221),
    .X(net4220));
 sg13g2_buf_1 fanout4221 (.A(net4222),
    .X(net4221));
 sg13g2_buf_1 fanout4222 (.A(net4224),
    .X(net4222));
 sg13g2_buf_8 fanout4223 (.A(net4224),
    .X(net4223));
 sg13g2_buf_1 fanout4224 (.A(net4225),
    .X(net4224));
 sg13g2_buf_2 fanout4225 (.A(net4231),
    .X(net4225));
 sg13g2_buf_8 fanout4226 (.A(net4228),
    .X(net4226));
 sg13g2_buf_1 fanout4227 (.A(net4228),
    .X(net4227));
 sg13g2_buf_2 fanout4228 (.A(net4229),
    .X(net4228));
 sg13g2_buf_8 fanout4229 (.A(net4231),
    .X(net4229));
 sg13g2_buf_8 fanout4230 (.A(net4231),
    .X(net4230));
 sg13g2_buf_8 fanout4231 (.A(_05699_),
    .X(net4231));
 sg13g2_buf_8 fanout4232 (.A(net4233),
    .X(net4232));
 sg13g2_buf_8 fanout4233 (.A(net4240),
    .X(net4233));
 sg13g2_buf_8 fanout4234 (.A(net4240),
    .X(net4234));
 sg13g2_buf_8 fanout4235 (.A(net4240),
    .X(net4235));
 sg13g2_buf_8 fanout4236 (.A(net4237),
    .X(net4236));
 sg13g2_buf_8 fanout4237 (.A(net4240),
    .X(net4237));
 sg13g2_buf_8 fanout4238 (.A(net4239),
    .X(net4238));
 sg13g2_buf_8 fanout4239 (.A(net4240),
    .X(net4239));
 sg13g2_buf_8 fanout4240 (.A(_12818_),
    .X(net4240));
 sg13g2_buf_8 fanout4241 (.A(_11054_),
    .X(net4241));
 sg13g2_buf_8 fanout4242 (.A(net4247),
    .X(net4242));
 sg13g2_buf_8 fanout4243 (.A(net4244),
    .X(net4243));
 sg13g2_buf_8 fanout4244 (.A(net4245),
    .X(net4244));
 sg13g2_buf_8 fanout4245 (.A(net4247),
    .X(net4245));
 sg13g2_buf_8 fanout4246 (.A(net4247),
    .X(net4246));
 sg13g2_buf_8 fanout4247 (.A(net4266),
    .X(net4247));
 sg13g2_buf_8 fanout4248 (.A(net4250),
    .X(net4248));
 sg13g2_buf_1 fanout4249 (.A(net4250),
    .X(net4249));
 sg13g2_buf_8 fanout4250 (.A(net4266),
    .X(net4250));
 sg13g2_buf_8 fanout4251 (.A(net4253),
    .X(net4251));
 sg13g2_buf_8 fanout4252 (.A(net4253),
    .X(net4252));
 sg13g2_buf_8 fanout4253 (.A(net4266),
    .X(net4253));
 sg13g2_buf_8 fanout4254 (.A(net4259),
    .X(net4254));
 sg13g2_buf_8 fanout4255 (.A(net4259),
    .X(net4255));
 sg13g2_buf_8 fanout4256 (.A(net4257),
    .X(net4256));
 sg13g2_buf_8 fanout4257 (.A(net4258),
    .X(net4257));
 sg13g2_buf_8 fanout4258 (.A(net4259),
    .X(net4258));
 sg13g2_buf_8 fanout4259 (.A(net4265),
    .X(net4259));
 sg13g2_buf_8 fanout4260 (.A(net4265),
    .X(net4260));
 sg13g2_buf_8 fanout4261 (.A(net4264),
    .X(net4261));
 sg13g2_buf_8 fanout4262 (.A(net4263),
    .X(net4262));
 sg13g2_buf_8 fanout4263 (.A(net4264),
    .X(net4263));
 sg13g2_buf_8 fanout4264 (.A(net4265),
    .X(net4264));
 sg13g2_buf_8 fanout4265 (.A(net4266),
    .X(net4265));
 sg13g2_buf_8 fanout4266 (.A(net4288),
    .X(net4266));
 sg13g2_buf_8 fanout4267 (.A(net4270),
    .X(net4267));
 sg13g2_buf_8 fanout4268 (.A(net4269),
    .X(net4268));
 sg13g2_buf_8 fanout4269 (.A(net4270),
    .X(net4269));
 sg13g2_buf_8 fanout4270 (.A(net4288),
    .X(net4270));
 sg13g2_buf_8 fanout4271 (.A(net4272),
    .X(net4271));
 sg13g2_buf_8 fanout4272 (.A(net4274),
    .X(net4272));
 sg13g2_buf_8 fanout4273 (.A(net4274),
    .X(net4273));
 sg13g2_buf_8 fanout4274 (.A(net4288),
    .X(net4274));
 sg13g2_buf_8 fanout4275 (.A(net4287),
    .X(net4275));
 sg13g2_buf_8 fanout4276 (.A(net4277),
    .X(net4276));
 sg13g2_buf_8 fanout4277 (.A(net4287),
    .X(net4277));
 sg13g2_buf_8 fanout4278 (.A(net4279),
    .X(net4278));
 sg13g2_buf_8 fanout4279 (.A(net4287),
    .X(net4279));
 sg13g2_buf_8 fanout4280 (.A(net4281),
    .X(net4280));
 sg13g2_buf_8 fanout4281 (.A(net4287),
    .X(net4281));
 sg13g2_buf_8 fanout4282 (.A(net4286),
    .X(net4282));
 sg13g2_buf_8 fanout4283 (.A(net4285),
    .X(net4283));
 sg13g2_buf_8 fanout4284 (.A(net4285),
    .X(net4284));
 sg13g2_buf_8 fanout4285 (.A(net4286),
    .X(net4285));
 sg13g2_buf_8 fanout4286 (.A(net4287),
    .X(net4286));
 sg13g2_buf_8 fanout4287 (.A(net4288),
    .X(net4287));
 sg13g2_buf_8 fanout4288 (.A(_10277_),
    .X(net4288));
 sg13g2_buf_8 fanout4289 (.A(net4290),
    .X(net4289));
 sg13g2_buf_8 fanout4290 (.A(net4291),
    .X(net4290));
 sg13g2_buf_8 fanout4291 (.A(net4294),
    .X(net4291));
 sg13g2_buf_8 fanout4292 (.A(net4293),
    .X(net4292));
 sg13g2_buf_8 fanout4293 (.A(net4294),
    .X(net4293));
 sg13g2_buf_8 fanout4294 (.A(_15658_),
    .X(net4294));
 sg13g2_buf_8 fanout4295 (.A(net4299),
    .X(net4295));
 sg13g2_buf_8 fanout4296 (.A(net4299),
    .X(net4296));
 sg13g2_buf_8 fanout4297 (.A(net4299),
    .X(net4297));
 sg13g2_buf_8 fanout4298 (.A(net4299),
    .X(net4298));
 sg13g2_buf_8 fanout4299 (.A(_15658_),
    .X(net4299));
 sg13g2_buf_8 fanout4300 (.A(net4308),
    .X(net4300));
 sg13g2_buf_8 fanout4301 (.A(net4308),
    .X(net4301));
 sg13g2_buf_8 fanout4302 (.A(net4304),
    .X(net4302));
 sg13g2_buf_1 fanout4303 (.A(net4304),
    .X(net4303));
 sg13g2_buf_8 fanout4304 (.A(net4308),
    .X(net4304));
 sg13g2_buf_8 fanout4305 (.A(net4307),
    .X(net4305));
 sg13g2_buf_1 fanout4306 (.A(net4307),
    .X(net4306));
 sg13g2_buf_8 fanout4307 (.A(net4308),
    .X(net4307));
 sg13g2_buf_8 fanout4308 (.A(net4333),
    .X(net4308));
 sg13g2_buf_8 fanout4309 (.A(net4311),
    .X(net4309));
 sg13g2_buf_1 fanout4310 (.A(net4311),
    .X(net4310));
 sg13g2_buf_8 fanout4311 (.A(net4317),
    .X(net4311));
 sg13g2_buf_8 fanout4312 (.A(net4314),
    .X(net4312));
 sg13g2_buf_1 fanout4313 (.A(net4314),
    .X(net4313));
 sg13g2_buf_8 fanout4314 (.A(net4317),
    .X(net4314));
 sg13g2_buf_8 fanout4315 (.A(net4316),
    .X(net4315));
 sg13g2_buf_8 fanout4316 (.A(net4317),
    .X(net4316));
 sg13g2_buf_8 fanout4317 (.A(net4333),
    .X(net4317));
 sg13g2_buf_8 fanout4318 (.A(net4319),
    .X(net4318));
 sg13g2_buf_8 fanout4319 (.A(net4323),
    .X(net4319));
 sg13g2_buf_8 fanout4320 (.A(net4321),
    .X(net4320));
 sg13g2_buf_8 fanout4321 (.A(net4322),
    .X(net4321));
 sg13g2_buf_8 fanout4322 (.A(net4323),
    .X(net4322));
 sg13g2_buf_2 fanout4323 (.A(net4333),
    .X(net4323));
 sg13g2_buf_8 fanout4324 (.A(net4326),
    .X(net4324));
 sg13g2_buf_1 fanout4325 (.A(net4326),
    .X(net4325));
 sg13g2_buf_8 fanout4326 (.A(net4327),
    .X(net4326));
 sg13g2_buf_8 fanout4327 (.A(net4332),
    .X(net4327));
 sg13g2_buf_8 fanout4328 (.A(net4330),
    .X(net4328));
 sg13g2_buf_8 fanout4329 (.A(net4330),
    .X(net4329));
 sg13g2_buf_8 fanout4330 (.A(net4332),
    .X(net4330));
 sg13g2_buf_8 fanout4331 (.A(net4332),
    .X(net4331));
 sg13g2_buf_8 fanout4332 (.A(net4333),
    .X(net4332));
 sg13g2_buf_8 fanout4333 (.A(_15657_),
    .X(net4333));
 sg13g2_buf_8 fanout4334 (.A(net4337),
    .X(net4334));
 sg13g2_buf_8 fanout4335 (.A(net4337),
    .X(net4335));
 sg13g2_buf_8 fanout4336 (.A(net4337),
    .X(net4336));
 sg13g2_buf_8 fanout4337 (.A(net4358),
    .X(net4337));
 sg13g2_buf_8 fanout4338 (.A(net4340),
    .X(net4338));
 sg13g2_buf_1 fanout4339 (.A(net4340),
    .X(net4339));
 sg13g2_buf_8 fanout4340 (.A(net4342),
    .X(net4340));
 sg13g2_buf_8 fanout4341 (.A(net4342),
    .X(net4341));
 sg13g2_buf_8 fanout4342 (.A(net4358),
    .X(net4342));
 sg13g2_buf_8 fanout4343 (.A(net4344),
    .X(net4343));
 sg13g2_buf_8 fanout4344 (.A(net4358),
    .X(net4344));
 sg13g2_buf_8 fanout4345 (.A(net4353),
    .X(net4345));
 sg13g2_buf_1 fanout4346 (.A(net4353),
    .X(net4346));
 sg13g2_buf_8 fanout4347 (.A(net4353),
    .X(net4347));
 sg13g2_buf_1 fanout4348 (.A(net4349),
    .X(net4348));
 sg13g2_buf_8 fanout4349 (.A(net4353),
    .X(net4349));
 sg13g2_buf_8 fanout4350 (.A(net4352),
    .X(net4350));
 sg13g2_buf_8 fanout4351 (.A(net4352),
    .X(net4351));
 sg13g2_buf_2 fanout4352 (.A(net4353),
    .X(net4352));
 sg13g2_buf_8 fanout4353 (.A(net4358),
    .X(net4353));
 sg13g2_buf_8 fanout4354 (.A(net4357),
    .X(net4354));
 sg13g2_buf_8 fanout4355 (.A(net4356),
    .X(net4355));
 sg13g2_buf_8 fanout4356 (.A(net4357),
    .X(net4356));
 sg13g2_buf_8 fanout4357 (.A(net4358),
    .X(net4357));
 sg13g2_buf_8 fanout4358 (.A(_15657_),
    .X(net4358));
 sg13g2_buf_8 fanout4359 (.A(net4360),
    .X(net4359));
 sg13g2_buf_8 fanout4360 (.A(net4364),
    .X(net4360));
 sg13g2_buf_8 fanout4361 (.A(net4362),
    .X(net4361));
 sg13g2_buf_8 fanout4362 (.A(net4363),
    .X(net4362));
 sg13g2_buf_8 fanout4363 (.A(net4364),
    .X(net4363));
 sg13g2_buf_8 fanout4364 (.A(net4377),
    .X(net4364));
 sg13g2_buf_8 fanout4365 (.A(net4367),
    .X(net4365));
 sg13g2_buf_2 fanout4366 (.A(net4367),
    .X(net4366));
 sg13g2_buf_8 fanout4367 (.A(net4377),
    .X(net4367));
 sg13g2_buf_8 fanout4368 (.A(net4370),
    .X(net4368));
 sg13g2_buf_8 fanout4369 (.A(net4370),
    .X(net4369));
 sg13g2_buf_8 fanout4370 (.A(net4377),
    .X(net4370));
 sg13g2_buf_8 fanout4371 (.A(net4372),
    .X(net4371));
 sg13g2_buf_8 fanout4372 (.A(net4377),
    .X(net4372));
 sg13g2_buf_8 fanout4373 (.A(net4376),
    .X(net4373));
 sg13g2_buf_1 fanout4374 (.A(net4376),
    .X(net4374));
 sg13g2_buf_8 fanout4375 (.A(net4376),
    .X(net4375));
 sg13g2_buf_8 fanout4376 (.A(net4377),
    .X(net4376));
 sg13g2_buf_8 fanout4377 (.A(_15657_),
    .X(net4377));
 sg13g2_buf_8 fanout4378 (.A(net4382),
    .X(net4378));
 sg13g2_buf_8 fanout4379 (.A(net4382),
    .X(net4379));
 sg13g2_buf_8 fanout4380 (.A(net4381),
    .X(net4380));
 sg13g2_buf_8 fanout4381 (.A(net4382),
    .X(net4381));
 sg13g2_buf_8 fanout4382 (.A(_11063_),
    .X(net4382));
 sg13g2_buf_8 fanout4383 (.A(net4386),
    .X(net4383));
 sg13g2_buf_8 fanout4384 (.A(net4385),
    .X(net4384));
 sg13g2_buf_8 fanout4385 (.A(net4386),
    .X(net4385));
 sg13g2_buf_8 fanout4386 (.A(_11063_),
    .X(net4386));
 sg13g2_buf_8 fanout4387 (.A(net4394),
    .X(net4387));
 sg13g2_buf_1 fanout4388 (.A(net4394),
    .X(net4388));
 sg13g2_buf_8 fanout4389 (.A(net4390),
    .X(net4389));
 sg13g2_buf_8 fanout4390 (.A(net4391),
    .X(net4390));
 sg13g2_buf_8 fanout4391 (.A(net4394),
    .X(net4391));
 sg13g2_buf_8 fanout4392 (.A(net4393),
    .X(net4392));
 sg13g2_buf_1 fanout4393 (.A(net4394),
    .X(net4393));
 sg13g2_buf_8 fanout4394 (.A(net4398),
    .X(net4394));
 sg13g2_buf_8 fanout4395 (.A(net4398),
    .X(net4395));
 sg13g2_buf_1 fanout4396 (.A(net4398),
    .X(net4396));
 sg13g2_buf_8 fanout4397 (.A(net4398),
    .X(net4397));
 sg13g2_buf_8 fanout4398 (.A(net4409),
    .X(net4398));
 sg13g2_buf_8 fanout4399 (.A(net4403),
    .X(net4399));
 sg13g2_buf_8 fanout4400 (.A(net4402),
    .X(net4400));
 sg13g2_buf_1 fanout4401 (.A(net4402),
    .X(net4401));
 sg13g2_buf_2 fanout4402 (.A(net4403),
    .X(net4402));
 sg13g2_buf_8 fanout4403 (.A(net4409),
    .X(net4403));
 sg13g2_buf_8 fanout4404 (.A(net4405),
    .X(net4404));
 sg13g2_buf_8 fanout4405 (.A(net4409),
    .X(net4405));
 sg13g2_buf_8 fanout4406 (.A(net4407),
    .X(net4406));
 sg13g2_buf_8 fanout4407 (.A(net4408),
    .X(net4407));
 sg13g2_buf_8 fanout4408 (.A(net4409),
    .X(net4408));
 sg13g2_buf_8 fanout4409 (.A(_11041_),
    .X(net4409));
 sg13g2_buf_8 fanout4410 (.A(net4412),
    .X(net4410));
 sg13g2_buf_8 fanout4411 (.A(net4412),
    .X(net4411));
 sg13g2_buf_8 fanout4412 (.A(net4413),
    .X(net4412));
 sg13g2_buf_8 fanout4413 (.A(net4418),
    .X(net4413));
 sg13g2_buf_8 fanout4414 (.A(net4418),
    .X(net4414));
 sg13g2_buf_1 fanout4415 (.A(net4418),
    .X(net4415));
 sg13g2_buf_8 fanout4416 (.A(net4417),
    .X(net4416));
 sg13g2_buf_2 fanout4417 (.A(net4418),
    .X(net4417));
 sg13g2_buf_8 fanout4418 (.A(_11041_),
    .X(net4418));
 sg13g2_buf_8 fanout4419 (.A(net4420),
    .X(net4419));
 sg13g2_buf_1 fanout4420 (.A(net4428),
    .X(net4420));
 sg13g2_buf_8 fanout4421 (.A(net4422),
    .X(net4421));
 sg13g2_buf_8 fanout4422 (.A(net4425),
    .X(net4422));
 sg13g2_buf_8 fanout4423 (.A(net4425),
    .X(net4423));
 sg13g2_buf_1 fanout4424 (.A(net4425),
    .X(net4424));
 sg13g2_buf_8 fanout4425 (.A(net4428),
    .X(net4425));
 sg13g2_buf_8 fanout4426 (.A(net4427),
    .X(net4426));
 sg13g2_buf_8 fanout4427 (.A(net4428),
    .X(net4427));
 sg13g2_buf_8 fanout4428 (.A(_11041_),
    .X(net4428));
 sg13g2_buf_8 fanout4429 (.A(_14840_),
    .X(net4429));
 sg13g2_buf_8 fanout4430 (.A(_14838_),
    .X(net4430));
 sg13g2_buf_8 fanout4431 (.A(_13825_),
    .X(net4431));
 sg13g2_buf_8 fanout4432 (.A(_11792_),
    .X(net4432));
 sg13g2_buf_8 fanout4433 (.A(_11763_),
    .X(net4433));
 sg13g2_buf_8 fanout4434 (.A(net4435),
    .X(net4434));
 sg13g2_buf_8 fanout4435 (.A(net4436),
    .X(net4435));
 sg13g2_buf_8 fanout4436 (.A(net4437),
    .X(net4436));
 sg13g2_buf_8 fanout4437 (.A(net4450),
    .X(net4437));
 sg13g2_buf_8 fanout4438 (.A(net4439),
    .X(net4438));
 sg13g2_buf_2 fanout4439 (.A(net4450),
    .X(net4439));
 sg13g2_buf_8 fanout4440 (.A(net4441),
    .X(net4440));
 sg13g2_buf_8 fanout4441 (.A(net4444),
    .X(net4441));
 sg13g2_buf_8 fanout4442 (.A(net4444),
    .X(net4442));
 sg13g2_buf_1 fanout4443 (.A(net4444),
    .X(net4443));
 sg13g2_buf_8 fanout4444 (.A(net4450),
    .X(net4444));
 sg13g2_buf_8 fanout4445 (.A(net4449),
    .X(net4445));
 sg13g2_buf_8 fanout4446 (.A(net4447),
    .X(net4446));
 sg13g2_buf_8 fanout4447 (.A(net4449),
    .X(net4447));
 sg13g2_buf_8 fanout4448 (.A(net4449),
    .X(net4448));
 sg13g2_buf_8 fanout4449 (.A(net4450),
    .X(net4449));
 sg13g2_buf_8 fanout4450 (.A(_11064_),
    .X(net4450));
 sg13g2_buf_8 fanout4451 (.A(net4452),
    .X(net4451));
 sg13g2_buf_8 fanout4452 (.A(net4454),
    .X(net4452));
 sg13g2_buf_8 fanout4453 (.A(net4454),
    .X(net4453));
 sg13g2_buf_8 fanout4454 (.A(net4472),
    .X(net4454));
 sg13g2_buf_8 fanout4455 (.A(net4456),
    .X(net4455));
 sg13g2_buf_8 fanout4456 (.A(net4457),
    .X(net4456));
 sg13g2_buf_8 fanout4457 (.A(net4472),
    .X(net4457));
 sg13g2_buf_8 fanout4458 (.A(net4460),
    .X(net4458));
 sg13g2_buf_1 fanout4459 (.A(net4460),
    .X(net4459));
 sg13g2_buf_1 fanout4460 (.A(net4472),
    .X(net4460));
 sg13g2_buf_8 fanout4461 (.A(net4465),
    .X(net4461));
 sg13g2_buf_1 fanout4462 (.A(net4465),
    .X(net4462));
 sg13g2_buf_8 fanout4463 (.A(net4465),
    .X(net4463));
 sg13g2_buf_2 fanout4464 (.A(net4465),
    .X(net4464));
 sg13g2_buf_8 fanout4465 (.A(net4472),
    .X(net4465));
 sg13g2_buf_2 fanout4466 (.A(net4468),
    .X(net4466));
 sg13g2_buf_1 fanout4467 (.A(net4468),
    .X(net4467));
 sg13g2_buf_8 fanout4468 (.A(net4471),
    .X(net4468));
 sg13g2_buf_2 fanout4469 (.A(net4470),
    .X(net4469));
 sg13g2_buf_8 fanout4470 (.A(net4471),
    .X(net4470));
 sg13g2_buf_8 fanout4471 (.A(net4472),
    .X(net4471));
 sg13g2_buf_8 fanout4472 (.A(_11042_),
    .X(net4472));
 sg13g2_buf_2 fanout4473 (.A(net4474),
    .X(net4473));
 sg13g2_buf_2 fanout4474 (.A(net4477),
    .X(net4474));
 sg13g2_buf_2 fanout4475 (.A(net4477),
    .X(net4475));
 sg13g2_buf_2 fanout4476 (.A(net4477),
    .X(net4476));
 sg13g2_buf_1 fanout4477 (.A(net4500),
    .X(net4477));
 sg13g2_buf_2 fanout4478 (.A(net4479),
    .X(net4478));
 sg13g2_buf_8 fanout4479 (.A(net4480),
    .X(net4479));
 sg13g2_buf_1 fanout4480 (.A(net4500),
    .X(net4480));
 sg13g2_buf_2 fanout4481 (.A(net4483),
    .X(net4481));
 sg13g2_buf_1 fanout4482 (.A(net4483),
    .X(net4482));
 sg13g2_buf_1 fanout4483 (.A(net4500),
    .X(net4483));
 sg13g2_buf_2 fanout4484 (.A(net4485),
    .X(net4484));
 sg13g2_buf_8 fanout4485 (.A(net4486),
    .X(net4485));
 sg13g2_buf_2 fanout4486 (.A(net4499),
    .X(net4486));
 sg13g2_buf_2 fanout4487 (.A(net4489),
    .X(net4487));
 sg13g2_buf_2 fanout4488 (.A(net4489),
    .X(net4488));
 sg13g2_buf_1 fanout4489 (.A(net4492),
    .X(net4489));
 sg13g2_buf_8 fanout4490 (.A(net4491),
    .X(net4490));
 sg13g2_buf_8 fanout4491 (.A(net4492),
    .X(net4491));
 sg13g2_buf_8 fanout4492 (.A(net4499),
    .X(net4492));
 sg13g2_buf_2 fanout4493 (.A(net4494),
    .X(net4493));
 sg13g2_buf_1 fanout4494 (.A(net4499),
    .X(net4494));
 sg13g2_buf_2 fanout4495 (.A(net4497),
    .X(net4495));
 sg13g2_buf_2 fanout4496 (.A(net4497),
    .X(net4496));
 sg13g2_buf_2 fanout4497 (.A(net4498),
    .X(net4497));
 sg13g2_buf_1 fanout4498 (.A(net4499),
    .X(net4498));
 sg13g2_buf_8 fanout4499 (.A(net4500),
    .X(net4499));
 sg13g2_buf_8 fanout4500 (.A(_11042_),
    .X(net4500));
 sg13g2_buf_8 fanout4501 (.A(net4502),
    .X(net4501));
 sg13g2_buf_8 fanout4502 (.A(net4503),
    .X(net4502));
 sg13g2_buf_8 fanout4503 (.A(_10634_),
    .X(net4503));
 sg13g2_buf_8 fanout4504 (.A(net4505),
    .X(net4504));
 sg13g2_buf_8 fanout4505 (.A(_10634_),
    .X(net4505));
 sg13g2_buf_8 fanout4506 (.A(net4510),
    .X(net4506));
 sg13g2_buf_1 fanout4507 (.A(net4510),
    .X(net4507));
 sg13g2_buf_8 fanout4508 (.A(net4510),
    .X(net4508));
 sg13g2_buf_8 fanout4509 (.A(net4510),
    .X(net4509));
 sg13g2_buf_8 fanout4510 (.A(_10634_),
    .X(net4510));
 sg13g2_buf_8 fanout4511 (.A(net4512),
    .X(net4511));
 sg13g2_buf_8 fanout4512 (.A(net4515),
    .X(net4512));
 sg13g2_buf_8 fanout4513 (.A(net4515),
    .X(net4513));
 sg13g2_buf_8 fanout4514 (.A(net4515),
    .X(net4514));
 sg13g2_buf_8 fanout4515 (.A(_10625_),
    .X(net4515));
 sg13g2_buf_8 fanout4516 (.A(net4518),
    .X(net4516));
 sg13g2_buf_2 fanout4517 (.A(net4518),
    .X(net4517));
 sg13g2_buf_8 fanout4518 (.A(_10625_),
    .X(net4518));
 sg13g2_buf_8 fanout4519 (.A(net4520),
    .X(net4519));
 sg13g2_buf_8 fanout4520 (.A(net4521),
    .X(net4520));
 sg13g2_buf_8 fanout4521 (.A(_10625_),
    .X(net4521));
 sg13g2_buf_8 fanout4522 (.A(net4523),
    .X(net4522));
 sg13g2_buf_8 fanout4523 (.A(net4524),
    .X(net4523));
 sg13g2_buf_8 fanout4524 (.A(net4529),
    .X(net4524));
 sg13g2_buf_8 fanout4525 (.A(net4529),
    .X(net4525));
 sg13g2_buf_8 fanout4526 (.A(net4528),
    .X(net4526));
 sg13g2_buf_8 fanout4527 (.A(net4528),
    .X(net4527));
 sg13g2_buf_8 fanout4528 (.A(net4529),
    .X(net4528));
 sg13g2_buf_8 fanout4529 (.A(net4558),
    .X(net4529));
 sg13g2_buf_8 fanout4530 (.A(net4531),
    .X(net4530));
 sg13g2_buf_8 fanout4531 (.A(net4539),
    .X(net4531));
 sg13g2_buf_8 fanout4532 (.A(net4535),
    .X(net4532));
 sg13g2_buf_8 fanout4533 (.A(net4535),
    .X(net4533));
 sg13g2_buf_1 fanout4534 (.A(net4535),
    .X(net4534));
 sg13g2_buf_8 fanout4535 (.A(net4539),
    .X(net4535));
 sg13g2_buf_8 fanout4536 (.A(net4538),
    .X(net4536));
 sg13g2_buf_8 fanout4537 (.A(net4538),
    .X(net4537));
 sg13g2_buf_8 fanout4538 (.A(net4539),
    .X(net4538));
 sg13g2_buf_8 fanout4539 (.A(net4558),
    .X(net4539));
 sg13g2_buf_8 fanout4540 (.A(net4542),
    .X(net4540));
 sg13g2_buf_2 fanout4541 (.A(net4542),
    .X(net4541));
 sg13g2_buf_8 fanout4542 (.A(net4547),
    .X(net4542));
 sg13g2_buf_8 fanout4543 (.A(net4545),
    .X(net4543));
 sg13g2_buf_1 fanout4544 (.A(net4545),
    .X(net4544));
 sg13g2_buf_8 fanout4545 (.A(net4547),
    .X(net4545));
 sg13g2_buf_8 fanout4546 (.A(net4547),
    .X(net4546));
 sg13g2_buf_8 fanout4547 (.A(net4558),
    .X(net4547));
 sg13g2_buf_8 fanout4548 (.A(net4549),
    .X(net4548));
 sg13g2_buf_8 fanout4549 (.A(net4557),
    .X(net4549));
 sg13g2_buf_8 fanout4550 (.A(net4551),
    .X(net4550));
 sg13g2_buf_8 fanout4551 (.A(net4554),
    .X(net4551));
 sg13g2_buf_8 fanout4552 (.A(net4554),
    .X(net4552));
 sg13g2_buf_1 fanout4553 (.A(net4554),
    .X(net4553));
 sg13g2_buf_8 fanout4554 (.A(net4557),
    .X(net4554));
 sg13g2_buf_8 fanout4555 (.A(net4557),
    .X(net4555));
 sg13g2_buf_8 fanout4556 (.A(net4557),
    .X(net4556));
 sg13g2_buf_8 fanout4557 (.A(net4558),
    .X(net4557));
 sg13g2_buf_8 fanout4558 (.A(_10577_),
    .X(net4558));
 sg13g2_buf_8 fanout4559 (.A(net4561),
    .X(net4559));
 sg13g2_buf_1 fanout4560 (.A(net4561),
    .X(net4560));
 sg13g2_buf_8 fanout4561 (.A(net4567),
    .X(net4561));
 sg13g2_buf_8 fanout4562 (.A(net4567),
    .X(net4562));
 sg13g2_buf_8 fanout4563 (.A(net4565),
    .X(net4563));
 sg13g2_buf_1 fanout4564 (.A(net4565),
    .X(net4564));
 sg13g2_buf_2 fanout4565 (.A(net4567),
    .X(net4565));
 sg13g2_buf_8 fanout4566 (.A(net4567),
    .X(net4566));
 sg13g2_buf_8 fanout4567 (.A(net4583),
    .X(net4567));
 sg13g2_buf_8 fanout4568 (.A(net4569),
    .X(net4568));
 sg13g2_buf_8 fanout4569 (.A(net4583),
    .X(net4569));
 sg13g2_buf_8 fanout4570 (.A(net4571),
    .X(net4570));
 sg13g2_buf_8 fanout4571 (.A(net4579),
    .X(net4571));
 sg13g2_buf_8 fanout4572 (.A(net4579),
    .X(net4572));
 sg13g2_buf_1 fanout4573 (.A(net4579),
    .X(net4573));
 sg13g2_buf_8 fanout4574 (.A(net4578),
    .X(net4574));
 sg13g2_buf_2 fanout4575 (.A(net4578),
    .X(net4575));
 sg13g2_buf_8 fanout4576 (.A(net4578),
    .X(net4576));
 sg13g2_buf_1 fanout4577 (.A(net4578),
    .X(net4577));
 sg13g2_buf_8 fanout4578 (.A(net4579),
    .X(net4578));
 sg13g2_buf_8 fanout4579 (.A(net4583),
    .X(net4579));
 sg13g2_buf_8 fanout4580 (.A(net4581),
    .X(net4580));
 sg13g2_buf_8 fanout4581 (.A(net4582),
    .X(net4581));
 sg13g2_buf_8 fanout4582 (.A(net4583),
    .X(net4582));
 sg13g2_buf_8 fanout4583 (.A(_10577_),
    .X(net4583));
 sg13g2_buf_8 fanout4584 (.A(net4585),
    .X(net4584));
 sg13g2_buf_8 fanout4585 (.A(net4586),
    .X(net4585));
 sg13g2_buf_8 fanout4586 (.A(net4600),
    .X(net4586));
 sg13g2_buf_8 fanout4587 (.A(net4589),
    .X(net4587));
 sg13g2_buf_8 fanout4588 (.A(net4589),
    .X(net4588));
 sg13g2_buf_8 fanout4589 (.A(net4600),
    .X(net4589));
 sg13g2_buf_8 fanout4590 (.A(net4593),
    .X(net4590));
 sg13g2_buf_1 fanout4591 (.A(net4593),
    .X(net4591));
 sg13g2_buf_8 fanout4592 (.A(net4593),
    .X(net4592));
 sg13g2_buf_8 fanout4593 (.A(net4600),
    .X(net4593));
 sg13g2_buf_8 fanout4594 (.A(net4595),
    .X(net4594));
 sg13g2_buf_8 fanout4595 (.A(net4596),
    .X(net4595));
 sg13g2_buf_8 fanout4596 (.A(net4600),
    .X(net4596));
 sg13g2_buf_8 fanout4597 (.A(net4599),
    .X(net4597));
 sg13g2_buf_1 fanout4598 (.A(net4599),
    .X(net4598));
 sg13g2_buf_2 fanout4599 (.A(net4600),
    .X(net4599));
 sg13g2_buf_8 fanout4600 (.A(_10577_),
    .X(net4600));
 sg13g2_buf_8 fanout4601 (.A(net4602),
    .X(net4601));
 sg13g2_buf_8 fanout4602 (.A(net4603),
    .X(net4602));
 sg13g2_buf_8 fanout4603 (.A(net4608),
    .X(net4603));
 sg13g2_buf_8 fanout4604 (.A(net4606),
    .X(net4604));
 sg13g2_buf_8 fanout4605 (.A(net4606),
    .X(net4605));
 sg13g2_buf_8 fanout4606 (.A(net4607),
    .X(net4606));
 sg13g2_buf_8 fanout4607 (.A(net4608),
    .X(net4607));
 sg13g2_buf_8 fanout4608 (.A(\u_inv.state[0] ),
    .X(net4608));
 sg13g2_buf_8 fanout4609 (.A(net4612),
    .X(net4609));
 sg13g2_buf_8 fanout4610 (.A(net4612),
    .X(net4610));
 sg13g2_buf_8 fanout4611 (.A(net4612),
    .X(net4611));
 sg13g2_buf_8 fanout4612 (.A(net4617),
    .X(net4612));
 sg13g2_buf_8 fanout4613 (.A(net4616),
    .X(net4613));
 sg13g2_buf_8 fanout4614 (.A(net4616),
    .X(net4614));
 sg13g2_buf_8 fanout4615 (.A(net4616),
    .X(net4615));
 sg13g2_buf_8 fanout4616 (.A(net4617),
    .X(net4616));
 sg13g2_buf_8 fanout4617 (.A(\u_inv.state[0] ),
    .X(net4617));
 sg13g2_buf_8 fanout4618 (.A(net4622),
    .X(net4618));
 sg13g2_buf_1 fanout4619 (.A(net4622),
    .X(net4619));
 sg13g2_buf_8 fanout4620 (.A(net4622),
    .X(net4620));
 sg13g2_buf_2 fanout4621 (.A(net4622),
    .X(net4621));
 sg13g2_buf_8 fanout4622 (.A(net4633),
    .X(net4622));
 sg13g2_buf_8 fanout4623 (.A(net4633),
    .X(net4623));
 sg13g2_buf_1 fanout4624 (.A(net4633),
    .X(net4624));
 sg13g2_buf_8 fanout4625 (.A(net4627),
    .X(net4625));
 sg13g2_buf_8 fanout4626 (.A(net4627),
    .X(net4626));
 sg13g2_buf_8 fanout4627 (.A(net4632),
    .X(net4627));
 sg13g2_buf_8 fanout4628 (.A(net4629),
    .X(net4628));
 sg13g2_buf_8 fanout4629 (.A(net4632),
    .X(net4629));
 sg13g2_buf_8 fanout4630 (.A(net4632),
    .X(net4630));
 sg13g2_buf_2 fanout4631 (.A(net4632),
    .X(net4631));
 sg13g2_buf_8 fanout4632 (.A(net4633),
    .X(net4632));
 sg13g2_buf_8 fanout4633 (.A(\u_inv.state[0] ),
    .X(net4633));
 sg13g2_buf_8 fanout4634 (.A(net4635),
    .X(net4634));
 sg13g2_buf_8 fanout4635 (.A(net4655),
    .X(net4635));
 sg13g2_buf_8 fanout4636 (.A(net4637),
    .X(net4636));
 sg13g2_buf_8 fanout4637 (.A(net4642),
    .X(net4637));
 sg13g2_buf_8 fanout4638 (.A(net4642),
    .X(net4638));
 sg13g2_buf_2 fanout4639 (.A(net4642),
    .X(net4639));
 sg13g2_buf_8 fanout4640 (.A(net4641),
    .X(net4640));
 sg13g2_buf_1 fanout4641 (.A(net4642),
    .X(net4641));
 sg13g2_buf_8 fanout4642 (.A(net4655),
    .X(net4642));
 sg13g2_buf_8 fanout4643 (.A(net4647),
    .X(net4643));
 sg13g2_buf_1 fanout4644 (.A(net4647),
    .X(net4644));
 sg13g2_buf_8 fanout4645 (.A(net4647),
    .X(net4645));
 sg13g2_buf_8 fanout4646 (.A(net4647),
    .X(net4646));
 sg13g2_buf_8 fanout4647 (.A(net4655),
    .X(net4647));
 sg13g2_buf_8 fanout4648 (.A(net4651),
    .X(net4648));
 sg13g2_buf_8 fanout4649 (.A(net4651),
    .X(net4649));
 sg13g2_buf_8 fanout4650 (.A(net4651),
    .X(net4650));
 sg13g2_buf_8 fanout4651 (.A(net4655),
    .X(net4651));
 sg13g2_buf_8 fanout4652 (.A(net4654),
    .X(net4652));
 sg13g2_buf_1 fanout4653 (.A(net4654),
    .X(net4653));
 sg13g2_buf_8 fanout4654 (.A(net4655),
    .X(net4654));
 sg13g2_buf_8 fanout4655 (.A(net4679),
    .X(net4655));
 sg13g2_buf_8 fanout4656 (.A(net4658),
    .X(net4656));
 sg13g2_buf_1 fanout4657 (.A(net4658),
    .X(net4657));
 sg13g2_buf_2 fanout4658 (.A(net4659),
    .X(net4658));
 sg13g2_buf_8 fanout4659 (.A(net4679),
    .X(net4659));
 sg13g2_buf_8 fanout4660 (.A(net4661),
    .X(net4660));
 sg13g2_buf_8 fanout4661 (.A(net4669),
    .X(net4661));
 sg13g2_buf_8 fanout4662 (.A(net4663),
    .X(net4662));
 sg13g2_buf_8 fanout4663 (.A(net4669),
    .X(net4663));
 sg13g2_buf_8 fanout4664 (.A(net4666),
    .X(net4664));
 sg13g2_buf_8 fanout4665 (.A(net4666),
    .X(net4665));
 sg13g2_buf_8 fanout4666 (.A(net4669),
    .X(net4666));
 sg13g2_buf_8 fanout4667 (.A(net4669),
    .X(net4667));
 sg13g2_buf_1 fanout4668 (.A(net4669),
    .X(net4668));
 sg13g2_buf_8 fanout4669 (.A(net4679),
    .X(net4669));
 sg13g2_buf_8 fanout4670 (.A(net4672),
    .X(net4670));
 sg13g2_buf_8 fanout4671 (.A(net4672),
    .X(net4671));
 sg13g2_buf_8 fanout4672 (.A(net4678),
    .X(net4672));
 sg13g2_buf_8 fanout4673 (.A(net4678),
    .X(net4673));
 sg13g2_buf_1 fanout4674 (.A(net4675),
    .X(net4674));
 sg13g2_buf_8 fanout4675 (.A(net4678),
    .X(net4675));
 sg13g2_buf_8 fanout4676 (.A(net4677),
    .X(net4676));
 sg13g2_buf_8 fanout4677 (.A(net4678),
    .X(net4677));
 sg13g2_buf_8 fanout4678 (.A(net4679),
    .X(net4678));
 sg13g2_buf_8 fanout4679 (.A(net4724),
    .X(net4679));
 sg13g2_buf_8 fanout4680 (.A(net4688),
    .X(net4680));
 sg13g2_buf_8 fanout4681 (.A(net4682),
    .X(net4681));
 sg13g2_buf_8 fanout4682 (.A(net4688),
    .X(net4682));
 sg13g2_buf_8 fanout4683 (.A(net4685),
    .X(net4683));
 sg13g2_buf_1 fanout4684 (.A(net4685),
    .X(net4684));
 sg13g2_buf_8 fanout4685 (.A(net4688),
    .X(net4685));
 sg13g2_buf_8 fanout4686 (.A(net4687),
    .X(net4686));
 sg13g2_buf_8 fanout4687 (.A(net4688),
    .X(net4687));
 sg13g2_buf_8 fanout4688 (.A(net4724),
    .X(net4688));
 sg13g2_buf_8 fanout4689 (.A(net4691),
    .X(net4689));
 sg13g2_buf_8 fanout4690 (.A(net4691),
    .X(net4690));
 sg13g2_buf_2 fanout4691 (.A(net4699),
    .X(net4691));
 sg13g2_buf_8 fanout4692 (.A(net4699),
    .X(net4692));
 sg13g2_buf_8 fanout4693 (.A(net4699),
    .X(net4693));
 sg13g2_buf_1 fanout4694 (.A(net4699),
    .X(net4694));
 sg13g2_buf_8 fanout4695 (.A(net4696),
    .X(net4695));
 sg13g2_buf_1 fanout4696 (.A(net4697),
    .X(net4696));
 sg13g2_buf_1 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_8 fanout4698 (.A(net4699),
    .X(net4698));
 sg13g2_buf_8 fanout4699 (.A(net4724),
    .X(net4699));
 sg13g2_buf_8 fanout4700 (.A(net4702),
    .X(net4700));
 sg13g2_buf_1 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_8 fanout4702 (.A(net4723),
    .X(net4702));
 sg13g2_buf_8 fanout4703 (.A(net4704),
    .X(net4703));
 sg13g2_buf_8 fanout4704 (.A(net4705),
    .X(net4704));
 sg13g2_buf_8 fanout4705 (.A(net4723),
    .X(net4705));
 sg13g2_buf_8 fanout4706 (.A(net4708),
    .X(net4706));
 sg13g2_buf_8 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_8 fanout4708 (.A(net4723),
    .X(net4708));
 sg13g2_buf_8 fanout4709 (.A(net4712),
    .X(net4709));
 sg13g2_buf_8 fanout4710 (.A(net4711),
    .X(net4710));
 sg13g2_buf_8 fanout4711 (.A(net4712),
    .X(net4711));
 sg13g2_buf_8 fanout4712 (.A(net4713),
    .X(net4712));
 sg13g2_buf_8 fanout4713 (.A(net4723),
    .X(net4713));
 sg13g2_buf_8 fanout4714 (.A(net4715),
    .X(net4714));
 sg13g2_buf_8 fanout4715 (.A(net4716),
    .X(net4715));
 sg13g2_buf_8 fanout4716 (.A(net4723),
    .X(net4716));
 sg13g2_buf_8 fanout4717 (.A(net4722),
    .X(net4717));
 sg13g2_buf_1 fanout4718 (.A(net4719),
    .X(net4718));
 sg13g2_buf_8 fanout4719 (.A(net4722),
    .X(net4719));
 sg13g2_buf_8 fanout4720 (.A(net4722),
    .X(net4720));
 sg13g2_buf_1 fanout4721 (.A(net4722),
    .X(net4721));
 sg13g2_buf_8 fanout4722 (.A(net4723),
    .X(net4722));
 sg13g2_buf_8 fanout4723 (.A(net4724),
    .X(net4723));
 sg13g2_buf_8 fanout4724 (.A(\u_inv.f_next[0] ),
    .X(net4724));
 sg13g2_buf_8 fanout4725 (.A(net4726),
    .X(net4725));
 sg13g2_buf_1 fanout4726 (.A(net4732),
    .X(net4726));
 sg13g2_buf_8 fanout4727 (.A(net4732),
    .X(net4727));
 sg13g2_buf_1 fanout4728 (.A(net4732),
    .X(net4728));
 sg13g2_buf_8 fanout4729 (.A(net4732),
    .X(net4729));
 sg13g2_buf_1 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(net4732),
    .X(net4731));
 sg13g2_buf_8 fanout4732 (.A(net4739),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(net4736),
    .X(net4733));
 sg13g2_buf_8 fanout4734 (.A(net4736),
    .X(net4734));
 sg13g2_buf_1 fanout4735 (.A(net4736),
    .X(net4735));
 sg13g2_buf_8 fanout4736 (.A(net4739),
    .X(net4736));
 sg13g2_buf_8 fanout4737 (.A(net4739),
    .X(net4737));
 sg13g2_buf_1 fanout4738 (.A(net4739),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(net4765),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(net4744),
    .X(net4740));
 sg13g2_buf_1 fanout4741 (.A(net4744),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(net4744),
    .X(net4742));
 sg13g2_buf_1 fanout4743 (.A(net4744),
    .X(net4743));
 sg13g2_buf_2 fanout4744 (.A(net4765),
    .X(net4744));
 sg13g2_buf_8 fanout4745 (.A(net4747),
    .X(net4745));
 sg13g2_buf_1 fanout4746 (.A(net4749),
    .X(net4746));
 sg13g2_buf_8 fanout4747 (.A(net4749),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(net4749),
    .X(net4748));
 sg13g2_buf_8 fanout4749 (.A(net4765),
    .X(net4749));
 sg13g2_buf_8 fanout4750 (.A(net4755),
    .X(net4750));
 sg13g2_buf_8 fanout4751 (.A(net4752),
    .X(net4751));
 sg13g2_buf_1 fanout4752 (.A(net4753),
    .X(net4752));
 sg13g2_buf_1 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(net4755),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(net4764),
    .X(net4755));
 sg13g2_buf_8 fanout4756 (.A(net4757),
    .X(net4756));
 sg13g2_buf_1 fanout4757 (.A(net4758),
    .X(net4757));
 sg13g2_buf_1 fanout4758 (.A(net4763),
    .X(net4758));
 sg13g2_buf_8 fanout4759 (.A(net4760),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(net4761),
    .X(net4760));
 sg13g2_buf_1 fanout4761 (.A(net4763),
    .X(net4761));
 sg13g2_buf_8 fanout4762 (.A(net4763),
    .X(net4762));
 sg13g2_buf_8 fanout4763 (.A(net4764),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(net4765),
    .X(net4764));
 sg13g2_buf_8 fanout4765 (.A(\u_inv.f_reg[256] ),
    .X(net4765));
 sg13g2_buf_8 fanout4766 (.A(net2904),
    .X(net4766));
 sg13g2_buf_8 fanout4767 (.A(net3188),
    .X(net4767));
 sg13g2_buf_8 fanout4768 (.A(\u_inv.d_reg[226] ),
    .X(net4768));
 sg13g2_buf_8 fanout4769 (.A(\u_inv.d_reg[209] ),
    .X(net4769));
 sg13g2_buf_8 fanout4770 (.A(\u_inv.d_reg[208] ),
    .X(net4770));
 sg13g2_buf_8 fanout4771 (.A(net3087),
    .X(net4771));
 sg13g2_buf_8 fanout4772 (.A(\u_inv.d_reg[197] ),
    .X(net4772));
 sg13g2_buf_8 fanout4773 (.A(net3239),
    .X(net4773));
 sg13g2_buf_8 fanout4774 (.A(\u_inv.d_reg[187] ),
    .X(net4774));
 sg13g2_buf_8 fanout4775 (.A(net4963),
    .X(net4775));
 sg13g2_buf_8 fanout4776 (.A(\u_inv.d_reg[150] ),
    .X(net4776));
 sg13g2_buf_8 fanout4777 (.A(net3307),
    .X(net4777));
 sg13g2_buf_8 fanout4778 (.A(net4962),
    .X(net4778));
 sg13g2_buf_8 fanout4779 (.A(net2978),
    .X(net4779));
 sg13g2_buf_8 fanout4780 (.A(net3016),
    .X(net4780));
 sg13g2_buf_8 fanout4781 (.A(\u_inv.d_reg[77] ),
    .X(net4781));
 sg13g2_buf_8 fanout4782 (.A(net3198),
    .X(net4782));
 sg13g2_buf_8 fanout4783 (.A(net3070),
    .X(net4783));
 sg13g2_buf_8 fanout4784 (.A(net3247),
    .X(net4784));
 sg13g2_buf_8 fanout4785 (.A(\u_inv.d_reg[58] ),
    .X(net4785));
 sg13g2_buf_8 fanout4786 (.A(\u_inv.d_reg[42] ),
    .X(net4786));
 sg13g2_buf_8 fanout4787 (.A(\u_inv.d_reg[26] ),
    .X(net4787));
 sg13g2_buf_8 fanout4788 (.A(net3062),
    .X(net4788));
 sg13g2_buf_8 fanout4789 (.A(net3222),
    .X(net4789));
 sg13g2_buf_8 fanout4790 (.A(\u_inv.d_reg[18] ),
    .X(net4790));
 sg13g2_buf_8 fanout4791 (.A(\u_inv.d_reg[17] ),
    .X(net4791));
 sg13g2_buf_8 fanout4792 (.A(\u_inv.d_reg[11] ),
    .X(net4792));
 sg13g2_buf_1 fanout4793 (.A(\u_inv.d_reg[11] ),
    .X(net4793));
 sg13g2_buf_8 fanout4794 (.A(\u_inv.d_reg[7] ),
    .X(net4794));
 sg13g2_buf_8 fanout4795 (.A(net1450),
    .X(net4795));
 sg13g2_buf_8 fanout4796 (.A(net3096),
    .X(net4796));
 sg13g2_buf_8 fanout4797 (.A(\u_inv.d_reg[1] ),
    .X(net4797));
 sg13g2_buf_1 fanout4798 (.A(\u_inv.d_reg[1] ),
    .X(net4798));
 sg13g2_buf_8 fanout4799 (.A(\u_inv.d_reg[0] ),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(\u_inv.d_reg[0] ),
    .X(net4800));
 sg13g2_buf_8 fanout4801 (.A(net3031),
    .X(net4801));
 sg13g2_buf_8 fanout4802 (.A(net3148),
    .X(net4802));
 sg13g2_buf_8 fanout4803 (.A(net1949),
    .X(net4803));
 sg13g2_buf_8 fanout4804 (.A(net3229),
    .X(net4804));
 sg13g2_buf_8 fanout4805 (.A(net4960),
    .X(net4805));
 sg13g2_buf_8 fanout4806 (.A(net2170),
    .X(net4806));
 sg13g2_buf_8 fanout4807 (.A(net4810),
    .X(net4807));
 sg13g2_buf_8 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_8 fanout4809 (.A(net4810),
    .X(net4809));
 sg13g2_buf_8 fanout4810 (.A(net4878),
    .X(net4810));
 sg13g2_buf_8 fanout4811 (.A(net4816),
    .X(net4811));
 sg13g2_buf_8 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_8 fanout4813 (.A(net4816),
    .X(net4813));
 sg13g2_buf_8 fanout4814 (.A(net4816),
    .X(net4814));
 sg13g2_buf_8 fanout4815 (.A(net4816),
    .X(net4815));
 sg13g2_buf_8 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_8 fanout4817 (.A(net4826),
    .X(net4817));
 sg13g2_buf_8 fanout4818 (.A(net4820),
    .X(net4818));
 sg13g2_buf_2 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_8 fanout4820 (.A(net4826),
    .X(net4820));
 sg13g2_buf_8 fanout4821 (.A(net4823),
    .X(net4821));
 sg13g2_buf_8 fanout4822 (.A(net4823),
    .X(net4822));
 sg13g2_buf_8 fanout4823 (.A(net4826),
    .X(net4823));
 sg13g2_buf_8 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_8 fanout4825 (.A(net4826),
    .X(net4825));
 sg13g2_buf_8 fanout4826 (.A(net4878),
    .X(net4826));
 sg13g2_buf_8 fanout4827 (.A(net4835),
    .X(net4827));
 sg13g2_buf_8 fanout4828 (.A(net4835),
    .X(net4828));
 sg13g2_buf_8 fanout4829 (.A(net4831),
    .X(net4829));
 sg13g2_buf_8 fanout4830 (.A(net4831),
    .X(net4830));
 sg13g2_buf_8 fanout4831 (.A(net4835),
    .X(net4831));
 sg13g2_buf_8 fanout4832 (.A(net4834),
    .X(net4832));
 sg13g2_buf_8 fanout4833 (.A(net4834),
    .X(net4833));
 sg13g2_buf_8 fanout4834 (.A(net4835),
    .X(net4834));
 sg13g2_buf_8 fanout4835 (.A(net4843),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(net4843),
    .X(net4836));
 sg13g2_buf_8 fanout4837 (.A(net4843),
    .X(net4837));
 sg13g2_buf_8 fanout4838 (.A(net4841),
    .X(net4838));
 sg13g2_buf_8 fanout4839 (.A(net4840),
    .X(net4839));
 sg13g2_buf_8 fanout4840 (.A(net4841),
    .X(net4840));
 sg13g2_buf_8 fanout4841 (.A(net4842),
    .X(net4841));
 sg13g2_buf_8 fanout4842 (.A(net4843),
    .X(net4842));
 sg13g2_buf_8 fanout4843 (.A(net4878),
    .X(net4843));
 sg13g2_buf_8 fanout4844 (.A(net4846),
    .X(net4844));
 sg13g2_buf_8 fanout4845 (.A(net4846),
    .X(net4845));
 sg13g2_buf_8 fanout4846 (.A(net4859),
    .X(net4846));
 sg13g2_buf_8 fanout4847 (.A(net4849),
    .X(net4847));
 sg13g2_buf_8 fanout4848 (.A(net4849),
    .X(net4848));
 sg13g2_buf_8 fanout4849 (.A(net4850),
    .X(net4849));
 sg13g2_buf_8 fanout4850 (.A(net4859),
    .X(net4850));
 sg13g2_buf_8 fanout4851 (.A(net4853),
    .X(net4851));
 sg13g2_buf_8 fanout4852 (.A(net4854),
    .X(net4852));
 sg13g2_buf_8 fanout4853 (.A(net4854),
    .X(net4853));
 sg13g2_buf_8 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_8 fanout4855 (.A(net4859),
    .X(net4855));
 sg13g2_buf_8 fanout4856 (.A(net4857),
    .X(net4856));
 sg13g2_buf_8 fanout4857 (.A(net4858),
    .X(net4857));
 sg13g2_buf_2 fanout4858 (.A(net4859),
    .X(net4858));
 sg13g2_buf_8 fanout4859 (.A(net4877),
    .X(net4859));
 sg13g2_buf_8 fanout4860 (.A(net4865),
    .X(net4860));
 sg13g2_buf_8 fanout4861 (.A(net4865),
    .X(net4861));
 sg13g2_buf_8 fanout4862 (.A(net4865),
    .X(net4862));
 sg13g2_buf_8 fanout4863 (.A(net4864),
    .X(net4863));
 sg13g2_buf_8 fanout4864 (.A(net4865),
    .X(net4864));
 sg13g2_buf_8 fanout4865 (.A(net4877),
    .X(net4865));
 sg13g2_buf_8 fanout4866 (.A(net4869),
    .X(net4866));
 sg13g2_buf_8 fanout4867 (.A(net4869),
    .X(net4867));
 sg13g2_buf_8 fanout4868 (.A(net4869),
    .X(net4868));
 sg13g2_buf_8 fanout4869 (.A(net4877),
    .X(net4869));
 sg13g2_buf_8 fanout4870 (.A(net4871),
    .X(net4870));
 sg13g2_buf_8 fanout4871 (.A(net4876),
    .X(net4871));
 sg13g2_buf_8 fanout4872 (.A(net4874),
    .X(net4872));
 sg13g2_buf_8 fanout4873 (.A(net4874),
    .X(net4873));
 sg13g2_buf_8 fanout4874 (.A(net4876),
    .X(net4874));
 sg13g2_buf_8 fanout4875 (.A(net4876),
    .X(net4875));
 sg13g2_buf_8 fanout4876 (.A(net4877),
    .X(net4876));
 sg13g2_buf_8 fanout4877 (.A(net4878),
    .X(net4877));
 sg13g2_buf_8 fanout4878 (.A(net4951),
    .X(net4878));
 sg13g2_buf_8 fanout4879 (.A(net4880),
    .X(net4879));
 sg13g2_buf_2 fanout4880 (.A(net4881),
    .X(net4880));
 sg13g2_buf_8 fanout4881 (.A(net4883),
    .X(net4881));
 sg13g2_buf_8 fanout4882 (.A(net4883),
    .X(net4882));
 sg13g2_buf_8 fanout4883 (.A(net4909),
    .X(net4883));
 sg13g2_buf_8 fanout4884 (.A(net4885),
    .X(net4884));
 sg13g2_buf_8 fanout4885 (.A(net4888),
    .X(net4885));
 sg13g2_buf_8 fanout4886 (.A(net4887),
    .X(net4886));
 sg13g2_buf_8 fanout4887 (.A(net4888),
    .X(net4887));
 sg13g2_buf_8 fanout4888 (.A(net4909),
    .X(net4888));
 sg13g2_buf_8 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_8 fanout4890 (.A(net4893),
    .X(net4890));
 sg13g2_buf_8 fanout4891 (.A(net4892),
    .X(net4891));
 sg13g2_buf_8 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_8 fanout4893 (.A(net4909),
    .X(net4893));
 sg13g2_buf_8 fanout4894 (.A(net4908),
    .X(net4894));
 sg13g2_buf_2 fanout4895 (.A(net4908),
    .X(net4895));
 sg13g2_buf_8 fanout4896 (.A(net4898),
    .X(net4896));
 sg13g2_buf_8 fanout4897 (.A(net4898),
    .X(net4897));
 sg13g2_buf_8 fanout4898 (.A(net4907),
    .X(net4898));
 sg13g2_buf_8 fanout4899 (.A(net4900),
    .X(net4899));
 sg13g2_buf_8 fanout4900 (.A(net4907),
    .X(net4900));
 sg13g2_buf_8 fanout4901 (.A(net4903),
    .X(net4901));
 sg13g2_buf_8 fanout4902 (.A(net4906),
    .X(net4902));
 sg13g2_buf_8 fanout4903 (.A(net4906),
    .X(net4903));
 sg13g2_buf_8 fanout4904 (.A(net4905),
    .X(net4904));
 sg13g2_buf_8 fanout4905 (.A(net4906),
    .X(net4905));
 sg13g2_buf_8 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_8 fanout4907 (.A(net4908),
    .X(net4907));
 sg13g2_buf_8 fanout4908 (.A(net4909),
    .X(net4908));
 sg13g2_buf_8 fanout4909 (.A(net4951),
    .X(net4909));
 sg13g2_buf_8 fanout4910 (.A(net4913),
    .X(net4910));
 sg13g2_buf_8 fanout4911 (.A(net4913),
    .X(net4911));
 sg13g2_buf_8 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_8 fanout4913 (.A(net4919),
    .X(net4913));
 sg13g2_buf_8 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_8 fanout4915 (.A(net4918),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4917),
    .X(net4916));
 sg13g2_buf_8 fanout4917 (.A(net4918),
    .X(net4917));
 sg13g2_buf_8 fanout4918 (.A(net4919),
    .X(net4918));
 sg13g2_buf_8 fanout4919 (.A(net4920),
    .X(net4919));
 sg13g2_buf_8 fanout4920 (.A(net4951),
    .X(net4920));
 sg13g2_buf_8 fanout4921 (.A(net4923),
    .X(net4921));
 sg13g2_buf_1 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_8 fanout4923 (.A(net4950),
    .X(net4923));
 sg13g2_buf_8 fanout4924 (.A(net4926),
    .X(net4924));
 sg13g2_buf_8 fanout4925 (.A(net4926),
    .X(net4925));
 sg13g2_buf_8 fanout4926 (.A(net4927),
    .X(net4926));
 sg13g2_buf_8 fanout4927 (.A(net4950),
    .X(net4927));
 sg13g2_buf_8 fanout4928 (.A(net4930),
    .X(net4928));
 sg13g2_buf_8 fanout4929 (.A(net4930),
    .X(net4929));
 sg13g2_buf_8 fanout4930 (.A(net4937),
    .X(net4930));
 sg13g2_buf_8 fanout4931 (.A(net4937),
    .X(net4931));
 sg13g2_buf_8 fanout4932 (.A(net4937),
    .X(net4932));
 sg13g2_buf_8 fanout4933 (.A(net4934),
    .X(net4933));
 sg13g2_buf_8 fanout4934 (.A(net4936),
    .X(net4934));
 sg13g2_buf_8 fanout4935 (.A(net4936),
    .X(net4935));
 sg13g2_buf_8 fanout4936 (.A(net4937),
    .X(net4936));
 sg13g2_buf_8 fanout4937 (.A(net4950),
    .X(net4937));
 sg13g2_buf_8 fanout4938 (.A(net4939),
    .X(net4938));
 sg13g2_buf_8 fanout4939 (.A(net4949),
    .X(net4939));
 sg13g2_buf_8 fanout4940 (.A(net4944),
    .X(net4940));
 sg13g2_buf_2 fanout4941 (.A(net4944),
    .X(net4941));
 sg13g2_buf_8 fanout4942 (.A(net4944),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_2 fanout4944 (.A(net4949),
    .X(net4944));
 sg13g2_buf_8 fanout4945 (.A(net4947),
    .X(net4945));
 sg13g2_buf_8 fanout4946 (.A(net4947),
    .X(net4946));
 sg13g2_buf_8 fanout4947 (.A(net4949),
    .X(net4947));
 sg13g2_buf_2 fanout4948 (.A(net4949),
    .X(net4948));
 sg13g2_buf_8 fanout4949 (.A(net4950),
    .X(net4949));
 sg13g2_buf_8 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_8 fanout4951 (.A(rst_n),
    .X(net4951));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_tielo tt_um_corey_11 (.L_LO(net11));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_8 clkbuf_5_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0_0_clk));
 sg13g2_buf_8 clkbuf_5_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1_0_clk));
 sg13g2_buf_8 clkbuf_5_2_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2_0_clk));
 sg13g2_buf_8 clkbuf_5_3_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3_0_clk));
 sg13g2_buf_8 clkbuf_5_4_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4_0_clk));
 sg13g2_buf_8 clkbuf_5_5_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5_0_clk));
 sg13g2_buf_8 clkbuf_5_6_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6_0_clk));
 sg13g2_buf_8 clkbuf_5_7_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7_0_clk));
 sg13g2_buf_8 clkbuf_5_8_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8_0_clk));
 sg13g2_buf_8 clkbuf_5_9_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9_0_clk));
 sg13g2_buf_8 clkbuf_5_10_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10_0_clk));
 sg13g2_buf_8 clkbuf_5_11_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11_0_clk));
 sg13g2_buf_8 clkbuf_5_12_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12_0_clk));
 sg13g2_buf_8 clkbuf_5_13_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13_0_clk));
 sg13g2_buf_8 clkbuf_5_14_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14_0_clk));
 sg13g2_buf_8 clkbuf_5_15_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15_0_clk));
 sg13g2_buf_8 clkbuf_5_16_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16_0_clk));
 sg13g2_buf_8 clkbuf_5_17_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17_0_clk));
 sg13g2_buf_8 clkbuf_5_18_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18_0_clk));
 sg13g2_buf_8 clkbuf_5_19_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19_0_clk));
 sg13g2_buf_8 clkbuf_5_20_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20_0_clk));
 sg13g2_buf_8 clkbuf_5_21_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21_0_clk));
 sg13g2_buf_8 clkbuf_5_22_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22_0_clk));
 sg13g2_buf_8 clkbuf_5_23_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23_0_clk));
 sg13g2_buf_8 clkbuf_5_24_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24_0_clk));
 sg13g2_buf_8 clkbuf_5_25_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25_0_clk));
 sg13g2_buf_8 clkbuf_5_26_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26_0_clk));
 sg13g2_buf_8 clkbuf_5_27_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27_0_clk));
 sg13g2_buf_8 clkbuf_5_28_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28_0_clk));
 sg13g2_buf_8 clkbuf_5_29_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29_0_clk));
 sg13g2_buf_8 clkbuf_5_30_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30_0_clk));
 sg13g2_buf_8 clkbuf_5_31_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31_0_clk));
 sg13g2_buf_8 clkbuf_6_0__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_8 clkbuf_6_1__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkbuf_6_2__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkbuf_6_3__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkbuf_6_4__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkbuf_6_5__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkbuf_6_6__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkbuf_6_7__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkbuf_6_8__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_8 clkbuf_6_9__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkbuf_6_10__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkbuf_6_11__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkbuf_6_12__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkbuf_6_13__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkbuf_6_14__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkbuf_6_15__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkbuf_6_16__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_8 clkbuf_6_17__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkbuf_6_18__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkbuf_6_19__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkbuf_6_20__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkbuf_6_21__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkbuf_6_22__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkbuf_6_23__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkbuf_6_24__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_8 clkbuf_6_25__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkbuf_6_26__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkbuf_6_27__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkbuf_6_28__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkbuf_6_29__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkbuf_6_30__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkbuf_6_31__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkbuf_6_32__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_8 clkbuf_6_33__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkbuf_6_34__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkbuf_6_35__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkbuf_6_36__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkbuf_6_37__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkbuf_6_38__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkbuf_6_39__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkbuf_6_40__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_8 clkbuf_6_41__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkbuf_6_42__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkbuf_6_43__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkbuf_6_44__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkbuf_6_45__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkbuf_6_46__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkbuf_6_47__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkbuf_6_48__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_8 clkbuf_6_49__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkbuf_6_50__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkbuf_6_51__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkbuf_6_52__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkbuf_6_53__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkbuf_6_54__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkbuf_6_55__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkbuf_6_56__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_8 clkbuf_6_57__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkbuf_6_58__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkbuf_6_59__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkbuf_6_60__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_8 clkbuf_6_61__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkbuf_6_62__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkbuf_6_63__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_53__leaf_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_78_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_leaf_222_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_223_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_215_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_leaf_18_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_0_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_233_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_196_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_194_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_208_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_213_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_176_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_117_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_124_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_inv.load_input ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00002_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_inv.d_next[184] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold4 (.A(_05619_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_inv.counter[9] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00276_),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold7 (.A(\byte_cnt[0] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00005_),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold9 (.A(\inv_result[230] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold10 (.A(\inv_result[37] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold11 (.A(\inv_result[224] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold12 (.A(\inv_result[35] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_inv.counter[7] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00274_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold15 (.A(\inv_result[43] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold16 (.A(\inv_result[42] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold17 (.A(\inv_result[227] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold18 (.A(\inv_result[56] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold19 (.A(\inv_result[202] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold20 (.A(\inv_result[114] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold21 (.A(\inv_result[222] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold22 (.A(\inv_result[193] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold23 (.A(\inv_result[172] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold24 (.A(\shift_reg[250] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold25 (.A(_00261_),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_inv.counter[3] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold27 (.A(_00270_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold28 (.A(\shift_reg[223] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold29 (.A(_00234_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold30 (.A(\inv_result[210] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold31 (.A(\inv_result[170] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold32 (.A(\inv_result[54] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold33 (.A(\inv_result[62] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold34 (.A(\inv_result[166] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold35 (.A(\shift_reg[249] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00260_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold37 (.A(\shift_reg[254] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold38 (.A(_00265_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold39 (.A(\inv_result[74] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold40 (.A(\byte_cnt[3] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold41 (.A(_11061_),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold42 (.A(_00008_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold43 (.A(\shift_reg[239] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold44 (.A(_00250_),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold45 (.A(\shift_reg[114] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold46 (.A(_00125_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold47 (.A(\shift_reg[255] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold48 (.A(_00266_),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold49 (.A(\inv_result[126] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold50 (.A(\shift_reg[127] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00138_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold52 (.A(\inv_result[221] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold53 (.A(\shift_reg[251] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold54 (.A(_00262_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold55 (.A(\inv_result[7] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold56 (.A(\shift_reg[237] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold57 (.A(_00248_),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold58 (.A(\inv_result[118] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold59 (.A(\shift_reg[253] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00264_),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold61 (.A(\shift_reg[51] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00062_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold63 (.A(\shift_reg[216] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold64 (.A(_00227_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold65 (.A(\shift_reg[248] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold66 (.A(_00259_),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold67 (.A(\shift_reg[234] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00245_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold69 (.A(\inv_result[205] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold70 (.A(\shift_reg[33] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold71 (.A(_00044_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold72 (.A(\inv_result[80] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold73 (.A(\inv_result[102] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold74 (.A(\shift_reg[215] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00226_),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold76 (.A(\shift_reg[241] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00252_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold78 (.A(\inv_result[171] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold79 (.A(\inv_result[48] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold80 (.A(\inv_result[243] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold81 (.A(\shift_reg[13] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold82 (.A(_00024_),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold83 (.A(\inv_result[195] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold84 (.A(\shift_reg[227] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00238_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold86 (.A(\shift_reg[31] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold87 (.A(_00042_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_inv.counter[0] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold89 (.A(\shift_reg[44] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold90 (.A(_00055_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold91 (.A(\shift_reg[252] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold92 (.A(_00263_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold93 (.A(\shift_reg[30] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00041_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold95 (.A(\shift_reg[69] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00080_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold97 (.A(\inv_result[229] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold98 (.A(\shift_reg[28] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold99 (.A(_00039_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold100 (.A(\shift_reg[35] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00046_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold102 (.A(\shift_reg[209] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold103 (.A(_00220_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold104 (.A(\inv_result[132] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold105 (.A(\shift_reg[183] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00194_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold107 (.A(\shift_reg[4] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold108 (.A(_00015_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold109 (.A(\inv_result[213] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold110 (.A(\inv_result[2] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold111 (.A(\shift_reg[105] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold112 (.A(_00116_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold113 (.A(\inv_result[192] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold114 (.A(\inv_result[134] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold115 (.A(\inv_result[91] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold116 (.A(\shift_reg[138] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00149_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold118 (.A(\shift_reg[124] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold119 (.A(_00135_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold120 (.A(\shift_reg[213] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold121 (.A(_00224_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold122 (.A(\inv_result[32] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold123 (.A(\inv_result[70] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold124 (.A(\inv_result[179] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold125 (.A(\inv_result[150] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold126 (.A(\shift_reg[232] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold127 (.A(_00243_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold128 (.A(\shift_reg[6] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold129 (.A(_01568_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold130 (.A(\shift_reg[229] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold131 (.A(_00240_),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold132 (.A(\shift_reg[236] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00247_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold134 (.A(\shift_reg[108] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold135 (.A(_00119_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold136 (.A(\shift_reg[50] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00061_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold138 (.A(\shift_reg[203] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold139 (.A(_00214_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold140 (.A(\shift_reg[230] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold141 (.A(_00241_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold142 (.A(\shift_reg[93] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold143 (.A(_00104_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold144 (.A(\inv_result[9] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold145 (.A(_01057_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold146 (.A(\shift_reg[72] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold147 (.A(_00083_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold148 (.A(\shift_reg[26] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold149 (.A(_00037_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold150 (.A(\shift_reg[12] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold151 (.A(_00023_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_inv.input_reg[4] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold153 (.A(\byte_cnt[4] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold154 (.A(_11048_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold155 (.A(_00000_),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold156 (.A(\shift_reg[132] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_inv.input_reg[159] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold158 (.A(_01463_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold159 (.A(\shift_reg[136] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold160 (.A(_00147_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold161 (.A(\inv_result[40] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold162 (.A(\inv_result[147] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold163 (.A(\inv_result[241] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold164 (.A(_01289_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_inv.counter[8] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold166 (.A(_13596_),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold167 (.A(_00275_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold168 (.A(\shift_reg[25] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold169 (.A(_00036_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold170 (.A(\shift_reg[55] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold171 (.A(_00066_),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold172 (.A(\shift_reg[139] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold173 (.A(_00150_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold174 (.A(\inv_result[65] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold175 (.A(\inv_result[237] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold176 (.A(\shift_reg[74] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold177 (.A(_00085_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold178 (.A(\inv_result[168] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold179 (.A(\shift_reg[11] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00022_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold181 (.A(\shift_reg[164] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold182 (.A(_00175_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold183 (.A(\inv_result[85] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold184 (.A(\inv_result[141] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold185 (.A(\shift_reg[87] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold186 (.A(_00098_),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold187 (.A(\shift_reg[9] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00020_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold189 (.A(\shift_reg[21] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold190 (.A(_00032_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold191 (.A(\shift_reg[85] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold192 (.A(_00096_),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold193 (.A(\inv_result[44] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold194 (.A(\inv_result[52] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold195 (.A(\shift_reg[71] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold196 (.A(_00082_),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold197 (.A(\shift_reg[117] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold198 (.A(_00128_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold199 (.A(\shift_reg[38] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold200 (.A(_00049_),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold201 (.A(\inv_result[140] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold202 (.A(\inv_result[106] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold203 (.A(\shift_reg[133] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold204 (.A(_00144_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_inv.input_reg[3] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold206 (.A(_01565_),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold207 (.A(\shift_reg[166] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00177_),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold209 (.A(\inv_result[137] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold210 (.A(\shift_reg[177] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold211 (.A(_00188_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold212 (.A(\shift_reg[42] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold213 (.A(_00053_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold214 (.A(\shift_reg[160] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold215 (.A(_00171_),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold216 (.A(\shift_reg[52] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold217 (.A(\inv_result[133] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold218 (.A(\shift_reg[193] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold219 (.A(_00204_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold220 (.A(\shift_reg[81] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00092_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold222 (.A(\shift_reg[54] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold223 (.A(_00065_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold224 (.A(\shift_reg[68] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00079_),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold226 (.A(\shift_reg[131] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold227 (.A(_00142_),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold228 (.A(\inv_result[190] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold229 (.A(\shift_reg[88] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold230 (.A(_00099_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold231 (.A(\inv_result[185] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold232 (.A(\byte_cnt[1] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold233 (.A(_11057_),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold234 (.A(_00006_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_inv.f_reg[0] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold236 (.A(\inv_result[93] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold237 (.A(\inv_result[59] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_inv.input_reg[5] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold239 (.A(_01567_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold240 (.A(\shift_reg[238] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold241 (.A(_00249_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold242 (.A(\shift_reg[175] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold243 (.A(_00186_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold244 (.A(\shift_reg[214] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00225_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold246 (.A(\inv_result[174] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold247 (.A(\inv_result[164] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold248 (.A(\shift_reg[41] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold249 (.A(_00052_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold250 (.A(\shift_reg[162] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold251 (.A(_00173_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold252 (.A(\inv_result[131] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold253 (.A(\shift_reg[204] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold254 (.A(_00215_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold255 (.A(\shift_reg[79] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold256 (.A(_00090_),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold257 (.A(\shift_reg[233] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold258 (.A(_00244_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold259 (.A(\inv_result[23] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold260 (.A(\inv_result[218] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold261 (.A(\shift_reg[207] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00218_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold263 (.A(\inv_result[109] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold264 (.A(\shift_reg[128] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold265 (.A(_00139_),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold266 (.A(\shift_reg[89] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00100_),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold268 (.A(\shift_reg[94] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00105_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold270 (.A(\shift_reg[62] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold271 (.A(\shift_reg[170] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold272 (.A(\inv_result[128] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold273 (.A(\inv_result[212] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold274 (.A(\shift_reg[40] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold275 (.A(_00051_),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold276 (.A(\inv_result[184] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold277 (.A(\shift_reg[80] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold278 (.A(\shift_reg[235] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold279 (.A(_00246_),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold280 (.A(\inv_result[20] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold281 (.A(\shift_reg[83] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold282 (.A(_00094_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold283 (.A(\shift_reg[191] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold284 (.A(_00202_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold285 (.A(\shift_reg[5] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold286 (.A(_00016_),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold287 (.A(\inv_result[198] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold288 (.A(\shift_reg[56] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00067_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold290 (.A(\inv_result[146] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold291 (.A(\shift_reg[112] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold292 (.A(_00123_),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold293 (.A(\shift_reg[37] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00048_),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold295 (.A(\shift_reg[202] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold296 (.A(_00213_),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold297 (.A(\shift_reg[22] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold298 (.A(_00033_),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold299 (.A(\shift_reg[97] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold300 (.A(_00108_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold301 (.A(\inv_result[136] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold302 (.A(\shift_reg[140] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold303 (.A(\shift_reg[161] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold304 (.A(_00172_),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold305 (.A(\inv_result[115] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold306 (.A(\inv_result[204] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold307 (.A(\shift_reg[1] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold308 (.A(_00012_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold309 (.A(\shift_reg[208] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00219_),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold311 (.A(\inv_result[160] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold312 (.A(\inv_result[200] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold313 (.A(\inv_result[244] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold314 (.A(_01292_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold315 (.A(\inv_result[61] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold316 (.A(\shift_reg[90] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00101_),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold318 (.A(\shift_reg[78] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold319 (.A(_00089_),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold320 (.A(\inv_result[225] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold321 (.A(\shift_reg[59] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold322 (.A(\shift_reg[32] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold323 (.A(_00043_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold324 (.A(\shift_reg[67] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold325 (.A(_00078_),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold326 (.A(\shift_reg[34] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00045_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold328 (.A(\inv_result[33] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold329 (.A(\inv_result[187] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold330 (.A(\inv_result[217] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold331 (.A(\inv_result[64] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold332 (.A(\shift_reg[135] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00146_),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold334 (.A(\shift_reg[106] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold335 (.A(_00117_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold336 (.A(\shift_reg[194] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold337 (.A(_00205_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold338 (.A(\inv_result[183] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold339 (.A(\inv_result[203] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold340 (.A(\shift_reg[75] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold341 (.A(_00086_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold342 (.A(\shift_reg[107] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold343 (.A(_00118_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold344 (.A(\shift_reg[171] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold345 (.A(_00182_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold346 (.A(\shift_reg[70] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold347 (.A(\inv_result[159] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold348 (.A(\inv_result[180] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold349 (.A(\inv_result[175] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_inv.f_next[234] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold351 (.A(_01538_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold352 (.A(\shift_reg[134] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold353 (.A(_00145_),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold354 (.A(\inv_result[182] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold355 (.A(\shift_reg[122] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold356 (.A(_00133_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold357 (.A(\shift_reg[20] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold358 (.A(\shift_reg[49] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00060_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold360 (.A(\shift_reg[181] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold361 (.A(_00192_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold362 (.A(\shift_reg[205] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00216_),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold364 (.A(\inv_result[6] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold365 (.A(\inv_result[0] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold366 (.A(_01048_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold367 (.A(\shift_reg[36] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold368 (.A(_00047_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold369 (.A(\inv_result[148] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold370 (.A(\inv_result[71] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold371 (.A(_01119_),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold372 (.A(\inv_result[86] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold373 (.A(\shift_reg[167] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold374 (.A(_00178_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold375 (.A(\inv_result[112] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold376 (.A(\inv_result[253] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold377 (.A(\u_inv.f_next[244] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold378 (.A(_01548_),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold379 (.A(\shift_reg[169] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold380 (.A(_00180_),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold381 (.A(\shift_reg[217] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold382 (.A(\shift_reg[86] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold383 (.A(\inv_result[167] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold384 (.A(\shift_reg[8] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold385 (.A(_00019_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold386 (.A(\inv_result[162] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold387 (.A(_01210_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold388 (.A(\u_inv.d_reg[6] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold389 (.A(_06172_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold390 (.A(\inv_result[251] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold391 (.A(\inv_result[16] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold392 (.A(\inv_result[231] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold393 (.A(\inv_result[208] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold394 (.A(_01256_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold395 (.A(\inv_result[158] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold396 (.A(\inv_result[138] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold397 (.A(\shift_reg[76] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold398 (.A(_00087_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold399 (.A(\shift_reg[29] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00040_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold401 (.A(\u_inv.f_next[222] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold402 (.A(_01526_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold403 (.A(\shift_reg[82] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold404 (.A(_00093_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold405 (.A(\inv_result[188] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold406 (.A(\inv_result[194] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold407 (.A(\shift_reg[99] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00110_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold409 (.A(\shift_reg[84] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00095_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold411 (.A(\shift_reg[65] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold412 (.A(_00076_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold413 (.A(\u_inv.f_next[158] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold414 (.A(_01462_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold415 (.A(\shift_reg[77] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold416 (.A(_00088_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold417 (.A(\shift_reg[39] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold418 (.A(_00050_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold419 (.A(\shift_reg[92] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold420 (.A(_00103_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold421 (.A(\shift_reg[43] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold422 (.A(\inv_result[152] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold423 (.A(\shift_reg[66] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold424 (.A(_00077_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold425 (.A(\shift_reg[23] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold426 (.A(_00034_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold427 (.A(\shift_reg[145] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold428 (.A(_00156_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold429 (.A(\shift_reg[0] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold430 (.A(_01562_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold431 (.A(\inv_result[34] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold432 (.A(\shift_reg[211] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold433 (.A(_00222_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold434 (.A(\shift_reg[148] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold435 (.A(\inv_result[196] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold436 (.A(\shift_reg[173] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00184_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold438 (.A(\shift_reg[121] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold439 (.A(_00132_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold440 (.A(\inv_result[46] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold441 (.A(\shift_reg[176] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold442 (.A(_00187_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold443 (.A(\inv_result[81] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold444 (.A(\inv_result[151] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold445 (.A(\inv_result[207] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold446 (.A(\inv_result[57] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold447 (.A(\inv_result[45] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold448 (.A(\inv_result[92] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold449 (.A(\inv_result[111] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold450 (.A(\shift_reg[231] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold451 (.A(\shift_reg[188] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00199_),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold453 (.A(\inv_result[53] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold454 (.A(\inv_result[189] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold455 (.A(\shift_reg[141] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold456 (.A(\inv_result[11] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold457 (.A(\shift_reg[63] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold458 (.A(_00074_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold459 (.A(\u_inv.delta_reg[6] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold460 (.A(_01824_),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold461 (.A(\inv_result[90] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold462 (.A(\shift_reg[149] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold463 (.A(_00160_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold464 (.A(\inv_result[87] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_inv.f_next[112] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold466 (.A(_01416_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold467 (.A(\u_inv.input_reg[1] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold468 (.A(\shift_reg[126] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold469 (.A(_00137_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold470 (.A(\inv_result[226] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold471 (.A(wr_prev),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold472 (.A(_11054_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold473 (.A(\inv_result[186] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold474 (.A(\shift_reg[144] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold475 (.A(_00155_),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold476 (.A(\inv_result[94] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_inv.f_next[70] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold478 (.A(_01374_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold479 (.A(\shift_reg[53] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00064_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold481 (.A(\inv_result[178] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold482 (.A(\shift_reg[225] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold483 (.A(\shift_reg[157] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold484 (.A(_00168_),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold485 (.A(\inv_result[8] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold486 (.A(\inv_result[1] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold487 (.A(\shift_reg[242] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold488 (.A(_00253_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold489 (.A(\inv_result[95] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold490 (.A(\inv_result[22] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold491 (.A(\inv_result[142] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold492 (.A(\shift_reg[168] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold493 (.A(\shift_reg[129] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold494 (.A(_00140_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold495 (.A(\shift_reg[210] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_inv.f_next[124] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold497 (.A(_01428_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold498 (.A(\inv_result[15] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold499 (.A(\inv_result[211] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold500 (.A(\u_inv.counter[1] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold501 (.A(_00268_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold502 (.A(\shift_reg[246] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold503 (.A(_00257_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold504 (.A(\inv_result[144] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold505 (.A(\shift_reg[201] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold506 (.A(_00212_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold507 (.A(\inv_result[233] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold508 (.A(\shift_reg[73] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00084_),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold510 (.A(\shift_reg[58] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold511 (.A(_00069_),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold512 (.A(\inv_result[104] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold513 (.A(\inv_result[215] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold514 (.A(\inv_result[139] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold515 (.A(\inv_result[214] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold516 (.A(\inv_result[68] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold517 (.A(\shift_reg[64] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold518 (.A(\inv_result[84] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold519 (.A(\inv_result[110] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold520 (.A(\shift_reg[7] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold521 (.A(\inv_result[242] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold522 (.A(\shift_reg[27] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold523 (.A(_00038_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold524 (.A(\inv_result[206] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold525 (.A(\shift_reg[219] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold526 (.A(_00230_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold527 (.A(\shift_reg[60] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold528 (.A(_00071_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold529 (.A(\inv_result[116] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold530 (.A(\shift_reg[142] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold531 (.A(\shift_reg[10] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold532 (.A(_00021_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold533 (.A(\inv_result[36] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold534 (.A(\shift_reg[182] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00193_),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold536 (.A(\inv_result[220] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold537 (.A(\u_inv.delta_reg[0] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold538 (.A(\shift_reg[151] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold539 (.A(_00162_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold540 (.A(\shift_reg[222] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_inv.delta_reg[1] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold542 (.A(_01819_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold543 (.A(\inv_result[100] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold544 (.A(\shift_reg[130] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold545 (.A(_00141_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold546 (.A(\inv_result[235] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold547 (.A(\inv_result[248] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold548 (.A(\inv_result[38] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold549 (.A(\inv_result[135] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold550 (.A(\shift_reg[147] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold551 (.A(\inv_result[154] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold552 (.A(_01202_),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold553 (.A(\shift_reg[91] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold554 (.A(\shift_reg[180] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold555 (.A(_00191_),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold556 (.A(\shift_reg[212] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_inv.input_reg[18] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold558 (.A(_01580_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold559 (.A(\u_inv.input_reg[2] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold560 (.A(_01564_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold561 (.A(\inv_result[75] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold562 (.A(\inv_result[83] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_inv.f_next[236] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold564 (.A(_01540_),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold565 (.A(\u_inv.f_next[198] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold566 (.A(_01502_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold567 (.A(\shift_reg[113] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold568 (.A(_00124_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_inv.counter[2] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold570 (.A(_00269_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold571 (.A(\shift_reg[24] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold572 (.A(_00035_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold573 (.A(\shift_reg[116] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold574 (.A(\inv_result[96] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_inv.input_reg[95] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold576 (.A(_01657_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold577 (.A(\shift_reg[245] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00256_),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold579 (.A(\inv_result[73] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold580 (.A(\shift_reg[218] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold581 (.A(\inv_result[228] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold582 (.A(\shift_reg[155] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold583 (.A(_00166_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold584 (.A(\inv_result[13] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold585 (.A(\inv_result[18] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold586 (.A(\shift_reg[143] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold587 (.A(_00154_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold588 (.A(\shift_reg[57] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold589 (.A(\shift_reg[165] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00176_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold591 (.A(\inv_result[66] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold592 (.A(\inv_result[199] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold593 (.A(\inv_result[163] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold594 (.A(\inv_result[191] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold595 (.A(\shift_reg[154] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold596 (.A(_00165_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold597 (.A(\shift_reg[192] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold598 (.A(_00203_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold599 (.A(\u_inv.f_next[246] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold600 (.A(_01550_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_inv.input_reg[31] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold602 (.A(\inv_result[130] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold603 (.A(\inv_result[77] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold604 (.A(\inv_result[123] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold605 (.A(\inv_result[82] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold606 (.A(\inv_result[19] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold607 (.A(_01067_),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold608 (.A(\u_inv.input_reg[7] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold609 (.A(\inv_result[117] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold610 (.A(\inv_result[129] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold611 (.A(\shift_reg[158] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00169_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold613 (.A(\shift_reg[179] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold614 (.A(\inv_result[234] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold615 (.A(\inv_result[10] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold616 (.A(\shift_reg[95] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold617 (.A(\shift_reg[159] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold618 (.A(\u_inv.delta_reg[7] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold619 (.A(_10316_),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold620 (.A(\u_inv.input_reg[90] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_inv.input_reg[16] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold622 (.A(_01578_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold623 (.A(\shift_reg[228] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold624 (.A(_00239_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold625 (.A(\shift_reg[186] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold626 (.A(_00197_),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold627 (.A(\inv_result[209] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold628 (.A(\inv_result[4] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold629 (.A(_01052_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold630 (.A(\inv_result[101] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold631 (.A(\inv_result[67] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold632 (.A(\u_inv.input_reg[32] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold633 (.A(\u_inv.input_reg[34] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold634 (.A(\u_inv.f_next[214] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold635 (.A(_01518_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold636 (.A(\shift_reg[123] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold637 (.A(_00134_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold638 (.A(\inv_result[63] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold639 (.A(\inv_result[21] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold640 (.A(\shift_reg[163] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold641 (.A(\inv_result[127] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold642 (.A(\u_inv.f_next[197] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold643 (.A(_01501_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold644 (.A(\shift_reg[247] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold645 (.A(_00258_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold646 (.A(\u_inv.input_reg[78] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold647 (.A(\u_inv.f_next[220] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold648 (.A(_01524_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold649 (.A(\shift_reg[47] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold650 (.A(_00058_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold651 (.A(\inv_result[72] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold652 (.A(\shift_reg[187] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold653 (.A(\u_inv.input_reg[76] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_inv.input_reg[187] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold655 (.A(\u_inv.input_reg[33] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold656 (.A(\u_inv.input_reg[48] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold657 (.A(_01610_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold658 (.A(\u_inv.input_reg[46] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold659 (.A(_01608_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold660 (.A(\u_inv.input_reg[30] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold661 (.A(\u_inv.input_reg[250] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold662 (.A(\inv_result[88] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_inv.input_reg[57] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold664 (.A(\shift_reg[172] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold665 (.A(\shift_reg[174] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold666 (.A(\u_inv.f_next[140] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold667 (.A(_01444_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold668 (.A(\shift_reg[220] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold669 (.A(\shift_reg[96] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_inv.input_reg[238] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold671 (.A(\u_inv.input_reg[91] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold672 (.A(\inv_result[14] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold673 (.A(\inv_result[99] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold674 (.A(\shift_reg[104] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold675 (.A(\u_inv.input_reg[25] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold676 (.A(\inv_result[153] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold677 (.A(\inv_result[216] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold678 (.A(\u_inv.input_reg[126] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_inv.input_reg[65] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold680 (.A(\u_inv.input_reg[228] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold681 (.A(\inv_result[124] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold682 (.A(\u_inv.f_next[17] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold683 (.A(_01321_),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold684 (.A(\inv_result[125] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold685 (.A(\u_inv.input_reg[29] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold686 (.A(\u_inv.f_next[156] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold687 (.A(_01460_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold688 (.A(\u_inv.input_reg[54] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold689 (.A(\u_inv.input_reg[137] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold690 (.A(_01699_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold691 (.A(\shift_reg[137] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_inv.f_next[24] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold693 (.A(_01328_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold694 (.A(\u_inv.input_reg[251] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold695 (.A(\inv_result[98] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold696 (.A(\u_inv.input_reg[26] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold697 (.A(\inv_result[156] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold698 (.A(\inv_result[76] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_inv.f_next[99] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold700 (.A(_01403_),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold701 (.A(\shift_reg[195] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold702 (.A(\u_inv.input_reg[61] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold703 (.A(_01623_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold704 (.A(\shift_reg[100] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_inv.input_reg[40] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold706 (.A(\inv_result[89] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold707 (.A(_01137_),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold708 (.A(\u_inv.f_next[196] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold709 (.A(_01500_),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold710 (.A(\u_inv.f_next[162] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold711 (.A(_01466_),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold712 (.A(\shift_reg[119] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00130_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold714 (.A(\shift_reg[110] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold715 (.A(_00121_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold716 (.A(\inv_result[47] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold717 (.A(\u_inv.input_reg[49] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold718 (.A(\u_inv.input_reg[53] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_inv.input_reg[206] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold720 (.A(_01768_),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold721 (.A(\u_inv.input_reg[246] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_inv.input_reg[28] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold723 (.A(\u_inv.input_reg[15] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold724 (.A(_01577_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold725 (.A(\u_inv.input_reg[136] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_inv.input_reg[244] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold727 (.A(_01806_),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold728 (.A(\u_inv.input_reg[185] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold729 (.A(_01747_),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold730 (.A(\u_inv.input_reg[219] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_inv.input_reg[113] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold732 (.A(\inv_result[60] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold733 (.A(\u_inv.input_reg[35] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_inv.input_reg[215] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold735 (.A(\u_inv.input_reg[209] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold736 (.A(\u_inv.input_reg[64] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold737 (.A(\u_inv.f_next[94] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold738 (.A(_01398_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold739 (.A(\u_inv.input_reg[58] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold740 (.A(\u_inv.input_reg[37] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold741 (.A(\u_inv.input_reg[47] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold742 (.A(\shift_reg[48] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold743 (.A(\shift_reg[206] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold744 (.A(_00217_),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold745 (.A(\u_inv.input_reg[220] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold746 (.A(\shift_reg[200] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold747 (.A(\shift_reg[178] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold748 (.A(\u_inv.input_reg[201] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold749 (.A(\u_inv.input_reg[14] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold750 (.A(_01576_),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold751 (.A(\u_inv.input_reg[66] ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold752 (.A(\u_inv.input_reg[38] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold753 (.A(\u_inv.input_reg[9] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold754 (.A(\inv_result[219] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold755 (.A(\u_inv.input_reg[130] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold756 (.A(\u_inv.input_reg[163] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold757 (.A(\u_inv.input_reg[153] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold758 (.A(_01715_),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold759 (.A(\inv_result[79] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold760 (.A(_01127_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold761 (.A(\u_inv.input_reg[207] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold762 (.A(\u_inv.input_reg[218] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold763 (.A(\u_inv.input_reg[222] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold764 (.A(\u_inv.f_next[242] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold765 (.A(_01546_),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold766 (.A(\u_inv.input_reg[236] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold767 (.A(\shift_reg[3] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold768 (.A(_00014_),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold769 (.A(\u_inv.input_reg[156] ),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold770 (.A(_01718_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold771 (.A(\u_inv.input_reg[197] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold772 (.A(_01759_),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold773 (.A(\u_inv.input_reg[224] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold774 (.A(_01786_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold775 (.A(\u_inv.input_reg[27] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold776 (.A(\u_inv.input_reg[50] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold777 (.A(\u_inv.input_reg[198] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold778 (.A(_01760_),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold779 (.A(\shift_reg[189] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold780 (.A(\shift_reg[46] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold781 (.A(\shift_reg[190] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold782 (.A(\u_inv.input_reg[189] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold783 (.A(\u_inv.input_reg[17] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold784 (.A(_01579_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold785 (.A(\u_inv.input_reg[79] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold786 (.A(\u_inv.input_reg[171] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold787 (.A(\u_inv.input_reg[242] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold788 (.A(\shift_reg[2] ),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold789 (.A(\u_inv.input_reg[168] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold790 (.A(\u_inv.input_reg[245] ),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold791 (.A(\u_inv.input_reg[129] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold792 (.A(\shift_reg[196] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold793 (.A(\u_inv.input_reg[19] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold794 (.A(_01581_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold795 (.A(\u_inv.counter[4] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold796 (.A(\u_inv.input_reg[83] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold797 (.A(\shift_reg[198] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold798 (.A(\u_inv.input_reg[42] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold799 (.A(\u_inv.input_reg[87] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold800 (.A(\u_inv.input_reg[12] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold801 (.A(\u_inv.input_reg[43] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold802 (.A(\shift_reg[109] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold803 (.A(_00120_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold804 (.A(\u_inv.input_reg[210] ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold805 (.A(\u_inv.f_reg[222] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold806 (.A(\u_inv.input_reg[188] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold807 (.A(\shift_reg[146] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold808 (.A(\u_inv.d_next[249] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold809 (.A(\shift_reg[19] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold810 (.A(\u_inv.input_reg[51] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold811 (.A(\u_inv.delta_reg[8] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold812 (.A(_01826_),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold813 (.A(\u_inv.input_reg[13] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold814 (.A(\u_inv.input_reg[101] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold815 (.A(_01663_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold816 (.A(\u_inv.f_next[129] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold817 (.A(_01433_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold818 (.A(\shift_reg[14] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold819 (.A(\inv_result[173] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold820 (.A(\u_inv.input_reg[165] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold821 (.A(\inv_result[26] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold822 (.A(\u_inv.input_reg[225] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold823 (.A(\u_inv.input_reg[167] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold824 (.A(\u_inv.input_reg[89] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold825 (.A(\u_inv.input_reg[161] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold826 (.A(\u_inv.input_reg[108] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold827 (.A(\shift_reg[120] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00131_),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold829 (.A(\u_inv.input_reg[184] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold830 (.A(_01746_),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold831 (.A(\inv_result[3] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold832 (.A(\u_inv.input_reg[116] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold833 (.A(\u_inv.input_reg[77] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold834 (.A(\u_inv.input_reg[164] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold835 (.A(\u_inv.input_reg[233] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold836 (.A(\u_inv.input_reg[175] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold837 (.A(\shift_reg[98] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold838 (.A(\u_inv.f_reg[86] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold839 (.A(_00877_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold840 (.A(\u_inv.input_reg[41] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold841 (.A(\u_inv.f_reg[70] ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold842 (.A(\u_inv.input_reg[123] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold843 (.A(\u_inv.f_next[41] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold844 (.A(_01345_),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold845 (.A(\shift_reg[101] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold846 (.A(\u_inv.f_next[163] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold847 (.A(_01467_),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold848 (.A(\shift_reg[224] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold849 (.A(\u_inv.input_reg[204] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold850 (.A(\u_inv.input_reg[23] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold851 (.A(\u_inv.input_reg[200] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold852 (.A(\inv_result[120] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold853 (.A(\u_inv.input_reg[199] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold854 (.A(_01761_),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold855 (.A(\shift_reg[150] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold856 (.A(\inv_result[143] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold857 (.A(\u_inv.input_reg[60] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold858 (.A(\u_inv.input_reg[92] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold859 (.A(\inv_result[103] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold860 (.A(\shift_reg[115] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold861 (.A(\u_inv.input_reg[75] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold862 (.A(\u_inv.f_reg[158] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold863 (.A(\u_inv.input_reg[144] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold864 (.A(\u_inv.f_reg[162] ),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold865 (.A(\shift_reg[226] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold866 (.A(\u_inv.input_reg[145] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold867 (.A(\u_inv.input_reg[98] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold868 (.A(\u_inv.input_reg[186] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold869 (.A(\inv_result[155] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold870 (.A(\u_inv.input_reg[243] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold871 (.A(_01805_),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold872 (.A(\u_inv.input_reg[133] ),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold873 (.A(\inv_result[223] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold874 (.A(\inv_result[250] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold875 (.A(\u_inv.input_reg[22] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold876 (.A(\u_inv.input_reg[134] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold877 (.A(\u_inv.input_reg[143] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold878 (.A(\u_inv.input_reg[36] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold879 (.A(\u_inv.f_reg[186] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold880 (.A(_00977_),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold881 (.A(\u_inv.input_reg[205] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold882 (.A(\inv_result[105] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold883 (.A(\shift_reg[153] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold884 (.A(\u_inv.input_reg[249] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold885 (.A(\u_inv.input_reg[160] ),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold886 (.A(\u_inv.input_reg[252] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold887 (.A(\u_inv.d_next[69] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold888 (.A(_05504_),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold889 (.A(\u_inv.input_reg[106] ),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold890 (.A(\u_inv.input_reg[253] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold891 (.A(\u_inv.input_reg[180] ),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold892 (.A(\inv_result[97] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold893 (.A(\u_inv.input_reg[73] ),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold894 (.A(\u_inv.f_reg[159] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold895 (.A(_00950_),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold896 (.A(\u_inv.input_reg[140] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold897 (.A(\u_inv.f_next[202] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold898 (.A(_01506_),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold899 (.A(\shift_reg[118] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold900 (.A(\u_inv.input_reg[21] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold901 (.A(\u_inv.input_reg[11] ),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold902 (.A(\inv_result[108] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold903 (.A(\u_inv.input_reg[247] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold904 (.A(\u_inv.input_reg[211] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold905 (.A(\u_inv.f_next[237] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold906 (.A(_01541_),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold907 (.A(\u_inv.f_next[62] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold908 (.A(_01366_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold909 (.A(\u_inv.f_reg[234] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold910 (.A(\u_inv.input_reg[162] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold911 (.A(\u_inv.input_reg[234] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold912 (.A(\u_inv.input_reg[80] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold913 (.A(\u_inv.input_reg[169] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold914 (.A(\u_inv.f_reg[102] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold915 (.A(_00893_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold916 (.A(\u_inv.input_reg[45] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold917 (.A(_01607_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold918 (.A(\u_inv.input_reg[100] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold919 (.A(\u_inv.input_reg[147] ),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold920 (.A(\u_inv.input_reg[190] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold921 (.A(\u_inv.input_reg[68] ),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold922 (.A(\u_inv.f_reg[2] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold923 (.A(_00793_),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold924 (.A(\shift_reg[125] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold925 (.A(\u_inv.input_reg[203] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold926 (.A(\u_inv.input_reg[217] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold927 (.A(\u_inv.input_reg[151] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold928 (.A(\u_inv.input_reg[196] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold929 (.A(\shift_reg[102] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold930 (.A(\u_inv.f_next[201] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold931 (.A(\u_inv.input_reg[39] ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold932 (.A(\inv_result[55] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold933 (.A(\u_inv.input_reg[176] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold934 (.A(\shift_reg[244] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold935 (.A(\u_inv.d_next[80] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold936 (.A(\u_inv.input_reg[105] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold937 (.A(\u_inv.input_reg[10] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold938 (.A(\u_inv.input_reg[166] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold939 (.A(\inv_result[201] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold940 (.A(\u_inv.f_reg[166] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold941 (.A(_00957_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold942 (.A(\u_inv.input_reg[240] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold943 (.A(_01802_),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold944 (.A(\u_inv.input_reg[178] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold945 (.A(\inv_result[232] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold946 (.A(\u_inv.input_reg[132] ),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold947 (.A(\u_inv.input_reg[24] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold948 (.A(\u_inv.input_reg[254] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold949 (.A(\byte_cnt[2] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold950 (.A(_00007_),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold951 (.A(\u_inv.d_next[221] ),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold952 (.A(_05656_),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold953 (.A(\u_inv.input_reg[44] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold954 (.A(\u_inv.input_reg[150] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold955 (.A(\inv_result[145] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold956 (.A(\u_inv.f_next[101] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold957 (.A(_01405_),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold958 (.A(\u_inv.input_reg[128] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold959 (.A(\u_inv.f_next[166] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold960 (.A(_01470_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold961 (.A(\u_inv.input_reg[179] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold962 (.A(\u_inv.f_reg[244] ),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold963 (.A(\u_inv.input_reg[85] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold964 (.A(\u_inv.input_reg[139] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold965 (.A(\u_inv.input_reg[72] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold966 (.A(\u_inv.d_next[16] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold967 (.A(\inv_result[78] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold968 (.A(\u_inv.d_next[126] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold969 (.A(\u_inv.input_reg[114] ),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold970 (.A(\inv_result[240] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01288_),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold972 (.A(\u_inv.f_reg[118] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold973 (.A(_00909_),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold974 (.A(\inv_result[236] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold975 (.A(\u_inv.input_reg[255] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold976 (.A(\shift_reg[17] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold977 (.A(_00028_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold978 (.A(\u_inv.input_reg[216] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold979 (.A(\u_inv.input_reg[202] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold980 (.A(\u_inv.input_reg[67] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold981 (.A(\inv_result[30] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold982 (.A(\u_inv.f_next[176] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold983 (.A(_01480_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold984 (.A(\u_inv.input_reg[59] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold985 (.A(\u_inv.f_reg[19] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold986 (.A(_00810_),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold987 (.A(\u_inv.f_next[224] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold988 (.A(\inv_result[29] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold989 (.A(\u_inv.f_next[65] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold990 (.A(_01369_),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold991 (.A(\u_inv.input_reg[208] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold992 (.A(\u_inv.input_reg[131] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold993 (.A(\inv_result[239] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold994 (.A(\u_inv.input_reg[172] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold995 (.A(\shift_reg[197] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold996 (.A(_00208_),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold997 (.A(\u_inv.input_reg[8] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold998 (.A(\u_inv.f_next[68] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold999 (.A(_01372_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\u_inv.input_reg[135] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\inv_result[17] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\u_inv.d_next[50] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\u_inv.input_reg[20] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\u_inv.d_next[10] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\u_inv.f_next[72] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1006 (.A(_01376_),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\inv_result[238] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\inv_result[5] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\u_inv.input_reg[94] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\state[1] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\u_inv.f_next[144] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_01448_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\u_inv.input_reg[102] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\u_inv.input_reg[181] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\u_inv.f_next[36] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold1016 (.A(_01340_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\u_inv.input_reg[125] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\inv_result[176] ),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\u_inv.input_reg[221] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_01783_),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\u_inv.f_next[169] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_01473_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\u_inv.input_reg[107] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\u_inv.f_next[98] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\inv_result[122] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\u_inv.d_next[241] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\inv_result[12] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\u_inv.f_reg[236] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\u_inv.f_reg[33] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_00824_),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\u_inv.input_reg[226] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\u_inv.d_next[60] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\inv_result[31] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\u_inv.input_reg[235] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\u_inv.f_next[132] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_01436_),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\u_inv.input_reg[81] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\u_inv.f_next[110] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold1039 (.A(_01414_),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\u_inv.f_reg[126] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold1041 (.A(_00917_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\u_inv.input_reg[56] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\u_inv.input_reg[124] ),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\inv_result[246] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_01294_),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\shift_reg[221] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\u_inv.f_next[218] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_01522_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\u_inv.input_reg[70] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\u_inv.d_next[56] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\u_inv.input_reg[223] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\u_inv.input_reg[63] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\u_inv.f_reg[214] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\inv_result[255] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\u_inv.input_reg[109] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\u_inv.input_reg[69] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\u_inv.counter[5] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold1058 (.A(_13587_),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\u_inv.input_reg[191] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\u_inv.f_next[5] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold1061 (.A(_00796_),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\u_inv.f_next[215] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_01519_),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\u_inv.input_reg[241] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\u_inv.d_next[244] ),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\u_inv.input_reg[212] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\u_inv.f_next[189] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_01493_),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\u_inv.input_reg[214] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\shift_reg[185] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\u_inv.d_next[168] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\u_inv.d_next[19] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\u_inv.input_reg[148] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\shift_reg[45] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\inv_result[247] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\shift_reg[18] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\u_inv.d_next[96] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\u_inv.f_next[161] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\u_inv.f_reg[81] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00872_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\u_inv.f_next[6] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_05693_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\u_inv.f_reg[238] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_01029_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\u_inv.f_next[64] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\u_inv.f_next[111] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_00902_),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\u_inv.d_next[144] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\u_inv.f_next[184] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold1090 (.A(_01488_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\u_inv.f_reg[38] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_00829_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\u_inv.d_next[4] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\u_inv.f_next[40] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\u_inv.input_reg[99] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\u_inv.f_reg[136] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_00927_),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\u_inv.input_reg[237] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\shift_reg[111] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1100 (.A(_00122_),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\shift_reg[240] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\u_inv.f_next[122] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_01426_),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\shift_reg[243] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\u_inv.f_reg[138] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_00929_),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\u_inv.f_reg[94] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\u_inv.d_next[6] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\u_inv.f_next[125] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1110 (.A(_00916_),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\u_inv.input_reg[173] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\inv_result[24] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\u_inv.f_next[185] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_01489_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\u_inv.f_next[207] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_01511_),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\u_inv.input_reg[117] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\u_inv.input_reg[248] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\u_inv.f_next[243] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\u_inv.input_reg[86] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\shift_reg[103] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\u_inv.input_reg[55] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\u_inv.input_reg[232] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\u_inv.f_next[3] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1125 (.A(_00794_),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\u_inv.f_next[188] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\u_inv.input_reg[183] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\inv_result[58] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\u_inv.f_next[175] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1130 (.A(_01479_),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\u_inv.f_next[233] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\u_inv.d_next[236] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\u_inv.f_next[216] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01520_),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\u_inv.f_next[245] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\u_inv.d_next[92] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\u_inv.f_reg[58] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_00849_),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\u_inv.input_reg[195] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\u_inv.f_next[173] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_00964_),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\u_inv.input_reg[88] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\u_inv.input_reg[239] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\u_inv.f_next[210] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1145 (.A(_01514_),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\inv_result[181] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_01229_),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\u_inv.d_next[94] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\u_inv.f_reg[202] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\u_inv.f_next[229] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_01533_),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\inv_result[41] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\u_inv.d_next[48] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\u_inv.input_reg[158] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\u_inv.f_next[66] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00857_),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\u_inv.f_reg[122] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\u_inv.input_reg[213] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1159 (.A(inv_done),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_00001_),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\u_inv.f_next[116] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_00907_),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\u_inv.input_reg[141] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\u_inv.f_reg[246] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\u_inv.f_reg[22] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1166 (.A(_00813_),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\inv_result[28] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\u_inv.d_next[240] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\u_inv.f_next[177] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1170 (.A(_01481_),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\inv_result[49] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\u_inv.f_next[50] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1173 (.A(_01354_),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\u_inv.f_next[219] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\u_inv.d_next[108] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\u_inv.input_reg[192] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\u_inv.input_reg[157] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\u_inv.counter[6] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\u_inv.d_next[81] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\u_inv.f_next[192] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_01496_),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\u_inv.f_next[252] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_01556_),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\inv_result[39] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\u_inv.f_reg[178] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1186 (.A(_00969_),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\inv_result[252] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\u_inv.f_next[21] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_00812_),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\u_inv.input_reg[120] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\inv_result[50] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\u_inv.f_reg[204] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00995_),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\u_inv.f_next[164] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_01468_),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\u_inv.f_next[217] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\u_inv.f_reg[44] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_00835_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\u_inv.f_reg[49] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_00840_),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\u_inv.d_next[101] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_05536_),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\u_inv.input_reg[71] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\u_inv.f_next[225] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1205 (.A(_01529_),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\u_inv.input_reg[84] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\u_inv.d_next[164] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_05599_),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\u_inv.f_next[78] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_00869_),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\u_inv.d_next[185] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_05620_),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\u_inv.d_next[245] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_05680_),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\u_inv.f_next[221] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\u_inv.f_reg[144] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\u_inv.f_reg[65] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\u_inv.f_next[32] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_01336_),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\u_inv.f_reg[132] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\shift_reg[16] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\inv_result[254] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\u_inv.f_reg[40] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\u_inv.input_reg[115] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\u_inv.f_reg[172] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_00963_),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\u_inv.input_reg[103] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\u_inv.f_next[18] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_00809_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\u_inv.d_next[107] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\u_inv.f_reg[50] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\u_inv.input_reg[229] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\u_inv.f_reg[15] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1234 (.A(_00806_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\u_inv.d_next[189] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_05624_),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\u_inv.input_reg[122] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\inv_result[119] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\u_inv.f_reg[156] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\u_inv.f_reg[76] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_00867_),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\u_inv.input_reg[52] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\u_inv.input_reg[193] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\u_inv.f_next[42] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_01346_),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\u_inv.f_next[73] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1247 (.A(_01377_),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\shift_reg[15] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\u_inv.d_next[159] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1250 (.A(_05594_),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\u_inv.f_next[55] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00846_),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\u_inv.d_next[73] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\u_inv.f_next[190] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\u_inv.f_next[71] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1256 (.A(_00862_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\u_inv.input_reg[138] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\u_inv.f_reg[212] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_01003_),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\u_inv.f_reg[252] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\u_inv.input_reg[127] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\u_inv.f_reg[98] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\u_inv.f_reg[190] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\u_inv.f_reg[32] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\u_inv.input_reg[231] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\u_inv.f_next[103] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_01407_),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\inv_result[169] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\u_inv.d_reg[10] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\u_inv.f_next[137] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1271 (.A(_01441_),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\u_inv.f_next[152] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_00943_),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\u_inv.f_next[247] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1275 (.A(_01551_),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\u_inv.f_next[223] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_01014_),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\u_inv.f_next[253] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_01044_),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\u_inv.d_next[173] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_05608_),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\u_inv.d_next[116] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\inv_result[245] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_01293_),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\u_inv.f_next[235] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1286 (.A(_01026_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\u_inv.f_next[67] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00858_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\u_inv.d_next[89] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_05524_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\u_inv.f_next[92] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_01396_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\u_inv.f_reg[60] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1294 (.A(_00851_),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\inv_result[51] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\u_inv.f_reg[194] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_00985_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\u_inv.d_reg[92] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\u_inv.f_reg[226] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_01017_),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\shift_reg[61] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\u_inv.d_next[151] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_05586_),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\u_inv.f_next[183] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\shift_reg[184] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\u_inv.input_reg[177] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\u_inv.d_reg[126] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\u_inv.f_reg[210] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\inv_result[27] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\u_inv.f_reg[106] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_00897_),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\u_inv.d_next[70] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\u_inv.f_next[81] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_01385_),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\u_inv.f_reg[88] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_00879_),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\u_inv.f_reg[242] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\u_inv.f_next[95] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_00886_),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\u_inv.f_next[82] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1321 (.A(_00873_),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\u_inv.d_reg[249] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\u_inv.input_reg[93] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\u_inv.f_reg[120] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00911_),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\u_inv.d_next[248] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_05683_),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\u_inv.d_next[237] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_05672_),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\u_inv.d_next[181] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_05616_),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\u_inv.f_next[9] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold1333 (.A(_01313_),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\u_inv.f_reg[137] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\u_inv.f_reg[73] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\u_inv.input_reg[96] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\u_inv.f_next[2] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\u_inv.f_next[133] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_01437_),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\u_inv.f_next[52] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_01356_),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\u_inv.f_next[114] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_00905_),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\u_inv.f_next[141] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold1345 (.A(_00932_),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\u_inv.input_reg[110] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\u_inv.f_reg[92] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\u_inv.f_reg[198] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\u_inv.f_next[154] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_00945_),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\u_inv.d_next[223] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\u_inv.f_reg[108] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_00899_),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\inv_result[25] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\u_inv.f_reg[225] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\inv_result[121] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\u_inv.f_next[143] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\u_inv.f_next[121] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_00912_),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\u_inv.d_reg[58] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_05493_),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\u_inv.f_reg[4] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_05692_),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\u_inv.input_reg[170] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\u_inv.f_reg[250] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1366 (.A(_01041_),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\u_inv.f_next[172] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\u_inv.f_next[23] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1369 (.A(_00814_),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\shift_reg[199] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\u_inv.input_reg[149] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\u_inv.f_reg[160] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_00951_),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\u_inv.d_next[174] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_05609_),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\u_inv.f_reg[201] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\shift_reg[152] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\u_inv.f_next[195] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_00986_),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\shift_reg[156] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\u_inv.input_reg[104] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\u_inv.f_reg[219] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\u_inv.d_next[106] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\u_inv.f_reg[216] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\u_inv.d_next[52] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\u_inv.input_reg[230] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\u_inv.d_next[224] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1388 (.A(_05659_),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\u_inv.input_reg[119] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\u_inv.d_next[255] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\u_inv.input_reg[62] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\u_inv.d_next[194] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_05629_),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\u_inv.f_reg[46] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1395 (.A(_00837_),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\u_inv.d_next[55] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1397 (.A(_05490_),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\u_inv.d_next[158] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\u_inv.input_reg[174] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\u_inv.input_reg[194] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\u_inv.input_reg[142] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\u_inv.f_reg[196] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\u_inv.d_next[25] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\u_inv.f_reg[42] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\u_inv.delta_reg[3] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1406 (.A(_10299_),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\u_inv.f_reg[119] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1408 (.A(_00910_),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\u_inv.f_reg[179] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_00970_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\u_inv.f_reg[61] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1412 (.A(_00852_),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\u_inv.f_reg[185] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\u_inv.d_reg[144] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\u_inv.f_next[213] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1416 (.A(_01004_),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\u_inv.d_next[0] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1418 (.A(_05435_),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\inv_result[107] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\u_inv.f_next[208] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_00999_),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\u_inv.f_reg[215] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\u_inv.f_next[48] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_00839_),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\u_inv.f_reg[129] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\u_inv.input_reg[152] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\u_inv.d_next[127] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1428 (.A(_05562_),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\inv_result[177] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\u_inv.d_next[11] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_05446_),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\u_inv.input_reg[227] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\u_inv.f_reg[217] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\u_inv.input_reg[74] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\u_inv.f_next[180] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1436 (.A(_00971_),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\u_inv.f_next[96] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1438 (.A(_00887_),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\u_inv.d_next[152] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\u_inv.f_reg[37] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_00828_),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\u_inv.f_next[167] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_00958_),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\inv_result[161] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\u_inv.d_next[182] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_05617_),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\u_inv.f_next[200] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\u_inv.d_reg[56] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\u_inv.d_next[12] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1450 (.A(_05447_),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\u_inv.f_next[39] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_00830_),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\u_inv.d_next[229] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\u_inv.d_next[8] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\u_inv.f_reg[28] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1456 (.A(_00819_),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\u_inv.d_next[232] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_05667_),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\u_inv.f_reg[90] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_00881_),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\u_inv.f_reg[224] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\u_inv.d_next[67] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1463 (.A(_05502_),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\u_inv.f_next[109] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_00900_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\u_inv.f_next[12] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1467 (.A(_01316_),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\u_inv.f_next[255] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1469 (.A(_01559_),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\u_inv.f_reg[84] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1471 (.A(_00875_),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\u_inv.input_reg[146] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\u_inv.f_next[254] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1474 (.A(_01045_),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\u_inv.d_reg[48] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\u_inv.d_next[202] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_05637_),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\u_inv.d_next[114] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\u_inv.input_reg[97] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\u_inv.f_next[138] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_01442_),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\u_inv.f_reg[220] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\u_inv.f_next[127] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_00918_),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\u_inv.d_next[7] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_05442_),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\u_inv.f_next[209] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\u_inv.input_reg[155] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\u_inv.f_reg[54] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_00845_),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\u_inv.f_reg[72] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\u_inv.f_next[69] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1493 (.A(_00860_),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\inv_result[149] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\u_inv.input_reg[112] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\u_inv.d_next[1] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_05436_),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\u_inv.f_next[255] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\u_inv.f_next[128] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\u_inv.f_reg[7] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_05694_),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\u_inv.d_reg[168] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\u_inv.d_next[136] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\u_inv.f_reg[200] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\u_inv.d_next[143] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\u_inv.f_next[79] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1507 (.A(_00870_),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\u_inv.d_next[256] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\u_inv.f_next[74] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1510 (.A(_00865_),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\u_inv.f_reg[13] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_00804_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\u_inv.f_reg[191] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1514 (.A(_00982_),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\inv_result[197] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\u_inv.f_reg[30] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_00821_),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\u_inv.d_next[128] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1519 (.A(_05563_),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\u_inv.d_reg[80] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\u_inv.f_reg[1] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_00792_),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\u_inv.f_next[107] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_00898_),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\u_inv.f_reg[20] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_00811_),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\u_inv.f_reg[99] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\u_inv.f_reg[128] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\u_inv.f_reg[175] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\u_inv.f_reg[124] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\u_inv.f_next[45] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1532 (.A(_00836_),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\u_inv.f_reg[104] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_00895_),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\u_inv.input_reg[82] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\u_inv.d_next[118] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\u_inv.d_reg[94] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\u_inv.delta_reg[4] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\u_inv.f_next[10] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_00801_),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\u_inv.f_reg[174] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_00965_),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\u_inv.d_next[28] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_05463_),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\u_inv.d_next[65] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_05500_),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\inv_result[165] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\u_inv.f_next[38] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1549 (.A(_01342_),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\u_inv.d_next[99] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\u_inv.f_reg[8] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_05695_),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\u_inv.d_next[84] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\u_inv.f_next[181] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1555 (.A(_00972_),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\u_inv.f_next[134] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_01438_),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\u_inv.f_reg[112] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\u_inv.input_reg[111] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\u_inv.f_next[20] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\u_inv.d_next[210] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_05645_),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\u_inv.d_next[51] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_05486_),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\u_inv.d_next[192] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_05627_),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\u_inv.f_reg[143] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\u_inv.f_next[174] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\u_inv.d_next[93] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_05528_),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\u_inv.f_reg[184] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\u_inv.f_reg[41] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\u_inv.d_next[177] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\u_inv.f_reg[17] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\u_inv.d_next[253] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_05688_),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\u_inv.f_reg[59] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_00850_),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\u_inv.d_next[142] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1580 (.A(_05577_),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\u_inv.f_next[22] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\u_inv.d_next[235] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_05670_),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\u_inv.f_reg[197] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\u_inv.d_next[61] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1586 (.A(_05496_),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\u_inv.d_next[29] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1588 (.A(_05464_),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\u_inv.input_reg[182] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\u_inv.d_reg[70] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\u_inv.f_reg[245] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\u_inv.input_reg[118] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\u_inv.f_next[59] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_01363_),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\u_inv.d_next[203] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_05638_),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\u_inv.d_reg[152] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\u_inv.f_reg[64] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\u_inv.f_next[113] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\u_inv.d_next[83] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_05518_),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\u_inv.f_next[206] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\u_inv.d_next[62] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1604 (.A(_05497_),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\u_inv.input_reg[121] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\inv_result[69] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\u_inv.d_next[238] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_05673_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\u_inv.f_next[179] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\u_inv.d_next[186] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_05621_),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\u_inv.d_next[176] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1613 (.A(_05611_),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\u_inv.f_reg[218] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\u_inv.f_reg[199] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_00990_),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\u_inv.f_reg[26] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_00817_),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\u_inv.f_reg[232] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_01023_),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\u_inv.f_reg[145] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1622 (.A(_00936_),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\u_inv.d_next[160] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\u_inv.f_reg[97] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_00888_),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\u_inv.f_reg[237] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\u_inv.f_next[56] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1628 (.A(_01360_),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\u_inv.f_reg[101] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\u_inv.d_reg[244] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\u_inv.d_reg[24] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1632 (.A(_05459_),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\u_inv.d_next[85] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\u_inv.f_next[240] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1635 (.A(_01544_),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\u_inv.input_reg[154] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\u_inv.d_reg[240] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\u_inv.f_next[226] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1639 (.A(_01530_),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\u_inv.f_next[51] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\u_inv.d_next[213] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1642 (.A(_05648_),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\u_inv.f_next[7] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1644 (.A(_01311_),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\u_inv.f_reg[68] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\u_inv.d_next[90] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\u_inv.f_reg[177] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\u_inv.f_reg[34] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1649 (.A(_00825_),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\u_inv.f_next[31] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1651 (.A(_00822_),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\u_inv.d_next[254] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\u_inv.f_reg[163] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\u_inv.d_next[76] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\u_inv.f_next[61] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\u_inv.f_reg[16] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1657 (.A(_00807_),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\u_inv.f_next[131] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\u_inv.d_next[198] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\u_inv.f_next[25] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1661 (.A(_01329_),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\u_inv.d_next[98] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1663 (.A(_05533_),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\u_inv.f_reg[176] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\u_inv.d_next[13] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1666 (.A(_05448_),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\u_inv.f_reg[24] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\u_inv.d_next[207] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1669 (.A(_05642_),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\u_inv.d_next[91] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1671 (.A(_05526_),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\u_inv.d_reg[150] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1673 (.A(_05585_),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\u_inv.f_reg[113] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\u_inv.d_reg[108] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\u_inv.f_next[145] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1677 (.A(_01449_),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\u_inv.d_reg[177] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\u_inv.f_reg[87] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_00878_),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\u_inv.d_next[252] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1682 (.A(_05687_),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\u_inv.d_next[193] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1684 (.A(_05628_),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\u_inv.d_next[154] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_05589_),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\u_inv.f_reg[233] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\u_inv.f_reg[170] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_00961_),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\u_inv.d_next[227] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_05662_),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\u_inv.f_reg[51] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\u_inv.f_reg[52] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\u_inv.d_next[121] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1695 (.A(_05556_),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\u_inv.d_next[242] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_05677_),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\u_inv.d_reg[241] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\u_inv.d_reg[16] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\u_inv.d_next[195] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1701 (.A(_05630_),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\u_inv.f_next[239] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1703 (.A(_01030_),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\u_inv.d_next[196] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\u_inv.f_next[119] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_01423_),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\u_inv.f_next[77] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00868_),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\u_inv.f_next[193] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1710 (.A(_00984_),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\u_inv.d_next[214] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1712 (.A(_05649_),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\u_inv.d_reg[81] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\u_inv.d_next[250] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1715 (.A(_05685_),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\u_inv.f_next[108] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\u_inv.f_reg[110] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\u_inv.d_next[27] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1719 (.A(_05462_),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\u_inv.d_next[97] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_05532_),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\u_inv.f_next[171] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_00962_),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\u_inv.f_reg[9] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\u_inv.d_next[71] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1726 (.A(_05506_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\u_inv.d_next[218] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1728 (.A(_05653_),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\u_inv.f_next[182] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\u_inv.f_next[149] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1731 (.A(_00940_),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\u_inv.d_next[167] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1733 (.A(_05602_),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\u_inv.d_next[104] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\u_inv.d_next[3] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1736 (.A(_05438_),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\u_inv.f_next[142] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\u_inv.d_reg[236] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\u_inv.f_next[35] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1740 (.A(_00826_),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\u_inv.d_reg[60] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\u_inv.d_next[209] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1743 (.A(_05644_),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\u_inv.d_next[105] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1745 (.A(_05540_),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\inv_result[157] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\u_inv.f_next[204] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\u_inv.d_next[220] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1749 (.A(_05655_),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\u_inv.f_next[19] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\u_inv.f_reg[130] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_00921_),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\u_inv.d_next[87] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\u_inv.d_next[5] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1755 (.A(_05440_),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\u_inv.f_next[168] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\u_inv.f_next[87] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1758 (.A(_01391_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\u_inv.f_next[126] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\u_inv.d_next[228] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\u_inv.d_next[188] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1762 (.A(_05623_),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\u_inv.d_next[132] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1764 (.A(_05567_),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\u_inv.f_reg[155] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1766 (.A(_00946_),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\u_inv.d_next[78] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1768 (.A(_05513_),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\u_inv.f_next[46] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\u_inv.f_next[211] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_01002_),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\u_inv.d_next[103] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1773 (.A(_05538_),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\u_inv.state[1] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\u_inv.d_next[148] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1776 (.A(_05583_),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\u_inv.f_reg[209] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\u_inv.d_next[22] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\u_inv.delta_reg[2] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\u_inv.f_next[93] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1781 (.A(_00884_),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\u_inv.d_next[35] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1783 (.A(_05470_),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\u_inv.d_next[175] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1785 (.A(_05610_),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\u_inv.d_next[79] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1787 (.A(_05514_),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\u_inv.d_next[243] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1789 (.A(_05678_),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\u_inv.d_next[140] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_05575_),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\u_inv.f_next[165] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\u_inv.d_next[161] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1794 (.A(_05596_),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\u_inv.f_next[53] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1796 (.A(_01357_),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\u_inv.d_reg[96] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\u_inv.f_reg[142] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\u_inv.f_reg[229] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\u_inv.d_next[82] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1801 (.A(_05517_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\u_inv.d_next[33] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\u_inv.f_next[89] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1804 (.A(_00880_),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\u_inv.d_reg[19] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\u_inv.f_next[135] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1807 (.A(_01439_),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\u_inv.d_next[153] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_05588_),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\u_inv.d_reg[106] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\u_inv.d_next[170] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_05605_),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\u_inv.d_reg[107] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\u_inv.d_next[112] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1815 (.A(_05547_),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\u_inv.f_next[153] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\u_inv.d_reg[50] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\u_inv.f_reg[247] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\u_inv.d_next[146] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1820 (.A(_05581_),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\state[0] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\u_inv.f_next[123] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_00914_),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\u_inv.f_reg[243] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\u_inv.f_reg[100] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_00891_),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\u_inv.d_next[34] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\u_inv.f_next[248] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1829 (.A(_01552_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\u_inv.d_reg[254] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\u_inv.d_next[178] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1832 (.A(_05613_),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\u_inv.d_next[225] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\u_inv.f_next[34] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\u_inv.d_next[200] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\inv_result[113] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\u_inv.d_next[141] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1838 (.A(_05576_),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\u_inv.d_next[9] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1840 (.A(_05444_),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\u_inv.f_reg[248] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\u_inv.d_reg[229] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\u_inv.d_next[204] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\u_inv.d_next[169] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1845 (.A(_05604_),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\u_inv.d_next[183] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\u_inv.d_next[133] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1848 (.A(_05568_),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\u_inv.d_next[20] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1850 (.A(_05455_),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\u_inv.d_next[211] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1852 (.A(_05646_),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\u_inv.f_reg[133] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\u_inv.f_reg[182] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\u_inv.d_next[113] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\u_inv.d_next[233] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1857 (.A(_05668_),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\u_inv.f_reg[47] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1859 (.A(_00838_),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\u_inv.d_next[37] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1861 (.A(_05472_),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\u_inv.d_next[134] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1863 (.A(_05569_),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\u_inv.d_next[119] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1865 (.A(_05554_),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\u_inv.f_reg[183] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\u_inv.d_next[215] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1868 (.A(_05650_),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\u_inv.d_next[217] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1870 (.A(_05652_),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\u_inv.f_next[4] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\u_inv.d_next[129] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\u_inv.d_next[165] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1874 (.A(_05600_),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\u_inv.f_next[37] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\u_inv.d_next[219] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1877 (.A(_05654_),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\u_inv.f_next[91] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\u_inv.f_reg[62] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\u_inv.f_reg[91] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\u_inv.f_next[205] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_00996_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\u_inv.d_next[14] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1884 (.A(_05449_),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\u_inv.f_next[232] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\u_inv.d_next[66] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1887 (.A(_05501_),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\u_inv.f_reg[168] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\u_inv.d_reg[155] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1890 (.A(_05590_),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\u_inv.delta_reg[5] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1892 (.A(_10306_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\u_inv.d_next[124] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1894 (.A(_05559_),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\u_inv.d_next[38] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1896 (.A(_05473_),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\u_inv.d_next[145] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_05580_),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\u_inv.f_next[23] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\u_inv.d_next[208] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1901 (.A(_05643_),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\u_inv.f_reg[230] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1903 (.A(_01021_),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\u_inv.d_next[155] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\u_inv.d_next[216] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1906 (.A(_05651_),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\u_inv.f_reg[36] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\u_inv.d_next[41] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1909 (.A(_05476_),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\u_inv.d_next[149] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1911 (.A(_05584_),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\u_inv.f_reg[25] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\u_inv.f_reg[134] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\u_inv.d_next[111] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1915 (.A(_05546_),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\u_inv.d_reg[129] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\u_inv.f_next[75] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1918 (.A(_00866_),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\u_inv.d_reg[84] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\u_inv.d_reg[4] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\u_inv.f_next[212] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\u_inv.f_next[187] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\u_inv.f_reg[105] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1924 (.A(_00896_),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\u_inv.d_next[172] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1926 (.A(_05607_),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\u_inv.f_next[117] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1928 (.A(_01421_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\u_inv.d_next[57] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1930 (.A(_05492_),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\u_inv.d_next[199] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1932 (.A(_05634_),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\u_inv.f_reg[188] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\u_inv.f_reg[255] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\u_inv.f_next[115] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\u_inv.d_next[201] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1937 (.A(_05636_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\u_inv.d_reg[116] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\u_inv.d_next[206] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1940 (.A(_05641_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\u_inv.f_reg[221] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\u_inv.d_reg[225] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\u_inv.f_next[194] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\u_inv.f_reg[189] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\u_inv.d_next[190] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1946 (.A(_05625_),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\u_inv.d_next[226] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1948 (.A(_05661_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\u_inv.f_reg[56] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\u_inv.f_reg[192] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\u_inv.f_next[44] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1952 (.A(_01348_),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\u_inv.f_next[49] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\u_inv.d_reg[104] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\u_inv.d_reg[183] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\u_inv.f_next[147] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1957 (.A(_00938_),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\u_inv.d_next[75] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_05510_),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\u_inv.d_reg[255] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\u_inv.d_next[45] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1962 (.A(_05480_),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\u_inv.f_next[8] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\u_inv.d_next[54] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1965 (.A(_05489_),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\u_inv.f_next[157] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1967 (.A(_00948_),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\u_inv.d_next[2] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\u_inv.d_next[162] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\u_inv.d_next[231] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1971 (.A(_05666_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\u_inv.d_reg[256] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\u_inv.d_next[234] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1974 (.A(_05669_),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\u_inv.f_next[76] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\u_inv.d_next[49] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1977 (.A(_05484_),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\u_inv.d_reg[85] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\u_inv.d_reg[223] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\u_inv.f_next[151] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1981 (.A(_00942_),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\u_inv.f_next[11] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\u_inv.d_next[239] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\u_inv.d_reg[160] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\u_inv.d_next[180] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1986 (.A(_05615_),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\u_inv.d_reg[52] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\u_inv.f_reg[207] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\u_inv.d_next[230] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1990 (.A(_05665_),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\u_inv.d_reg[8] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\u_inv.f_reg[53] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\u_inv.d_reg[143] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\u_inv.d_next[251] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_05686_),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\u_inv.d_next[72] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\u_inv.d_reg[204] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\u_inv.d_next[120] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1999 (.A(_05555_),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\u_inv.d_reg[25] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\u_inv.f_reg[115] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\u_inv.f_next[15] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold2003 (.A(_01319_),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\u_inv.d_next[100] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold2005 (.A(_05535_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\u_inv.d_next[102] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold2007 (.A(_05537_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\u_inv.d_reg[72] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\u_inv.f_next[80] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold2010 (.A(_00871_),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\u_inv.d_next[246] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold2012 (.A(_05681_),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\u_inv.f_reg[251] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold2014 (.A(_01042_),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\u_inv.f_reg[150] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold2016 (.A(_00941_),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\u_inv.d_next[53] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold2018 (.A(_05488_),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\u_inv.d_next[117] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold2020 (.A(_05552_),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\u_inv.f_next[100] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\u_inv.f_next[83] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\u_inv.d_next[21] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold2024 (.A(_05456_),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\u_inv.d_reg[198] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\u_inv.f_reg[14] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold2027 (.A(_00805_),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\u_inv.d_next[135] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\u_inv.f_reg[249] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold2030 (.A(_01040_),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\u_inv.f_next[150] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\u_inv.d_next[42] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold2033 (.A(_05477_),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\u_inv.d_reg[2] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\u_inv.d_reg[99] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\u_inv.d_next[88] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\u_inv.f_reg[74] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\u_inv.f_reg[146] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold2039 (.A(_00937_),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\u_inv.f_reg[153] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\u_inv.f_reg[135] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\u_inv.d_next[32] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_05467_),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\u_inv.d_next[157] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold2045 (.A(_05592_),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\u_inv.d_reg[200] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\u_inv.f_reg[117] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\u_inv.f_reg[103] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\u_inv.f_next[90] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\u_inv.d_next[212] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_05647_),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\u_inv.d_next[63] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\u_inv.d_next[24] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\u_inv.f_reg[187] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\u_inv.d_next[40] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold2056 (.A(_05475_),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\u_inv.f_next[29] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold2058 (.A(_01333_),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\u_inv.f_reg[12] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\u_inv.d_next[36] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold2061 (.A(_05471_),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\u_inv.f_next[60] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold2063 (.A(_01364_),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\u_inv.d_next[125] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\u_inv.d_reg[73] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\u_inv.f_reg[169] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\u_inv.f_reg[63] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold2068 (.A(_00854_),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\u_inv.d_next[247] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold2070 (.A(_05682_),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\u_inv.f_next[27] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_00818_),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\u_inv.f_next[47] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\u_inv.d_reg[158] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\u_inv.f_next[170] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\u_inv.d_next[187] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold2077 (.A(_05622_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\u_inv.f_next[118] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\u_inv.f_next[139] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold2080 (.A(_00930_),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\u_inv.d_next[26] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold2082 (.A(_05461_),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\u_inv.f_reg[140] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\u_inv.d_next[44] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_05479_),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\u_inv.d_next[130] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\u_inv.d_reg[135] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\u_inv.d_next[68] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold2089 (.A(_05503_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\u_inv.d_next[150] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\u_inv.f_next[84] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold2092 (.A(_01388_),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\u_inv.d_reg[239] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\u_inv.f_next[85] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_00876_),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\u_inv.d_next[166] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold2097 (.A(_05601_),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\u_inv.delta_reg[9] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\u_inv.d_reg[87] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\u_inv.f_next[104] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_01408_),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\u_inv.d_next[171] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold2103 (.A(_05606_),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\u_inv.d_reg[136] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\u_inv.d_next[191] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\u_inv.d_next[39] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\u_inv.f_next[54] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\inv_result[249] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\u_inv.f_next[249] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold2110 (.A(_01553_),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\u_inv.d_reg[90] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\u_inv.d_next[86] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold2113 (.A(_05521_),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\u_inv.d_reg[191] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\u_inv.f_reg[240] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\u_inv.f_next[57] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold2117 (.A(_00848_),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\u_inv.f_next[250] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold2119 (.A(_01554_),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\u_inv.d_next[46] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\u_inv.f_reg[131] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\u_inv.f_reg[241] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold2123 (.A(_01032_),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\u_inv.f_reg[83] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\u_inv.f_reg[161] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\u_inv.d_reg[228] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\u_inv.f_next[16] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\u_inv.d_next[156] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\u_inv.d_next[18] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold2130 (.A(_05453_),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\u_inv.f_reg[227] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold2132 (.A(_01018_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\u_inv.d_reg[125] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\u_inv.d_reg[114] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\u_inv.d_next[147] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\u_inv.d_reg[76] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\u_inv.f_next[155] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\u_inv.f_reg[29] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\u_inv.d_next[115] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold2140 (.A(_05550_),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\u_inv.d_reg[34] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\u_inv.f_next[97] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\u_inv.d_next[197] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold2144 (.A(_05632_),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\u_inv.d_next[139] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold2146 (.A(_05574_),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\u_inv.f_next[28] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold2148 (.A(\u_inv.d_reg[63] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\u_inv.d_next[74] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold2150 (.A(_05509_),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\u_inv.d_reg[31] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold2152 (.A(_05466_),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\u_inv.d_next[15] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\u_inv.d_next[179] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\u_inv.d_next[110] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold2156 (.A(_05545_),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\u_inv.d_next[59] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold2158 (.A(_05494_),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\u_inv.f_next[102] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\u_inv.d_reg[22] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\u_inv.d_reg[23] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold2162 (.A(_05458_),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\u_inv.d_next[47] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold2164 (.A(_05482_),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\u_inv.f_next[86] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\u_inv.f_next[33] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\u_inv.d_next[58] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\u_inv.d_next[122] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold2169 (.A(_05557_),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\u_inv.f_next[238] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\u_inv.input_reg[0] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\u_inv.d_reg[179] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\u_inv.d_next[123] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold2174 (.A(_05558_),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\u_inv.d_reg[46] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\u_inv.d_reg[118] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\u_inv.d_reg[196] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\u_inv.d_next[222] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\u_inv.d_next[64] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\u_inv.f_next[148] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\u_inv.d_reg[15] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\u_inv.d_next[205] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\u_inv.f_next[88] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\u_inv.f_next[26] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\u_inv.d_reg[64] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\u_inv.f_next[58] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\u_inv.f_next[231] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold2188 (.A(_01022_),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\u_inv.f_reg[165] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\u_inv.d_reg[222] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\u_inv.f_reg[43] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold2192 (.A(_00834_),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\u_inv.d_next[163] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold2194 (.A(_05598_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\u_inv.input_reg[6] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\u_inv.d_next[23] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\u_inv.f_reg[203] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold2198 (.A(_00994_),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\u_inv.f_reg[11] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\u_inv.d_reg[147] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\u_inv.f_next[230] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold2202 (.A(_01534_),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\u_inv.f_next[186] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\u_inv.d_reg[33] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\u_inv.d_next[77] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_05512_),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\u_inv.d_reg[88] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\u_inv.f_reg[206] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\u_inv.f_next[160] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold2210 (.A(_01464_),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\u_inv.d_next[43] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\u_inv.d_next[131] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold2213 (.A(_05566_),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\u_inv.f_next[191] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\u_inv.f_next[228] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold2216 (.A(_01019_),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\u_inv.f_next[130] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\u_inv.f_reg[164] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\u_inv.d_next[30] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\u_inv.f_next[251] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\u_inv.f_next[136] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\u_inv.f_next[106] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold2223 (.A(_01410_),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\u_inv.d_reg[205] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\u_inv.d_reg[30] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\u_inv.d_reg[43] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\u_inv.d_reg[113] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\u_inv.f_next[1] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\u_inv.d_next[138] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\u_inv.d_next[137] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\u_inv.d_next[109] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\u_inv.d_reg[109] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\u_inv.f_next[178] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\u_inv.f_reg[148] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\u_inv.f_next[14] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold2236 (.A(inv_done),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\u_inv.f_next[120] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\u_inv.d_reg[156] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\u_inv.f_next[63] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\u_inv.d_reg[39] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\u_inv.d_next[31] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\u_inv.f_next[199] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\u_inv.f_next[146] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\u_inv.f_next[43] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\u_inv.d_reg[138] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\u_inv.f_next[30] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\u_inv.f_next[241] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\u_inv.d_reg[137] ),
    .X(net4952));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\u_inv.f_next[203] ),
    .X(net4953));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\u_inv.f_next[227] ),
    .X(net4954));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\u_inv.d_next[95] ),
    .X(net4955));
 sg13g2_dlygate4sd3_1 hold2252 (.A(_05530_),
    .X(net4956));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\u_inv.f_next[105] ),
    .X(net4957));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\u_inv.f_next[13] ),
    .X(net4958));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\u_inv.f_next[256] ),
    .X(net4959));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\u_inv.d_next[17] ),
    .X(net4960));
 sg13g2_dlygate4sd3_1 hold2257 (.A(_05452_),
    .X(net4961));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\u_inv.d_reg[130] ),
    .X(net4962));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\u_inv.d_reg[162] ),
    .X(net4963));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\u_inv.input_valid ),
    .X(net4964));
 sg13g2_dlygate4sd3_1 hold2261 (.A(_11045_),
    .X(net4965));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\state[0] ),
    .X(net4966));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\u_inv.f_next[225] ),
    .X(net4967));
 sg13g2_antennanp ANTENNA_1 (.A(rst_n));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_fill_2 FILLER_0_714 ();
 sg13g2_fill_1 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_8 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_0_1032 ();
 sg13g2_decap_8 FILLER_0_1039 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_8 FILLER_0_1053 ();
 sg13g2_decap_8 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1067 ();
 sg13g2_decap_8 FILLER_0_1074 ();
 sg13g2_decap_8 FILLER_0_1081 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_8 FILLER_0_1095 ();
 sg13g2_decap_8 FILLER_0_1102 ();
 sg13g2_decap_8 FILLER_0_1109 ();
 sg13g2_decap_8 FILLER_0_1116 ();
 sg13g2_decap_8 FILLER_0_1123 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1158 ();
 sg13g2_decap_8 FILLER_0_1165 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_8 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1186 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_fill_2 FILLER_0_1235 ();
 sg13g2_fill_1 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1245 ();
 sg13g2_fill_1 FILLER_0_1252 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_8 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1290 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_decap_8 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_0_1332 ();
 sg13g2_decap_8 FILLER_0_1339 ();
 sg13g2_decap_8 FILLER_0_1346 ();
 sg13g2_decap_8 FILLER_0_1353 ();
 sg13g2_decap_8 FILLER_0_1360 ();
 sg13g2_decap_8 FILLER_0_1367 ();
 sg13g2_decap_8 FILLER_0_1374 ();
 sg13g2_decap_8 FILLER_0_1381 ();
 sg13g2_decap_8 FILLER_0_1388 ();
 sg13g2_decap_8 FILLER_0_1395 ();
 sg13g2_decap_8 FILLER_0_1402 ();
 sg13g2_decap_8 FILLER_0_1409 ();
 sg13g2_decap_8 FILLER_0_1416 ();
 sg13g2_decap_8 FILLER_0_1423 ();
 sg13g2_decap_8 FILLER_0_1430 ();
 sg13g2_decap_8 FILLER_0_1437 ();
 sg13g2_decap_8 FILLER_0_1444 ();
 sg13g2_decap_8 FILLER_0_1451 ();
 sg13g2_decap_8 FILLER_0_1458 ();
 sg13g2_decap_8 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1472 ();
 sg13g2_decap_8 FILLER_0_1479 ();
 sg13g2_decap_8 FILLER_0_1486 ();
 sg13g2_decap_8 FILLER_0_1493 ();
 sg13g2_decap_8 FILLER_0_1500 ();
 sg13g2_decap_8 FILLER_0_1507 ();
 sg13g2_decap_8 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_8 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_decap_8 FILLER_0_1563 ();
 sg13g2_decap_8 FILLER_0_1570 ();
 sg13g2_decap_8 FILLER_0_1577 ();
 sg13g2_decap_8 FILLER_0_1584 ();
 sg13g2_decap_8 FILLER_0_1591 ();
 sg13g2_decap_8 FILLER_0_1598 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_4 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1658 ();
 sg13g2_decap_8 FILLER_0_1665 ();
 sg13g2_decap_8 FILLER_0_1672 ();
 sg13g2_fill_2 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1688 ();
 sg13g2_decap_8 FILLER_0_1695 ();
 sg13g2_decap_8 FILLER_0_1702 ();
 sg13g2_decap_4 FILLER_0_1709 ();
 sg13g2_fill_2 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1718 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1739 ();
 sg13g2_decap_8 FILLER_0_1746 ();
 sg13g2_decap_8 FILLER_0_1753 ();
 sg13g2_decap_8 FILLER_0_1760 ();
 sg13g2_decap_8 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_0_1774 ();
 sg13g2_decap_8 FILLER_0_1781 ();
 sg13g2_decap_8 FILLER_0_1788 ();
 sg13g2_decap_8 FILLER_0_1795 ();
 sg13g2_decap_8 FILLER_0_1802 ();
 sg13g2_decap_8 FILLER_0_1809 ();
 sg13g2_decap_8 FILLER_0_1816 ();
 sg13g2_decap_4 FILLER_0_1823 ();
 sg13g2_fill_1 FILLER_0_1827 ();
 sg13g2_decap_8 FILLER_0_1832 ();
 sg13g2_decap_4 FILLER_0_1839 ();
 sg13g2_fill_1 FILLER_0_1843 ();
 sg13g2_decap_4 FILLER_0_1871 ();
 sg13g2_fill_2 FILLER_0_1875 ();
 sg13g2_decap_8 FILLER_0_1881 ();
 sg13g2_decap_8 FILLER_0_1888 ();
 sg13g2_decap_8 FILLER_0_1895 ();
 sg13g2_fill_2 FILLER_0_1902 ();
 sg13g2_fill_1 FILLER_0_1904 ();
 sg13g2_decap_4 FILLER_0_1936 ();
 sg13g2_fill_1 FILLER_0_1940 ();
 sg13g2_fill_1 FILLER_0_1946 ();
 sg13g2_fill_2 FILLER_0_1957 ();
 sg13g2_decap_8 FILLER_0_1970 ();
 sg13g2_fill_1 FILLER_0_1977 ();
 sg13g2_fill_1 FILLER_0_1985 ();
 sg13g2_fill_2 FILLER_0_2014 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_fill_2 FILLER_0_2058 ();
 sg13g2_fill_1 FILLER_0_2060 ();
 sg13g2_decap_8 FILLER_0_2089 ();
 sg13g2_decap_8 FILLER_0_2096 ();
 sg13g2_decap_8 FILLER_0_2103 ();
 sg13g2_decap_8 FILLER_0_2110 ();
 sg13g2_decap_8 FILLER_0_2117 ();
 sg13g2_decap_8 FILLER_0_2124 ();
 sg13g2_decap_4 FILLER_0_2131 ();
 sg13g2_fill_1 FILLER_0_2135 ();
 sg13g2_decap_8 FILLER_0_2164 ();
 sg13g2_decap_8 FILLER_0_2171 ();
 sg13g2_decap_8 FILLER_0_2178 ();
 sg13g2_decap_8 FILLER_0_2185 ();
 sg13g2_decap_8 FILLER_0_2192 ();
 sg13g2_decap_8 FILLER_0_2199 ();
 sg13g2_decap_8 FILLER_0_2206 ();
 sg13g2_decap_8 FILLER_0_2213 ();
 sg13g2_decap_8 FILLER_0_2220 ();
 sg13g2_decap_8 FILLER_0_2227 ();
 sg13g2_decap_8 FILLER_0_2234 ();
 sg13g2_decap_8 FILLER_0_2241 ();
 sg13g2_decap_8 FILLER_0_2248 ();
 sg13g2_decap_8 FILLER_0_2255 ();
 sg13g2_decap_8 FILLER_0_2262 ();
 sg13g2_decap_8 FILLER_0_2269 ();
 sg13g2_decap_8 FILLER_0_2276 ();
 sg13g2_decap_8 FILLER_0_2283 ();
 sg13g2_decap_8 FILLER_0_2290 ();
 sg13g2_decap_8 FILLER_0_2297 ();
 sg13g2_decap_8 FILLER_0_2304 ();
 sg13g2_decap_8 FILLER_0_2311 ();
 sg13g2_decap_8 FILLER_0_2318 ();
 sg13g2_decap_8 FILLER_0_2325 ();
 sg13g2_decap_8 FILLER_0_2332 ();
 sg13g2_decap_8 FILLER_0_2339 ();
 sg13g2_decap_8 FILLER_0_2346 ();
 sg13g2_decap_8 FILLER_0_2353 ();
 sg13g2_decap_8 FILLER_0_2360 ();
 sg13g2_decap_8 FILLER_0_2367 ();
 sg13g2_decap_8 FILLER_0_2374 ();
 sg13g2_decap_8 FILLER_0_2381 ();
 sg13g2_decap_8 FILLER_0_2388 ();
 sg13g2_decap_8 FILLER_0_2395 ();
 sg13g2_decap_8 FILLER_0_2402 ();
 sg13g2_fill_2 FILLER_0_2409 ();
 sg13g2_fill_1 FILLER_0_2411 ();
 sg13g2_fill_2 FILLER_0_2440 ();
 sg13g2_decap_4 FILLER_0_2449 ();
 sg13g2_fill_1 FILLER_0_2453 ();
 sg13g2_decap_8 FILLER_0_2458 ();
 sg13g2_decap_8 FILLER_0_2465 ();
 sg13g2_decap_8 FILLER_0_2472 ();
 sg13g2_decap_8 FILLER_0_2479 ();
 sg13g2_decap_8 FILLER_0_2486 ();
 sg13g2_decap_8 FILLER_0_2493 ();
 sg13g2_decap_8 FILLER_0_2500 ();
 sg13g2_decap_4 FILLER_0_2507 ();
 sg13g2_decap_8 FILLER_0_2531 ();
 sg13g2_decap_8 FILLER_0_2538 ();
 sg13g2_fill_2 FILLER_0_2545 ();
 sg13g2_fill_2 FILLER_0_2552 ();
 sg13g2_decap_8 FILLER_0_2564 ();
 sg13g2_decap_8 FILLER_0_2578 ();
 sg13g2_fill_1 FILLER_0_2585 ();
 sg13g2_fill_1 FILLER_0_2592 ();
 sg13g2_fill_1 FILLER_0_2596 ();
 sg13g2_fill_1 FILLER_0_2600 ();
 sg13g2_decap_8 FILLER_0_2629 ();
 sg13g2_decap_8 FILLER_0_2636 ();
 sg13g2_fill_2 FILLER_0_2643 ();
 sg13g2_fill_1 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_decap_8 FILLER_0_2667 ();
 sg13g2_decap_8 FILLER_0_2674 ();
 sg13g2_decap_8 FILLER_0_2681 ();
 sg13g2_decap_8 FILLER_0_2688 ();
 sg13g2_decap_8 FILLER_0_2695 ();
 sg13g2_decap_8 FILLER_0_2702 ();
 sg13g2_decap_8 FILLER_0_2709 ();
 sg13g2_decap_8 FILLER_0_2716 ();
 sg13g2_decap_8 FILLER_0_2723 ();
 sg13g2_decap_8 FILLER_0_2730 ();
 sg13g2_decap_8 FILLER_0_2737 ();
 sg13g2_decap_8 FILLER_0_2744 ();
 sg13g2_decap_8 FILLER_0_2751 ();
 sg13g2_decap_8 FILLER_0_2758 ();
 sg13g2_decap_8 FILLER_0_2765 ();
 sg13g2_decap_8 FILLER_0_2772 ();
 sg13g2_decap_8 FILLER_0_2779 ();
 sg13g2_decap_8 FILLER_0_2786 ();
 sg13g2_decap_8 FILLER_0_2793 ();
 sg13g2_decap_8 FILLER_0_2800 ();
 sg13g2_decap_8 FILLER_0_2807 ();
 sg13g2_fill_2 FILLER_0_2814 ();
 sg13g2_decap_8 FILLER_0_2820 ();
 sg13g2_decap_8 FILLER_0_2827 ();
 sg13g2_decap_8 FILLER_0_2834 ();
 sg13g2_fill_1 FILLER_0_2841 ();
 sg13g2_decap_8 FILLER_0_2849 ();
 sg13g2_decap_4 FILLER_0_2856 ();
 sg13g2_decap_4 FILLER_0_2888 ();
 sg13g2_fill_2 FILLER_0_2892 ();
 sg13g2_decap_8 FILLER_0_2898 ();
 sg13g2_decap_8 FILLER_0_2905 ();
 sg13g2_decap_8 FILLER_0_2912 ();
 sg13g2_decap_8 FILLER_0_2919 ();
 sg13g2_fill_2 FILLER_0_2926 ();
 sg13g2_decap_8 FILLER_0_2935 ();
 sg13g2_decap_8 FILLER_0_2942 ();
 sg13g2_decap_8 FILLER_0_2949 ();
 sg13g2_decap_8 FILLER_0_2956 ();
 sg13g2_decap_8 FILLER_0_2963 ();
 sg13g2_decap_8 FILLER_0_2970 ();
 sg13g2_decap_8 FILLER_0_2977 ();
 sg13g2_decap_8 FILLER_0_2984 ();
 sg13g2_decap_8 FILLER_0_2991 ();
 sg13g2_decap_8 FILLER_0_2998 ();
 sg13g2_decap_8 FILLER_0_3005 ();
 sg13g2_decap_8 FILLER_0_3012 ();
 sg13g2_decap_8 FILLER_0_3019 ();
 sg13g2_decap_8 FILLER_0_3026 ();
 sg13g2_decap_8 FILLER_0_3033 ();
 sg13g2_decap_8 FILLER_0_3040 ();
 sg13g2_decap_8 FILLER_0_3047 ();
 sg13g2_decap_8 FILLER_0_3054 ();
 sg13g2_decap_8 FILLER_0_3061 ();
 sg13g2_decap_8 FILLER_0_3068 ();
 sg13g2_decap_8 FILLER_0_3075 ();
 sg13g2_decap_8 FILLER_0_3082 ();
 sg13g2_decap_8 FILLER_0_3089 ();
 sg13g2_decap_8 FILLER_0_3096 ();
 sg13g2_decap_8 FILLER_0_3103 ();
 sg13g2_decap_8 FILLER_0_3110 ();
 sg13g2_decap_8 FILLER_0_3117 ();
 sg13g2_decap_8 FILLER_0_3124 ();
 sg13g2_decap_8 FILLER_0_3131 ();
 sg13g2_decap_8 FILLER_0_3138 ();
 sg13g2_decap_8 FILLER_0_3145 ();
 sg13g2_decap_8 FILLER_0_3152 ();
 sg13g2_decap_8 FILLER_0_3159 ();
 sg13g2_decap_8 FILLER_0_3166 ();
 sg13g2_decap_8 FILLER_0_3173 ();
 sg13g2_decap_8 FILLER_0_3180 ();
 sg13g2_decap_8 FILLER_0_3187 ();
 sg13g2_decap_8 FILLER_0_3194 ();
 sg13g2_decap_8 FILLER_0_3201 ();
 sg13g2_decap_8 FILLER_0_3208 ();
 sg13g2_decap_8 FILLER_0_3215 ();
 sg13g2_decap_8 FILLER_0_3222 ();
 sg13g2_decap_8 FILLER_0_3229 ();
 sg13g2_decap_8 FILLER_0_3236 ();
 sg13g2_decap_8 FILLER_0_3243 ();
 sg13g2_decap_8 FILLER_0_3250 ();
 sg13g2_decap_8 FILLER_0_3257 ();
 sg13g2_decap_8 FILLER_0_3264 ();
 sg13g2_decap_8 FILLER_0_3271 ();
 sg13g2_decap_8 FILLER_0_3278 ();
 sg13g2_decap_8 FILLER_0_3285 ();
 sg13g2_decap_8 FILLER_0_3292 ();
 sg13g2_decap_8 FILLER_0_3299 ();
 sg13g2_decap_8 FILLER_0_3306 ();
 sg13g2_decap_8 FILLER_0_3313 ();
 sg13g2_decap_8 FILLER_0_3320 ();
 sg13g2_decap_8 FILLER_0_3327 ();
 sg13g2_decap_8 FILLER_0_3334 ();
 sg13g2_decap_8 FILLER_0_3341 ();
 sg13g2_decap_8 FILLER_0_3348 ();
 sg13g2_decap_8 FILLER_0_3355 ();
 sg13g2_decap_8 FILLER_0_3362 ();
 sg13g2_decap_8 FILLER_0_3369 ();
 sg13g2_decap_8 FILLER_0_3376 ();
 sg13g2_decap_8 FILLER_0_3383 ();
 sg13g2_decap_8 FILLER_0_3390 ();
 sg13g2_decap_8 FILLER_0_3397 ();
 sg13g2_decap_8 FILLER_0_3404 ();
 sg13g2_decap_8 FILLER_0_3411 ();
 sg13g2_decap_8 FILLER_0_3418 ();
 sg13g2_decap_8 FILLER_0_3425 ();
 sg13g2_decap_8 FILLER_0_3432 ();
 sg13g2_decap_8 FILLER_0_3439 ();
 sg13g2_decap_8 FILLER_0_3446 ();
 sg13g2_decap_8 FILLER_0_3453 ();
 sg13g2_decap_8 FILLER_0_3460 ();
 sg13g2_decap_8 FILLER_0_3467 ();
 sg13g2_decap_8 FILLER_0_3474 ();
 sg13g2_decap_8 FILLER_0_3481 ();
 sg13g2_decap_8 FILLER_0_3488 ();
 sg13g2_decap_8 FILLER_0_3495 ();
 sg13g2_decap_8 FILLER_0_3502 ();
 sg13g2_decap_8 FILLER_0_3509 ();
 sg13g2_decap_8 FILLER_0_3516 ();
 sg13g2_decap_8 FILLER_0_3523 ();
 sg13g2_decap_8 FILLER_0_3530 ();
 sg13g2_decap_8 FILLER_0_3537 ();
 sg13g2_decap_8 FILLER_0_3544 ();
 sg13g2_decap_8 FILLER_0_3551 ();
 sg13g2_decap_8 FILLER_0_3558 ();
 sg13g2_decap_8 FILLER_0_3565 ();
 sg13g2_decap_8 FILLER_0_3572 ();
 sg13g2_fill_1 FILLER_0_3579 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_fill_2 FILLER_1_623 ();
 sg13g2_fill_1 FILLER_1_625 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_692 ();
 sg13g2_decap_8 FILLER_1_699 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_8 FILLER_1_720 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_fill_2 FILLER_1_734 ();
 sg13g2_fill_1 FILLER_1_736 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_fill_2 FILLER_1_772 ();
 sg13g2_fill_1 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_780 ();
 sg13g2_decap_8 FILLER_1_787 ();
 sg13g2_decap_8 FILLER_1_794 ();
 sg13g2_decap_4 FILLER_1_801 ();
 sg13g2_fill_2 FILLER_1_805 ();
 sg13g2_decap_4 FILLER_1_812 ();
 sg13g2_fill_2 FILLER_1_816 ();
 sg13g2_fill_2 FILLER_1_822 ();
 sg13g2_fill_1 FILLER_1_824 ();
 sg13g2_decap_8 FILLER_1_834 ();
 sg13g2_decap_8 FILLER_1_841 ();
 sg13g2_decap_8 FILLER_1_848 ();
 sg13g2_decap_8 FILLER_1_855 ();
 sg13g2_decap_8 FILLER_1_862 ();
 sg13g2_decap_8 FILLER_1_869 ();
 sg13g2_decap_8 FILLER_1_876 ();
 sg13g2_decap_8 FILLER_1_883 ();
 sg13g2_decap_8 FILLER_1_890 ();
 sg13g2_decap_8 FILLER_1_897 ();
 sg13g2_decap_8 FILLER_1_904 ();
 sg13g2_decap_8 FILLER_1_911 ();
 sg13g2_decap_8 FILLER_1_918 ();
 sg13g2_decap_8 FILLER_1_925 ();
 sg13g2_decap_8 FILLER_1_932 ();
 sg13g2_decap_8 FILLER_1_939 ();
 sg13g2_decap_8 FILLER_1_946 ();
 sg13g2_decap_8 FILLER_1_953 ();
 sg13g2_decap_8 FILLER_1_960 ();
 sg13g2_decap_8 FILLER_1_967 ();
 sg13g2_decap_8 FILLER_1_974 ();
 sg13g2_decap_8 FILLER_1_981 ();
 sg13g2_decap_8 FILLER_1_988 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1002 ();
 sg13g2_decap_8 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1016 ();
 sg13g2_decap_8 FILLER_1_1023 ();
 sg13g2_decap_8 FILLER_1_1030 ();
 sg13g2_decap_8 FILLER_1_1037 ();
 sg13g2_decap_8 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1051 ();
 sg13g2_decap_8 FILLER_1_1058 ();
 sg13g2_decap_8 FILLER_1_1065 ();
 sg13g2_decap_8 FILLER_1_1072 ();
 sg13g2_decap_8 FILLER_1_1079 ();
 sg13g2_decap_8 FILLER_1_1086 ();
 sg13g2_decap_8 FILLER_1_1093 ();
 sg13g2_decap_8 FILLER_1_1100 ();
 sg13g2_decap_8 FILLER_1_1107 ();
 sg13g2_decap_8 FILLER_1_1114 ();
 sg13g2_decap_8 FILLER_1_1121 ();
 sg13g2_decap_8 FILLER_1_1128 ();
 sg13g2_decap_8 FILLER_1_1135 ();
 sg13g2_decap_8 FILLER_1_1142 ();
 sg13g2_decap_8 FILLER_1_1149 ();
 sg13g2_decap_8 FILLER_1_1156 ();
 sg13g2_decap_8 FILLER_1_1163 ();
 sg13g2_decap_8 FILLER_1_1170 ();
 sg13g2_decap_8 FILLER_1_1177 ();
 sg13g2_decap_8 FILLER_1_1184 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1198 ();
 sg13g2_fill_2 FILLER_1_1205 ();
 sg13g2_fill_1 FILLER_1_1207 ();
 sg13g2_decap_8 FILLER_1_1219 ();
 sg13g2_decap_4 FILLER_1_1226 ();
 sg13g2_fill_2 FILLER_1_1230 ();
 sg13g2_decap_8 FILLER_1_1264 ();
 sg13g2_decap_8 FILLER_1_1271 ();
 sg13g2_decap_8 FILLER_1_1278 ();
 sg13g2_decap_8 FILLER_1_1285 ();
 sg13g2_decap_8 FILLER_1_1292 ();
 sg13g2_decap_8 FILLER_1_1299 ();
 sg13g2_decap_8 FILLER_1_1306 ();
 sg13g2_decap_8 FILLER_1_1313 ();
 sg13g2_decap_8 FILLER_1_1320 ();
 sg13g2_decap_8 FILLER_1_1327 ();
 sg13g2_decap_8 FILLER_1_1334 ();
 sg13g2_decap_8 FILLER_1_1341 ();
 sg13g2_decap_8 FILLER_1_1348 ();
 sg13g2_decap_8 FILLER_1_1355 ();
 sg13g2_decap_8 FILLER_1_1362 ();
 sg13g2_decap_8 FILLER_1_1369 ();
 sg13g2_decap_8 FILLER_1_1376 ();
 sg13g2_decap_8 FILLER_1_1383 ();
 sg13g2_decap_8 FILLER_1_1390 ();
 sg13g2_decap_8 FILLER_1_1397 ();
 sg13g2_decap_8 FILLER_1_1404 ();
 sg13g2_decap_8 FILLER_1_1411 ();
 sg13g2_decap_8 FILLER_1_1418 ();
 sg13g2_decap_8 FILLER_1_1425 ();
 sg13g2_decap_8 FILLER_1_1432 ();
 sg13g2_decap_8 FILLER_1_1439 ();
 sg13g2_decap_8 FILLER_1_1446 ();
 sg13g2_fill_2 FILLER_1_1453 ();
 sg13g2_fill_1 FILLER_1_1455 ();
 sg13g2_fill_1 FILLER_1_1459 ();
 sg13g2_decap_8 FILLER_1_1464 ();
 sg13g2_decap_8 FILLER_1_1471 ();
 sg13g2_decap_8 FILLER_1_1478 ();
 sg13g2_decap_8 FILLER_1_1485 ();
 sg13g2_decap_8 FILLER_1_1492 ();
 sg13g2_decap_8 FILLER_1_1499 ();
 sg13g2_decap_8 FILLER_1_1506 ();
 sg13g2_fill_2 FILLER_1_1513 ();
 sg13g2_decap_8 FILLER_1_1519 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1561 ();
 sg13g2_decap_8 FILLER_1_1568 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_8 FILLER_1_1582 ();
 sg13g2_decap_8 FILLER_1_1589 ();
 sg13g2_decap_8 FILLER_1_1596 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_decap_8 FILLER_1_1610 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_4 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1639 ();
 sg13g2_decap_4 FILLER_1_1646 ();
 sg13g2_decap_8 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1741 ();
 sg13g2_decap_8 FILLER_1_1748 ();
 sg13g2_decap_8 FILLER_1_1755 ();
 sg13g2_decap_8 FILLER_1_1762 ();
 sg13g2_decap_8 FILLER_1_1769 ();
 sg13g2_decap_8 FILLER_1_1776 ();
 sg13g2_decap_8 FILLER_1_1783 ();
 sg13g2_decap_8 FILLER_1_1790 ();
 sg13g2_decap_8 FILLER_1_1797 ();
 sg13g2_decap_8 FILLER_1_1804 ();
 sg13g2_fill_2 FILLER_1_1811 ();
 sg13g2_fill_1 FILLER_1_1813 ();
 sg13g2_decap_4 FILLER_1_1818 ();
 sg13g2_fill_1 FILLER_1_1822 ();
 sg13g2_decap_8 FILLER_1_1926 ();
 sg13g2_fill_2 FILLER_1_1933 ();
 sg13g2_decap_8 FILLER_1_1955 ();
 sg13g2_fill_2 FILLER_1_1975 ();
 sg13g2_fill_2 FILLER_1_1993 ();
 sg13g2_fill_1 FILLER_1_1995 ();
 sg13g2_fill_2 FILLER_1_2009 ();
 sg13g2_fill_1 FILLER_1_2011 ();
 sg13g2_decap_8 FILLER_1_2038 ();
 sg13g2_decap_8 FILLER_1_2045 ();
 sg13g2_decap_8 FILLER_1_2052 ();
 sg13g2_decap_4 FILLER_1_2059 ();
 sg13g2_fill_2 FILLER_1_2070 ();
 sg13g2_decap_8 FILLER_1_2091 ();
 sg13g2_decap_8 FILLER_1_2098 ();
 sg13g2_decap_4 FILLER_1_2105 ();
 sg13g2_fill_2 FILLER_1_2109 ();
 sg13g2_decap_8 FILLER_1_2115 ();
 sg13g2_decap_4 FILLER_1_2122 ();
 sg13g2_decap_8 FILLER_1_2148 ();
 sg13g2_decap_8 FILLER_1_2155 ();
 sg13g2_decap_4 FILLER_1_2162 ();
 sg13g2_fill_2 FILLER_1_2166 ();
 sg13g2_decap_8 FILLER_1_2209 ();
 sg13g2_decap_8 FILLER_1_2216 ();
 sg13g2_fill_2 FILLER_1_2223 ();
 sg13g2_fill_1 FILLER_1_2225 ();
 sg13g2_decap_8 FILLER_1_2229 ();
 sg13g2_decap_8 FILLER_1_2236 ();
 sg13g2_decap_8 FILLER_1_2243 ();
 sg13g2_decap_8 FILLER_1_2250 ();
 sg13g2_fill_1 FILLER_1_2257 ();
 sg13g2_decap_8 FILLER_1_2265 ();
 sg13g2_decap_8 FILLER_1_2272 ();
 sg13g2_decap_8 FILLER_1_2279 ();
 sg13g2_decap_4 FILLER_1_2286 ();
 sg13g2_fill_2 FILLER_1_2290 ();
 sg13g2_decap_8 FILLER_1_2299 ();
 sg13g2_decap_8 FILLER_1_2306 ();
 sg13g2_decap_8 FILLER_1_2313 ();
 sg13g2_decap_8 FILLER_1_2320 ();
 sg13g2_decap_8 FILLER_1_2327 ();
 sg13g2_decap_8 FILLER_1_2334 ();
 sg13g2_decap_8 FILLER_1_2341 ();
 sg13g2_fill_2 FILLER_1_2348 ();
 sg13g2_decap_8 FILLER_1_2354 ();
 sg13g2_decap_8 FILLER_1_2361 ();
 sg13g2_decap_8 FILLER_1_2368 ();
 sg13g2_decap_8 FILLER_1_2375 ();
 sg13g2_decap_8 FILLER_1_2382 ();
 sg13g2_decap_8 FILLER_1_2389 ();
 sg13g2_decap_4 FILLER_1_2396 ();
 sg13g2_fill_1 FILLER_1_2400 ();
 sg13g2_fill_1 FILLER_1_2416 ();
 sg13g2_decap_4 FILLER_1_2421 ();
 sg13g2_fill_1 FILLER_1_2425 ();
 sg13g2_decap_4 FILLER_1_2430 ();
 sg13g2_fill_2 FILLER_1_2447 ();
 sg13g2_decap_8 FILLER_1_2477 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_fill_1 FILLER_1_2491 ();
 sg13g2_decap_4 FILLER_1_2497 ();
 sg13g2_fill_2 FILLER_1_2505 ();
 sg13g2_fill_1 FILLER_1_2532 ();
 sg13g2_fill_2 FILLER_1_2567 ();
 sg13g2_fill_1 FILLER_1_2597 ();
 sg13g2_fill_2 FILLER_1_2606 ();
 sg13g2_fill_1 FILLER_1_2608 ();
 sg13g2_decap_8 FILLER_1_2618 ();
 sg13g2_decap_8 FILLER_1_2625 ();
 sg13g2_decap_4 FILLER_1_2632 ();
 sg13g2_fill_1 FILLER_1_2636 ();
 sg13g2_decap_8 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_1_2676 ();
 sg13g2_decap_8 FILLER_1_2683 ();
 sg13g2_decap_8 FILLER_1_2690 ();
 sg13g2_decap_8 FILLER_1_2697 ();
 sg13g2_decap_8 FILLER_1_2704 ();
 sg13g2_decap_4 FILLER_1_2711 ();
 sg13g2_decap_4 FILLER_1_2719 ();
 sg13g2_fill_2 FILLER_1_2723 ();
 sg13g2_decap_8 FILLER_1_2732 ();
 sg13g2_decap_8 FILLER_1_2739 ();
 sg13g2_decap_8 FILLER_1_2746 ();
 sg13g2_decap_8 FILLER_1_2753 ();
 sg13g2_decap_8 FILLER_1_2760 ();
 sg13g2_decap_8 FILLER_1_2767 ();
 sg13g2_decap_8 FILLER_1_2774 ();
 sg13g2_decap_8 FILLER_1_2781 ();
 sg13g2_decap_8 FILLER_1_2788 ();
 sg13g2_decap_8 FILLER_1_2795 ();
 sg13g2_decap_8 FILLER_1_2802 ();
 sg13g2_fill_1 FILLER_1_2809 ();
 sg13g2_fill_2 FILLER_1_2838 ();
 sg13g2_fill_1 FILLER_1_2840 ();
 sg13g2_decap_8 FILLER_1_2873 ();
 sg13g2_fill_2 FILLER_1_2880 ();
 sg13g2_fill_2 FILLER_1_2917 ();
 sg13g2_fill_1 FILLER_1_2919 ();
 sg13g2_decap_8 FILLER_1_2948 ();
 sg13g2_decap_8 FILLER_1_2955 ();
 sg13g2_decap_8 FILLER_1_2962 ();
 sg13g2_decap_8 FILLER_1_2969 ();
 sg13g2_decap_8 FILLER_1_2976 ();
 sg13g2_decap_8 FILLER_1_2983 ();
 sg13g2_decap_8 FILLER_1_2990 ();
 sg13g2_decap_8 FILLER_1_2997 ();
 sg13g2_decap_8 FILLER_1_3004 ();
 sg13g2_decap_8 FILLER_1_3011 ();
 sg13g2_decap_8 FILLER_1_3018 ();
 sg13g2_decap_8 FILLER_1_3025 ();
 sg13g2_decap_8 FILLER_1_3032 ();
 sg13g2_decap_8 FILLER_1_3039 ();
 sg13g2_decap_8 FILLER_1_3046 ();
 sg13g2_decap_8 FILLER_1_3053 ();
 sg13g2_decap_8 FILLER_1_3060 ();
 sg13g2_decap_8 FILLER_1_3067 ();
 sg13g2_decap_8 FILLER_1_3074 ();
 sg13g2_decap_8 FILLER_1_3081 ();
 sg13g2_decap_8 FILLER_1_3088 ();
 sg13g2_decap_8 FILLER_1_3095 ();
 sg13g2_decap_8 FILLER_1_3102 ();
 sg13g2_decap_8 FILLER_1_3109 ();
 sg13g2_decap_8 FILLER_1_3116 ();
 sg13g2_decap_8 FILLER_1_3123 ();
 sg13g2_decap_8 FILLER_1_3130 ();
 sg13g2_decap_8 FILLER_1_3137 ();
 sg13g2_decap_8 FILLER_1_3144 ();
 sg13g2_decap_8 FILLER_1_3151 ();
 sg13g2_decap_8 FILLER_1_3158 ();
 sg13g2_decap_8 FILLER_1_3165 ();
 sg13g2_decap_8 FILLER_1_3172 ();
 sg13g2_decap_8 FILLER_1_3179 ();
 sg13g2_decap_8 FILLER_1_3186 ();
 sg13g2_decap_8 FILLER_1_3193 ();
 sg13g2_decap_8 FILLER_1_3200 ();
 sg13g2_decap_8 FILLER_1_3207 ();
 sg13g2_decap_8 FILLER_1_3214 ();
 sg13g2_decap_8 FILLER_1_3221 ();
 sg13g2_decap_8 FILLER_1_3228 ();
 sg13g2_decap_8 FILLER_1_3235 ();
 sg13g2_decap_8 FILLER_1_3242 ();
 sg13g2_decap_8 FILLER_1_3249 ();
 sg13g2_decap_8 FILLER_1_3256 ();
 sg13g2_decap_8 FILLER_1_3263 ();
 sg13g2_decap_8 FILLER_1_3270 ();
 sg13g2_decap_8 FILLER_1_3277 ();
 sg13g2_decap_8 FILLER_1_3284 ();
 sg13g2_decap_8 FILLER_1_3291 ();
 sg13g2_decap_8 FILLER_1_3298 ();
 sg13g2_decap_8 FILLER_1_3305 ();
 sg13g2_decap_8 FILLER_1_3312 ();
 sg13g2_decap_8 FILLER_1_3319 ();
 sg13g2_decap_8 FILLER_1_3326 ();
 sg13g2_decap_8 FILLER_1_3333 ();
 sg13g2_decap_8 FILLER_1_3340 ();
 sg13g2_decap_8 FILLER_1_3347 ();
 sg13g2_decap_8 FILLER_1_3354 ();
 sg13g2_decap_8 FILLER_1_3361 ();
 sg13g2_decap_8 FILLER_1_3368 ();
 sg13g2_decap_8 FILLER_1_3375 ();
 sg13g2_decap_8 FILLER_1_3382 ();
 sg13g2_decap_8 FILLER_1_3389 ();
 sg13g2_decap_8 FILLER_1_3396 ();
 sg13g2_decap_8 FILLER_1_3403 ();
 sg13g2_decap_8 FILLER_1_3410 ();
 sg13g2_decap_8 FILLER_1_3417 ();
 sg13g2_decap_8 FILLER_1_3424 ();
 sg13g2_decap_8 FILLER_1_3431 ();
 sg13g2_decap_8 FILLER_1_3438 ();
 sg13g2_decap_8 FILLER_1_3445 ();
 sg13g2_decap_8 FILLER_1_3452 ();
 sg13g2_decap_8 FILLER_1_3459 ();
 sg13g2_decap_8 FILLER_1_3466 ();
 sg13g2_decap_8 FILLER_1_3473 ();
 sg13g2_decap_8 FILLER_1_3480 ();
 sg13g2_decap_8 FILLER_1_3487 ();
 sg13g2_decap_8 FILLER_1_3494 ();
 sg13g2_decap_8 FILLER_1_3501 ();
 sg13g2_decap_8 FILLER_1_3508 ();
 sg13g2_decap_8 FILLER_1_3515 ();
 sg13g2_decap_8 FILLER_1_3522 ();
 sg13g2_decap_8 FILLER_1_3529 ();
 sg13g2_decap_8 FILLER_1_3536 ();
 sg13g2_decap_8 FILLER_1_3543 ();
 sg13g2_decap_8 FILLER_1_3550 ();
 sg13g2_decap_8 FILLER_1_3557 ();
 sg13g2_decap_8 FILLER_1_3564 ();
 sg13g2_decap_8 FILLER_1_3571 ();
 sg13g2_fill_2 FILLER_1_3578 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_fill_2 FILLER_2_511 ();
 sg13g2_fill_1 FILLER_2_513 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_fill_2 FILLER_2_560 ();
 sg13g2_fill_2 FILLER_2_590 ();
 sg13g2_fill_1 FILLER_2_592 ();
 sg13g2_fill_2 FILLER_2_621 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_4 FILLER_2_693 ();
 sg13g2_fill_1 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_705 ();
 sg13g2_decap_4 FILLER_2_712 ();
 sg13g2_fill_2 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_729 ();
 sg13g2_decap_4 FILLER_2_736 ();
 sg13g2_fill_2 FILLER_2_740 ();
 sg13g2_fill_1 FILLER_2_746 ();
 sg13g2_decap_4 FILLER_2_754 ();
 sg13g2_fill_2 FILLER_2_758 ();
 sg13g2_decap_4 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_785 ();
 sg13g2_decap_8 FILLER_2_792 ();
 sg13g2_decap_4 FILLER_2_799 ();
 sg13g2_fill_1 FILLER_2_803 ();
 sg13g2_decap_8 FILLER_2_841 ();
 sg13g2_decap_8 FILLER_2_848 ();
 sg13g2_decap_8 FILLER_2_855 ();
 sg13g2_decap_8 FILLER_2_862 ();
 sg13g2_decap_4 FILLER_2_869 ();
 sg13g2_fill_1 FILLER_2_873 ();
 sg13g2_decap_4 FILLER_2_885 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_4 FILLER_2_900 ();
 sg13g2_fill_1 FILLER_2_904 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_4 FILLER_2_928 ();
 sg13g2_fill_1 FILLER_2_932 ();
 sg13g2_fill_2 FILLER_2_941 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1036 ();
 sg13g2_decap_8 FILLER_2_1043 ();
 sg13g2_decap_8 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1057 ();
 sg13g2_decap_8 FILLER_2_1064 ();
 sg13g2_decap_8 FILLER_2_1071 ();
 sg13g2_decap_8 FILLER_2_1078 ();
 sg13g2_decap_8 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1092 ();
 sg13g2_decap_8 FILLER_2_1099 ();
 sg13g2_decap_8 FILLER_2_1106 ();
 sg13g2_decap_8 FILLER_2_1113 ();
 sg13g2_decap_8 FILLER_2_1120 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_4 FILLER_2_1162 ();
 sg13g2_fill_1 FILLER_2_1166 ();
 sg13g2_decap_4 FILLER_2_1180 ();
 sg13g2_decap_8 FILLER_2_1197 ();
 sg13g2_decap_4 FILLER_2_1204 ();
 sg13g2_decap_8 FILLER_2_1226 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_fill_2 FILLER_2_1240 ();
 sg13g2_fill_1 FILLER_2_1242 ();
 sg13g2_fill_2 FILLER_2_1248 ();
 sg13g2_fill_1 FILLER_2_1250 ();
 sg13g2_decap_4 FILLER_2_1255 ();
 sg13g2_fill_2 FILLER_2_1259 ();
 sg13g2_fill_2 FILLER_2_1292 ();
 sg13g2_fill_1 FILLER_2_1294 ();
 sg13g2_fill_2 FILLER_2_1323 ();
 sg13g2_fill_1 FILLER_2_1325 ();
 sg13g2_decap_8 FILLER_2_1354 ();
 sg13g2_decap_8 FILLER_2_1361 ();
 sg13g2_decap_8 FILLER_2_1368 ();
 sg13g2_decap_8 FILLER_2_1375 ();
 sg13g2_decap_8 FILLER_2_1382 ();
 sg13g2_decap_8 FILLER_2_1389 ();
 sg13g2_decap_8 FILLER_2_1396 ();
 sg13g2_decap_8 FILLER_2_1403 ();
 sg13g2_decap_8 FILLER_2_1410 ();
 sg13g2_decap_8 FILLER_2_1417 ();
 sg13g2_fill_2 FILLER_2_1424 ();
 sg13g2_fill_1 FILLER_2_1426 ();
 sg13g2_fill_2 FILLER_2_1483 ();
 sg13g2_fill_1 FILLER_2_1485 ();
 sg13g2_fill_2 FILLER_2_1490 ();
 sg13g2_fill_1 FILLER_2_1492 ();
 sg13g2_decap_8 FILLER_2_1500 ();
 sg13g2_fill_2 FILLER_2_1507 ();
 sg13g2_fill_1 FILLER_2_1509 ();
 sg13g2_decap_8 FILLER_2_1538 ();
 sg13g2_decap_8 FILLER_2_1545 ();
 sg13g2_decap_8 FILLER_2_1552 ();
 sg13g2_decap_8 FILLER_2_1559 ();
 sg13g2_decap_8 FILLER_2_1566 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_decap_8 FILLER_2_1580 ();
 sg13g2_decap_8 FILLER_2_1587 ();
 sg13g2_decap_8 FILLER_2_1594 ();
 sg13g2_decap_8 FILLER_2_1601 ();
 sg13g2_fill_2 FILLER_2_1608 ();
 sg13g2_decap_8 FILLER_2_1614 ();
 sg13g2_decap_8 FILLER_2_1621 ();
 sg13g2_decap_4 FILLER_2_1628 ();
 sg13g2_fill_1 FILLER_2_1632 ();
 sg13g2_decap_4 FILLER_2_1636 ();
 sg13g2_fill_1 FILLER_2_1662 ();
 sg13g2_fill_2 FILLER_2_1667 ();
 sg13g2_fill_1 FILLER_2_1669 ();
 sg13g2_fill_2 FILLER_2_1727 ();
 sg13g2_decap_8 FILLER_2_1742 ();
 sg13g2_decap_8 FILLER_2_1749 ();
 sg13g2_decap_8 FILLER_2_1756 ();
 sg13g2_decap_8 FILLER_2_1763 ();
 sg13g2_decap_8 FILLER_2_1770 ();
 sg13g2_fill_2 FILLER_2_1777 ();
 sg13g2_fill_1 FILLER_2_1779 ();
 sg13g2_decap_8 FILLER_2_1784 ();
 sg13g2_decap_8 FILLER_2_1791 ();
 sg13g2_decap_8 FILLER_2_1798 ();
 sg13g2_decap_4 FILLER_2_1805 ();
 sg13g2_fill_2 FILLER_2_1841 ();
 sg13g2_decap_8 FILLER_2_1862 ();
 sg13g2_decap_8 FILLER_2_1869 ();
 sg13g2_fill_2 FILLER_2_1881 ();
 sg13g2_fill_1 FILLER_2_1883 ();
 sg13g2_decap_4 FILLER_2_1935 ();
 sg13g2_decap_8 FILLER_2_1952 ();
 sg13g2_fill_1 FILLER_2_1959 ();
 sg13g2_fill_1 FILLER_2_1985 ();
 sg13g2_decap_8 FILLER_2_1998 ();
 sg13g2_decap_8 FILLER_2_2005 ();
 sg13g2_decap_8 FILLER_2_2012 ();
 sg13g2_decap_4 FILLER_2_2019 ();
 sg13g2_fill_2 FILLER_2_2023 ();
 sg13g2_decap_8 FILLER_2_2058 ();
 sg13g2_fill_1 FILLER_2_2065 ();
 sg13g2_fill_2 FILLER_2_2072 ();
 sg13g2_fill_1 FILLER_2_2102 ();
 sg13g2_fill_2 FILLER_2_2134 ();
 sg13g2_fill_1 FILLER_2_2177 ();
 sg13g2_fill_2 FILLER_2_2189 ();
 sg13g2_decap_4 FILLER_2_2284 ();
 sg13g2_fill_1 FILLER_2_2288 ();
 sg13g2_decap_8 FILLER_2_2321 ();
 sg13g2_decap_8 FILLER_2_2328 ();
 sg13g2_decap_8 FILLER_2_2335 ();
 sg13g2_fill_2 FILLER_2_2342 ();
 sg13g2_fill_1 FILLER_2_2344 ();
 sg13g2_decap_8 FILLER_2_2358 ();
 sg13g2_fill_2 FILLER_2_2365 ();
 sg13g2_decap_4 FILLER_2_2374 ();
 sg13g2_fill_1 FILLER_2_2378 ();
 sg13g2_decap_4 FILLER_2_2384 ();
 sg13g2_fill_2 FILLER_2_2388 ();
 sg13g2_decap_4 FILLER_2_2420 ();
 sg13g2_fill_2 FILLER_2_2437 ();
 sg13g2_decap_8 FILLER_2_2449 ();
 sg13g2_decap_4 FILLER_2_2456 ();
 sg13g2_decap_4 FILLER_2_2464 ();
 sg13g2_decap_4 FILLER_2_2472 ();
 sg13g2_fill_2 FILLER_2_2485 ();
 sg13g2_fill_1 FILLER_2_2487 ();
 sg13g2_decap_8 FILLER_2_2507 ();
 sg13g2_fill_2 FILLER_2_2514 ();
 sg13g2_fill_1 FILLER_2_2516 ();
 sg13g2_fill_2 FILLER_2_2527 ();
 sg13g2_fill_1 FILLER_2_2529 ();
 sg13g2_fill_1 FILLER_2_2544 ();
 sg13g2_fill_1 FILLER_2_2549 ();
 sg13g2_fill_1 FILLER_2_2555 ();
 sg13g2_decap_8 FILLER_2_2561 ();
 sg13g2_fill_2 FILLER_2_2568 ();
 sg13g2_fill_1 FILLER_2_2600 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_fill_2 FILLER_2_2636 ();
 sg13g2_fill_1 FILLER_2_2638 ();
 sg13g2_fill_2 FILLER_2_2652 ();
 sg13g2_fill_1 FILLER_2_2654 ();
 sg13g2_decap_8 FILLER_2_2665 ();
 sg13g2_fill_2 FILLER_2_2680 ();
 sg13g2_decap_8 FILLER_2_2695 ();
 sg13g2_fill_2 FILLER_2_2702 ();
 sg13g2_fill_1 FILLER_2_2704 ();
 sg13g2_fill_1 FILLER_2_2709 ();
 sg13g2_decap_8 FILLER_2_2738 ();
 sg13g2_fill_1 FILLER_2_2750 ();
 sg13g2_decap_8 FILLER_2_2761 ();
 sg13g2_decap_8 FILLER_2_2768 ();
 sg13g2_decap_8 FILLER_2_2775 ();
 sg13g2_decap_8 FILLER_2_2795 ();
 sg13g2_decap_8 FILLER_2_2802 ();
 sg13g2_decap_4 FILLER_2_2809 ();
 sg13g2_fill_2 FILLER_2_2813 ();
 sg13g2_fill_2 FILLER_2_2835 ();
 sg13g2_fill_1 FILLER_2_2837 ();
 sg13g2_fill_1 FILLER_2_2851 ();
 sg13g2_decap_4 FILLER_2_2874 ();
 sg13g2_decap_8 FILLER_2_2892 ();
 sg13g2_fill_1 FILLER_2_2899 ();
 sg13g2_fill_2 FILLER_2_2909 ();
 sg13g2_fill_1 FILLER_2_2924 ();
 sg13g2_decap_8 FILLER_2_2929 ();
 sg13g2_decap_8 FILLER_2_2943 ();
 sg13g2_decap_4 FILLER_2_2950 ();
 sg13g2_decap_4 FILLER_2_2959 ();
 sg13g2_fill_2 FILLER_2_2963 ();
 sg13g2_decap_8 FILLER_2_2993 ();
 sg13g2_decap_8 FILLER_2_3000 ();
 sg13g2_decap_8 FILLER_2_3007 ();
 sg13g2_decap_8 FILLER_2_3014 ();
 sg13g2_decap_8 FILLER_2_3021 ();
 sg13g2_decap_8 FILLER_2_3028 ();
 sg13g2_decap_8 FILLER_2_3035 ();
 sg13g2_decap_8 FILLER_2_3042 ();
 sg13g2_decap_8 FILLER_2_3049 ();
 sg13g2_decap_8 FILLER_2_3056 ();
 sg13g2_decap_8 FILLER_2_3063 ();
 sg13g2_decap_8 FILLER_2_3070 ();
 sg13g2_decap_8 FILLER_2_3077 ();
 sg13g2_decap_8 FILLER_2_3084 ();
 sg13g2_decap_8 FILLER_2_3091 ();
 sg13g2_decap_8 FILLER_2_3098 ();
 sg13g2_decap_8 FILLER_2_3105 ();
 sg13g2_decap_8 FILLER_2_3112 ();
 sg13g2_decap_8 FILLER_2_3119 ();
 sg13g2_decap_8 FILLER_2_3126 ();
 sg13g2_decap_8 FILLER_2_3133 ();
 sg13g2_decap_8 FILLER_2_3140 ();
 sg13g2_decap_8 FILLER_2_3147 ();
 sg13g2_decap_8 FILLER_2_3154 ();
 sg13g2_decap_8 FILLER_2_3161 ();
 sg13g2_decap_8 FILLER_2_3168 ();
 sg13g2_decap_8 FILLER_2_3175 ();
 sg13g2_decap_8 FILLER_2_3182 ();
 sg13g2_decap_8 FILLER_2_3189 ();
 sg13g2_decap_8 FILLER_2_3196 ();
 sg13g2_decap_8 FILLER_2_3203 ();
 sg13g2_decap_8 FILLER_2_3210 ();
 sg13g2_decap_8 FILLER_2_3217 ();
 sg13g2_decap_8 FILLER_2_3224 ();
 sg13g2_decap_8 FILLER_2_3231 ();
 sg13g2_decap_8 FILLER_2_3238 ();
 sg13g2_decap_8 FILLER_2_3245 ();
 sg13g2_decap_8 FILLER_2_3252 ();
 sg13g2_decap_8 FILLER_2_3259 ();
 sg13g2_decap_8 FILLER_2_3266 ();
 sg13g2_decap_8 FILLER_2_3273 ();
 sg13g2_decap_8 FILLER_2_3280 ();
 sg13g2_decap_8 FILLER_2_3287 ();
 sg13g2_decap_8 FILLER_2_3294 ();
 sg13g2_decap_8 FILLER_2_3301 ();
 sg13g2_decap_8 FILLER_2_3308 ();
 sg13g2_decap_8 FILLER_2_3315 ();
 sg13g2_decap_8 FILLER_2_3322 ();
 sg13g2_decap_8 FILLER_2_3329 ();
 sg13g2_decap_8 FILLER_2_3336 ();
 sg13g2_decap_8 FILLER_2_3343 ();
 sg13g2_decap_8 FILLER_2_3350 ();
 sg13g2_decap_8 FILLER_2_3357 ();
 sg13g2_decap_8 FILLER_2_3364 ();
 sg13g2_decap_8 FILLER_2_3371 ();
 sg13g2_decap_8 FILLER_2_3378 ();
 sg13g2_decap_8 FILLER_2_3385 ();
 sg13g2_decap_8 FILLER_2_3392 ();
 sg13g2_decap_8 FILLER_2_3399 ();
 sg13g2_decap_8 FILLER_2_3406 ();
 sg13g2_decap_8 FILLER_2_3413 ();
 sg13g2_decap_8 FILLER_2_3420 ();
 sg13g2_decap_8 FILLER_2_3427 ();
 sg13g2_decap_8 FILLER_2_3434 ();
 sg13g2_decap_8 FILLER_2_3441 ();
 sg13g2_decap_8 FILLER_2_3448 ();
 sg13g2_decap_8 FILLER_2_3455 ();
 sg13g2_decap_8 FILLER_2_3462 ();
 sg13g2_decap_8 FILLER_2_3469 ();
 sg13g2_decap_8 FILLER_2_3476 ();
 sg13g2_decap_8 FILLER_2_3483 ();
 sg13g2_decap_8 FILLER_2_3490 ();
 sg13g2_decap_8 FILLER_2_3497 ();
 sg13g2_decap_8 FILLER_2_3504 ();
 sg13g2_decap_8 FILLER_2_3511 ();
 sg13g2_decap_8 FILLER_2_3518 ();
 sg13g2_decap_8 FILLER_2_3525 ();
 sg13g2_decap_8 FILLER_2_3532 ();
 sg13g2_decap_8 FILLER_2_3539 ();
 sg13g2_decap_8 FILLER_2_3546 ();
 sg13g2_decap_8 FILLER_2_3553 ();
 sg13g2_decap_8 FILLER_2_3560 ();
 sg13g2_decap_8 FILLER_2_3567 ();
 sg13g2_decap_4 FILLER_2_3574 ();
 sg13g2_fill_2 FILLER_2_3578 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_4 FILLER_3_504 ();
 sg13g2_fill_1 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_544 ();
 sg13g2_decap_8 FILLER_3_551 ();
 sg13g2_fill_1 FILLER_3_558 ();
 sg13g2_decap_4 FILLER_3_591 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_4 FILLER_3_620 ();
 sg13g2_fill_1 FILLER_3_624 ();
 sg13g2_decap_8 FILLER_3_635 ();
 sg13g2_decap_8 FILLER_3_642 ();
 sg13g2_decap_4 FILLER_3_649 ();
 sg13g2_fill_1 FILLER_3_653 ();
 sg13g2_fill_1 FILLER_3_673 ();
 sg13g2_decap_8 FILLER_3_687 ();
 sg13g2_fill_1 FILLER_3_694 ();
 sg13g2_decap_4 FILLER_3_723 ();
 sg13g2_fill_1 FILLER_3_727 ();
 sg13g2_decap_8 FILLER_3_741 ();
 sg13g2_fill_1 FILLER_3_766 ();
 sg13g2_fill_1 FILLER_3_785 ();
 sg13g2_decap_4 FILLER_3_794 ();
 sg13g2_fill_2 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_820 ();
 sg13g2_decap_8 FILLER_3_827 ();
 sg13g2_decap_8 FILLER_3_834 ();
 sg13g2_decap_8 FILLER_3_841 ();
 sg13g2_decap_8 FILLER_3_848 ();
 sg13g2_decap_8 FILLER_3_855 ();
 sg13g2_decap_8 FILLER_3_862 ();
 sg13g2_fill_1 FILLER_3_869 ();
 sg13g2_fill_2 FILLER_3_1010 ();
 sg13g2_decap_4 FILLER_3_1040 ();
 sg13g2_fill_2 FILLER_3_1044 ();
 sg13g2_decap_8 FILLER_3_1059 ();
 sg13g2_fill_2 FILLER_3_1066 ();
 sg13g2_decap_8 FILLER_3_1071 ();
 sg13g2_decap_8 FILLER_3_1078 ();
 sg13g2_decap_8 FILLER_3_1085 ();
 sg13g2_decap_8 FILLER_3_1092 ();
 sg13g2_decap_8 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1113 ();
 sg13g2_decap_8 FILLER_3_1124 ();
 sg13g2_fill_1 FILLER_3_1148 ();
 sg13g2_decap_4 FILLER_3_1161 ();
 sg13g2_fill_2 FILLER_3_1165 ();
 sg13g2_decap_4 FILLER_3_1206 ();
 sg13g2_fill_1 FILLER_3_1210 ();
 sg13g2_fill_2 FILLER_3_1228 ();
 sg13g2_decap_8 FILLER_3_1283 ();
 sg13g2_decap_4 FILLER_3_1290 ();
 sg13g2_fill_2 FILLER_3_1294 ();
 sg13g2_decap_8 FILLER_3_1307 ();
 sg13g2_decap_8 FILLER_3_1314 ();
 sg13g2_decap_4 FILLER_3_1321 ();
 sg13g2_fill_1 FILLER_3_1341 ();
 sg13g2_decap_8 FILLER_3_1361 ();
 sg13g2_decap_8 FILLER_3_1368 ();
 sg13g2_decap_4 FILLER_3_1375 ();
 sg13g2_fill_1 FILLER_3_1379 ();
 sg13g2_fill_1 FILLER_3_1408 ();
 sg13g2_decap_8 FILLER_3_1416 ();
 sg13g2_decap_4 FILLER_3_1423 ();
 sg13g2_fill_2 FILLER_3_1427 ();
 sg13g2_decap_4 FILLER_3_1436 ();
 sg13g2_decap_8 FILLER_3_1468 ();
 sg13g2_decap_4 FILLER_3_1475 ();
 sg13g2_fill_1 FILLER_3_1479 ();
 sg13g2_fill_2 FILLER_3_1524 ();
 sg13g2_decap_8 FILLER_3_1562 ();
 sg13g2_decap_8 FILLER_3_1569 ();
 sg13g2_decap_8 FILLER_3_1576 ();
 sg13g2_decap_8 FILLER_3_1590 ();
 sg13g2_decap_8 FILLER_3_1597 ();
 sg13g2_fill_1 FILLER_3_1604 ();
 sg13g2_fill_2 FILLER_3_1633 ();
 sg13g2_decap_4 FILLER_3_1665 ();
 sg13g2_fill_2 FILLER_3_1673 ();
 sg13g2_fill_1 FILLER_3_1675 ();
 sg13g2_decap_8 FILLER_3_1689 ();
 sg13g2_fill_2 FILLER_3_1730 ();
 sg13g2_decap_4 FILLER_3_1745 ();
 sg13g2_fill_2 FILLER_3_1749 ();
 sg13g2_decap_8 FILLER_3_1755 ();
 sg13g2_decap_8 FILLER_3_1762 ();
 sg13g2_fill_2 FILLER_3_1769 ();
 sg13g2_fill_1 FILLER_3_1771 ();
 sg13g2_fill_2 FILLER_3_1803 ();
 sg13g2_fill_1 FILLER_3_1805 ();
 sg13g2_fill_1 FILLER_3_1812 ();
 sg13g2_fill_1 FILLER_3_1823 ();
 sg13g2_fill_2 FILLER_3_1834 ();
 sg13g2_decap_8 FILLER_3_1858 ();
 sg13g2_fill_1 FILLER_3_1865 ();
 sg13g2_fill_2 FILLER_3_1876 ();
 sg13g2_fill_1 FILLER_3_1878 ();
 sg13g2_fill_1 FILLER_3_1888 ();
 sg13g2_fill_1 FILLER_3_1905 ();
 sg13g2_fill_2 FILLER_3_1924 ();
 sg13g2_fill_1 FILLER_3_1926 ();
 sg13g2_fill_1 FILLER_3_1938 ();
 sg13g2_fill_1 FILLER_3_1949 ();
 sg13g2_decap_8 FILLER_3_1958 ();
 sg13g2_decap_8 FILLER_3_1965 ();
 sg13g2_fill_2 FILLER_3_1972 ();
 sg13g2_fill_1 FILLER_3_1974 ();
 sg13g2_fill_1 FILLER_3_1980 ();
 sg13g2_fill_2 FILLER_3_1986 ();
 sg13g2_fill_1 FILLER_3_1988 ();
 sg13g2_decap_8 FILLER_3_1996 ();
 sg13g2_decap_8 FILLER_3_2003 ();
 sg13g2_decap_8 FILLER_3_2027 ();
 sg13g2_decap_4 FILLER_3_2065 ();
 sg13g2_fill_2 FILLER_3_2069 ();
 sg13g2_decap_8 FILLER_3_2083 ();
 sg13g2_decap_8 FILLER_3_2118 ();
 sg13g2_decap_8 FILLER_3_2125 ();
 sg13g2_decap_4 FILLER_3_2132 ();
 sg13g2_fill_1 FILLER_3_2136 ();
 sg13g2_fill_1 FILLER_3_2143 ();
 sg13g2_fill_1 FILLER_3_2183 ();
 sg13g2_decap_8 FILLER_3_2189 ();
 sg13g2_fill_1 FILLER_3_2196 ();
 sg13g2_decap_4 FILLER_3_2200 ();
 sg13g2_fill_1 FILLER_3_2204 ();
 sg13g2_fill_2 FILLER_3_2220 ();
 sg13g2_fill_1 FILLER_3_2222 ();
 sg13g2_fill_2 FILLER_3_2229 ();
 sg13g2_fill_2 FILLER_3_2258 ();
 sg13g2_fill_1 FILLER_3_2260 ();
 sg13g2_decap_4 FILLER_3_2265 ();
 sg13g2_fill_1 FILLER_3_2269 ();
 sg13g2_decap_8 FILLER_3_2278 ();
 sg13g2_decap_8 FILLER_3_2285 ();
 sg13g2_fill_2 FILLER_3_2292 ();
 sg13g2_fill_1 FILLER_3_2294 ();
 sg13g2_fill_2 FILLER_3_2299 ();
 sg13g2_fill_2 FILLER_3_2310 ();
 sg13g2_decap_4 FILLER_3_2340 ();
 sg13g2_fill_1 FILLER_3_2344 ();
 sg13g2_fill_1 FILLER_3_2373 ();
 sg13g2_fill_2 FILLER_3_2395 ();
 sg13g2_fill_1 FILLER_3_2397 ();
 sg13g2_decap_8 FILLER_3_2416 ();
 sg13g2_fill_1 FILLER_3_2423 ();
 sg13g2_fill_2 FILLER_3_2450 ();
 sg13g2_decap_4 FILLER_3_2490 ();
 sg13g2_decap_4 FILLER_3_2505 ();
 sg13g2_fill_2 FILLER_3_2509 ();
 sg13g2_fill_2 FILLER_3_2523 ();
 sg13g2_decap_8 FILLER_3_2535 ();
 sg13g2_fill_2 FILLER_3_2542 ();
 sg13g2_decap_4 FILLER_3_2583 ();
 sg13g2_fill_1 FILLER_3_2587 ();
 sg13g2_decap_4 FILLER_3_2616 ();
 sg13g2_fill_1 FILLER_3_2620 ();
 sg13g2_fill_2 FILLER_3_2671 ();
 sg13g2_fill_1 FILLER_3_2673 ();
 sg13g2_fill_2 FILLER_3_2705 ();
 sg13g2_fill_2 FILLER_3_2719 ();
 sg13g2_fill_1 FILLER_3_2721 ();
 sg13g2_fill_1 FILLER_3_2735 ();
 sg13g2_fill_2 FILLER_3_2745 ();
 sg13g2_decap_8 FILLER_3_2763 ();
 sg13g2_decap_4 FILLER_3_2770 ();
 sg13g2_fill_1 FILLER_3_2774 ();
 sg13g2_decap_4 FILLER_3_2788 ();
 sg13g2_fill_2 FILLER_3_2792 ();
 sg13g2_decap_8 FILLER_3_2812 ();
 sg13g2_fill_2 FILLER_3_2819 ();
 sg13g2_fill_1 FILLER_3_2821 ();
 sg13g2_fill_2 FILLER_3_2844 ();
 sg13g2_fill_2 FILLER_3_2855 ();
 sg13g2_fill_1 FILLER_3_2862 ();
 sg13g2_fill_2 FILLER_3_2871 ();
 sg13g2_fill_1 FILLER_3_2873 ();
 sg13g2_decap_8 FILLER_3_2899 ();
 sg13g2_fill_1 FILLER_3_2927 ();
 sg13g2_fill_2 FILLER_3_2959 ();
 sg13g2_fill_2 FILLER_3_2968 ();
 sg13g2_fill_1 FILLER_3_2970 ();
 sg13g2_decap_8 FILLER_3_2975 ();
 sg13g2_decap_8 FILLER_3_2982 ();
 sg13g2_decap_8 FILLER_3_2989 ();
 sg13g2_decap_8 FILLER_3_2996 ();
 sg13g2_decap_8 FILLER_3_3003 ();
 sg13g2_decap_8 FILLER_3_3010 ();
 sg13g2_decap_8 FILLER_3_3017 ();
 sg13g2_decap_8 FILLER_3_3024 ();
 sg13g2_decap_8 FILLER_3_3031 ();
 sg13g2_decap_8 FILLER_3_3038 ();
 sg13g2_decap_8 FILLER_3_3045 ();
 sg13g2_decap_8 FILLER_3_3052 ();
 sg13g2_decap_8 FILLER_3_3059 ();
 sg13g2_decap_8 FILLER_3_3066 ();
 sg13g2_decap_8 FILLER_3_3073 ();
 sg13g2_decap_8 FILLER_3_3080 ();
 sg13g2_decap_8 FILLER_3_3087 ();
 sg13g2_decap_8 FILLER_3_3094 ();
 sg13g2_decap_8 FILLER_3_3101 ();
 sg13g2_decap_8 FILLER_3_3108 ();
 sg13g2_decap_8 FILLER_3_3115 ();
 sg13g2_decap_8 FILLER_3_3122 ();
 sg13g2_decap_8 FILLER_3_3129 ();
 sg13g2_decap_8 FILLER_3_3136 ();
 sg13g2_decap_8 FILLER_3_3143 ();
 sg13g2_decap_8 FILLER_3_3150 ();
 sg13g2_decap_8 FILLER_3_3157 ();
 sg13g2_decap_8 FILLER_3_3164 ();
 sg13g2_decap_8 FILLER_3_3171 ();
 sg13g2_decap_8 FILLER_3_3178 ();
 sg13g2_decap_8 FILLER_3_3185 ();
 sg13g2_decap_8 FILLER_3_3192 ();
 sg13g2_decap_8 FILLER_3_3199 ();
 sg13g2_decap_8 FILLER_3_3206 ();
 sg13g2_decap_8 FILLER_3_3213 ();
 sg13g2_decap_8 FILLER_3_3220 ();
 sg13g2_decap_8 FILLER_3_3227 ();
 sg13g2_decap_8 FILLER_3_3234 ();
 sg13g2_decap_8 FILLER_3_3241 ();
 sg13g2_decap_8 FILLER_3_3248 ();
 sg13g2_decap_8 FILLER_3_3255 ();
 sg13g2_decap_8 FILLER_3_3262 ();
 sg13g2_decap_8 FILLER_3_3269 ();
 sg13g2_decap_8 FILLER_3_3276 ();
 sg13g2_decap_8 FILLER_3_3283 ();
 sg13g2_decap_8 FILLER_3_3290 ();
 sg13g2_decap_8 FILLER_3_3297 ();
 sg13g2_decap_8 FILLER_3_3304 ();
 sg13g2_decap_8 FILLER_3_3311 ();
 sg13g2_decap_8 FILLER_3_3318 ();
 sg13g2_decap_8 FILLER_3_3325 ();
 sg13g2_decap_8 FILLER_3_3332 ();
 sg13g2_decap_8 FILLER_3_3339 ();
 sg13g2_decap_8 FILLER_3_3346 ();
 sg13g2_decap_8 FILLER_3_3353 ();
 sg13g2_decap_8 FILLER_3_3360 ();
 sg13g2_decap_8 FILLER_3_3367 ();
 sg13g2_decap_8 FILLER_3_3374 ();
 sg13g2_decap_8 FILLER_3_3381 ();
 sg13g2_decap_8 FILLER_3_3388 ();
 sg13g2_decap_8 FILLER_3_3395 ();
 sg13g2_decap_8 FILLER_3_3402 ();
 sg13g2_decap_8 FILLER_3_3409 ();
 sg13g2_decap_8 FILLER_3_3416 ();
 sg13g2_decap_8 FILLER_3_3423 ();
 sg13g2_decap_8 FILLER_3_3430 ();
 sg13g2_decap_8 FILLER_3_3437 ();
 sg13g2_decap_8 FILLER_3_3444 ();
 sg13g2_decap_8 FILLER_3_3451 ();
 sg13g2_decap_8 FILLER_3_3458 ();
 sg13g2_decap_8 FILLER_3_3465 ();
 sg13g2_decap_8 FILLER_3_3472 ();
 sg13g2_decap_8 FILLER_3_3479 ();
 sg13g2_decap_8 FILLER_3_3486 ();
 sg13g2_decap_8 FILLER_3_3493 ();
 sg13g2_decap_8 FILLER_3_3500 ();
 sg13g2_decap_8 FILLER_3_3507 ();
 sg13g2_decap_8 FILLER_3_3514 ();
 sg13g2_decap_8 FILLER_3_3521 ();
 sg13g2_decap_8 FILLER_3_3528 ();
 sg13g2_decap_8 FILLER_3_3535 ();
 sg13g2_decap_8 FILLER_3_3542 ();
 sg13g2_decap_8 FILLER_3_3549 ();
 sg13g2_decap_8 FILLER_3_3556 ();
 sg13g2_decap_8 FILLER_3_3563 ();
 sg13g2_decap_8 FILLER_3_3570 ();
 sg13g2_fill_2 FILLER_3_3577 ();
 sg13g2_fill_1 FILLER_3_3579 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_4 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_440 ();
 sg13g2_decap_8 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_461 ();
 sg13g2_decap_8 FILLER_4_468 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_482 ();
 sg13g2_decap_8 FILLER_4_489 ();
 sg13g2_decap_8 FILLER_4_496 ();
 sg13g2_decap_8 FILLER_4_503 ();
 sg13g2_decap_8 FILLER_4_510 ();
 sg13g2_decap_8 FILLER_4_517 ();
 sg13g2_fill_2 FILLER_4_524 ();
 sg13g2_fill_1 FILLER_4_526 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_fill_1 FILLER_4_557 ();
 sg13g2_decap_8 FILLER_4_578 ();
 sg13g2_fill_2 FILLER_4_585 ();
 sg13g2_fill_2 FILLER_4_608 ();
 sg13g2_fill_1 FILLER_4_610 ();
 sg13g2_fill_2 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_4 FILLER_4_677 ();
 sg13g2_fill_1 FILLER_4_681 ();
 sg13g2_fill_1 FILLER_4_722 ();
 sg13g2_fill_2 FILLER_4_754 ();
 sg13g2_fill_2 FILLER_4_761 ();
 sg13g2_fill_1 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_4 FILLER_4_825 ();
 sg13g2_fill_1 FILLER_4_842 ();
 sg13g2_decap_4 FILLER_4_856 ();
 sg13g2_fill_1 FILLER_4_860 ();
 sg13g2_fill_2 FILLER_4_874 ();
 sg13g2_fill_2 FILLER_4_889 ();
 sg13g2_fill_1 FILLER_4_891 ();
 sg13g2_fill_2 FILLER_4_907 ();
 sg13g2_fill_1 FILLER_4_909 ();
 sg13g2_fill_1 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_943 ();
 sg13g2_decap_4 FILLER_4_950 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_fill_1 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_4 FILLER_4_1005 ();
 sg13g2_fill_1 FILLER_4_1016 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_fill_2 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_4_1043 ();
 sg13g2_fill_1 FILLER_4_1050 ();
 sg13g2_fill_2 FILLER_4_1079 ();
 sg13g2_fill_1 FILLER_4_1081 ();
 sg13g2_decap_8 FILLER_4_1086 ();
 sg13g2_decap_8 FILLER_4_1093 ();
 sg13g2_decap_8 FILLER_4_1100 ();
 sg13g2_fill_2 FILLER_4_1107 ();
 sg13g2_fill_1 FILLER_4_1109 ();
 sg13g2_fill_1 FILLER_4_1114 ();
 sg13g2_fill_2 FILLER_4_1151 ();
 sg13g2_fill_1 FILLER_4_1153 ();
 sg13g2_fill_1 FILLER_4_1175 ();
 sg13g2_decap_4 FILLER_4_1181 ();
 sg13g2_fill_1 FILLER_4_1185 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_4 FILLER_4_1206 ();
 sg13g2_fill_2 FILLER_4_1210 ();
 sg13g2_fill_2 FILLER_4_1229 ();
 sg13g2_fill_2 FILLER_4_1255 ();
 sg13g2_decap_4 FILLER_4_1285 ();
 sg13g2_fill_2 FILLER_4_1315 ();
 sg13g2_fill_1 FILLER_4_1338 ();
 sg13g2_decap_4 FILLER_4_1376 ();
 sg13g2_fill_1 FILLER_4_1380 ();
 sg13g2_decap_8 FILLER_4_1392 ();
 sg13g2_decap_8 FILLER_4_1399 ();
 sg13g2_fill_2 FILLER_4_1447 ();
 sg13g2_fill_2 FILLER_4_1472 ();
 sg13g2_decap_8 FILLER_4_1491 ();
 sg13g2_decap_8 FILLER_4_1498 ();
 sg13g2_fill_2 FILLER_4_1505 ();
 sg13g2_fill_1 FILLER_4_1507 ();
 sg13g2_decap_4 FILLER_4_1515 ();
 sg13g2_fill_1 FILLER_4_1529 ();
 sg13g2_decap_8 FILLER_4_1539 ();
 sg13g2_fill_2 FILLER_4_1546 ();
 sg13g2_fill_2 FILLER_4_1573 ();
 sg13g2_fill_1 FILLER_4_1607 ();
 sg13g2_fill_1 FILLER_4_1674 ();
 sg13g2_decap_4 FILLER_4_1685 ();
 sg13g2_fill_2 FILLER_4_1689 ();
 sg13g2_fill_2 FILLER_4_1706 ();
 sg13g2_fill_2 FILLER_4_1717 ();
 sg13g2_decap_4 FILLER_4_1728 ();
 sg13g2_fill_2 FILLER_4_1737 ();
 sg13g2_decap_4 FILLER_4_1774 ();
 sg13g2_fill_2 FILLER_4_1778 ();
 sg13g2_decap_8 FILLER_4_1838 ();
 sg13g2_decap_4 FILLER_4_1845 ();
 sg13g2_fill_1 FILLER_4_1854 ();
 sg13g2_fill_1 FILLER_4_1864 ();
 sg13g2_decap_8 FILLER_4_1889 ();
 sg13g2_decap_8 FILLER_4_1896 ();
 sg13g2_fill_2 FILLER_4_1903 ();
 sg13g2_fill_1 FILLER_4_1905 ();
 sg13g2_fill_2 FILLER_4_1914 ();
 sg13g2_fill_1 FILLER_4_1916 ();
 sg13g2_decap_8 FILLER_4_1927 ();
 sg13g2_fill_2 FILLER_4_1934 ();
 sg13g2_fill_1 FILLER_4_1936 ();
 sg13g2_decap_4 FILLER_4_1969 ();
 sg13g2_decap_4 FILLER_4_1982 ();
 sg13g2_fill_2 FILLER_4_1986 ();
 sg13g2_decap_8 FILLER_4_1998 ();
 sg13g2_fill_2 FILLER_4_2005 ();
 sg13g2_decap_8 FILLER_4_2031 ();
 sg13g2_fill_1 FILLER_4_2038 ();
 sg13g2_fill_2 FILLER_4_2049 ();
 sg13g2_fill_1 FILLER_4_2056 ();
 sg13g2_decap_4 FILLER_4_2065 ();
 sg13g2_fill_1 FILLER_4_2069 ();
 sg13g2_fill_2 FILLER_4_2078 ();
 sg13g2_decap_4 FILLER_4_2143 ();
 sg13g2_fill_1 FILLER_4_2147 ();
 sg13g2_fill_1 FILLER_4_2160 ();
 sg13g2_decap_8 FILLER_4_2171 ();
 sg13g2_fill_2 FILLER_4_2178 ();
 sg13g2_decap_8 FILLER_4_2197 ();
 sg13g2_decap_8 FILLER_4_2204 ();
 sg13g2_fill_1 FILLER_4_2211 ();
 sg13g2_decap_8 FILLER_4_2232 ();
 sg13g2_fill_1 FILLER_4_2257 ();
 sg13g2_decap_8 FILLER_4_2289 ();
 sg13g2_fill_2 FILLER_4_2296 ();
 sg13g2_decap_8 FILLER_4_2313 ();
 sg13g2_fill_1 FILLER_4_2320 ();
 sg13g2_fill_1 FILLER_4_2330 ();
 sg13g2_decap_4 FILLER_4_2357 ();
 sg13g2_fill_1 FILLER_4_2361 ();
 sg13g2_decap_4 FILLER_4_2375 ();
 sg13g2_fill_1 FILLER_4_2379 ();
 sg13g2_decap_8 FILLER_4_2385 ();
 sg13g2_decap_8 FILLER_4_2392 ();
 sg13g2_decap_4 FILLER_4_2399 ();
 sg13g2_decap_8 FILLER_4_2408 ();
 sg13g2_decap_8 FILLER_4_2415 ();
 sg13g2_decap_8 FILLER_4_2422 ();
 sg13g2_decap_4 FILLER_4_2429 ();
 sg13g2_fill_1 FILLER_4_2433 ();
 sg13g2_fill_2 FILLER_4_2443 ();
 sg13g2_fill_1 FILLER_4_2445 ();
 sg13g2_decap_8 FILLER_4_2451 ();
 sg13g2_fill_1 FILLER_4_2458 ();
 sg13g2_decap_4 FILLER_4_2464 ();
 sg13g2_fill_2 FILLER_4_2490 ();
 sg13g2_fill_1 FILLER_4_2492 ();
 sg13g2_decap_8 FILLER_4_2502 ();
 sg13g2_fill_2 FILLER_4_2509 ();
 sg13g2_fill_1 FILLER_4_2511 ();
 sg13g2_fill_1 FILLER_4_2540 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_fill_1 FILLER_4_2577 ();
 sg13g2_decap_8 FILLER_4_2597 ();
 sg13g2_decap_8 FILLER_4_2604 ();
 sg13g2_decap_8 FILLER_4_2611 ();
 sg13g2_decap_8 FILLER_4_2618 ();
 sg13g2_fill_1 FILLER_4_2625 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_4 FILLER_4_2644 ();
 sg13g2_fill_1 FILLER_4_2648 ();
 sg13g2_fill_1 FILLER_4_2656 ();
 sg13g2_fill_2 FILLER_4_2684 ();
 sg13g2_fill_1 FILLER_4_2686 ();
 sg13g2_fill_2 FILLER_4_2694 ();
 sg13g2_fill_1 FILLER_4_2696 ();
 sg13g2_decap_8 FILLER_4_2705 ();
 sg13g2_decap_8 FILLER_4_2712 ();
 sg13g2_fill_2 FILLER_4_2719 ();
 sg13g2_fill_1 FILLER_4_2721 ();
 sg13g2_decap_8 FILLER_4_2735 ();
 sg13g2_decap_8 FILLER_4_2767 ();
 sg13g2_decap_4 FILLER_4_2774 ();
 sg13g2_fill_1 FILLER_4_2790 ();
 sg13g2_decap_8 FILLER_4_2820 ();
 sg13g2_fill_2 FILLER_4_2827 ();
 sg13g2_decap_4 FILLER_4_2859 ();
 sg13g2_fill_1 FILLER_4_2868 ();
 sg13g2_decap_4 FILLER_4_2873 ();
 sg13g2_fill_1 FILLER_4_2877 ();
 sg13g2_decap_4 FILLER_4_2903 ();
 sg13g2_fill_1 FILLER_4_2907 ();
 sg13g2_decap_8 FILLER_4_2920 ();
 sg13g2_decap_8 FILLER_4_2927 ();
 sg13g2_fill_2 FILLER_4_2934 ();
 sg13g2_fill_1 FILLER_4_2936 ();
 sg13g2_decap_8 FILLER_4_2954 ();
 sg13g2_fill_2 FILLER_4_2961 ();
 sg13g2_fill_1 FILLER_4_2963 ();
 sg13g2_decap_8 FILLER_4_2990 ();
 sg13g2_fill_2 FILLER_4_2997 ();
 sg13g2_fill_1 FILLER_4_2999 ();
 sg13g2_decap_8 FILLER_4_3004 ();
 sg13g2_decap_8 FILLER_4_3011 ();
 sg13g2_decap_8 FILLER_4_3018 ();
 sg13g2_decap_8 FILLER_4_3025 ();
 sg13g2_decap_8 FILLER_4_3032 ();
 sg13g2_decap_8 FILLER_4_3039 ();
 sg13g2_decap_8 FILLER_4_3046 ();
 sg13g2_decap_8 FILLER_4_3053 ();
 sg13g2_decap_8 FILLER_4_3060 ();
 sg13g2_decap_8 FILLER_4_3067 ();
 sg13g2_decap_8 FILLER_4_3074 ();
 sg13g2_decap_8 FILLER_4_3081 ();
 sg13g2_decap_8 FILLER_4_3088 ();
 sg13g2_decap_8 FILLER_4_3095 ();
 sg13g2_decap_8 FILLER_4_3102 ();
 sg13g2_decap_8 FILLER_4_3109 ();
 sg13g2_decap_8 FILLER_4_3116 ();
 sg13g2_decap_8 FILLER_4_3123 ();
 sg13g2_decap_8 FILLER_4_3130 ();
 sg13g2_decap_8 FILLER_4_3137 ();
 sg13g2_decap_8 FILLER_4_3144 ();
 sg13g2_decap_8 FILLER_4_3151 ();
 sg13g2_decap_8 FILLER_4_3158 ();
 sg13g2_decap_8 FILLER_4_3165 ();
 sg13g2_decap_8 FILLER_4_3172 ();
 sg13g2_decap_8 FILLER_4_3179 ();
 sg13g2_decap_8 FILLER_4_3186 ();
 sg13g2_decap_8 FILLER_4_3193 ();
 sg13g2_decap_8 FILLER_4_3200 ();
 sg13g2_decap_8 FILLER_4_3207 ();
 sg13g2_decap_8 FILLER_4_3214 ();
 sg13g2_decap_8 FILLER_4_3221 ();
 sg13g2_decap_8 FILLER_4_3228 ();
 sg13g2_decap_8 FILLER_4_3235 ();
 sg13g2_decap_8 FILLER_4_3242 ();
 sg13g2_decap_8 FILLER_4_3249 ();
 sg13g2_decap_8 FILLER_4_3256 ();
 sg13g2_decap_8 FILLER_4_3263 ();
 sg13g2_decap_8 FILLER_4_3270 ();
 sg13g2_decap_8 FILLER_4_3277 ();
 sg13g2_decap_8 FILLER_4_3284 ();
 sg13g2_decap_8 FILLER_4_3291 ();
 sg13g2_decap_8 FILLER_4_3298 ();
 sg13g2_decap_8 FILLER_4_3305 ();
 sg13g2_decap_8 FILLER_4_3312 ();
 sg13g2_decap_8 FILLER_4_3319 ();
 sg13g2_decap_8 FILLER_4_3326 ();
 sg13g2_decap_8 FILLER_4_3333 ();
 sg13g2_decap_8 FILLER_4_3340 ();
 sg13g2_decap_8 FILLER_4_3347 ();
 sg13g2_decap_8 FILLER_4_3354 ();
 sg13g2_decap_8 FILLER_4_3361 ();
 sg13g2_decap_8 FILLER_4_3368 ();
 sg13g2_decap_8 FILLER_4_3375 ();
 sg13g2_decap_8 FILLER_4_3382 ();
 sg13g2_decap_8 FILLER_4_3389 ();
 sg13g2_decap_8 FILLER_4_3396 ();
 sg13g2_decap_8 FILLER_4_3403 ();
 sg13g2_decap_8 FILLER_4_3410 ();
 sg13g2_decap_8 FILLER_4_3417 ();
 sg13g2_decap_8 FILLER_4_3424 ();
 sg13g2_decap_8 FILLER_4_3431 ();
 sg13g2_decap_8 FILLER_4_3438 ();
 sg13g2_decap_8 FILLER_4_3445 ();
 sg13g2_decap_8 FILLER_4_3452 ();
 sg13g2_decap_8 FILLER_4_3459 ();
 sg13g2_decap_8 FILLER_4_3466 ();
 sg13g2_decap_8 FILLER_4_3473 ();
 sg13g2_decap_8 FILLER_4_3480 ();
 sg13g2_decap_8 FILLER_4_3487 ();
 sg13g2_decap_8 FILLER_4_3494 ();
 sg13g2_decap_8 FILLER_4_3501 ();
 sg13g2_decap_8 FILLER_4_3508 ();
 sg13g2_decap_8 FILLER_4_3515 ();
 sg13g2_decap_8 FILLER_4_3522 ();
 sg13g2_decap_8 FILLER_4_3529 ();
 sg13g2_decap_8 FILLER_4_3536 ();
 sg13g2_decap_8 FILLER_4_3543 ();
 sg13g2_decap_8 FILLER_4_3550 ();
 sg13g2_decap_8 FILLER_4_3557 ();
 sg13g2_decap_8 FILLER_4_3564 ();
 sg13g2_decap_8 FILLER_4_3571 ();
 sg13g2_fill_2 FILLER_4_3578 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_fill_1 FILLER_5_473 ();
 sg13g2_decap_4 FILLER_5_482 ();
 sg13g2_fill_2 FILLER_5_486 ();
 sg13g2_fill_2 FILLER_5_493 ();
 sg13g2_fill_1 FILLER_5_495 ();
 sg13g2_decap_4 FILLER_5_503 ();
 sg13g2_fill_1 FILLER_5_507 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_1 FILLER_5_523 ();
 sg13g2_fill_2 FILLER_5_532 ();
 sg13g2_fill_1 FILLER_5_534 ();
 sg13g2_fill_2 FILLER_5_551 ();
 sg13g2_fill_2 FILLER_5_565 ();
 sg13g2_fill_1 FILLER_5_583 ();
 sg13g2_fill_1 FILLER_5_589 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_fill_1 FILLER_5_623 ();
 sg13g2_fill_2 FILLER_5_638 ();
 sg13g2_decap_4 FILLER_5_656 ();
 sg13g2_fill_1 FILLER_5_660 ();
 sg13g2_decap_4 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_fill_2 FILLER_5_725 ();
 sg13g2_fill_1 FILLER_5_727 ();
 sg13g2_fill_2 FILLER_5_760 ();
 sg13g2_fill_1 FILLER_5_762 ();
 sg13g2_fill_1 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_778 ();
 sg13g2_fill_2 FILLER_5_785 ();
 sg13g2_fill_2 FILLER_5_800 ();
 sg13g2_decap_4 FILLER_5_822 ();
 sg13g2_fill_1 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_fill_2 FILLER_5_878 ();
 sg13g2_fill_1 FILLER_5_893 ();
 sg13g2_fill_1 FILLER_5_922 ();
 sg13g2_fill_1 FILLER_5_928 ();
 sg13g2_fill_1 FILLER_5_947 ();
 sg13g2_decap_4 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_960 ();
 sg13g2_decap_4 FILLER_5_967 ();
 sg13g2_fill_1 FILLER_5_971 ();
 sg13g2_decap_4 FILLER_5_990 ();
 sg13g2_decap_4 FILLER_5_998 ();
 sg13g2_fill_2 FILLER_5_1017 ();
 sg13g2_fill_1 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1055 ();
 sg13g2_decap_4 FILLER_5_1133 ();
 sg13g2_fill_2 FILLER_5_1137 ();
 sg13g2_fill_2 FILLER_5_1160 ();
 sg13g2_fill_1 FILLER_5_1162 ();
 sg13g2_decap_8 FILLER_5_1167 ();
 sg13g2_decap_8 FILLER_5_1174 ();
 sg13g2_fill_1 FILLER_5_1186 ();
 sg13g2_decap_4 FILLER_5_1204 ();
 sg13g2_decap_8 FILLER_5_1213 ();
 sg13g2_decap_4 FILLER_5_1220 ();
 sg13g2_fill_1 FILLER_5_1224 ();
 sg13g2_fill_2 FILLER_5_1237 ();
 sg13g2_fill_1 FILLER_5_1239 ();
 sg13g2_fill_1 FILLER_5_1259 ();
 sg13g2_decap_8 FILLER_5_1269 ();
 sg13g2_decap_8 FILLER_5_1276 ();
 sg13g2_fill_2 FILLER_5_1296 ();
 sg13g2_fill_1 FILLER_5_1298 ();
 sg13g2_fill_1 FILLER_5_1309 ();
 sg13g2_decap_4 FILLER_5_1334 ();
 sg13g2_fill_1 FILLER_5_1338 ();
 sg13g2_decap_8 FILLER_5_1342 ();
 sg13g2_decap_4 FILLER_5_1349 ();
 sg13g2_fill_2 FILLER_5_1353 ();
 sg13g2_decap_8 FILLER_5_1363 ();
 sg13g2_decap_4 FILLER_5_1370 ();
 sg13g2_fill_2 FILLER_5_1374 ();
 sg13g2_decap_8 FILLER_5_1398 ();
 sg13g2_fill_2 FILLER_5_1405 ();
 sg13g2_decap_4 FILLER_5_1416 ();
 sg13g2_fill_2 FILLER_5_1433 ();
 sg13g2_fill_1 FILLER_5_1435 ();
 sg13g2_decap_8 FILLER_5_1471 ();
 sg13g2_fill_1 FILLER_5_1478 ();
 sg13g2_fill_2 FILLER_5_1520 ();
 sg13g2_decap_4 FILLER_5_1531 ();
 sg13g2_fill_2 FILLER_5_1542 ();
 sg13g2_fill_1 FILLER_5_1544 ();
 sg13g2_decap_8 FILLER_5_1563 ();
 sg13g2_decap_8 FILLER_5_1570 ();
 sg13g2_fill_2 FILLER_5_1577 ();
 sg13g2_decap_8 FILLER_5_1592 ();
 sg13g2_decap_4 FILLER_5_1607 ();
 sg13g2_fill_2 FILLER_5_1616 ();
 sg13g2_fill_1 FILLER_5_1618 ();
 sg13g2_decap_8 FILLER_5_1637 ();
 sg13g2_fill_1 FILLER_5_1644 ();
 sg13g2_decap_4 FILLER_5_1666 ();
 sg13g2_fill_2 FILLER_5_1670 ();
 sg13g2_decap_4 FILLER_5_1690 ();
 sg13g2_fill_2 FILLER_5_1694 ();
 sg13g2_fill_2 FILLER_5_1733 ();
 sg13g2_fill_1 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1746 ();
 sg13g2_decap_8 FILLER_5_1753 ();
 sg13g2_decap_4 FILLER_5_1760 ();
 sg13g2_fill_2 FILLER_5_1764 ();
 sg13g2_decap_8 FILLER_5_1770 ();
 sg13g2_decap_8 FILLER_5_1777 ();
 sg13g2_fill_2 FILLER_5_1784 ();
 sg13g2_fill_2 FILLER_5_1790 ();
 sg13g2_decap_4 FILLER_5_1842 ();
 sg13g2_fill_2 FILLER_5_1846 ();
 sg13g2_fill_2 FILLER_5_1860 ();
 sg13g2_fill_1 FILLER_5_1880 ();
 sg13g2_decap_8 FILLER_5_1885 ();
 sg13g2_decap_4 FILLER_5_1892 ();
 sg13g2_decap_4 FILLER_5_1938 ();
 sg13g2_fill_2 FILLER_5_1942 ();
 sg13g2_fill_2 FILLER_5_1949 ();
 sg13g2_fill_1 FILLER_5_1951 ();
 sg13g2_decap_8 FILLER_5_1963 ();
 sg13g2_fill_2 FILLER_5_1970 ();
 sg13g2_fill_1 FILLER_5_1972 ();
 sg13g2_fill_2 FILLER_5_1986 ();
 sg13g2_decap_4 FILLER_5_2008 ();
 sg13g2_fill_1 FILLER_5_2022 ();
 sg13g2_decap_8 FILLER_5_2033 ();
 sg13g2_fill_2 FILLER_5_2040 ();
 sg13g2_fill_1 FILLER_5_2042 ();
 sg13g2_fill_1 FILLER_5_2059 ();
 sg13g2_decap_4 FILLER_5_2086 ();
 sg13g2_fill_2 FILLER_5_2090 ();
 sg13g2_decap_8 FILLER_5_2105 ();
 sg13g2_fill_1 FILLER_5_2112 ();
 sg13g2_fill_1 FILLER_5_2118 ();
 sg13g2_decap_8 FILLER_5_2127 ();
 sg13g2_fill_1 FILLER_5_2143 ();
 sg13g2_fill_1 FILLER_5_2157 ();
 sg13g2_decap_4 FILLER_5_2176 ();
 sg13g2_fill_2 FILLER_5_2180 ();
 sg13g2_fill_2 FILLER_5_2211 ();
 sg13g2_fill_1 FILLER_5_2213 ();
 sg13g2_decap_4 FILLER_5_2222 ();
 sg13g2_fill_2 FILLER_5_2239 ();
 sg13g2_decap_8 FILLER_5_2252 ();
 sg13g2_decap_4 FILLER_5_2259 ();
 sg13g2_fill_2 FILLER_5_2263 ();
 sg13g2_decap_8 FILLER_5_2285 ();
 sg13g2_decap_8 FILLER_5_2320 ();
 sg13g2_fill_2 FILLER_5_2327 ();
 sg13g2_fill_2 FILLER_5_2355 ();
 sg13g2_decap_8 FILLER_5_2379 ();
 sg13g2_fill_2 FILLER_5_2386 ();
 sg13g2_fill_2 FILLER_5_2398 ();
 sg13g2_decap_8 FILLER_5_2412 ();
 sg13g2_fill_1 FILLER_5_2419 ();
 sg13g2_fill_2 FILLER_5_2433 ();
 sg13g2_fill_1 FILLER_5_2435 ();
 sg13g2_fill_2 FILLER_5_2440 ();
 sg13g2_fill_2 FILLER_5_2454 ();
 sg13g2_fill_1 FILLER_5_2456 ();
 sg13g2_fill_1 FILLER_5_2463 ();
 sg13g2_decap_8 FILLER_5_2479 ();
 sg13g2_decap_4 FILLER_5_2509 ();
 sg13g2_fill_2 FILLER_5_2517 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_fill_1 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2557 ();
 sg13g2_fill_1 FILLER_5_2564 ();
 sg13g2_fill_2 FILLER_5_2571 ();
 sg13g2_fill_2 FILLER_5_2619 ();
 sg13g2_fill_1 FILLER_5_2621 ();
 sg13g2_decap_8 FILLER_5_2635 ();
 sg13g2_decap_8 FILLER_5_2642 ();
 sg13g2_fill_2 FILLER_5_2664 ();
 sg13g2_fill_1 FILLER_5_2683 ();
 sg13g2_decap_8 FILLER_5_2700 ();
 sg13g2_fill_2 FILLER_5_2707 ();
 sg13g2_decap_8 FILLER_5_2714 ();
 sg13g2_fill_2 FILLER_5_2721 ();
 sg13g2_fill_1 FILLER_5_2723 ();
 sg13g2_decap_4 FILLER_5_2737 ();
 sg13g2_fill_2 FILLER_5_2751 ();
 sg13g2_fill_1 FILLER_5_2753 ();
 sg13g2_fill_2 FILLER_5_2770 ();
 sg13g2_fill_1 FILLER_5_2795 ();
 sg13g2_fill_2 FILLER_5_2804 ();
 sg13g2_fill_1 FILLER_5_2806 ();
 sg13g2_decap_8 FILLER_5_2819 ();
 sg13g2_decap_4 FILLER_5_2845 ();
 sg13g2_fill_1 FILLER_5_2849 ();
 sg13g2_decap_4 FILLER_5_2863 ();
 sg13g2_fill_2 FILLER_5_2867 ();
 sg13g2_decap_4 FILLER_5_2882 ();
 sg13g2_fill_2 FILLER_5_2886 ();
 sg13g2_decap_8 FILLER_5_2897 ();
 sg13g2_decap_8 FILLER_5_2904 ();
 sg13g2_decap_4 FILLER_5_2911 ();
 sg13g2_decap_4 FILLER_5_2923 ();
 sg13g2_fill_2 FILLER_5_2927 ();
 sg13g2_fill_2 FILLER_5_2936 ();
 sg13g2_fill_1 FILLER_5_2938 ();
 sg13g2_fill_1 FILLER_5_2958 ();
 sg13g2_fill_1 FILLER_5_2972 ();
 sg13g2_fill_1 FILLER_5_2987 ();
 sg13g2_decap_8 FILLER_5_3023 ();
 sg13g2_decap_8 FILLER_5_3030 ();
 sg13g2_decap_8 FILLER_5_3037 ();
 sg13g2_decap_8 FILLER_5_3044 ();
 sg13g2_decap_8 FILLER_5_3051 ();
 sg13g2_decap_8 FILLER_5_3058 ();
 sg13g2_decap_8 FILLER_5_3065 ();
 sg13g2_decap_8 FILLER_5_3072 ();
 sg13g2_decap_8 FILLER_5_3079 ();
 sg13g2_decap_8 FILLER_5_3086 ();
 sg13g2_decap_8 FILLER_5_3093 ();
 sg13g2_decap_8 FILLER_5_3100 ();
 sg13g2_decap_8 FILLER_5_3107 ();
 sg13g2_decap_8 FILLER_5_3114 ();
 sg13g2_decap_8 FILLER_5_3121 ();
 sg13g2_decap_8 FILLER_5_3128 ();
 sg13g2_decap_8 FILLER_5_3135 ();
 sg13g2_decap_8 FILLER_5_3142 ();
 sg13g2_decap_8 FILLER_5_3149 ();
 sg13g2_decap_8 FILLER_5_3156 ();
 sg13g2_decap_8 FILLER_5_3163 ();
 sg13g2_decap_8 FILLER_5_3170 ();
 sg13g2_decap_8 FILLER_5_3177 ();
 sg13g2_decap_8 FILLER_5_3184 ();
 sg13g2_decap_8 FILLER_5_3191 ();
 sg13g2_decap_8 FILLER_5_3198 ();
 sg13g2_decap_8 FILLER_5_3205 ();
 sg13g2_decap_8 FILLER_5_3212 ();
 sg13g2_decap_8 FILLER_5_3219 ();
 sg13g2_decap_8 FILLER_5_3226 ();
 sg13g2_decap_8 FILLER_5_3233 ();
 sg13g2_decap_8 FILLER_5_3240 ();
 sg13g2_decap_8 FILLER_5_3247 ();
 sg13g2_decap_8 FILLER_5_3254 ();
 sg13g2_decap_8 FILLER_5_3261 ();
 sg13g2_decap_8 FILLER_5_3268 ();
 sg13g2_decap_8 FILLER_5_3275 ();
 sg13g2_decap_8 FILLER_5_3282 ();
 sg13g2_decap_8 FILLER_5_3289 ();
 sg13g2_decap_8 FILLER_5_3296 ();
 sg13g2_decap_8 FILLER_5_3303 ();
 sg13g2_decap_8 FILLER_5_3310 ();
 sg13g2_decap_8 FILLER_5_3317 ();
 sg13g2_decap_8 FILLER_5_3324 ();
 sg13g2_decap_8 FILLER_5_3331 ();
 sg13g2_decap_8 FILLER_5_3338 ();
 sg13g2_decap_8 FILLER_5_3345 ();
 sg13g2_decap_8 FILLER_5_3352 ();
 sg13g2_decap_8 FILLER_5_3359 ();
 sg13g2_decap_8 FILLER_5_3366 ();
 sg13g2_decap_8 FILLER_5_3373 ();
 sg13g2_decap_8 FILLER_5_3380 ();
 sg13g2_decap_8 FILLER_5_3387 ();
 sg13g2_decap_8 FILLER_5_3394 ();
 sg13g2_decap_8 FILLER_5_3401 ();
 sg13g2_decap_8 FILLER_5_3408 ();
 sg13g2_decap_8 FILLER_5_3415 ();
 sg13g2_decap_8 FILLER_5_3422 ();
 sg13g2_decap_8 FILLER_5_3429 ();
 sg13g2_decap_8 FILLER_5_3436 ();
 sg13g2_decap_8 FILLER_5_3443 ();
 sg13g2_decap_8 FILLER_5_3450 ();
 sg13g2_decap_8 FILLER_5_3457 ();
 sg13g2_decap_8 FILLER_5_3464 ();
 sg13g2_decap_8 FILLER_5_3471 ();
 sg13g2_decap_8 FILLER_5_3478 ();
 sg13g2_decap_8 FILLER_5_3485 ();
 sg13g2_decap_8 FILLER_5_3492 ();
 sg13g2_decap_8 FILLER_5_3499 ();
 sg13g2_decap_8 FILLER_5_3506 ();
 sg13g2_decap_8 FILLER_5_3513 ();
 sg13g2_decap_8 FILLER_5_3520 ();
 sg13g2_decap_8 FILLER_5_3527 ();
 sg13g2_decap_8 FILLER_5_3534 ();
 sg13g2_decap_8 FILLER_5_3541 ();
 sg13g2_decap_8 FILLER_5_3548 ();
 sg13g2_decap_8 FILLER_5_3555 ();
 sg13g2_decap_8 FILLER_5_3562 ();
 sg13g2_decap_8 FILLER_5_3569 ();
 sg13g2_decap_4 FILLER_5_3576 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_4 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_6_414 ();
 sg13g2_fill_2 FILLER_6_420 ();
 sg13g2_fill_1 FILLER_6_422 ();
 sg13g2_fill_2 FILLER_6_436 ();
 sg13g2_fill_2 FILLER_6_455 ();
 sg13g2_fill_2 FILLER_6_462 ();
 sg13g2_fill_1 FILLER_6_481 ();
 sg13g2_fill_1 FILLER_6_523 ();
 sg13g2_fill_1 FILLER_6_564 ();
 sg13g2_fill_1 FILLER_6_570 ();
 sg13g2_decap_8 FILLER_6_576 ();
 sg13g2_decap_8 FILLER_6_583 ();
 sg13g2_decap_8 FILLER_6_590 ();
 sg13g2_decap_8 FILLER_6_597 ();
 sg13g2_fill_1 FILLER_6_604 ();
 sg13g2_decap_4 FILLER_6_618 ();
 sg13g2_fill_2 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_629 ();
 sg13g2_fill_1 FILLER_6_640 ();
 sg13g2_decap_4 FILLER_6_644 ();
 sg13g2_fill_2 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_664 ();
 sg13g2_decap_8 FILLER_6_675 ();
 sg13g2_decap_8 FILLER_6_682 ();
 sg13g2_decap_8 FILLER_6_689 ();
 sg13g2_decap_8 FILLER_6_696 ();
 sg13g2_decap_4 FILLER_6_707 ();
 sg13g2_fill_2 FILLER_6_711 ();
 sg13g2_fill_1 FILLER_6_733 ();
 sg13g2_fill_2 FILLER_6_751 ();
 sg13g2_decap_8 FILLER_6_771 ();
 sg13g2_fill_1 FILLER_6_778 ();
 sg13g2_fill_2 FILLER_6_784 ();
 sg13g2_fill_2 FILLER_6_796 ();
 sg13g2_fill_1 FILLER_6_798 ();
 sg13g2_fill_2 FILLER_6_807 ();
 sg13g2_decap_8 FILLER_6_822 ();
 sg13g2_decap_4 FILLER_6_829 ();
 sg13g2_fill_2 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_856 ();
 sg13g2_decap_8 FILLER_6_863 ();
 sg13g2_fill_2 FILLER_6_870 ();
 sg13g2_fill_1 FILLER_6_872 ();
 sg13g2_decap_4 FILLER_6_895 ();
 sg13g2_decap_4 FILLER_6_904 ();
 sg13g2_fill_1 FILLER_6_913 ();
 sg13g2_fill_1 FILLER_6_927 ();
 sg13g2_fill_2 FILLER_6_946 ();
 sg13g2_fill_1 FILLER_6_965 ();
 sg13g2_fill_2 FILLER_6_987 ();
 sg13g2_fill_2 FILLER_6_1007 ();
 sg13g2_fill_2 FILLER_6_1018 ();
 sg13g2_fill_1 FILLER_6_1020 ();
 sg13g2_fill_1 FILLER_6_1024 ();
 sg13g2_decap_8 FILLER_6_1029 ();
 sg13g2_fill_2 FILLER_6_1036 ();
 sg13g2_fill_1 FILLER_6_1051 ();
 sg13g2_decap_8 FILLER_6_1086 ();
 sg13g2_decap_8 FILLER_6_1093 ();
 sg13g2_decap_4 FILLER_6_1104 ();
 sg13g2_decap_8 FILLER_6_1111 ();
 sg13g2_decap_8 FILLER_6_1118 ();
 sg13g2_fill_2 FILLER_6_1125 ();
 sg13g2_fill_2 FILLER_6_1155 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_fill_2 FILLER_6_1177 ();
 sg13g2_fill_1 FILLER_6_1179 ();
 sg13g2_decap_8 FILLER_6_1201 ();
 sg13g2_decap_4 FILLER_6_1208 ();
 sg13g2_fill_2 FILLER_6_1212 ();
 sg13g2_fill_2 FILLER_6_1222 ();
 sg13g2_fill_2 FILLER_6_1269 ();
 sg13g2_decap_8 FILLER_6_1309 ();
 sg13g2_fill_1 FILLER_6_1316 ();
 sg13g2_fill_1 FILLER_6_1322 ();
 sg13g2_decap_8 FILLER_6_1344 ();
 sg13g2_fill_2 FILLER_6_1351 ();
 sg13g2_fill_1 FILLER_6_1353 ();
 sg13g2_fill_2 FILLER_6_1374 ();
 sg13g2_fill_1 FILLER_6_1376 ();
 sg13g2_fill_2 FILLER_6_1414 ();
 sg13g2_fill_1 FILLER_6_1416 ();
 sg13g2_decap_4 FILLER_6_1441 ();
 sg13g2_fill_2 FILLER_6_1445 ();
 sg13g2_fill_1 FILLER_6_1452 ();
 sg13g2_fill_1 FILLER_6_1463 ();
 sg13g2_fill_1 FILLER_6_1469 ();
 sg13g2_fill_1 FILLER_6_1482 ();
 sg13g2_decap_8 FILLER_6_1492 ();
 sg13g2_decap_4 FILLER_6_1499 ();
 sg13g2_fill_2 FILLER_6_1503 ();
 sg13g2_fill_1 FILLER_6_1520 ();
 sg13g2_decap_4 FILLER_6_1545 ();
 sg13g2_fill_1 FILLER_6_1549 ();
 sg13g2_fill_2 FILLER_6_1559 ();
 sg13g2_fill_1 FILLER_6_1561 ();
 sg13g2_decap_8 FILLER_6_1581 ();
 sg13g2_decap_8 FILLER_6_1623 ();
 sg13g2_decap_8 FILLER_6_1630 ();
 sg13g2_decap_4 FILLER_6_1637 ();
 sg13g2_fill_1 FILLER_6_1641 ();
 sg13g2_fill_1 FILLER_6_1655 ();
 sg13g2_fill_2 FILLER_6_1666 ();
 sg13g2_decap_8 FILLER_6_1673 ();
 sg13g2_fill_2 FILLER_6_1685 ();
 sg13g2_fill_1 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1697 ();
 sg13g2_decap_4 FILLER_6_1704 ();
 sg13g2_fill_2 FILLER_6_1718 ();
 sg13g2_fill_2 FILLER_6_1751 ();
 sg13g2_decap_4 FILLER_6_1828 ();
 sg13g2_fill_2 FILLER_6_1832 ();
 sg13g2_decap_4 FILLER_6_1839 ();
 sg13g2_fill_2 FILLER_6_1865 ();
 sg13g2_fill_1 FILLER_6_1867 ();
 sg13g2_fill_2 FILLER_6_1872 ();
 sg13g2_fill_1 FILLER_6_1874 ();
 sg13g2_decap_8 FILLER_6_1891 ();
 sg13g2_fill_1 FILLER_6_1898 ();
 sg13g2_fill_1 FILLER_6_1904 ();
 sg13g2_decap_4 FILLER_6_1910 ();
 sg13g2_fill_1 FILLER_6_1927 ();
 sg13g2_fill_2 FILLER_6_1956 ();
 sg13g2_decap_4 FILLER_6_1976 ();
 sg13g2_decap_8 FILLER_6_1985 ();
 sg13g2_decap_4 FILLER_6_2018 ();
 sg13g2_fill_1 FILLER_6_2022 ();
 sg13g2_decap_4 FILLER_6_2036 ();
 sg13g2_fill_1 FILLER_6_2040 ();
 sg13g2_decap_8 FILLER_6_2055 ();
 sg13g2_fill_2 FILLER_6_2065 ();
 sg13g2_fill_1 FILLER_6_2067 ();
 sg13g2_decap_8 FILLER_6_2078 ();
 sg13g2_decap_8 FILLER_6_2085 ();
 sg13g2_decap_4 FILLER_6_2092 ();
 sg13g2_fill_1 FILLER_6_2096 ();
 sg13g2_decap_4 FILLER_6_2122 ();
 sg13g2_decap_8 FILLER_6_2136 ();
 sg13g2_fill_2 FILLER_6_2151 ();
 sg13g2_decap_4 FILLER_6_2176 ();
 sg13g2_fill_2 FILLER_6_2180 ();
 sg13g2_decap_8 FILLER_6_2196 ();
 sg13g2_decap_8 FILLER_6_2203 ();
 sg13g2_decap_4 FILLER_6_2210 ();
 sg13g2_fill_2 FILLER_6_2219 ();
 sg13g2_fill_1 FILLER_6_2221 ();
 sg13g2_decap_8 FILLER_6_2241 ();
 sg13g2_fill_1 FILLER_6_2248 ();
 sg13g2_decap_8 FILLER_6_2262 ();
 sg13g2_fill_2 FILLER_6_2269 ();
 sg13g2_decap_8 FILLER_6_2288 ();
 sg13g2_fill_2 FILLER_6_2295 ();
 sg13g2_decap_8 FILLER_6_2315 ();
 sg13g2_decap_8 FILLER_6_2322 ();
 sg13g2_decap_4 FILLER_6_2329 ();
 sg13g2_fill_2 FILLER_6_2341 ();
 sg13g2_fill_1 FILLER_6_2343 ();
 sg13g2_decap_8 FILLER_6_2352 ();
 sg13g2_decap_4 FILLER_6_2382 ();
 sg13g2_fill_2 FILLER_6_2386 ();
 sg13g2_fill_2 FILLER_6_2393 ();
 sg13g2_fill_1 FILLER_6_2432 ();
 sg13g2_decap_8 FILLER_6_2450 ();
 sg13g2_fill_2 FILLER_6_2457 ();
 sg13g2_fill_2 FILLER_6_2466 ();
 sg13g2_decap_4 FILLER_6_2485 ();
 sg13g2_decap_8 FILLER_6_2498 ();
 sg13g2_fill_2 FILLER_6_2505 ();
 sg13g2_fill_2 FILLER_6_2517 ();
 sg13g2_decap_8 FILLER_6_2524 ();
 sg13g2_decap_8 FILLER_6_2531 ();
 sg13g2_decap_4 FILLER_6_2538 ();
 sg13g2_fill_1 FILLER_6_2542 ();
 sg13g2_fill_1 FILLER_6_2548 ();
 sg13g2_fill_1 FILLER_6_2559 ();
 sg13g2_fill_2 FILLER_6_2569 ();
 sg13g2_decap_8 FILLER_6_2609 ();
 sg13g2_fill_2 FILLER_6_2674 ();
 sg13g2_fill_1 FILLER_6_2676 ();
 sg13g2_decap_8 FILLER_6_2688 ();
 sg13g2_fill_2 FILLER_6_2695 ();
 sg13g2_fill_1 FILLER_6_2705 ();
 sg13g2_decap_8 FILLER_6_2717 ();
 sg13g2_decap_8 FILLER_6_2724 ();
 sg13g2_decap_4 FILLER_6_2768 ();
 sg13g2_fill_2 FILLER_6_2772 ();
 sg13g2_decap_8 FILLER_6_2781 ();
 sg13g2_decap_4 FILLER_6_2793 ();
 sg13g2_fill_1 FILLER_6_2797 ();
 sg13g2_decap_8 FILLER_6_2816 ();
 sg13g2_decap_8 FILLER_6_2823 ();
 sg13g2_fill_2 FILLER_6_2830 ();
 sg13g2_fill_1 FILLER_6_2832 ();
 sg13g2_fill_2 FILLER_6_2837 ();
 sg13g2_fill_1 FILLER_6_2844 ();
 sg13g2_fill_1 FILLER_6_2873 ();
 sg13g2_fill_2 FILLER_6_2894 ();
 sg13g2_decap_8 FILLER_6_2901 ();
 sg13g2_decap_8 FILLER_6_2939 ();
 sg13g2_decap_4 FILLER_6_2946 ();
 sg13g2_decap_8 FILLER_6_2954 ();
 sg13g2_decap_4 FILLER_6_2961 ();
 sg13g2_fill_2 FILLER_6_2969 ();
 sg13g2_fill_1 FILLER_6_2984 ();
 sg13g2_decap_8 FILLER_6_3005 ();
 sg13g2_decap_8 FILLER_6_3012 ();
 sg13g2_decap_8 FILLER_6_3019 ();
 sg13g2_decap_8 FILLER_6_3026 ();
 sg13g2_decap_8 FILLER_6_3033 ();
 sg13g2_decap_8 FILLER_6_3040 ();
 sg13g2_decap_8 FILLER_6_3047 ();
 sg13g2_decap_8 FILLER_6_3054 ();
 sg13g2_decap_8 FILLER_6_3061 ();
 sg13g2_decap_8 FILLER_6_3068 ();
 sg13g2_decap_8 FILLER_6_3075 ();
 sg13g2_decap_8 FILLER_6_3082 ();
 sg13g2_decap_8 FILLER_6_3089 ();
 sg13g2_decap_8 FILLER_6_3096 ();
 sg13g2_decap_8 FILLER_6_3103 ();
 sg13g2_decap_8 FILLER_6_3110 ();
 sg13g2_decap_8 FILLER_6_3117 ();
 sg13g2_decap_8 FILLER_6_3124 ();
 sg13g2_decap_8 FILLER_6_3131 ();
 sg13g2_decap_8 FILLER_6_3138 ();
 sg13g2_decap_8 FILLER_6_3145 ();
 sg13g2_decap_8 FILLER_6_3152 ();
 sg13g2_decap_8 FILLER_6_3159 ();
 sg13g2_decap_8 FILLER_6_3166 ();
 sg13g2_decap_8 FILLER_6_3173 ();
 sg13g2_decap_8 FILLER_6_3180 ();
 sg13g2_decap_8 FILLER_6_3187 ();
 sg13g2_decap_8 FILLER_6_3194 ();
 sg13g2_decap_8 FILLER_6_3201 ();
 sg13g2_decap_8 FILLER_6_3208 ();
 sg13g2_decap_8 FILLER_6_3215 ();
 sg13g2_decap_8 FILLER_6_3222 ();
 sg13g2_decap_8 FILLER_6_3229 ();
 sg13g2_decap_8 FILLER_6_3236 ();
 sg13g2_decap_8 FILLER_6_3243 ();
 sg13g2_decap_8 FILLER_6_3250 ();
 sg13g2_decap_8 FILLER_6_3257 ();
 sg13g2_decap_8 FILLER_6_3264 ();
 sg13g2_decap_8 FILLER_6_3271 ();
 sg13g2_decap_8 FILLER_6_3278 ();
 sg13g2_decap_8 FILLER_6_3285 ();
 sg13g2_decap_8 FILLER_6_3292 ();
 sg13g2_decap_8 FILLER_6_3299 ();
 sg13g2_decap_8 FILLER_6_3306 ();
 sg13g2_decap_8 FILLER_6_3313 ();
 sg13g2_decap_8 FILLER_6_3320 ();
 sg13g2_decap_8 FILLER_6_3327 ();
 sg13g2_decap_8 FILLER_6_3334 ();
 sg13g2_decap_8 FILLER_6_3341 ();
 sg13g2_decap_8 FILLER_6_3348 ();
 sg13g2_decap_8 FILLER_6_3355 ();
 sg13g2_decap_8 FILLER_6_3362 ();
 sg13g2_decap_8 FILLER_6_3369 ();
 sg13g2_decap_8 FILLER_6_3376 ();
 sg13g2_decap_8 FILLER_6_3383 ();
 sg13g2_decap_8 FILLER_6_3390 ();
 sg13g2_decap_8 FILLER_6_3397 ();
 sg13g2_decap_8 FILLER_6_3404 ();
 sg13g2_decap_8 FILLER_6_3411 ();
 sg13g2_decap_8 FILLER_6_3418 ();
 sg13g2_decap_8 FILLER_6_3425 ();
 sg13g2_decap_8 FILLER_6_3432 ();
 sg13g2_decap_8 FILLER_6_3439 ();
 sg13g2_decap_8 FILLER_6_3446 ();
 sg13g2_decap_8 FILLER_6_3453 ();
 sg13g2_decap_8 FILLER_6_3460 ();
 sg13g2_decap_8 FILLER_6_3467 ();
 sg13g2_decap_8 FILLER_6_3474 ();
 sg13g2_decap_8 FILLER_6_3481 ();
 sg13g2_decap_8 FILLER_6_3488 ();
 sg13g2_decap_8 FILLER_6_3495 ();
 sg13g2_decap_8 FILLER_6_3502 ();
 sg13g2_decap_8 FILLER_6_3509 ();
 sg13g2_decap_8 FILLER_6_3516 ();
 sg13g2_decap_8 FILLER_6_3523 ();
 sg13g2_decap_8 FILLER_6_3530 ();
 sg13g2_decap_8 FILLER_6_3537 ();
 sg13g2_decap_8 FILLER_6_3544 ();
 sg13g2_decap_8 FILLER_6_3551 ();
 sg13g2_decap_8 FILLER_6_3558 ();
 sg13g2_decap_8 FILLER_6_3565 ();
 sg13g2_decap_8 FILLER_6_3572 ();
 sg13g2_fill_1 FILLER_6_3579 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_4 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_347 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_2 FILLER_7_413 ();
 sg13g2_fill_1 FILLER_7_415 ();
 sg13g2_fill_1 FILLER_7_442 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_fill_2 FILLER_7_497 ();
 sg13g2_fill_1 FILLER_7_499 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_fill_2 FILLER_7_511 ();
 sg13g2_fill_1 FILLER_7_513 ();
 sg13g2_fill_1 FILLER_7_529 ();
 sg13g2_decap_8 FILLER_7_535 ();
 sg13g2_fill_2 FILLER_7_542 ();
 sg13g2_decap_4 FILLER_7_553 ();
 sg13g2_decap_4 FILLER_7_562 ();
 sg13g2_decap_4 FILLER_7_580 ();
 sg13g2_fill_2 FILLER_7_584 ();
 sg13g2_decap_8 FILLER_7_597 ();
 sg13g2_decap_4 FILLER_7_638 ();
 sg13g2_fill_1 FILLER_7_642 ();
 sg13g2_decap_4 FILLER_7_654 ();
 sg13g2_fill_2 FILLER_7_658 ();
 sg13g2_fill_1 FILLER_7_664 ();
 sg13g2_fill_2 FILLER_7_693 ();
 sg13g2_fill_1 FILLER_7_695 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_fill_2 FILLER_7_725 ();
 sg13g2_fill_1 FILLER_7_727 ();
 sg13g2_fill_2 FILLER_7_741 ();
 sg13g2_fill_1 FILLER_7_743 ();
 sg13g2_decap_4 FILLER_7_753 ();
 sg13g2_fill_2 FILLER_7_757 ();
 sg13g2_fill_1 FILLER_7_766 ();
 sg13g2_fill_2 FILLER_7_772 ();
 sg13g2_fill_1 FILLER_7_774 ();
 sg13g2_decap_4 FILLER_7_794 ();
 sg13g2_fill_1 FILLER_7_798 ();
 sg13g2_fill_1 FILLER_7_808 ();
 sg13g2_decap_8 FILLER_7_834 ();
 sg13g2_fill_1 FILLER_7_841 ();
 sg13g2_fill_2 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_fill_2 FILLER_7_919 ();
 sg13g2_fill_1 FILLER_7_921 ();
 sg13g2_decap_8 FILLER_7_930 ();
 sg13g2_decap_8 FILLER_7_937 ();
 sg13g2_decap_8 FILLER_7_944 ();
 sg13g2_decap_4 FILLER_7_951 ();
 sg13g2_fill_1 FILLER_7_955 ();
 sg13g2_fill_2 FILLER_7_960 ();
 sg13g2_fill_1 FILLER_7_962 ();
 sg13g2_fill_2 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_991 ();
 sg13g2_fill_1 FILLER_7_998 ();
 sg13g2_fill_2 FILLER_7_1009 ();
 sg13g2_decap_4 FILLER_7_1014 ();
 sg13g2_fill_1 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_fill_1 FILLER_7_1029 ();
 sg13g2_fill_2 FILLER_7_1049 ();
 sg13g2_fill_2 FILLER_7_1064 ();
 sg13g2_fill_1 FILLER_7_1066 ();
 sg13g2_fill_2 FILLER_7_1075 ();
 sg13g2_fill_1 FILLER_7_1077 ();
 sg13g2_fill_1 FILLER_7_1091 ();
 sg13g2_fill_2 FILLER_7_1175 ();
 sg13g2_fill_1 FILLER_7_1177 ();
 sg13g2_fill_2 FILLER_7_1203 ();
 sg13g2_decap_8 FILLER_7_1230 ();
 sg13g2_decap_4 FILLER_7_1237 ();
 sg13g2_decap_8 FILLER_7_1246 ();
 sg13g2_decap_8 FILLER_7_1253 ();
 sg13g2_fill_1 FILLER_7_1260 ();
 sg13g2_decap_4 FILLER_7_1266 ();
 sg13g2_fill_1 FILLER_7_1270 ();
 sg13g2_decap_8 FILLER_7_1276 ();
 sg13g2_decap_4 FILLER_7_1283 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_4 FILLER_7_1309 ();
 sg13g2_fill_2 FILLER_7_1313 ();
 sg13g2_fill_1 FILLER_7_1325 ();
 sg13g2_fill_2 FILLER_7_1331 ();
 sg13g2_decap_8 FILLER_7_1338 ();
 sg13g2_decap_8 FILLER_7_1371 ();
 sg13g2_fill_2 FILLER_7_1378 ();
 sg13g2_fill_1 FILLER_7_1384 ();
 sg13g2_decap_4 FILLER_7_1390 ();
 sg13g2_fill_1 FILLER_7_1394 ();
 sg13g2_fill_2 FILLER_7_1400 ();
 sg13g2_fill_1 FILLER_7_1402 ();
 sg13g2_decap_4 FILLER_7_1408 ();
 sg13g2_fill_2 FILLER_7_1412 ();
 sg13g2_decap_4 FILLER_7_1446 ();
 sg13g2_fill_1 FILLER_7_1450 ();
 sg13g2_decap_8 FILLER_7_1479 ();
 sg13g2_decap_8 FILLER_7_1486 ();
 sg13g2_decap_4 FILLER_7_1493 ();
 sg13g2_fill_2 FILLER_7_1509 ();
 sg13g2_fill_1 FILLER_7_1511 ();
 sg13g2_decap_8 FILLER_7_1542 ();
 sg13g2_fill_2 FILLER_7_1549 ();
 sg13g2_fill_1 FILLER_7_1551 ();
 sg13g2_decap_8 FILLER_7_1566 ();
 sg13g2_fill_2 FILLER_7_1573 ();
 sg13g2_fill_2 FILLER_7_1580 ();
 sg13g2_decap_8 FILLER_7_1591 ();
 sg13g2_fill_1 FILLER_7_1598 ();
 sg13g2_decap_4 FILLER_7_1631 ();
 sg13g2_decap_8 FILLER_7_1665 ();
 sg13g2_fill_1 FILLER_7_1672 ();
 sg13g2_decap_4 FILLER_7_1699 ();
 sg13g2_decap_8 FILLER_7_1713 ();
 sg13g2_decap_4 FILLER_7_1720 ();
 sg13g2_fill_1 FILLER_7_1724 ();
 sg13g2_decap_8 FILLER_7_1748 ();
 sg13g2_decap_4 FILLER_7_1755 ();
 sg13g2_fill_2 FILLER_7_1759 ();
 sg13g2_decap_8 FILLER_7_1774 ();
 sg13g2_fill_2 FILLER_7_1793 ();
 sg13g2_fill_1 FILLER_7_1795 ();
 sg13g2_fill_2 FILLER_7_1813 ();
 sg13g2_fill_1 FILLER_7_1815 ();
 sg13g2_decap_8 FILLER_7_1838 ();
 sg13g2_fill_1 FILLER_7_1845 ();
 sg13g2_decap_4 FILLER_7_1859 ();
 sg13g2_fill_1 FILLER_7_1863 ();
 sg13g2_decap_8 FILLER_7_1878 ();
 sg13g2_decap_8 FILLER_7_1885 ();
 sg13g2_decap_4 FILLER_7_1892 ();
 sg13g2_decap_4 FILLER_7_1902 ();
 sg13g2_decap_8 FILLER_7_1914 ();
 sg13g2_decap_4 FILLER_7_1921 ();
 sg13g2_decap_8 FILLER_7_1933 ();
 sg13g2_fill_1 FILLER_7_1940 ();
 sg13g2_decap_8 FILLER_7_1950 ();
 sg13g2_fill_2 FILLER_7_1961 ();
 sg13g2_fill_1 FILLER_7_1963 ();
 sg13g2_decap_4 FILLER_7_1969 ();
 sg13g2_fill_2 FILLER_7_1973 ();
 sg13g2_decap_8 FILLER_7_1988 ();
 sg13g2_fill_2 FILLER_7_1995 ();
 sg13g2_decap_8 FILLER_7_2001 ();
 sg13g2_fill_2 FILLER_7_2008 ();
 sg13g2_fill_1 FILLER_7_2010 ();
 sg13g2_fill_2 FILLER_7_2023 ();
 sg13g2_fill_2 FILLER_7_2057 ();
 sg13g2_decap_8 FILLER_7_2087 ();
 sg13g2_fill_2 FILLER_7_2094 ();
 sg13g2_fill_2 FILLER_7_2101 ();
 sg13g2_decap_4 FILLER_7_2115 ();
 sg13g2_fill_2 FILLER_7_2119 ();
 sg13g2_decap_8 FILLER_7_2140 ();
 sg13g2_decap_4 FILLER_7_2147 ();
 sg13g2_decap_8 FILLER_7_2164 ();
 sg13g2_decap_8 FILLER_7_2171 ();
 sg13g2_fill_2 FILLER_7_2178 ();
 sg13g2_decap_4 FILLER_7_2185 ();
 sg13g2_fill_2 FILLER_7_2209 ();
 sg13g2_fill_1 FILLER_7_2211 ();
 sg13g2_fill_2 FILLER_7_2235 ();
 sg13g2_fill_1 FILLER_7_2237 ();
 sg13g2_fill_1 FILLER_7_2250 ();
 sg13g2_decap_8 FILLER_7_2265 ();
 sg13g2_fill_1 FILLER_7_2289 ();
 sg13g2_fill_2 FILLER_7_2319 ();
 sg13g2_fill_1 FILLER_7_2321 ();
 sg13g2_decap_8 FILLER_7_2329 ();
 sg13g2_fill_1 FILLER_7_2336 ();
 sg13g2_fill_1 FILLER_7_2374 ();
 sg13g2_decap_4 FILLER_7_2388 ();
 sg13g2_fill_2 FILLER_7_2392 ();
 sg13g2_decap_8 FILLER_7_2399 ();
 sg13g2_fill_2 FILLER_7_2406 ();
 sg13g2_fill_1 FILLER_7_2408 ();
 sg13g2_decap_8 FILLER_7_2414 ();
 sg13g2_decap_8 FILLER_7_2421 ();
 sg13g2_decap_4 FILLER_7_2428 ();
 sg13g2_fill_1 FILLER_7_2432 ();
 sg13g2_decap_4 FILLER_7_2445 ();
 sg13g2_fill_2 FILLER_7_2449 ();
 sg13g2_decap_8 FILLER_7_2456 ();
 sg13g2_fill_2 FILLER_7_2463 ();
 sg13g2_decap_8 FILLER_7_2480 ();
 sg13g2_fill_2 FILLER_7_2490 ();
 sg13g2_decap_4 FILLER_7_2504 ();
 sg13g2_decap_8 FILLER_7_2529 ();
 sg13g2_fill_2 FILLER_7_2536 ();
 sg13g2_fill_1 FILLER_7_2538 ();
 sg13g2_decap_8 FILLER_7_2543 ();
 sg13g2_decap_8 FILLER_7_2550 ();
 sg13g2_fill_2 FILLER_7_2557 ();
 sg13g2_fill_1 FILLER_7_2559 ();
 sg13g2_decap_8 FILLER_7_2586 ();
 sg13g2_fill_2 FILLER_7_2593 ();
 sg13g2_fill_1 FILLER_7_2595 ();
 sg13g2_decap_8 FILLER_7_2613 ();
 sg13g2_fill_1 FILLER_7_2620 ();
 sg13g2_decap_4 FILLER_7_2625 ();
 sg13g2_fill_1 FILLER_7_2667 ();
 sg13g2_decap_4 FILLER_7_2698 ();
 sg13g2_decap_8 FILLER_7_2719 ();
 sg13g2_fill_1 FILLER_7_2726 ();
 sg13g2_fill_1 FILLER_7_2747 ();
 sg13g2_decap_8 FILLER_7_2771 ();
 sg13g2_fill_2 FILLER_7_2778 ();
 sg13g2_decap_8 FILLER_7_2793 ();
 sg13g2_decap_4 FILLER_7_2800 ();
 sg13g2_decap_8 FILLER_7_2827 ();
 sg13g2_decap_4 FILLER_7_2839 ();
 sg13g2_decap_4 FILLER_7_2861 ();
 sg13g2_decap_8 FILLER_7_2874 ();
 sg13g2_fill_2 FILLER_7_2881 ();
 sg13g2_fill_1 FILLER_7_2883 ();
 sg13g2_fill_2 FILLER_7_2895 ();
 sg13g2_fill_1 FILLER_7_2897 ();
 sg13g2_decap_8 FILLER_7_2911 ();
 sg13g2_decap_8 FILLER_7_2918 ();
 sg13g2_decap_8 FILLER_7_2936 ();
 sg13g2_fill_2 FILLER_7_2943 ();
 sg13g2_fill_1 FILLER_7_2945 ();
 sg13g2_decap_8 FILLER_7_2962 ();
 sg13g2_fill_1 FILLER_7_2969 ();
 sg13g2_fill_2 FILLER_7_2991 ();
 sg13g2_fill_1 FILLER_7_2993 ();
 sg13g2_decap_8 FILLER_7_3050 ();
 sg13g2_decap_8 FILLER_7_3057 ();
 sg13g2_decap_8 FILLER_7_3064 ();
 sg13g2_decap_8 FILLER_7_3071 ();
 sg13g2_decap_8 FILLER_7_3078 ();
 sg13g2_decap_8 FILLER_7_3085 ();
 sg13g2_decap_8 FILLER_7_3092 ();
 sg13g2_decap_8 FILLER_7_3099 ();
 sg13g2_decap_8 FILLER_7_3106 ();
 sg13g2_decap_8 FILLER_7_3113 ();
 sg13g2_decap_8 FILLER_7_3120 ();
 sg13g2_decap_8 FILLER_7_3127 ();
 sg13g2_decap_8 FILLER_7_3134 ();
 sg13g2_decap_8 FILLER_7_3141 ();
 sg13g2_decap_8 FILLER_7_3148 ();
 sg13g2_decap_8 FILLER_7_3155 ();
 sg13g2_decap_8 FILLER_7_3162 ();
 sg13g2_decap_8 FILLER_7_3169 ();
 sg13g2_decap_8 FILLER_7_3176 ();
 sg13g2_decap_8 FILLER_7_3183 ();
 sg13g2_decap_8 FILLER_7_3190 ();
 sg13g2_decap_8 FILLER_7_3197 ();
 sg13g2_decap_8 FILLER_7_3204 ();
 sg13g2_decap_8 FILLER_7_3211 ();
 sg13g2_decap_8 FILLER_7_3218 ();
 sg13g2_decap_8 FILLER_7_3225 ();
 sg13g2_decap_8 FILLER_7_3232 ();
 sg13g2_decap_8 FILLER_7_3239 ();
 sg13g2_decap_8 FILLER_7_3246 ();
 sg13g2_decap_8 FILLER_7_3253 ();
 sg13g2_decap_8 FILLER_7_3260 ();
 sg13g2_decap_8 FILLER_7_3267 ();
 sg13g2_decap_8 FILLER_7_3274 ();
 sg13g2_decap_8 FILLER_7_3281 ();
 sg13g2_decap_8 FILLER_7_3288 ();
 sg13g2_decap_8 FILLER_7_3295 ();
 sg13g2_decap_8 FILLER_7_3302 ();
 sg13g2_decap_8 FILLER_7_3309 ();
 sg13g2_decap_8 FILLER_7_3316 ();
 sg13g2_decap_8 FILLER_7_3323 ();
 sg13g2_decap_8 FILLER_7_3330 ();
 sg13g2_decap_8 FILLER_7_3337 ();
 sg13g2_decap_8 FILLER_7_3344 ();
 sg13g2_decap_8 FILLER_7_3351 ();
 sg13g2_decap_8 FILLER_7_3358 ();
 sg13g2_decap_8 FILLER_7_3365 ();
 sg13g2_decap_8 FILLER_7_3372 ();
 sg13g2_decap_8 FILLER_7_3379 ();
 sg13g2_decap_8 FILLER_7_3386 ();
 sg13g2_decap_8 FILLER_7_3393 ();
 sg13g2_decap_8 FILLER_7_3400 ();
 sg13g2_decap_8 FILLER_7_3407 ();
 sg13g2_decap_8 FILLER_7_3414 ();
 sg13g2_decap_8 FILLER_7_3421 ();
 sg13g2_decap_8 FILLER_7_3428 ();
 sg13g2_decap_8 FILLER_7_3435 ();
 sg13g2_decap_8 FILLER_7_3442 ();
 sg13g2_decap_8 FILLER_7_3449 ();
 sg13g2_decap_8 FILLER_7_3456 ();
 sg13g2_decap_8 FILLER_7_3463 ();
 sg13g2_decap_8 FILLER_7_3470 ();
 sg13g2_decap_8 FILLER_7_3477 ();
 sg13g2_decap_8 FILLER_7_3484 ();
 sg13g2_decap_8 FILLER_7_3491 ();
 sg13g2_decap_8 FILLER_7_3498 ();
 sg13g2_decap_8 FILLER_7_3505 ();
 sg13g2_decap_8 FILLER_7_3512 ();
 sg13g2_decap_8 FILLER_7_3519 ();
 sg13g2_decap_8 FILLER_7_3526 ();
 sg13g2_decap_8 FILLER_7_3533 ();
 sg13g2_decap_8 FILLER_7_3540 ();
 sg13g2_decap_8 FILLER_7_3547 ();
 sg13g2_decap_8 FILLER_7_3554 ();
 sg13g2_decap_8 FILLER_7_3561 ();
 sg13g2_decap_8 FILLER_7_3568 ();
 sg13g2_decap_4 FILLER_7_3575 ();
 sg13g2_fill_1 FILLER_7_3579 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_4 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_340 ();
 sg13g2_decap_4 FILLER_8_363 ();
 sg13g2_decap_4 FILLER_8_397 ();
 sg13g2_fill_2 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_410 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_fill_2 FILLER_8_460 ();
 sg13g2_fill_2 FILLER_8_471 ();
 sg13g2_decap_4 FILLER_8_521 ();
 sg13g2_fill_2 FILLER_8_560 ();
 sg13g2_fill_1 FILLER_8_562 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_4 FILLER_8_606 ();
 sg13g2_fill_2 FILLER_8_628 ();
 sg13g2_decap_8 FILLER_8_657 ();
 sg13g2_fill_2 FILLER_8_675 ();
 sg13g2_fill_2 FILLER_8_686 ();
 sg13g2_fill_1 FILLER_8_719 ();
 sg13g2_fill_1 FILLER_8_729 ();
 sg13g2_fill_1 FILLER_8_743 ();
 sg13g2_decap_8 FILLER_8_748 ();
 sg13g2_fill_2 FILLER_8_755 ();
 sg13g2_fill_1 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_fill_2 FILLER_8_770 ();
 sg13g2_fill_1 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_782 ();
 sg13g2_fill_2 FILLER_8_789 ();
 sg13g2_fill_2 FILLER_8_796 ();
 sg13g2_decap_4 FILLER_8_824 ();
 sg13g2_fill_2 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_fill_2 FILLER_8_879 ();
 sg13g2_decap_4 FILLER_8_889 ();
 sg13g2_decap_4 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_8_928 ();
 sg13g2_decap_4 FILLER_8_935 ();
 sg13g2_fill_1 FILLER_8_948 ();
 sg13g2_decap_4 FILLER_8_964 ();
 sg13g2_decap_8 FILLER_8_985 ();
 sg13g2_fill_2 FILLER_8_992 ();
 sg13g2_fill_1 FILLER_8_994 ();
 sg13g2_fill_2 FILLER_8_1051 ();
 sg13g2_fill_1 FILLER_8_1053 ();
 sg13g2_decap_4 FILLER_8_1072 ();
 sg13g2_decap_8 FILLER_8_1109 ();
 sg13g2_fill_2 FILLER_8_1120 ();
 sg13g2_fill_1 FILLER_8_1122 ();
 sg13g2_decap_8 FILLER_8_1132 ();
 sg13g2_fill_2 FILLER_8_1139 ();
 sg13g2_decap_8 FILLER_8_1165 ();
 sg13g2_decap_8 FILLER_8_1172 ();
 sg13g2_fill_2 FILLER_8_1179 ();
 sg13g2_fill_1 FILLER_8_1186 ();
 sg13g2_decap_8 FILLER_8_1196 ();
 sg13g2_decap_4 FILLER_8_1203 ();
 sg13g2_fill_1 FILLER_8_1207 ();
 sg13g2_decap_4 FILLER_8_1216 ();
 sg13g2_fill_2 FILLER_8_1220 ();
 sg13g2_decap_4 FILLER_8_1235 ();
 sg13g2_fill_1 FILLER_8_1244 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_decap_4 FILLER_8_1267 ();
 sg13g2_fill_1 FILLER_8_1271 ();
 sg13g2_decap_8 FILLER_8_1295 ();
 sg13g2_fill_2 FILLER_8_1302 ();
 sg13g2_fill_1 FILLER_8_1304 ();
 sg13g2_fill_2 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_8_1337 ();
 sg13g2_decap_8 FILLER_8_1344 ();
 sg13g2_fill_2 FILLER_8_1351 ();
 sg13g2_fill_1 FILLER_8_1353 ();
 sg13g2_fill_2 FILLER_8_1359 ();
 sg13g2_fill_1 FILLER_8_1365 ();
 sg13g2_decap_8 FILLER_8_1379 ();
 sg13g2_decap_8 FILLER_8_1386 ();
 sg13g2_fill_2 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1399 ();
 sg13g2_fill_2 FILLER_8_1406 ();
 sg13g2_fill_1 FILLER_8_1408 ();
 sg13g2_fill_2 FILLER_8_1418 ();
 sg13g2_decap_8 FILLER_8_1427 ();
 sg13g2_decap_4 FILLER_8_1434 ();
 sg13g2_fill_2 FILLER_8_1438 ();
 sg13g2_decap_8 FILLER_8_1447 ();
 sg13g2_decap_4 FILLER_8_1454 ();
 sg13g2_fill_2 FILLER_8_1458 ();
 sg13g2_fill_2 FILLER_8_1487 ();
 sg13g2_decap_4 FILLER_8_1516 ();
 sg13g2_fill_2 FILLER_8_1520 ();
 sg13g2_fill_2 FILLER_8_1569 ();
 sg13g2_fill_1 FILLER_8_1571 ();
 sg13g2_decap_8 FILLER_8_1595 ();
 sg13g2_fill_2 FILLER_8_1602 ();
 sg13g2_decap_8 FILLER_8_1612 ();
 sg13g2_decap_4 FILLER_8_1619 ();
 sg13g2_fill_1 FILLER_8_1623 ();
 sg13g2_decap_8 FILLER_8_1629 ();
 sg13g2_fill_1 FILLER_8_1636 ();
 sg13g2_decap_4 FILLER_8_1664 ();
 sg13g2_fill_2 FILLER_8_1668 ();
 sg13g2_decap_8 FILLER_8_1677 ();
 sg13g2_decap_8 FILLER_8_1684 ();
 sg13g2_decap_4 FILLER_8_1691 ();
 sg13g2_decap_8 FILLER_8_1714 ();
 sg13g2_decap_8 FILLER_8_1721 ();
 sg13g2_fill_1 FILLER_8_1728 ();
 sg13g2_fill_2 FILLER_8_1734 ();
 sg13g2_decap_4 FILLER_8_1759 ();
 sg13g2_fill_1 FILLER_8_1763 ();
 sg13g2_decap_8 FILLER_8_1851 ();
 sg13g2_fill_1 FILLER_8_1858 ();
 sg13g2_fill_2 FILLER_8_1882 ();
 sg13g2_decap_8 FILLER_8_1922 ();
 sg13g2_decap_8 FILLER_8_1951 ();
 sg13g2_decap_8 FILLER_8_1958 ();
 sg13g2_decap_4 FILLER_8_1965 ();
 sg13g2_fill_1 FILLER_8_1969 ();
 sg13g2_decap_4 FILLER_8_1980 ();
 sg13g2_fill_2 FILLER_8_1984 ();
 sg13g2_decap_4 FILLER_8_2005 ();
 sg13g2_fill_2 FILLER_8_2009 ();
 sg13g2_decap_8 FILLER_8_2028 ();
 sg13g2_decap_8 FILLER_8_2035 ();
 sg13g2_decap_8 FILLER_8_2042 ();
 sg13g2_fill_1 FILLER_8_2058 ();
 sg13g2_fill_1 FILLER_8_2070 ();
 sg13g2_decap_8 FILLER_8_2079 ();
 sg13g2_decap_4 FILLER_8_2086 ();
 sg13g2_fill_2 FILLER_8_2090 ();
 sg13g2_decap_8 FILLER_8_2112 ();
 sg13g2_decap_8 FILLER_8_2136 ();
 sg13g2_decap_8 FILLER_8_2143 ();
 sg13g2_fill_2 FILLER_8_2150 ();
 sg13g2_fill_2 FILLER_8_2156 ();
 sg13g2_decap_4 FILLER_8_2165 ();
 sg13g2_fill_1 FILLER_8_2169 ();
 sg13g2_decap_4 FILLER_8_2175 ();
 sg13g2_fill_2 FILLER_8_2179 ();
 sg13g2_fill_2 FILLER_8_2198 ();
 sg13g2_fill_1 FILLER_8_2200 ();
 sg13g2_decap_4 FILLER_8_2206 ();
 sg13g2_fill_2 FILLER_8_2215 ();
 sg13g2_fill_1 FILLER_8_2217 ();
 sg13g2_decap_4 FILLER_8_2227 ();
 sg13g2_fill_1 FILLER_8_2231 ();
 sg13g2_decap_8 FILLER_8_2237 ();
 sg13g2_decap_4 FILLER_8_2244 ();
 sg13g2_decap_4 FILLER_8_2257 ();
 sg13g2_fill_1 FILLER_8_2261 ();
 sg13g2_fill_2 FILLER_8_2267 ();
 sg13g2_fill_1 FILLER_8_2269 ();
 sg13g2_fill_2 FILLER_8_2275 ();
 sg13g2_fill_1 FILLER_8_2277 ();
 sg13g2_fill_2 FILLER_8_2295 ();
 sg13g2_decap_8 FILLER_8_2302 ();
 sg13g2_decap_8 FILLER_8_2309 ();
 sg13g2_decap_4 FILLER_8_2316 ();
 sg13g2_decap_8 FILLER_8_2348 ();
 sg13g2_fill_1 FILLER_8_2363 ();
 sg13g2_fill_2 FILLER_8_2373 ();
 sg13g2_fill_2 FILLER_8_2383 ();
 sg13g2_fill_1 FILLER_8_2385 ();
 sg13g2_fill_1 FILLER_8_2399 ();
 sg13g2_fill_1 FILLER_8_2435 ();
 sg13g2_fill_1 FILLER_8_2446 ();
 sg13g2_decap_4 FILLER_8_2465 ();
 sg13g2_fill_2 FILLER_8_2469 ();
 sg13g2_fill_1 FILLER_8_2484 ();
 sg13g2_decap_8 FILLER_8_2502 ();
 sg13g2_decap_8 FILLER_8_2509 ();
 sg13g2_fill_2 FILLER_8_2516 ();
 sg13g2_fill_1 FILLER_8_2518 ();
 sg13g2_decap_4 FILLER_8_2529 ();
 sg13g2_fill_1 FILLER_8_2533 ();
 sg13g2_fill_1 FILLER_8_2562 ();
 sg13g2_decap_8 FILLER_8_2594 ();
 sg13g2_fill_1 FILLER_8_2650 ();
 sg13g2_decap_4 FILLER_8_2676 ();
 sg13g2_decap_4 FILLER_8_2685 ();
 sg13g2_fill_1 FILLER_8_2689 ();
 sg13g2_fill_2 FILLER_8_2695 ();
 sg13g2_fill_1 FILLER_8_2697 ();
 sg13g2_decap_8 FILLER_8_2720 ();
 sg13g2_decap_8 FILLER_8_2727 ();
 sg13g2_fill_1 FILLER_8_2734 ();
 sg13g2_decap_8 FILLER_8_2751 ();
 sg13g2_decap_8 FILLER_8_2763 ();
 sg13g2_decap_4 FILLER_8_2770 ();
 sg13g2_decap_8 FILLER_8_2818 ();
 sg13g2_decap_8 FILLER_8_2825 ();
 sg13g2_fill_1 FILLER_8_2832 ();
 sg13g2_fill_1 FILLER_8_2839 ();
 sg13g2_fill_2 FILLER_8_2845 ();
 sg13g2_fill_1 FILLER_8_2847 ();
 sg13g2_decap_8 FILLER_8_2865 ();
 sg13g2_decap_8 FILLER_8_2872 ();
 sg13g2_fill_1 FILLER_8_2879 ();
 sg13g2_fill_1 FILLER_8_2888 ();
 sg13g2_fill_1 FILLER_8_2917 ();
 sg13g2_fill_2 FILLER_8_2953 ();
 sg13g2_fill_1 FILLER_8_2970 ();
 sg13g2_fill_1 FILLER_8_2984 ();
 sg13g2_fill_1 FILLER_8_2990 ();
 sg13g2_decap_4 FILLER_8_3000 ();
 sg13g2_decap_8 FILLER_8_3035 ();
 sg13g2_decap_8 FILLER_8_3042 ();
 sg13g2_decap_8 FILLER_8_3049 ();
 sg13g2_decap_8 FILLER_8_3056 ();
 sg13g2_decap_8 FILLER_8_3063 ();
 sg13g2_decap_8 FILLER_8_3070 ();
 sg13g2_decap_8 FILLER_8_3077 ();
 sg13g2_decap_8 FILLER_8_3084 ();
 sg13g2_decap_8 FILLER_8_3091 ();
 sg13g2_decap_8 FILLER_8_3098 ();
 sg13g2_decap_8 FILLER_8_3105 ();
 sg13g2_decap_8 FILLER_8_3112 ();
 sg13g2_decap_8 FILLER_8_3119 ();
 sg13g2_decap_8 FILLER_8_3126 ();
 sg13g2_decap_8 FILLER_8_3133 ();
 sg13g2_decap_8 FILLER_8_3140 ();
 sg13g2_decap_8 FILLER_8_3147 ();
 sg13g2_decap_8 FILLER_8_3154 ();
 sg13g2_decap_8 FILLER_8_3161 ();
 sg13g2_decap_8 FILLER_8_3168 ();
 sg13g2_decap_8 FILLER_8_3175 ();
 sg13g2_decap_8 FILLER_8_3182 ();
 sg13g2_decap_8 FILLER_8_3189 ();
 sg13g2_decap_8 FILLER_8_3196 ();
 sg13g2_decap_8 FILLER_8_3203 ();
 sg13g2_decap_8 FILLER_8_3210 ();
 sg13g2_decap_8 FILLER_8_3217 ();
 sg13g2_decap_8 FILLER_8_3224 ();
 sg13g2_decap_8 FILLER_8_3231 ();
 sg13g2_decap_8 FILLER_8_3238 ();
 sg13g2_decap_8 FILLER_8_3245 ();
 sg13g2_decap_8 FILLER_8_3252 ();
 sg13g2_decap_8 FILLER_8_3259 ();
 sg13g2_decap_8 FILLER_8_3266 ();
 sg13g2_decap_8 FILLER_8_3273 ();
 sg13g2_decap_8 FILLER_8_3280 ();
 sg13g2_decap_8 FILLER_8_3287 ();
 sg13g2_decap_8 FILLER_8_3294 ();
 sg13g2_decap_8 FILLER_8_3301 ();
 sg13g2_decap_8 FILLER_8_3308 ();
 sg13g2_decap_8 FILLER_8_3315 ();
 sg13g2_decap_8 FILLER_8_3322 ();
 sg13g2_decap_8 FILLER_8_3329 ();
 sg13g2_decap_8 FILLER_8_3336 ();
 sg13g2_decap_8 FILLER_8_3343 ();
 sg13g2_decap_8 FILLER_8_3350 ();
 sg13g2_decap_8 FILLER_8_3357 ();
 sg13g2_decap_8 FILLER_8_3364 ();
 sg13g2_decap_8 FILLER_8_3371 ();
 sg13g2_decap_8 FILLER_8_3378 ();
 sg13g2_decap_8 FILLER_8_3385 ();
 sg13g2_decap_8 FILLER_8_3392 ();
 sg13g2_decap_8 FILLER_8_3399 ();
 sg13g2_decap_8 FILLER_8_3406 ();
 sg13g2_decap_8 FILLER_8_3413 ();
 sg13g2_decap_8 FILLER_8_3420 ();
 sg13g2_decap_8 FILLER_8_3427 ();
 sg13g2_decap_8 FILLER_8_3434 ();
 sg13g2_decap_8 FILLER_8_3441 ();
 sg13g2_decap_8 FILLER_8_3448 ();
 sg13g2_decap_8 FILLER_8_3455 ();
 sg13g2_decap_8 FILLER_8_3462 ();
 sg13g2_decap_8 FILLER_8_3469 ();
 sg13g2_decap_8 FILLER_8_3476 ();
 sg13g2_decap_8 FILLER_8_3483 ();
 sg13g2_decap_8 FILLER_8_3490 ();
 sg13g2_decap_8 FILLER_8_3497 ();
 sg13g2_decap_8 FILLER_8_3504 ();
 sg13g2_decap_8 FILLER_8_3511 ();
 sg13g2_decap_8 FILLER_8_3518 ();
 sg13g2_decap_8 FILLER_8_3525 ();
 sg13g2_decap_8 FILLER_8_3532 ();
 sg13g2_decap_8 FILLER_8_3539 ();
 sg13g2_decap_8 FILLER_8_3546 ();
 sg13g2_decap_8 FILLER_8_3553 ();
 sg13g2_decap_8 FILLER_8_3560 ();
 sg13g2_decap_8 FILLER_8_3567 ();
 sg13g2_decap_4 FILLER_8_3574 ();
 sg13g2_fill_2 FILLER_8_3578 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_4 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_decap_4 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_9_432 ();
 sg13g2_decap_8 FILLER_9_450 ();
 sg13g2_decap_4 FILLER_9_457 ();
 sg13g2_decap_8 FILLER_9_475 ();
 sg13g2_fill_2 FILLER_9_482 ();
 sg13g2_fill_1 FILLER_9_484 ();
 sg13g2_decap_4 FILLER_9_489 ();
 sg13g2_decap_8 FILLER_9_498 ();
 sg13g2_decap_8 FILLER_9_505 ();
 sg13g2_decap_8 FILLER_9_512 ();
 sg13g2_fill_2 FILLER_9_519 ();
 sg13g2_fill_1 FILLER_9_521 ();
 sg13g2_fill_1 FILLER_9_537 ();
 sg13g2_decap_8 FILLER_9_548 ();
 sg13g2_decap_8 FILLER_9_555 ();
 sg13g2_fill_1 FILLER_9_562 ();
 sg13g2_fill_2 FILLER_9_567 ();
 sg13g2_fill_1 FILLER_9_569 ();
 sg13g2_fill_2 FILLER_9_579 ();
 sg13g2_fill_1 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_4 FILLER_9_594 ();
 sg13g2_fill_1 FILLER_9_598 ();
 sg13g2_fill_2 FILLER_9_654 ();
 sg13g2_decap_4 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_671 ();
 sg13g2_fill_2 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_691 ();
 sg13g2_fill_1 FILLER_9_705 ();
 sg13g2_decap_4 FILLER_9_719 ();
 sg13g2_fill_2 FILLER_9_723 ();
 sg13g2_fill_1 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_789 ();
 sg13g2_decap_8 FILLER_9_796 ();
 sg13g2_fill_1 FILLER_9_816 ();
 sg13g2_fill_2 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_865 ();
 sg13g2_fill_2 FILLER_9_874 ();
 sg13g2_decap_8 FILLER_9_892 ();
 sg13g2_fill_1 FILLER_9_917 ();
 sg13g2_fill_1 FILLER_9_936 ();
 sg13g2_decap_4 FILLER_9_956 ();
 sg13g2_decap_8 FILLER_9_1011 ();
 sg13g2_fill_1 FILLER_9_1018 ();
 sg13g2_decap_8 FILLER_9_1023 ();
 sg13g2_decap_4 FILLER_9_1030 ();
 sg13g2_fill_2 FILLER_9_1051 ();
 sg13g2_fill_1 FILLER_9_1053 ();
 sg13g2_decap_8 FILLER_9_1060 ();
 sg13g2_fill_1 FILLER_9_1067 ();
 sg13g2_fill_1 FILLER_9_1085 ();
 sg13g2_decap_8 FILLER_9_1090 ();
 sg13g2_fill_1 FILLER_9_1101 ();
 sg13g2_fill_2 FILLER_9_1146 ();
 sg13g2_fill_1 FILLER_9_1153 ();
 sg13g2_fill_2 FILLER_9_1161 ();
 sg13g2_fill_1 FILLER_9_1163 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1191 ();
 sg13g2_decap_4 FILLER_9_1198 ();
 sg13g2_fill_1 FILLER_9_1202 ();
 sg13g2_fill_1 FILLER_9_1215 ();
 sg13g2_fill_2 FILLER_9_1224 ();
 sg13g2_fill_2 FILLER_9_1249 ();
 sg13g2_fill_1 FILLER_9_1251 ();
 sg13g2_decap_8 FILLER_9_1270 ();
 sg13g2_decap_8 FILLER_9_1277 ();
 sg13g2_fill_2 FILLER_9_1284 ();
 sg13g2_fill_1 FILLER_9_1286 ();
 sg13g2_decap_8 FILLER_9_1292 ();
 sg13g2_fill_2 FILLER_9_1299 ();
 sg13g2_fill_2 FILLER_9_1322 ();
 sg13g2_decap_8 FILLER_9_1335 ();
 sg13g2_decap_8 FILLER_9_1357 ();
 sg13g2_fill_2 FILLER_9_1375 ();
 sg13g2_fill_1 FILLER_9_1382 ();
 sg13g2_fill_2 FILLER_9_1446 ();
 sg13g2_fill_1 FILLER_9_1448 ();
 sg13g2_fill_2 FILLER_9_1470 ();
 sg13g2_fill_1 FILLER_9_1472 ();
 sg13g2_decap_4 FILLER_9_1488 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_fill_2 FILLER_9_1526 ();
 sg13g2_decap_4 FILLER_9_1533 ();
 sg13g2_fill_2 FILLER_9_1537 ();
 sg13g2_fill_2 FILLER_9_1544 ();
 sg13g2_fill_1 FILLER_9_1546 ();
 sg13g2_fill_1 FILLER_9_1556 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_fill_2 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1590 ();
 sg13g2_decap_8 FILLER_9_1597 ();
 sg13g2_fill_2 FILLER_9_1604 ();
 sg13g2_decap_4 FILLER_9_1620 ();
 sg13g2_fill_1 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1630 ();
 sg13g2_decap_8 FILLER_9_1637 ();
 sg13g2_fill_2 FILLER_9_1644 ();
 sg13g2_fill_1 FILLER_9_1646 ();
 sg13g2_fill_2 FILLER_9_1652 ();
 sg13g2_fill_1 FILLER_9_1654 ();
 sg13g2_decap_8 FILLER_9_1668 ();
 sg13g2_fill_1 FILLER_9_1675 ();
 sg13g2_decap_8 FILLER_9_1689 ();
 sg13g2_decap_4 FILLER_9_1701 ();
 sg13g2_fill_1 FILLER_9_1710 ();
 sg13g2_decap_8 FILLER_9_1716 ();
 sg13g2_decap_8 FILLER_9_1731 ();
 sg13g2_decap_8 FILLER_9_1738 ();
 sg13g2_fill_1 FILLER_9_1745 ();
 sg13g2_decap_8 FILLER_9_1786 ();
 sg13g2_decap_8 FILLER_9_1793 ();
 sg13g2_decap_4 FILLER_9_1810 ();
 sg13g2_fill_2 FILLER_9_1814 ();
 sg13g2_decap_8 FILLER_9_1842 ();
 sg13g2_decap_4 FILLER_9_1849 ();
 sg13g2_fill_2 FILLER_9_1869 ();
 sg13g2_decap_8 FILLER_9_1884 ();
 sg13g2_fill_1 FILLER_9_1891 ();
 sg13g2_decap_4 FILLER_9_1909 ();
 sg13g2_fill_1 FILLER_9_1913 ();
 sg13g2_fill_2 FILLER_9_1924 ();
 sg13g2_fill_1 FILLER_9_1926 ();
 sg13g2_decap_4 FILLER_9_1950 ();
 sg13g2_fill_2 FILLER_9_1954 ();
 sg13g2_fill_1 FILLER_9_1963 ();
 sg13g2_decap_8 FILLER_9_1984 ();
 sg13g2_fill_1 FILLER_9_1991 ();
 sg13g2_decap_4 FILLER_9_1997 ();
 sg13g2_fill_1 FILLER_9_2001 ();
 sg13g2_decap_8 FILLER_9_2031 ();
 sg13g2_fill_1 FILLER_9_2054 ();
 sg13g2_decap_4 FILLER_9_2063 ();
 sg13g2_fill_2 FILLER_9_2084 ();
 sg13g2_decap_8 FILLER_9_2104 ();
 sg13g2_fill_1 FILLER_9_2121 ();
 sg13g2_fill_2 FILLER_9_2127 ();
 sg13g2_fill_1 FILLER_9_2129 ();
 sg13g2_decap_8 FILLER_9_2138 ();
 sg13g2_fill_2 FILLER_9_2145 ();
 sg13g2_fill_2 FILLER_9_2157 ();
 sg13g2_fill_2 FILLER_9_2170 ();
 sg13g2_fill_1 FILLER_9_2172 ();
 sg13g2_fill_2 FILLER_9_2179 ();
 sg13g2_fill_1 FILLER_9_2181 ();
 sg13g2_decap_4 FILLER_9_2186 ();
 sg13g2_fill_2 FILLER_9_2190 ();
 sg13g2_decap_8 FILLER_9_2205 ();
 sg13g2_fill_1 FILLER_9_2212 ();
 sg13g2_fill_1 FILLER_9_2216 ();
 sg13g2_fill_2 FILLER_9_2225 ();
 sg13g2_fill_1 FILLER_9_2227 ();
 sg13g2_decap_4 FILLER_9_2231 ();
 sg13g2_decap_8 FILLER_9_2239 ();
 sg13g2_decap_8 FILLER_9_2246 ();
 sg13g2_decap_4 FILLER_9_2253 ();
 sg13g2_fill_1 FILLER_9_2257 ();
 sg13g2_fill_2 FILLER_9_2274 ();
 sg13g2_decap_8 FILLER_9_2294 ();
 sg13g2_fill_2 FILLER_9_2301 ();
 sg13g2_fill_1 FILLER_9_2303 ();
 sg13g2_decap_8 FILLER_9_2321 ();
 sg13g2_decap_8 FILLER_9_2328 ();
 sg13g2_decap_8 FILLER_9_2335 ();
 sg13g2_fill_2 FILLER_9_2342 ();
 sg13g2_fill_1 FILLER_9_2344 ();
 sg13g2_fill_2 FILLER_9_2363 ();
 sg13g2_fill_2 FILLER_9_2373 ();
 sg13g2_fill_2 FILLER_9_2380 ();
 sg13g2_fill_1 FILLER_9_2382 ();
 sg13g2_fill_2 FILLER_9_2403 ();
 sg13g2_fill_1 FILLER_9_2405 ();
 sg13g2_decap_8 FILLER_9_2410 ();
 sg13g2_decap_8 FILLER_9_2417 ();
 sg13g2_fill_2 FILLER_9_2424 ();
 sg13g2_fill_1 FILLER_9_2426 ();
 sg13g2_fill_1 FILLER_9_2434 ();
 sg13g2_decap_4 FILLER_9_2444 ();
 sg13g2_fill_1 FILLER_9_2448 ();
 sg13g2_decap_8 FILLER_9_2477 ();
 sg13g2_decap_4 FILLER_9_2484 ();
 sg13g2_decap_8 FILLER_9_2511 ();
 sg13g2_fill_1 FILLER_9_2518 ();
 sg13g2_decap_8 FILLER_9_2527 ();
 sg13g2_decap_8 FILLER_9_2534 ();
 sg13g2_fill_2 FILLER_9_2541 ();
 sg13g2_decap_8 FILLER_9_2563 ();
 sg13g2_fill_1 FILLER_9_2570 ();
 sg13g2_decap_4 FILLER_9_2588 ();
 sg13g2_fill_1 FILLER_9_2592 ();
 sg13g2_decap_8 FILLER_9_2606 ();
 sg13g2_decap_8 FILLER_9_2613 ();
 sg13g2_decap_8 FILLER_9_2620 ();
 sg13g2_decap_8 FILLER_9_2627 ();
 sg13g2_decap_4 FILLER_9_2634 ();
 sg13g2_fill_2 FILLER_9_2661 ();
 sg13g2_fill_1 FILLER_9_2663 ();
 sg13g2_fill_2 FILLER_9_2688 ();
 sg13g2_fill_1 FILLER_9_2690 ();
 sg13g2_decap_8 FILLER_9_2719 ();
 sg13g2_fill_2 FILLER_9_2726 ();
 sg13g2_decap_8 FILLER_9_2748 ();
 sg13g2_fill_2 FILLER_9_2755 ();
 sg13g2_decap_8 FILLER_9_2769 ();
 sg13g2_fill_2 FILLER_9_2776 ();
 sg13g2_fill_1 FILLER_9_2778 ();
 sg13g2_decap_8 FILLER_9_2792 ();
 sg13g2_fill_1 FILLER_9_2799 ();
 sg13g2_decap_8 FILLER_9_2819 ();
 sg13g2_decap_8 FILLER_9_2826 ();
 sg13g2_fill_2 FILLER_9_2833 ();
 sg13g2_fill_1 FILLER_9_2835 ();
 sg13g2_fill_1 FILLER_9_2848 ();
 sg13g2_fill_2 FILLER_9_2854 ();
 sg13g2_fill_1 FILLER_9_2856 ();
 sg13g2_fill_1 FILLER_9_2862 ();
 sg13g2_fill_1 FILLER_9_2873 ();
 sg13g2_decap_8 FILLER_9_2882 ();
 sg13g2_decap_8 FILLER_9_2889 ();
 sg13g2_fill_1 FILLER_9_2896 ();
 sg13g2_decap_8 FILLER_9_2916 ();
 sg13g2_decap_4 FILLER_9_2923 ();
 sg13g2_fill_1 FILLER_9_2927 ();
 sg13g2_fill_2 FILLER_9_2937 ();
 sg13g2_fill_1 FILLER_9_2939 ();
 sg13g2_fill_1 FILLER_9_2948 ();
 sg13g2_fill_2 FILLER_9_2968 ();
 sg13g2_fill_1 FILLER_9_2970 ();
 sg13g2_decap_4 FILLER_9_2975 ();
 sg13g2_decap_4 FILLER_9_2985 ();
 sg13g2_fill_1 FILLER_9_3039 ();
 sg13g2_decap_8 FILLER_9_3057 ();
 sg13g2_decap_8 FILLER_9_3064 ();
 sg13g2_decap_8 FILLER_9_3071 ();
 sg13g2_decap_8 FILLER_9_3078 ();
 sg13g2_decap_8 FILLER_9_3085 ();
 sg13g2_decap_8 FILLER_9_3092 ();
 sg13g2_decap_8 FILLER_9_3099 ();
 sg13g2_decap_8 FILLER_9_3106 ();
 sg13g2_decap_8 FILLER_9_3113 ();
 sg13g2_decap_8 FILLER_9_3120 ();
 sg13g2_decap_8 FILLER_9_3127 ();
 sg13g2_decap_8 FILLER_9_3134 ();
 sg13g2_decap_8 FILLER_9_3141 ();
 sg13g2_decap_8 FILLER_9_3148 ();
 sg13g2_decap_8 FILLER_9_3155 ();
 sg13g2_decap_8 FILLER_9_3162 ();
 sg13g2_decap_8 FILLER_9_3169 ();
 sg13g2_decap_8 FILLER_9_3176 ();
 sg13g2_decap_8 FILLER_9_3183 ();
 sg13g2_decap_8 FILLER_9_3190 ();
 sg13g2_decap_8 FILLER_9_3197 ();
 sg13g2_decap_8 FILLER_9_3204 ();
 sg13g2_decap_8 FILLER_9_3211 ();
 sg13g2_decap_8 FILLER_9_3218 ();
 sg13g2_decap_8 FILLER_9_3225 ();
 sg13g2_decap_8 FILLER_9_3232 ();
 sg13g2_decap_8 FILLER_9_3239 ();
 sg13g2_decap_8 FILLER_9_3246 ();
 sg13g2_decap_8 FILLER_9_3253 ();
 sg13g2_decap_8 FILLER_9_3260 ();
 sg13g2_decap_8 FILLER_9_3267 ();
 sg13g2_decap_8 FILLER_9_3274 ();
 sg13g2_decap_8 FILLER_9_3281 ();
 sg13g2_decap_8 FILLER_9_3288 ();
 sg13g2_decap_8 FILLER_9_3295 ();
 sg13g2_decap_8 FILLER_9_3302 ();
 sg13g2_decap_8 FILLER_9_3309 ();
 sg13g2_decap_8 FILLER_9_3316 ();
 sg13g2_decap_8 FILLER_9_3323 ();
 sg13g2_decap_8 FILLER_9_3330 ();
 sg13g2_decap_8 FILLER_9_3337 ();
 sg13g2_decap_8 FILLER_9_3344 ();
 sg13g2_decap_8 FILLER_9_3351 ();
 sg13g2_decap_8 FILLER_9_3358 ();
 sg13g2_decap_8 FILLER_9_3365 ();
 sg13g2_decap_8 FILLER_9_3372 ();
 sg13g2_decap_8 FILLER_9_3379 ();
 sg13g2_decap_8 FILLER_9_3386 ();
 sg13g2_decap_8 FILLER_9_3393 ();
 sg13g2_decap_8 FILLER_9_3400 ();
 sg13g2_decap_8 FILLER_9_3407 ();
 sg13g2_decap_8 FILLER_9_3414 ();
 sg13g2_decap_8 FILLER_9_3421 ();
 sg13g2_decap_8 FILLER_9_3428 ();
 sg13g2_decap_8 FILLER_9_3435 ();
 sg13g2_decap_8 FILLER_9_3442 ();
 sg13g2_decap_8 FILLER_9_3449 ();
 sg13g2_decap_8 FILLER_9_3456 ();
 sg13g2_decap_8 FILLER_9_3463 ();
 sg13g2_decap_8 FILLER_9_3470 ();
 sg13g2_decap_8 FILLER_9_3477 ();
 sg13g2_decap_8 FILLER_9_3484 ();
 sg13g2_decap_8 FILLER_9_3491 ();
 sg13g2_decap_8 FILLER_9_3498 ();
 sg13g2_decap_8 FILLER_9_3505 ();
 sg13g2_decap_8 FILLER_9_3512 ();
 sg13g2_decap_8 FILLER_9_3519 ();
 sg13g2_decap_8 FILLER_9_3526 ();
 sg13g2_decap_8 FILLER_9_3533 ();
 sg13g2_decap_8 FILLER_9_3540 ();
 sg13g2_decap_8 FILLER_9_3547 ();
 sg13g2_decap_8 FILLER_9_3554 ();
 sg13g2_decap_8 FILLER_9_3561 ();
 sg13g2_decap_8 FILLER_9_3568 ();
 sg13g2_decap_4 FILLER_9_3575 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_301 ();
 sg13g2_fill_1 FILLER_10_303 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_4 FILLER_10_369 ();
 sg13g2_fill_2 FILLER_10_373 ();
 sg13g2_fill_2 FILLER_10_403 ();
 sg13g2_decap_4 FILLER_10_424 ();
 sg13g2_decap_4 FILLER_10_456 ();
 sg13g2_fill_1 FILLER_10_460 ();
 sg13g2_decap_4 FILLER_10_481 ();
 sg13g2_fill_2 FILLER_10_485 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_508 ();
 sg13g2_fill_2 FILLER_10_534 ();
 sg13g2_fill_1 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_545 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_2 FILLER_10_557 ();
 sg13g2_fill_2 FILLER_10_564 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_4 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_621 ();
 sg13g2_decap_8 FILLER_10_628 ();
 sg13g2_decap_4 FILLER_10_635 ();
 sg13g2_fill_1 FILLER_10_639 ();
 sg13g2_fill_1 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_4 FILLER_10_722 ();
 sg13g2_fill_1 FILLER_10_740 ();
 sg13g2_decap_8 FILLER_10_745 ();
 sg13g2_fill_1 FILLER_10_756 ();
 sg13g2_decap_4 FILLER_10_762 ();
 sg13g2_fill_1 FILLER_10_766 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_4 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_834 ();
 sg13g2_fill_2 FILLER_10_841 ();
 sg13g2_fill_1 FILLER_10_872 ();
 sg13g2_fill_2 FILLER_10_878 ();
 sg13g2_fill_1 FILLER_10_880 ();
 sg13g2_decap_4 FILLER_10_898 ();
 sg13g2_fill_2 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_fill_2 FILLER_10_938 ();
 sg13g2_fill_2 FILLER_10_948 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_4 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_4 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_decap_8 FILLER_10_1069 ();
 sg13g2_decap_8 FILLER_10_1076 ();
 sg13g2_fill_1 FILLER_10_1111 ();
 sg13g2_fill_2 FILLER_10_1184 ();
 sg13g2_fill_1 FILLER_10_1186 ();
 sg13g2_decap_4 FILLER_10_1197 ();
 sg13g2_fill_2 FILLER_10_1201 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_fill_2 FILLER_10_1239 ();
 sg13g2_fill_1 FILLER_10_1241 ();
 sg13g2_decap_8 FILLER_10_1257 ();
 sg13g2_decap_8 FILLER_10_1264 ();
 sg13g2_decap_8 FILLER_10_1271 ();
 sg13g2_decap_4 FILLER_10_1278 ();
 sg13g2_fill_2 FILLER_10_1300 ();
 sg13g2_decap_4 FILLER_10_1321 ();
 sg13g2_fill_2 FILLER_10_1341 ();
 sg13g2_fill_1 FILLER_10_1343 ();
 sg13g2_fill_1 FILLER_10_1349 ();
 sg13g2_decap_8 FILLER_10_1360 ();
 sg13g2_decap_8 FILLER_10_1367 ();
 sg13g2_fill_1 FILLER_10_1374 ();
 sg13g2_decap_8 FILLER_10_1380 ();
 sg13g2_decap_4 FILLER_10_1387 ();
 sg13g2_fill_1 FILLER_10_1391 ();
 sg13g2_decap_8 FILLER_10_1406 ();
 sg13g2_decap_8 FILLER_10_1413 ();
 sg13g2_decap_4 FILLER_10_1420 ();
 sg13g2_decap_8 FILLER_10_1430 ();
 sg13g2_decap_8 FILLER_10_1437 ();
 sg13g2_decap_8 FILLER_10_1451 ();
 sg13g2_decap_4 FILLER_10_1458 ();
 sg13g2_fill_2 FILLER_10_1462 ();
 sg13g2_fill_2 FILLER_10_1505 ();
 sg13g2_fill_1 FILLER_10_1507 ();
 sg13g2_decap_4 FILLER_10_1521 ();
 sg13g2_fill_1 FILLER_10_1525 ();
 sg13g2_fill_2 FILLER_10_1547 ();
 sg13g2_decap_8 FILLER_10_1567 ();
 sg13g2_decap_4 FILLER_10_1574 ();
 sg13g2_fill_1 FILLER_10_1578 ();
 sg13g2_decap_8 FILLER_10_1587 ();
 sg13g2_fill_2 FILLER_10_1594 ();
 sg13g2_fill_2 FILLER_10_1609 ();
 sg13g2_decap_8 FILLER_10_1628 ();
 sg13g2_fill_1 FILLER_10_1635 ();
 sg13g2_fill_1 FILLER_10_1649 ();
 sg13g2_decap_4 FILLER_10_1655 ();
 sg13g2_fill_1 FILLER_10_1670 ();
 sg13g2_fill_1 FILLER_10_1716 ();
 sg13g2_decap_8 FILLER_10_1750 ();
 sg13g2_fill_2 FILLER_10_1757 ();
 sg13g2_decap_8 FILLER_10_1763 ();
 sg13g2_fill_2 FILLER_10_1770 ();
 sg13g2_fill_1 FILLER_10_1772 ();
 sg13g2_decap_8 FILLER_10_1777 ();
 sg13g2_fill_2 FILLER_10_1784 ();
 sg13g2_fill_1 FILLER_10_1786 ();
 sg13g2_decap_4 FILLER_10_1804 ();
 sg13g2_fill_1 FILLER_10_1821 ();
 sg13g2_fill_2 FILLER_10_1833 ();
 sg13g2_fill_1 FILLER_10_1835 ();
 sg13g2_fill_2 FILLER_10_1848 ();
 sg13g2_fill_1 FILLER_10_1850 ();
 sg13g2_decap_4 FILLER_10_1882 ();
 sg13g2_fill_1 FILLER_10_1886 ();
 sg13g2_fill_1 FILLER_10_1913 ();
 sg13g2_fill_2 FILLER_10_1919 ();
 sg13g2_fill_1 FILLER_10_1921 ();
 sg13g2_decap_8 FILLER_10_1926 ();
 sg13g2_decap_8 FILLER_10_1933 ();
 sg13g2_decap_8 FILLER_10_1940 ();
 sg13g2_decap_4 FILLER_10_1947 ();
 sg13g2_fill_1 FILLER_10_1951 ();
 sg13g2_fill_2 FILLER_10_1960 ();
 sg13g2_fill_1 FILLER_10_1962 ();
 sg13g2_fill_1 FILLER_10_1966 ();
 sg13g2_decap_8 FILLER_10_1975 ();
 sg13g2_decap_8 FILLER_10_1982 ();
 sg13g2_decap_4 FILLER_10_1989 ();
 sg13g2_fill_1 FILLER_10_1993 ();
 sg13g2_decap_8 FILLER_10_1998 ();
 sg13g2_decap_8 FILLER_10_2005 ();
 sg13g2_fill_1 FILLER_10_2012 ();
 sg13g2_decap_4 FILLER_10_2023 ();
 sg13g2_decap_8 FILLER_10_2036 ();
 sg13g2_fill_1 FILLER_10_2051 ();
 sg13g2_decap_4 FILLER_10_2057 ();
 sg13g2_fill_2 FILLER_10_2061 ();
 sg13g2_decap_8 FILLER_10_2072 ();
 sg13g2_decap_8 FILLER_10_2079 ();
 sg13g2_fill_1 FILLER_10_2086 ();
 sg13g2_fill_2 FILLER_10_2092 ();
 sg13g2_decap_8 FILLER_10_2104 ();
 sg13g2_fill_1 FILLER_10_2111 ();
 sg13g2_fill_2 FILLER_10_2120 ();
 sg13g2_fill_1 FILLER_10_2131 ();
 sg13g2_decap_4 FILLER_10_2142 ();
 sg13g2_decap_8 FILLER_10_2150 ();
 sg13g2_fill_1 FILLER_10_2157 ();
 sg13g2_decap_4 FILLER_10_2172 ();
 sg13g2_fill_1 FILLER_10_2176 ();
 sg13g2_decap_8 FILLER_10_2190 ();
 sg13g2_decap_8 FILLER_10_2197 ();
 sg13g2_fill_2 FILLER_10_2204 ();
 sg13g2_fill_2 FILLER_10_2216 ();
 sg13g2_fill_2 FILLER_10_2268 ();
 sg13g2_fill_1 FILLER_10_2270 ();
 sg13g2_decap_8 FILLER_10_2297 ();
 sg13g2_fill_2 FILLER_10_2304 ();
 sg13g2_fill_1 FILLER_10_2306 ();
 sg13g2_decap_4 FILLER_10_2353 ();
 sg13g2_decap_4 FILLER_10_2365 ();
 sg13g2_fill_2 FILLER_10_2369 ();
 sg13g2_decap_4 FILLER_10_2412 ();
 sg13g2_fill_1 FILLER_10_2416 ();
 sg13g2_fill_1 FILLER_10_2449 ();
 sg13g2_decap_8 FILLER_10_2481 ();
 sg13g2_decap_8 FILLER_10_2488 ();
 sg13g2_decap_8 FILLER_10_2508 ();
 sg13g2_fill_2 FILLER_10_2515 ();
 sg13g2_fill_1 FILLER_10_2517 ();
 sg13g2_fill_1 FILLER_10_2530 ();
 sg13g2_fill_1 FILLER_10_2556 ();
 sg13g2_decap_4 FILLER_10_2566 ();
 sg13g2_fill_1 FILLER_10_2570 ();
 sg13g2_fill_2 FILLER_10_2630 ();
 sg13g2_fill_1 FILLER_10_2632 ();
 sg13g2_fill_2 FILLER_10_2641 ();
 sg13g2_fill_1 FILLER_10_2643 ();
 sg13g2_fill_1 FILLER_10_2660 ();
 sg13g2_fill_2 FILLER_10_2674 ();
 sg13g2_fill_1 FILLER_10_2676 ();
 sg13g2_fill_1 FILLER_10_2695 ();
 sg13g2_fill_1 FILLER_10_2700 ();
 sg13g2_decap_4 FILLER_10_2711 ();
 sg13g2_decap_8 FILLER_10_2727 ();
 sg13g2_decap_8 FILLER_10_2734 ();
 sg13g2_fill_1 FILLER_10_2741 ();
 sg13g2_fill_2 FILLER_10_2747 ();
 sg13g2_fill_1 FILLER_10_2762 ();
 sg13g2_fill_2 FILLER_10_2781 ();
 sg13g2_fill_1 FILLER_10_2783 ();
 sg13g2_decap_8 FILLER_10_2800 ();
 sg13g2_decap_8 FILLER_10_2811 ();
 sg13g2_decap_8 FILLER_10_2826 ();
 sg13g2_fill_1 FILLER_10_2833 ();
 sg13g2_fill_2 FILLER_10_2852 ();
 sg13g2_fill_1 FILLER_10_2854 ();
 sg13g2_fill_1 FILLER_10_2860 ();
 sg13g2_fill_1 FILLER_10_2866 ();
 sg13g2_decap_4 FILLER_10_2884 ();
 sg13g2_fill_2 FILLER_10_2888 ();
 sg13g2_fill_2 FILLER_10_2900 ();
 sg13g2_decap_4 FILLER_10_2913 ();
 sg13g2_fill_2 FILLER_10_2917 ();
 sg13g2_decap_8 FILLER_10_2931 ();
 sg13g2_fill_1 FILLER_10_2938 ();
 sg13g2_decap_4 FILLER_10_2952 ();
 sg13g2_fill_1 FILLER_10_2956 ();
 sg13g2_decap_4 FILLER_10_2975 ();
 sg13g2_decap_8 FILLER_10_2992 ();
 sg13g2_decap_4 FILLER_10_2999 ();
 sg13g2_fill_1 FILLER_10_3003 ();
 sg13g2_fill_2 FILLER_10_3008 ();
 sg13g2_decap_8 FILLER_10_3058 ();
 sg13g2_decap_8 FILLER_10_3065 ();
 sg13g2_decap_8 FILLER_10_3072 ();
 sg13g2_decap_8 FILLER_10_3079 ();
 sg13g2_decap_8 FILLER_10_3086 ();
 sg13g2_decap_8 FILLER_10_3093 ();
 sg13g2_decap_8 FILLER_10_3100 ();
 sg13g2_decap_8 FILLER_10_3107 ();
 sg13g2_decap_8 FILLER_10_3114 ();
 sg13g2_decap_8 FILLER_10_3121 ();
 sg13g2_decap_8 FILLER_10_3128 ();
 sg13g2_decap_8 FILLER_10_3135 ();
 sg13g2_decap_8 FILLER_10_3142 ();
 sg13g2_decap_8 FILLER_10_3149 ();
 sg13g2_decap_8 FILLER_10_3156 ();
 sg13g2_decap_8 FILLER_10_3163 ();
 sg13g2_decap_8 FILLER_10_3170 ();
 sg13g2_decap_8 FILLER_10_3177 ();
 sg13g2_decap_8 FILLER_10_3184 ();
 sg13g2_decap_8 FILLER_10_3191 ();
 sg13g2_decap_8 FILLER_10_3198 ();
 sg13g2_decap_8 FILLER_10_3205 ();
 sg13g2_decap_8 FILLER_10_3212 ();
 sg13g2_decap_8 FILLER_10_3219 ();
 sg13g2_decap_8 FILLER_10_3226 ();
 sg13g2_decap_8 FILLER_10_3233 ();
 sg13g2_decap_8 FILLER_10_3240 ();
 sg13g2_decap_8 FILLER_10_3247 ();
 sg13g2_decap_8 FILLER_10_3254 ();
 sg13g2_decap_8 FILLER_10_3261 ();
 sg13g2_decap_8 FILLER_10_3268 ();
 sg13g2_decap_8 FILLER_10_3275 ();
 sg13g2_decap_8 FILLER_10_3282 ();
 sg13g2_decap_8 FILLER_10_3289 ();
 sg13g2_decap_8 FILLER_10_3296 ();
 sg13g2_decap_8 FILLER_10_3303 ();
 sg13g2_decap_8 FILLER_10_3310 ();
 sg13g2_decap_8 FILLER_10_3317 ();
 sg13g2_decap_8 FILLER_10_3324 ();
 sg13g2_decap_8 FILLER_10_3331 ();
 sg13g2_decap_8 FILLER_10_3338 ();
 sg13g2_decap_8 FILLER_10_3345 ();
 sg13g2_decap_8 FILLER_10_3352 ();
 sg13g2_decap_8 FILLER_10_3359 ();
 sg13g2_decap_8 FILLER_10_3366 ();
 sg13g2_decap_8 FILLER_10_3373 ();
 sg13g2_decap_8 FILLER_10_3380 ();
 sg13g2_decap_8 FILLER_10_3387 ();
 sg13g2_decap_8 FILLER_10_3394 ();
 sg13g2_decap_8 FILLER_10_3401 ();
 sg13g2_decap_8 FILLER_10_3408 ();
 sg13g2_decap_8 FILLER_10_3415 ();
 sg13g2_decap_8 FILLER_10_3422 ();
 sg13g2_decap_8 FILLER_10_3429 ();
 sg13g2_decap_8 FILLER_10_3436 ();
 sg13g2_decap_8 FILLER_10_3443 ();
 sg13g2_decap_8 FILLER_10_3450 ();
 sg13g2_decap_8 FILLER_10_3457 ();
 sg13g2_decap_8 FILLER_10_3464 ();
 sg13g2_decap_8 FILLER_10_3471 ();
 sg13g2_decap_8 FILLER_10_3478 ();
 sg13g2_decap_8 FILLER_10_3485 ();
 sg13g2_decap_8 FILLER_10_3492 ();
 sg13g2_decap_8 FILLER_10_3499 ();
 sg13g2_decap_8 FILLER_10_3506 ();
 sg13g2_decap_8 FILLER_10_3513 ();
 sg13g2_decap_8 FILLER_10_3520 ();
 sg13g2_decap_8 FILLER_10_3527 ();
 sg13g2_decap_8 FILLER_10_3534 ();
 sg13g2_decap_8 FILLER_10_3541 ();
 sg13g2_decap_8 FILLER_10_3548 ();
 sg13g2_decap_8 FILLER_10_3555 ();
 sg13g2_decap_8 FILLER_10_3562 ();
 sg13g2_decap_8 FILLER_10_3569 ();
 sg13g2_decap_4 FILLER_10_3576 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_fill_2 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_4 FILLER_11_371 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_2 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_11_415 ();
 sg13g2_decap_4 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_425 ();
 sg13g2_decap_4 FILLER_11_436 ();
 sg13g2_fill_1 FILLER_11_440 ();
 sg13g2_decap_8 FILLER_11_450 ();
 sg13g2_fill_1 FILLER_11_457 ();
 sg13g2_fill_1 FILLER_11_472 ();
 sg13g2_decap_4 FILLER_11_503 ();
 sg13g2_fill_2 FILLER_11_507 ();
 sg13g2_fill_2 FILLER_11_529 ();
 sg13g2_fill_1 FILLER_11_531 ();
 sg13g2_fill_1 FILLER_11_546 ();
 sg13g2_fill_1 FILLER_11_555 ();
 sg13g2_decap_4 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_569 ();
 sg13g2_fill_2 FILLER_11_583 ();
 sg13g2_fill_1 FILLER_11_594 ();
 sg13g2_decap_8 FILLER_11_605 ();
 sg13g2_fill_1 FILLER_11_618 ();
 sg13g2_decap_8 FILLER_11_639 ();
 sg13g2_fill_1 FILLER_11_646 ();
 sg13g2_decap_4 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_677 ();
 sg13g2_fill_2 FILLER_11_684 ();
 sg13g2_decap_8 FILLER_11_691 ();
 sg13g2_fill_2 FILLER_11_698 ();
 sg13g2_fill_1 FILLER_11_700 ();
 sg13g2_fill_1 FILLER_11_731 ();
 sg13g2_fill_2 FILLER_11_737 ();
 sg13g2_fill_1 FILLER_11_739 ();
 sg13g2_fill_2 FILLER_11_745 ();
 sg13g2_fill_2 FILLER_11_751 ();
 sg13g2_fill_1 FILLER_11_753 ();
 sg13g2_fill_2 FILLER_11_758 ();
 sg13g2_decap_8 FILLER_11_765 ();
 sg13g2_decap_4 FILLER_11_772 ();
 sg13g2_fill_1 FILLER_11_776 ();
 sg13g2_decap_4 FILLER_11_786 ();
 sg13g2_fill_1 FILLER_11_790 ();
 sg13g2_decap_8 FILLER_11_796 ();
 sg13g2_decap_8 FILLER_11_803 ();
 sg13g2_decap_4 FILLER_11_810 ();
 sg13g2_fill_1 FILLER_11_814 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_4 FILLER_11_840 ();
 sg13g2_fill_2 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_857 ();
 sg13g2_decap_4 FILLER_11_880 ();
 sg13g2_fill_2 FILLER_11_884 ();
 sg13g2_decap_4 FILLER_11_902 ();
 sg13g2_fill_1 FILLER_11_906 ();
 sg13g2_decap_8 FILLER_11_912 ();
 sg13g2_decap_4 FILLER_11_963 ();
 sg13g2_fill_2 FILLER_11_967 ();
 sg13g2_decap_4 FILLER_11_990 ();
 sg13g2_decap_4 FILLER_11_1029 ();
 sg13g2_fill_2 FILLER_11_1033 ();
 sg13g2_decap_8 FILLER_11_1050 ();
 sg13g2_decap_8 FILLER_11_1057 ();
 sg13g2_decap_8 FILLER_11_1064 ();
 sg13g2_fill_1 FILLER_11_1071 ();
 sg13g2_decap_8 FILLER_11_1076 ();
 sg13g2_decap_4 FILLER_11_1083 ();
 sg13g2_fill_1 FILLER_11_1087 ();
 sg13g2_fill_2 FILLER_11_1140 ();
 sg13g2_fill_1 FILLER_11_1142 ();
 sg13g2_fill_1 FILLER_11_1148 ();
 sg13g2_decap_8 FILLER_11_1157 ();
 sg13g2_decap_8 FILLER_11_1169 ();
 sg13g2_fill_1 FILLER_11_1176 ();
 sg13g2_fill_2 FILLER_11_1182 ();
 sg13g2_decap_8 FILLER_11_1200 ();
 sg13g2_decap_8 FILLER_11_1215 ();
 sg13g2_decap_8 FILLER_11_1222 ();
 sg13g2_decap_4 FILLER_11_1229 ();
 sg13g2_fill_1 FILLER_11_1233 ();
 sg13g2_decap_8 FILLER_11_1237 ();
 sg13g2_fill_2 FILLER_11_1244 ();
 sg13g2_decap_4 FILLER_11_1267 ();
 sg13g2_fill_1 FILLER_11_1288 ();
 sg13g2_decap_4 FILLER_11_1307 ();
 sg13g2_fill_1 FILLER_11_1311 ();
 sg13g2_fill_1 FILLER_11_1331 ();
 sg13g2_decap_4 FILLER_11_1336 ();
 sg13g2_fill_2 FILLER_11_1349 ();
 sg13g2_decap_8 FILLER_11_1363 ();
 sg13g2_fill_2 FILLER_11_1370 ();
 sg13g2_fill_1 FILLER_11_1372 ();
 sg13g2_decap_4 FILLER_11_1381 ();
 sg13g2_decap_8 FILLER_11_1412 ();
 sg13g2_fill_2 FILLER_11_1419 ();
 sg13g2_fill_2 FILLER_11_1449 ();
 sg13g2_fill_2 FILLER_11_1464 ();
 sg13g2_fill_2 FILLER_11_1479 ();
 sg13g2_decap_8 FILLER_11_1485 ();
 sg13g2_decap_8 FILLER_11_1511 ();
 sg13g2_fill_2 FILLER_11_1518 ();
 sg13g2_fill_1 FILLER_11_1520 ();
 sg13g2_fill_2 FILLER_11_1529 ();
 sg13g2_fill_1 FILLER_11_1531 ();
 sg13g2_decap_8 FILLER_11_1537 ();
 sg13g2_fill_1 FILLER_11_1544 ();
 sg13g2_decap_8 FILLER_11_1571 ();
 sg13g2_decap_4 FILLER_11_1578 ();
 sg13g2_fill_2 FILLER_11_1608 ();
 sg13g2_fill_1 FILLER_11_1610 ();
 sg13g2_decap_8 FILLER_11_1633 ();
 sg13g2_decap_4 FILLER_11_1640 ();
 sg13g2_fill_1 FILLER_11_1644 ();
 sg13g2_decap_8 FILLER_11_1660 ();
 sg13g2_decap_4 FILLER_11_1667 ();
 sg13g2_fill_1 FILLER_11_1671 ();
 sg13g2_fill_1 FILLER_11_1677 ();
 sg13g2_decap_8 FILLER_11_1685 ();
 sg13g2_fill_2 FILLER_11_1692 ();
 sg13g2_fill_1 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1700 ();
 sg13g2_fill_2 FILLER_11_1707 ();
 sg13g2_fill_1 FILLER_11_1709 ();
 sg13g2_fill_2 FILLER_11_1735 ();
 sg13g2_fill_1 FILLER_11_1737 ();
 sg13g2_decap_8 FILLER_11_1751 ();
 sg13g2_decap_8 FILLER_11_1758 ();
 sg13g2_fill_2 FILLER_11_1765 ();
 sg13g2_fill_1 FILLER_11_1767 ();
 sg13g2_fill_2 FILLER_11_1810 ();
 sg13g2_decap_8 FILLER_11_1842 ();
 sg13g2_decap_8 FILLER_11_1849 ();
 sg13g2_fill_1 FILLER_11_1863 ();
 sg13g2_decap_8 FILLER_11_1872 ();
 sg13g2_decap_8 FILLER_11_1879 ();
 sg13g2_fill_2 FILLER_11_1886 ();
 sg13g2_fill_1 FILLER_11_1888 ();
 sg13g2_decap_8 FILLER_11_1899 ();
 sg13g2_fill_1 FILLER_11_1947 ();
 sg13g2_decap_8 FILLER_11_1968 ();
 sg13g2_decap_8 FILLER_11_1975 ();
 sg13g2_decap_8 FILLER_11_2017 ();
 sg13g2_decap_8 FILLER_11_2024 ();
 sg13g2_decap_8 FILLER_11_2031 ();
 sg13g2_decap_4 FILLER_11_2038 ();
 sg13g2_fill_1 FILLER_11_2042 ();
 sg13g2_decap_4 FILLER_11_2047 ();
 sg13g2_fill_2 FILLER_11_2051 ();
 sg13g2_decap_8 FILLER_11_2062 ();
 sg13g2_decap_8 FILLER_11_2069 ();
 sg13g2_fill_1 FILLER_11_2096 ();
 sg13g2_decap_4 FILLER_11_2110 ();
 sg13g2_fill_1 FILLER_11_2122 ();
 sg13g2_fill_2 FILLER_11_2129 ();
 sg13g2_fill_2 FILLER_11_2144 ();
 sg13g2_fill_1 FILLER_11_2146 ();
 sg13g2_fill_2 FILLER_11_2162 ();
 sg13g2_fill_1 FILLER_11_2164 ();
 sg13g2_fill_2 FILLER_11_2181 ();
 sg13g2_decap_4 FILLER_11_2192 ();
 sg13g2_fill_1 FILLER_11_2206 ();
 sg13g2_decap_4 FILLER_11_2220 ();
 sg13g2_decap_8 FILLER_11_2230 ();
 sg13g2_decap_8 FILLER_11_2237 ();
 sg13g2_decap_4 FILLER_11_2244 ();
 sg13g2_fill_1 FILLER_11_2248 ();
 sg13g2_fill_2 FILLER_11_2266 ();
 sg13g2_fill_1 FILLER_11_2268 ();
 sg13g2_fill_2 FILLER_11_2304 ();
 sg13g2_decap_8 FILLER_11_2314 ();
 sg13g2_decap_4 FILLER_11_2321 ();
 sg13g2_decap_8 FILLER_11_2343 ();
 sg13g2_decap_4 FILLER_11_2350 ();
 sg13g2_fill_1 FILLER_11_2354 ();
 sg13g2_fill_2 FILLER_11_2363 ();
 sg13g2_fill_1 FILLER_11_2365 ();
 sg13g2_fill_1 FILLER_11_2379 ();
 sg13g2_decap_8 FILLER_11_2403 ();
 sg13g2_decap_8 FILLER_11_2410 ();
 sg13g2_fill_1 FILLER_11_2417 ();
 sg13g2_decap_8 FILLER_11_2446 ();
 sg13g2_decap_8 FILLER_11_2470 ();
 sg13g2_fill_2 FILLER_11_2477 ();
 sg13g2_fill_1 FILLER_11_2479 ();
 sg13g2_fill_2 FILLER_11_2484 ();
 sg13g2_fill_1 FILLER_11_2486 ();
 sg13g2_fill_1 FILLER_11_2498 ();
 sg13g2_decap_8 FILLER_11_2504 ();
 sg13g2_fill_2 FILLER_11_2511 ();
 sg13g2_fill_2 FILLER_11_2543 ();
 sg13g2_fill_1 FILLER_11_2545 ();
 sg13g2_decap_4 FILLER_11_2567 ();
 sg13g2_decap_8 FILLER_11_2582 ();
 sg13g2_fill_2 FILLER_11_2589 ();
 sg13g2_decap_8 FILLER_11_2619 ();
 sg13g2_decap_8 FILLER_11_2626 ();
 sg13g2_decap_8 FILLER_11_2633 ();
 sg13g2_fill_2 FILLER_11_2640 ();
 sg13g2_fill_1 FILLER_11_2642 ();
 sg13g2_decap_8 FILLER_11_2653 ();
 sg13g2_decap_8 FILLER_11_2660 ();
 sg13g2_decap_4 FILLER_11_2667 ();
 sg13g2_fill_2 FILLER_11_2671 ();
 sg13g2_decap_8 FILLER_11_2686 ();
 sg13g2_decap_4 FILLER_11_2693 ();
 sg13g2_fill_2 FILLER_11_2697 ();
 sg13g2_fill_1 FILLER_11_2717 ();
 sg13g2_decap_4 FILLER_11_2723 ();
 sg13g2_decap_4 FILLER_11_2731 ();
 sg13g2_fill_1 FILLER_11_2735 ();
 sg13g2_fill_2 FILLER_11_2748 ();
 sg13g2_fill_2 FILLER_11_2761 ();
 sg13g2_fill_1 FILLER_11_2778 ();
 sg13g2_fill_2 FILLER_11_2787 ();
 sg13g2_fill_1 FILLER_11_2816 ();
 sg13g2_fill_2 FILLER_11_2830 ();
 sg13g2_decap_8 FILLER_11_2837 ();
 sg13g2_fill_1 FILLER_11_2844 ();
 sg13g2_fill_2 FILLER_11_2863 ();
 sg13g2_fill_1 FILLER_11_2865 ();
 sg13g2_decap_4 FILLER_11_2874 ();
 sg13g2_fill_2 FILLER_11_2878 ();
 sg13g2_decap_4 FILLER_11_2884 ();
 sg13g2_fill_2 FILLER_11_2888 ();
 sg13g2_decap_8 FILLER_11_2918 ();
 sg13g2_decap_4 FILLER_11_2932 ();
 sg13g2_fill_1 FILLER_11_2936 ();
 sg13g2_fill_1 FILLER_11_2949 ();
 sg13g2_decap_4 FILLER_11_2966 ();
 sg13g2_fill_2 FILLER_11_2970 ();
 sg13g2_fill_2 FILLER_11_2985 ();
 sg13g2_decap_4 FILLER_11_2995 ();
 sg13g2_fill_2 FILLER_11_3009 ();
 sg13g2_fill_1 FILLER_11_3011 ();
 sg13g2_decap_8 FILLER_11_3034 ();
 sg13g2_fill_1 FILLER_11_3041 ();
 sg13g2_decap_8 FILLER_11_3070 ();
 sg13g2_decap_8 FILLER_11_3077 ();
 sg13g2_decap_8 FILLER_11_3084 ();
 sg13g2_decap_8 FILLER_11_3091 ();
 sg13g2_decap_8 FILLER_11_3098 ();
 sg13g2_fill_2 FILLER_11_3105 ();
 sg13g2_fill_1 FILLER_11_3107 ();
 sg13g2_decap_8 FILLER_11_3112 ();
 sg13g2_decap_8 FILLER_11_3119 ();
 sg13g2_decap_8 FILLER_11_3126 ();
 sg13g2_decap_8 FILLER_11_3133 ();
 sg13g2_decap_4 FILLER_11_3140 ();
 sg13g2_decap_8 FILLER_11_3148 ();
 sg13g2_decap_8 FILLER_11_3155 ();
 sg13g2_decap_8 FILLER_11_3162 ();
 sg13g2_decap_8 FILLER_11_3169 ();
 sg13g2_decap_8 FILLER_11_3176 ();
 sg13g2_decap_8 FILLER_11_3183 ();
 sg13g2_decap_8 FILLER_11_3190 ();
 sg13g2_decap_8 FILLER_11_3197 ();
 sg13g2_decap_8 FILLER_11_3204 ();
 sg13g2_decap_8 FILLER_11_3211 ();
 sg13g2_decap_8 FILLER_11_3218 ();
 sg13g2_decap_8 FILLER_11_3225 ();
 sg13g2_decap_8 FILLER_11_3232 ();
 sg13g2_decap_8 FILLER_11_3239 ();
 sg13g2_decap_8 FILLER_11_3246 ();
 sg13g2_decap_8 FILLER_11_3253 ();
 sg13g2_decap_8 FILLER_11_3260 ();
 sg13g2_decap_8 FILLER_11_3267 ();
 sg13g2_decap_8 FILLER_11_3274 ();
 sg13g2_decap_8 FILLER_11_3281 ();
 sg13g2_decap_8 FILLER_11_3288 ();
 sg13g2_decap_8 FILLER_11_3295 ();
 sg13g2_decap_8 FILLER_11_3302 ();
 sg13g2_decap_8 FILLER_11_3309 ();
 sg13g2_decap_8 FILLER_11_3316 ();
 sg13g2_decap_8 FILLER_11_3323 ();
 sg13g2_decap_8 FILLER_11_3330 ();
 sg13g2_decap_8 FILLER_11_3337 ();
 sg13g2_decap_8 FILLER_11_3344 ();
 sg13g2_decap_8 FILLER_11_3351 ();
 sg13g2_decap_8 FILLER_11_3358 ();
 sg13g2_decap_8 FILLER_11_3365 ();
 sg13g2_decap_8 FILLER_11_3372 ();
 sg13g2_decap_8 FILLER_11_3379 ();
 sg13g2_decap_8 FILLER_11_3386 ();
 sg13g2_decap_8 FILLER_11_3393 ();
 sg13g2_decap_8 FILLER_11_3400 ();
 sg13g2_decap_8 FILLER_11_3407 ();
 sg13g2_decap_8 FILLER_11_3414 ();
 sg13g2_decap_8 FILLER_11_3421 ();
 sg13g2_decap_8 FILLER_11_3428 ();
 sg13g2_decap_8 FILLER_11_3435 ();
 sg13g2_decap_8 FILLER_11_3442 ();
 sg13g2_decap_8 FILLER_11_3449 ();
 sg13g2_decap_8 FILLER_11_3456 ();
 sg13g2_decap_8 FILLER_11_3463 ();
 sg13g2_decap_8 FILLER_11_3470 ();
 sg13g2_decap_8 FILLER_11_3477 ();
 sg13g2_decap_8 FILLER_11_3484 ();
 sg13g2_decap_8 FILLER_11_3491 ();
 sg13g2_decap_8 FILLER_11_3498 ();
 sg13g2_decap_8 FILLER_11_3505 ();
 sg13g2_decap_8 FILLER_11_3512 ();
 sg13g2_decap_8 FILLER_11_3519 ();
 sg13g2_decap_8 FILLER_11_3526 ();
 sg13g2_decap_8 FILLER_11_3533 ();
 sg13g2_decap_8 FILLER_11_3540 ();
 sg13g2_decap_8 FILLER_11_3547 ();
 sg13g2_decap_8 FILLER_11_3554 ();
 sg13g2_decap_8 FILLER_11_3561 ();
 sg13g2_decap_8 FILLER_11_3568 ();
 sg13g2_decap_4 FILLER_11_3575 ();
 sg13g2_fill_1 FILLER_11_3579 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_fill_2 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_335 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_436 ();
 sg13g2_fill_2 FILLER_12_443 ();
 sg13g2_fill_2 FILLER_12_451 ();
 sg13g2_decap_8 FILLER_12_457 ();
 sg13g2_fill_1 FILLER_12_464 ();
 sg13g2_decap_8 FILLER_12_484 ();
 sg13g2_fill_2 FILLER_12_491 ();
 sg13g2_fill_1 FILLER_12_493 ();
 sg13g2_decap_4 FILLER_12_503 ();
 sg13g2_fill_2 FILLER_12_507 ();
 sg13g2_decap_4 FILLER_12_518 ();
 sg13g2_fill_2 FILLER_12_522 ();
 sg13g2_fill_2 FILLER_12_528 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_4 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_566 ();
 sg13g2_decap_4 FILLER_12_573 ();
 sg13g2_fill_1 FILLER_12_577 ();
 sg13g2_fill_1 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_fill_2 FILLER_12_597 ();
 sg13g2_fill_1 FILLER_12_599 ();
 sg13g2_fill_1 FILLER_12_603 ();
 sg13g2_fill_2 FILLER_12_626 ();
 sg13g2_decap_4 FILLER_12_642 ();
 sg13g2_fill_1 FILLER_12_646 ();
 sg13g2_decap_8 FILLER_12_673 ();
 sg13g2_fill_2 FILLER_12_680 ();
 sg13g2_fill_1 FILLER_12_682 ();
 sg13g2_decap_4 FILLER_12_691 ();
 sg13g2_fill_1 FILLER_12_695 ();
 sg13g2_decap_8 FILLER_12_724 ();
 sg13g2_decap_4 FILLER_12_731 ();
 sg13g2_decap_8 FILLER_12_764 ();
 sg13g2_decap_8 FILLER_12_771 ();
 sg13g2_fill_2 FILLER_12_778 ();
 sg13g2_fill_1 FILLER_12_799 ();
 sg13g2_decap_4 FILLER_12_808 ();
 sg13g2_fill_1 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_fill_2 FILLER_12_838 ();
 sg13g2_fill_1 FILLER_12_840 ();
 sg13g2_decap_4 FILLER_12_860 ();
 sg13g2_fill_2 FILLER_12_864 ();
 sg13g2_fill_2 FILLER_12_881 ();
 sg13g2_decap_4 FILLER_12_908 ();
 sg13g2_fill_1 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_8 FILLER_12_940 ();
 sg13g2_fill_1 FILLER_12_947 ();
 sg13g2_fill_2 FILLER_12_955 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_decap_4 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_fill_2 FILLER_12_989 ();
 sg13g2_decap_8 FILLER_12_1021 ();
 sg13g2_decap_8 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_12_1035 ();
 sg13g2_fill_2 FILLER_12_1042 ();
 sg13g2_decap_4 FILLER_12_1051 ();
 sg13g2_decap_8 FILLER_12_1060 ();
 sg13g2_decap_4 FILLER_12_1095 ();
 sg13g2_fill_2 FILLER_12_1099 ();
 sg13g2_decap_8 FILLER_12_1132 ();
 sg13g2_fill_2 FILLER_12_1147 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1185 ();
 sg13g2_fill_1 FILLER_12_1192 ();
 sg13g2_fill_1 FILLER_12_1207 ();
 sg13g2_decap_4 FILLER_12_1213 ();
 sg13g2_decap_4 FILLER_12_1245 ();
 sg13g2_fill_1 FILLER_12_1249 ();
 sg13g2_decap_8 FILLER_12_1255 ();
 sg13g2_decap_4 FILLER_12_1262 ();
 sg13g2_fill_2 FILLER_12_1266 ();
 sg13g2_fill_1 FILLER_12_1275 ();
 sg13g2_decap_4 FILLER_12_1281 ();
 sg13g2_fill_1 FILLER_12_1285 ();
 sg13g2_decap_4 FILLER_12_1303 ();
 sg13g2_fill_1 FILLER_12_1307 ();
 sg13g2_decap_4 FILLER_12_1312 ();
 sg13g2_fill_1 FILLER_12_1316 ();
 sg13g2_decap_8 FILLER_12_1322 ();
 sg13g2_decap_8 FILLER_12_1329 ();
 sg13g2_decap_8 FILLER_12_1336 ();
 sg13g2_decap_8 FILLER_12_1343 ();
 sg13g2_fill_1 FILLER_12_1355 ();
 sg13g2_decap_8 FILLER_12_1361 ();
 sg13g2_fill_2 FILLER_12_1368 ();
 sg13g2_decap_4 FILLER_12_1386 ();
 sg13g2_decap_8 FILLER_12_1416 ();
 sg13g2_decap_4 FILLER_12_1423 ();
 sg13g2_fill_2 FILLER_12_1431 ();
 sg13g2_fill_1 FILLER_12_1438 ();
 sg13g2_decap_4 FILLER_12_1444 ();
 sg13g2_fill_2 FILLER_12_1465 ();
 sg13g2_fill_1 FILLER_12_1467 ();
 sg13g2_fill_1 FILLER_12_1484 ();
 sg13g2_decap_4 FILLER_12_1490 ();
 sg13g2_fill_2 FILLER_12_1494 ();
 sg13g2_decap_4 FILLER_12_1500 ();
 sg13g2_decap_4 FILLER_12_1509 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_4 FILLER_12_1540 ();
 sg13g2_fill_2 FILLER_12_1544 ();
 sg13g2_decap_8 FILLER_12_1551 ();
 sg13g2_decap_4 FILLER_12_1558 ();
 sg13g2_fill_2 FILLER_12_1562 ();
 sg13g2_decap_4 FILLER_12_1576 ();
 sg13g2_fill_1 FILLER_12_1586 ();
 sg13g2_decap_4 FILLER_12_1612 ();
 sg13g2_decap_8 FILLER_12_1628 ();
 sg13g2_decap_4 FILLER_12_1635 ();
 sg13g2_fill_2 FILLER_12_1639 ();
 sg13g2_decap_4 FILLER_12_1656 ();
 sg13g2_decap_4 FILLER_12_1684 ();
 sg13g2_fill_1 FILLER_12_1688 ();
 sg13g2_decap_4 FILLER_12_1723 ();
 sg13g2_decap_4 FILLER_12_1732 ();
 sg13g2_fill_2 FILLER_12_1736 ();
 sg13g2_decap_4 FILLER_12_1751 ();
 sg13g2_fill_2 FILLER_12_1755 ();
 sg13g2_decap_8 FILLER_12_1783 ();
 sg13g2_decap_8 FILLER_12_1790 ();
 sg13g2_fill_2 FILLER_12_1797 ();
 sg13g2_decap_8 FILLER_12_1804 ();
 sg13g2_fill_2 FILLER_12_1824 ();
 sg13g2_fill_1 FILLER_12_1826 ();
 sg13g2_decap_4 FILLER_12_1840 ();
 sg13g2_decap_4 FILLER_12_1849 ();
 sg13g2_fill_1 FILLER_12_1853 ();
 sg13g2_decap_8 FILLER_12_1872 ();
 sg13g2_fill_2 FILLER_12_1879 ();
 sg13g2_fill_1 FILLER_12_1881 ();
 sg13g2_fill_1 FILLER_12_1910 ();
 sg13g2_decap_4 FILLER_12_1916 ();
 sg13g2_fill_2 FILLER_12_1950 ();
 sg13g2_fill_2 FILLER_12_1957 ();
 sg13g2_fill_2 FILLER_12_1969 ();
 sg13g2_decap_8 FILLER_12_1984 ();
 sg13g2_fill_1 FILLER_12_2100 ();
 sg13g2_decap_4 FILLER_12_2133 ();
 sg13g2_fill_2 FILLER_12_2137 ();
 sg13g2_decap_8 FILLER_12_2146 ();
 sg13g2_decap_4 FILLER_12_2153 ();
 sg13g2_fill_2 FILLER_12_2180 ();
 sg13g2_fill_2 FILLER_12_2195 ();
 sg13g2_fill_1 FILLER_12_2197 ();
 sg13g2_fill_2 FILLER_12_2201 ();
 sg13g2_decap_4 FILLER_12_2211 ();
 sg13g2_fill_1 FILLER_12_2215 ();
 sg13g2_decap_8 FILLER_12_2241 ();
 sg13g2_decap_4 FILLER_12_2283 ();
 sg13g2_decap_4 FILLER_12_2300 ();
 sg13g2_fill_2 FILLER_12_2304 ();
 sg13g2_fill_2 FILLER_12_2319 ();
 sg13g2_fill_1 FILLER_12_2321 ();
 sg13g2_decap_4 FILLER_12_2334 ();
 sg13g2_fill_2 FILLER_12_2356 ();
 sg13g2_decap_4 FILLER_12_2371 ();
 sg13g2_fill_1 FILLER_12_2375 ();
 sg13g2_decap_8 FILLER_12_2385 ();
 sg13g2_decap_4 FILLER_12_2413 ();
 sg13g2_fill_1 FILLER_12_2417 ();
 sg13g2_fill_1 FILLER_12_2431 ();
 sg13g2_decap_4 FILLER_12_2440 ();
 sg13g2_fill_1 FILLER_12_2444 ();
 sg13g2_fill_1 FILLER_12_2450 ();
 sg13g2_decap_4 FILLER_12_2459 ();
 sg13g2_fill_1 FILLER_12_2463 ();
 sg13g2_fill_2 FILLER_12_2473 ();
 sg13g2_fill_1 FILLER_12_2475 ();
 sg13g2_decap_8 FILLER_12_2486 ();
 sg13g2_fill_1 FILLER_12_2493 ();
 sg13g2_decap_4 FILLER_12_2499 ();
 sg13g2_fill_2 FILLER_12_2503 ();
 sg13g2_decap_8 FILLER_12_2536 ();
 sg13g2_fill_1 FILLER_12_2549 ();
 sg13g2_decap_8 FILLER_12_2557 ();
 sg13g2_fill_2 FILLER_12_2564 ();
 sg13g2_fill_1 FILLER_12_2566 ();
 sg13g2_decap_4 FILLER_12_2583 ();
 sg13g2_fill_2 FILLER_12_2587 ();
 sg13g2_decap_8 FILLER_12_2617 ();
 sg13g2_decap_8 FILLER_12_2624 ();
 sg13g2_fill_2 FILLER_12_2631 ();
 sg13g2_fill_1 FILLER_12_2633 ();
 sg13g2_decap_8 FILLER_12_2658 ();
 sg13g2_decap_4 FILLER_12_2665 ();
 sg13g2_fill_2 FILLER_12_2706 ();
 sg13g2_fill_1 FILLER_12_2708 ();
 sg13g2_decap_8 FILLER_12_2715 ();
 sg13g2_fill_2 FILLER_12_2763 ();
 sg13g2_fill_1 FILLER_12_2765 ();
 sg13g2_fill_2 FILLER_12_2770 ();
 sg13g2_decap_4 FILLER_12_2800 ();
 sg13g2_fill_1 FILLER_12_2804 ();
 sg13g2_decap_4 FILLER_12_2831 ();
 sg13g2_fill_1 FILLER_12_2835 ();
 sg13g2_decap_8 FILLER_12_2842 ();
 sg13g2_decap_4 FILLER_12_2849 ();
 sg13g2_decap_4 FILLER_12_2865 ();
 sg13g2_fill_2 FILLER_12_2869 ();
 sg13g2_fill_2 FILLER_12_2887 ();
 sg13g2_fill_1 FILLER_12_2889 ();
 sg13g2_fill_2 FILLER_12_2905 ();
 sg13g2_fill_1 FILLER_12_2907 ();
 sg13g2_decap_8 FILLER_12_2913 ();
 sg13g2_decap_4 FILLER_12_2920 ();
 sg13g2_fill_1 FILLER_12_2924 ();
 sg13g2_fill_1 FILLER_12_2934 ();
 sg13g2_decap_8 FILLER_12_2960 ();
 sg13g2_decap_4 FILLER_12_2967 ();
 sg13g2_decap_4 FILLER_12_2994 ();
 sg13g2_fill_1 FILLER_12_2998 ();
 sg13g2_fill_2 FILLER_12_3012 ();
 sg13g2_fill_1 FILLER_12_3014 ();
 sg13g2_decap_8 FILLER_12_3052 ();
 sg13g2_decap_8 FILLER_12_3059 ();
 sg13g2_decap_8 FILLER_12_3083 ();
 sg13g2_decap_8 FILLER_12_3090 ();
 sg13g2_fill_2 FILLER_12_3097 ();
 sg13g2_fill_1 FILLER_12_3099 ();
 sg13g2_decap_8 FILLER_12_3131 ();
 sg13g2_fill_1 FILLER_12_3138 ();
 sg13g2_decap_8 FILLER_12_3170 ();
 sg13g2_decap_8 FILLER_12_3181 ();
 sg13g2_decap_8 FILLER_12_3188 ();
 sg13g2_decap_8 FILLER_12_3195 ();
 sg13g2_decap_8 FILLER_12_3202 ();
 sg13g2_decap_8 FILLER_12_3209 ();
 sg13g2_decap_8 FILLER_12_3216 ();
 sg13g2_decap_8 FILLER_12_3223 ();
 sg13g2_decap_8 FILLER_12_3230 ();
 sg13g2_decap_8 FILLER_12_3237 ();
 sg13g2_decap_8 FILLER_12_3244 ();
 sg13g2_decap_8 FILLER_12_3251 ();
 sg13g2_decap_8 FILLER_12_3258 ();
 sg13g2_decap_8 FILLER_12_3265 ();
 sg13g2_decap_8 FILLER_12_3272 ();
 sg13g2_decap_8 FILLER_12_3279 ();
 sg13g2_decap_8 FILLER_12_3286 ();
 sg13g2_decap_8 FILLER_12_3293 ();
 sg13g2_decap_8 FILLER_12_3300 ();
 sg13g2_decap_8 FILLER_12_3307 ();
 sg13g2_decap_8 FILLER_12_3314 ();
 sg13g2_decap_8 FILLER_12_3321 ();
 sg13g2_decap_8 FILLER_12_3328 ();
 sg13g2_decap_8 FILLER_12_3335 ();
 sg13g2_decap_8 FILLER_12_3342 ();
 sg13g2_decap_8 FILLER_12_3349 ();
 sg13g2_decap_8 FILLER_12_3356 ();
 sg13g2_decap_8 FILLER_12_3363 ();
 sg13g2_decap_8 FILLER_12_3370 ();
 sg13g2_decap_8 FILLER_12_3377 ();
 sg13g2_decap_8 FILLER_12_3384 ();
 sg13g2_decap_8 FILLER_12_3391 ();
 sg13g2_decap_8 FILLER_12_3398 ();
 sg13g2_decap_8 FILLER_12_3405 ();
 sg13g2_decap_8 FILLER_12_3412 ();
 sg13g2_decap_8 FILLER_12_3419 ();
 sg13g2_decap_8 FILLER_12_3426 ();
 sg13g2_decap_8 FILLER_12_3433 ();
 sg13g2_decap_8 FILLER_12_3440 ();
 sg13g2_decap_8 FILLER_12_3447 ();
 sg13g2_decap_8 FILLER_12_3454 ();
 sg13g2_decap_8 FILLER_12_3461 ();
 sg13g2_decap_8 FILLER_12_3468 ();
 sg13g2_decap_8 FILLER_12_3475 ();
 sg13g2_decap_8 FILLER_12_3482 ();
 sg13g2_decap_8 FILLER_12_3489 ();
 sg13g2_decap_8 FILLER_12_3496 ();
 sg13g2_decap_8 FILLER_12_3503 ();
 sg13g2_decap_8 FILLER_12_3510 ();
 sg13g2_decap_8 FILLER_12_3517 ();
 sg13g2_decap_8 FILLER_12_3524 ();
 sg13g2_decap_8 FILLER_12_3531 ();
 sg13g2_decap_8 FILLER_12_3538 ();
 sg13g2_decap_8 FILLER_12_3545 ();
 sg13g2_decap_8 FILLER_12_3552 ();
 sg13g2_decap_8 FILLER_12_3559 ();
 sg13g2_decap_8 FILLER_12_3566 ();
 sg13g2_decap_8 FILLER_12_3573 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_4 FILLER_13_301 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_fill_2 FILLER_13_394 ();
 sg13g2_fill_1 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_fill_2 FILLER_13_409 ();
 sg13g2_decap_4 FILLER_13_431 ();
 sg13g2_fill_1 FILLER_13_435 ();
 sg13g2_fill_2 FILLER_13_456 ();
 sg13g2_fill_1 FILLER_13_458 ();
 sg13g2_fill_2 FILLER_13_472 ();
 sg13g2_fill_1 FILLER_13_474 ();
 sg13g2_decap_4 FILLER_13_496 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_fill_2 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_593 ();
 sg13g2_fill_1 FILLER_13_600 ();
 sg13g2_decap_4 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_656 ();
 sg13g2_fill_1 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_673 ();
 sg13g2_decap_4 FILLER_13_689 ();
 sg13g2_fill_2 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_730 ();
 sg13g2_fill_1 FILLER_13_732 ();
 sg13g2_fill_1 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_768 ();
 sg13g2_fill_1 FILLER_13_775 ();
 sg13g2_fill_2 FILLER_13_794 ();
 sg13g2_fill_1 FILLER_13_796 ();
 sg13g2_decap_4 FILLER_13_807 ();
 sg13g2_fill_1 FILLER_13_829 ();
 sg13g2_fill_2 FILLER_13_837 ();
 sg13g2_fill_1 FILLER_13_839 ();
 sg13g2_fill_2 FILLER_13_847 ();
 sg13g2_fill_1 FILLER_13_849 ();
 sg13g2_decap_8 FILLER_13_862 ();
 sg13g2_decap_8 FILLER_13_869 ();
 sg13g2_decap_8 FILLER_13_876 ();
 sg13g2_fill_2 FILLER_13_910 ();
 sg13g2_fill_1 FILLER_13_912 ();
 sg13g2_decap_4 FILLER_13_938 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_fill_1 FILLER_13_1007 ();
 sg13g2_decap_8 FILLER_13_1064 ();
 sg13g2_fill_1 FILLER_13_1071 ();
 sg13g2_fill_1 FILLER_13_1075 ();
 sg13g2_decap_8 FILLER_13_1129 ();
 sg13g2_fill_2 FILLER_13_1136 ();
 sg13g2_decap_8 FILLER_13_1151 ();
 sg13g2_fill_2 FILLER_13_1158 ();
 sg13g2_fill_1 FILLER_13_1160 ();
 sg13g2_fill_1 FILLER_13_1180 ();
 sg13g2_fill_2 FILLER_13_1191 ();
 sg13g2_fill_1 FILLER_13_1199 ();
 sg13g2_decap_4 FILLER_13_1208 ();
 sg13g2_fill_2 FILLER_13_1212 ();
 sg13g2_decap_8 FILLER_13_1242 ();
 sg13g2_fill_1 FILLER_13_1249 ();
 sg13g2_fill_2 FILLER_13_1278 ();
 sg13g2_fill_1 FILLER_13_1280 ();
 sg13g2_decap_4 FILLER_13_1289 ();
 sg13g2_decap_4 FILLER_13_1315 ();
 sg13g2_fill_1 FILLER_13_1344 ();
 sg13g2_fill_2 FILLER_13_1350 ();
 sg13g2_fill_1 FILLER_13_1352 ();
 sg13g2_decap_4 FILLER_13_1358 ();
 sg13g2_fill_2 FILLER_13_1378 ();
 sg13g2_fill_1 FILLER_13_1380 ();
 sg13g2_fill_2 FILLER_13_1425 ();
 sg13g2_decap_4 FILLER_13_1437 ();
 sg13g2_fill_2 FILLER_13_1455 ();
 sg13g2_decap_8 FILLER_13_1487 ();
 sg13g2_decap_8 FILLER_13_1504 ();
 sg13g2_decap_4 FILLER_13_1511 ();
 sg13g2_decap_8 FILLER_13_1531 ();
 sg13g2_fill_2 FILLER_13_1538 ();
 sg13g2_fill_1 FILLER_13_1540 ();
 sg13g2_fill_2 FILLER_13_1554 ();
 sg13g2_fill_1 FILLER_13_1556 ();
 sg13g2_decap_4 FILLER_13_1564 ();
 sg13g2_fill_2 FILLER_13_1568 ();
 sg13g2_decap_8 FILLER_13_1587 ();
 sg13g2_fill_1 FILLER_13_1603 ();
 sg13g2_decap_8 FILLER_13_1660 ();
 sg13g2_fill_1 FILLER_13_1667 ();
 sg13g2_decap_4 FILLER_13_1677 ();
 sg13g2_fill_2 FILLER_13_1681 ();
 sg13g2_decap_4 FILLER_13_1705 ();
 sg13g2_fill_1 FILLER_13_1723 ();
 sg13g2_fill_2 FILLER_13_1737 ();
 sg13g2_fill_1 FILLER_13_1742 ();
 sg13g2_fill_2 FILLER_13_1746 ();
 sg13g2_fill_1 FILLER_13_1794 ();
 sg13g2_decap_8 FILLER_13_1802 ();
 sg13g2_decap_4 FILLER_13_1824 ();
 sg13g2_fill_2 FILLER_13_1828 ();
 sg13g2_fill_2 FILLER_13_1849 ();
 sg13g2_decap_8 FILLER_13_1856 ();
 sg13g2_fill_1 FILLER_13_1863 ();
 sg13g2_decap_8 FILLER_13_1869 ();
 sg13g2_decap_8 FILLER_13_1876 ();
 sg13g2_decap_8 FILLER_13_1883 ();
 sg13g2_fill_1 FILLER_13_1890 ();
 sg13g2_fill_2 FILLER_13_1909 ();
 sg13g2_decap_4 FILLER_13_1915 ();
 sg13g2_fill_2 FILLER_13_1919 ();
 sg13g2_fill_2 FILLER_13_1927 ();
 sg13g2_fill_1 FILLER_13_1937 ();
 sg13g2_fill_1 FILLER_13_1955 ();
 sg13g2_fill_2 FILLER_13_1964 ();
 sg13g2_fill_1 FILLER_13_1977 ();
 sg13g2_decap_4 FILLER_13_1986 ();
 sg13g2_fill_2 FILLER_13_1990 ();
 sg13g2_fill_2 FILLER_13_1997 ();
 sg13g2_fill_1 FILLER_13_2012 ();
 sg13g2_decap_4 FILLER_13_2026 ();
 sg13g2_fill_2 FILLER_13_2030 ();
 sg13g2_decap_4 FILLER_13_2041 ();
 sg13g2_fill_2 FILLER_13_2045 ();
 sg13g2_fill_1 FILLER_13_2051 ();
 sg13g2_decap_8 FILLER_13_2061 ();
 sg13g2_fill_2 FILLER_13_2068 ();
 sg13g2_fill_1 FILLER_13_2070 ();
 sg13g2_decap_8 FILLER_13_2075 ();
 sg13g2_decap_4 FILLER_13_2082 ();
 sg13g2_fill_2 FILLER_13_2086 ();
 sg13g2_fill_1 FILLER_13_2094 ();
 sg13g2_decap_8 FILLER_13_2123 ();
 sg13g2_fill_1 FILLER_13_2130 ();
 sg13g2_fill_1 FILLER_13_2135 ();
 sg13g2_decap_4 FILLER_13_2193 ();
 sg13g2_fill_2 FILLER_13_2197 ();
 sg13g2_decap_4 FILLER_13_2217 ();
 sg13g2_fill_2 FILLER_13_2221 ();
 sg13g2_decap_8 FILLER_13_2231 ();
 sg13g2_decap_8 FILLER_13_2238 ();
 sg13g2_fill_1 FILLER_13_2245 ();
 sg13g2_fill_2 FILLER_13_2255 ();
 sg13g2_fill_1 FILLER_13_2262 ();
 sg13g2_decap_4 FILLER_13_2269 ();
 sg13g2_decap_4 FILLER_13_2296 ();
 sg13g2_fill_2 FILLER_13_2300 ();
 sg13g2_decap_4 FILLER_13_2315 ();
 sg13g2_decap_8 FILLER_13_2345 ();
 sg13g2_fill_2 FILLER_13_2352 ();
 sg13g2_decap_8 FILLER_13_2360 ();
 sg13g2_fill_2 FILLER_13_2367 ();
 sg13g2_fill_1 FILLER_13_2369 ();
 sg13g2_fill_2 FILLER_13_2378 ();
 sg13g2_decap_4 FILLER_13_2394 ();
 sg13g2_decap_8 FILLER_13_2414 ();
 sg13g2_fill_1 FILLER_13_2421 ();
 sg13g2_fill_1 FILLER_13_2434 ();
 sg13g2_fill_2 FILLER_13_2446 ();
 sg13g2_fill_1 FILLER_13_2448 ();
 sg13g2_fill_2 FILLER_13_2459 ();
 sg13g2_decap_8 FILLER_13_2486 ();
 sg13g2_decap_8 FILLER_13_2493 ();
 sg13g2_fill_1 FILLER_13_2500 ();
 sg13g2_decap_4 FILLER_13_2512 ();
 sg13g2_fill_1 FILLER_13_2516 ();
 sg13g2_decap_8 FILLER_13_2528 ();
 sg13g2_fill_2 FILLER_13_2535 ();
 sg13g2_fill_1 FILLER_13_2537 ();
 sg13g2_fill_2 FILLER_13_2563 ();
 sg13g2_decap_8 FILLER_13_2587 ();
 sg13g2_fill_2 FILLER_13_2598 ();
 sg13g2_fill_2 FILLER_13_2614 ();
 sg13g2_decap_8 FILLER_13_2623 ();
 sg13g2_fill_2 FILLER_13_2630 ();
 sg13g2_fill_2 FILLER_13_2696 ();
 sg13g2_decap_4 FILLER_13_2706 ();
 sg13g2_fill_2 FILLER_13_2710 ();
 sg13g2_decap_4 FILLER_13_2751 ();
 sg13g2_decap_4 FILLER_13_2782 ();
 sg13g2_decap_8 FILLER_13_2795 ();
 sg13g2_decap_8 FILLER_13_2807 ();
 sg13g2_decap_4 FILLER_13_2814 ();
 sg13g2_fill_2 FILLER_13_2818 ();
 sg13g2_decap_4 FILLER_13_2826 ();
 sg13g2_fill_1 FILLER_13_2830 ();
 sg13g2_decap_4 FILLER_13_2874 ();
 sg13g2_fill_1 FILLER_13_2878 ();
 sg13g2_fill_2 FILLER_13_2884 ();
 sg13g2_fill_1 FILLER_13_2886 ();
 sg13g2_decap_8 FILLER_13_2898 ();
 sg13g2_decap_8 FILLER_13_2905 ();
 sg13g2_decap_8 FILLER_13_2925 ();
 sg13g2_fill_1 FILLER_13_2932 ();
 sg13g2_decap_8 FILLER_13_2937 ();
 sg13g2_fill_1 FILLER_13_2947 ();
 sg13g2_fill_2 FILLER_13_2952 ();
 sg13g2_decap_4 FILLER_13_2959 ();
 sg13g2_fill_2 FILLER_13_2963 ();
 sg13g2_decap_8 FILLER_13_2988 ();
 sg13g2_decap_8 FILLER_13_2995 ();
 sg13g2_decap_4 FILLER_13_3002 ();
 sg13g2_fill_1 FILLER_13_3013 ();
 sg13g2_fill_2 FILLER_13_3030 ();
 sg13g2_fill_1 FILLER_13_3032 ();
 sg13g2_decap_8 FILLER_13_3036 ();
 sg13g2_fill_1 FILLER_13_3043 ();
 sg13g2_fill_1 FILLER_13_3057 ();
 sg13g2_fill_1 FILLER_13_3068 ();
 sg13g2_decap_4 FILLER_13_3097 ();
 sg13g2_fill_1 FILLER_13_3101 ();
 sg13g2_decap_4 FILLER_13_3145 ();
 sg13g2_fill_1 FILLER_13_3149 ();
 sg13g2_fill_2 FILLER_13_3154 ();
 sg13g2_fill_1 FILLER_13_3165 ();
 sg13g2_fill_2 FILLER_13_3200 ();
 sg13g2_decap_8 FILLER_13_3206 ();
 sg13g2_decap_8 FILLER_13_3213 ();
 sg13g2_decap_8 FILLER_13_3220 ();
 sg13g2_decap_8 FILLER_13_3227 ();
 sg13g2_decap_8 FILLER_13_3234 ();
 sg13g2_decap_8 FILLER_13_3241 ();
 sg13g2_decap_8 FILLER_13_3248 ();
 sg13g2_decap_8 FILLER_13_3255 ();
 sg13g2_decap_8 FILLER_13_3262 ();
 sg13g2_decap_8 FILLER_13_3269 ();
 sg13g2_decap_8 FILLER_13_3276 ();
 sg13g2_decap_8 FILLER_13_3283 ();
 sg13g2_decap_8 FILLER_13_3290 ();
 sg13g2_decap_8 FILLER_13_3297 ();
 sg13g2_decap_8 FILLER_13_3304 ();
 sg13g2_decap_8 FILLER_13_3311 ();
 sg13g2_decap_8 FILLER_13_3318 ();
 sg13g2_decap_8 FILLER_13_3325 ();
 sg13g2_decap_8 FILLER_13_3332 ();
 sg13g2_decap_8 FILLER_13_3339 ();
 sg13g2_decap_8 FILLER_13_3346 ();
 sg13g2_decap_8 FILLER_13_3353 ();
 sg13g2_decap_8 FILLER_13_3360 ();
 sg13g2_decap_8 FILLER_13_3367 ();
 sg13g2_decap_8 FILLER_13_3374 ();
 sg13g2_decap_8 FILLER_13_3381 ();
 sg13g2_decap_8 FILLER_13_3388 ();
 sg13g2_decap_8 FILLER_13_3395 ();
 sg13g2_decap_8 FILLER_13_3402 ();
 sg13g2_decap_8 FILLER_13_3409 ();
 sg13g2_decap_8 FILLER_13_3416 ();
 sg13g2_decap_8 FILLER_13_3423 ();
 sg13g2_decap_8 FILLER_13_3430 ();
 sg13g2_decap_8 FILLER_13_3437 ();
 sg13g2_decap_8 FILLER_13_3444 ();
 sg13g2_decap_8 FILLER_13_3451 ();
 sg13g2_decap_8 FILLER_13_3458 ();
 sg13g2_decap_8 FILLER_13_3465 ();
 sg13g2_decap_8 FILLER_13_3472 ();
 sg13g2_decap_8 FILLER_13_3479 ();
 sg13g2_decap_8 FILLER_13_3486 ();
 sg13g2_decap_8 FILLER_13_3493 ();
 sg13g2_decap_8 FILLER_13_3500 ();
 sg13g2_decap_8 FILLER_13_3507 ();
 sg13g2_decap_8 FILLER_13_3514 ();
 sg13g2_decap_8 FILLER_13_3521 ();
 sg13g2_decap_8 FILLER_13_3528 ();
 sg13g2_decap_8 FILLER_13_3535 ();
 sg13g2_decap_8 FILLER_13_3542 ();
 sg13g2_decap_8 FILLER_13_3549 ();
 sg13g2_decap_8 FILLER_13_3556 ();
 sg13g2_decap_8 FILLER_13_3563 ();
 sg13g2_decap_8 FILLER_13_3570 ();
 sg13g2_fill_2 FILLER_13_3577 ();
 sg13g2_fill_1 FILLER_13_3579 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_fill_2 FILLER_14_338 ();
 sg13g2_fill_1 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_4 FILLER_14_413 ();
 sg13g2_fill_1 FILLER_14_417 ();
 sg13g2_fill_2 FILLER_14_426 ();
 sg13g2_fill_1 FILLER_14_428 ();
 sg13g2_fill_2 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_446 ();
 sg13g2_decap_4 FILLER_14_453 ();
 sg13g2_fill_1 FILLER_14_494 ();
 sg13g2_fill_2 FILLER_14_523 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_decap_8 FILLER_14_552 ();
 sg13g2_decap_4 FILLER_14_559 ();
 sg13g2_fill_2 FILLER_14_563 ();
 sg13g2_decap_4 FILLER_14_569 ();
 sg13g2_fill_2 FILLER_14_573 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_fill_2 FILLER_14_656 ();
 sg13g2_decap_4 FILLER_14_693 ();
 sg13g2_fill_2 FILLER_14_697 ();
 sg13g2_fill_2 FILLER_14_707 ();
 sg13g2_fill_2 FILLER_14_713 ();
 sg13g2_fill_1 FILLER_14_715 ();
 sg13g2_decap_8 FILLER_14_723 ();
 sg13g2_decap_4 FILLER_14_730 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_fill_2 FILLER_14_758 ();
 sg13g2_decap_4 FILLER_14_770 ();
 sg13g2_fill_2 FILLER_14_779 ();
 sg13g2_fill_1 FILLER_14_804 ();
 sg13g2_fill_2 FILLER_14_824 ();
 sg13g2_fill_2 FILLER_14_888 ();
 sg13g2_decap_8 FILLER_14_902 ();
 sg13g2_decap_8 FILLER_14_909 ();
 sg13g2_decap_8 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_fill_2 FILLER_14_945 ();
 sg13g2_fill_1 FILLER_14_947 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_decap_8 FILLER_14_967 ();
 sg13g2_fill_1 FILLER_14_1043 ();
 sg13g2_fill_2 FILLER_14_1065 ();
 sg13g2_fill_1 FILLER_14_1067 ();
 sg13g2_fill_2 FILLER_14_1090 ();
 sg13g2_fill_2 FILLER_14_1129 ();
 sg13g2_fill_1 FILLER_14_1170 ();
 sg13g2_decap_4 FILLER_14_1178 ();
 sg13g2_fill_1 FILLER_14_1182 ();
 sg13g2_decap_8 FILLER_14_1196 ();
 sg13g2_decap_4 FILLER_14_1203 ();
 sg13g2_fill_1 FILLER_14_1207 ();
 sg13g2_fill_2 FILLER_14_1213 ();
 sg13g2_decap_8 FILLER_14_1224 ();
 sg13g2_fill_2 FILLER_14_1231 ();
 sg13g2_fill_2 FILLER_14_1237 ();
 sg13g2_decap_8 FILLER_14_1244 ();
 sg13g2_fill_2 FILLER_14_1251 ();
 sg13g2_decap_8 FILLER_14_1264 ();
 sg13g2_fill_2 FILLER_14_1271 ();
 sg13g2_fill_1 FILLER_14_1273 ();
 sg13g2_fill_1 FILLER_14_1282 ();
 sg13g2_fill_2 FILLER_14_1288 ();
 sg13g2_fill_1 FILLER_14_1290 ();
 sg13g2_decap_8 FILLER_14_1305 ();
 sg13g2_fill_1 FILLER_14_1312 ();
 sg13g2_fill_2 FILLER_14_1331 ();
 sg13g2_decap_8 FILLER_14_1363 ();
 sg13g2_fill_1 FILLER_14_1370 ();
 sg13g2_fill_2 FILLER_14_1389 ();
 sg13g2_fill_2 FILLER_14_1409 ();
 sg13g2_decap_8 FILLER_14_1421 ();
 sg13g2_decap_4 FILLER_14_1428 ();
 sg13g2_fill_1 FILLER_14_1432 ();
 sg13g2_fill_2 FILLER_14_1440 ();
 sg13g2_fill_1 FILLER_14_1442 ();
 sg13g2_fill_2 FILLER_14_1451 ();
 sg13g2_fill_1 FILLER_14_1453 ();
 sg13g2_fill_2 FILLER_14_1467 ();
 sg13g2_fill_1 FILLER_14_1469 ();
 sg13g2_decap_4 FILLER_14_1487 ();
 sg13g2_fill_1 FILLER_14_1491 ();
 sg13g2_decap_4 FILLER_14_1534 ();
 sg13g2_fill_2 FILLER_14_1538 ();
 sg13g2_decap_4 FILLER_14_1572 ();
 sg13g2_fill_1 FILLER_14_1576 ();
 sg13g2_decap_8 FILLER_14_1605 ();
 sg13g2_decap_4 FILLER_14_1612 ();
 sg13g2_fill_1 FILLER_14_1616 ();
 sg13g2_fill_2 FILLER_14_1657 ();
 sg13g2_fill_1 FILLER_14_1659 ();
 sg13g2_decap_8 FILLER_14_1681 ();
 sg13g2_fill_2 FILLER_14_1688 ();
 sg13g2_decap_4 FILLER_14_1698 ();
 sg13g2_fill_1 FILLER_14_1730 ();
 sg13g2_fill_2 FILLER_14_1759 ();
 sg13g2_fill_2 FILLER_14_1860 ();
 sg13g2_fill_1 FILLER_14_1862 ();
 sg13g2_decap_8 FILLER_14_1884 ();
 sg13g2_decap_8 FILLER_14_1891 ();
 sg13g2_decap_8 FILLER_14_1916 ();
 sg13g2_fill_1 FILLER_14_1923 ();
 sg13g2_fill_2 FILLER_14_1947 ();
 sg13g2_fill_1 FILLER_14_1949 ();
 sg13g2_fill_1 FILLER_14_1954 ();
 sg13g2_fill_2 FILLER_14_1967 ();
 sg13g2_fill_1 FILLER_14_1985 ();
 sg13g2_decap_8 FILLER_14_1991 ();
 sg13g2_fill_2 FILLER_14_1998 ();
 sg13g2_fill_1 FILLER_14_2040 ();
 sg13g2_fill_2 FILLER_14_2069 ();
 sg13g2_fill_1 FILLER_14_2071 ();
 sg13g2_fill_1 FILLER_14_2097 ();
 sg13g2_fill_2 FILLER_14_2108 ();
 sg13g2_fill_1 FILLER_14_2134 ();
 sg13g2_decap_4 FILLER_14_2166 ();
 sg13g2_decap_8 FILLER_14_2230 ();
 sg13g2_fill_2 FILLER_14_2237 ();
 sg13g2_fill_1 FILLER_14_2257 ();
 sg13g2_decap_8 FILLER_14_2276 ();
 sg13g2_decap_4 FILLER_14_2283 ();
 sg13g2_decap_4 FILLER_14_2297 ();
 sg13g2_fill_2 FILLER_14_2319 ();
 sg13g2_decap_4 FILLER_14_2383 ();
 sg13g2_fill_1 FILLER_14_2387 ();
 sg13g2_fill_2 FILLER_14_2396 ();
 sg13g2_fill_1 FILLER_14_2398 ();
 sg13g2_decap_4 FILLER_14_2425 ();
 sg13g2_fill_2 FILLER_14_2429 ();
 sg13g2_fill_2 FILLER_14_2444 ();
 sg13g2_fill_1 FILLER_14_2446 ();
 sg13g2_decap_4 FILLER_14_2459 ();
 sg13g2_fill_2 FILLER_14_2477 ();
 sg13g2_fill_1 FILLER_14_2479 ();
 sg13g2_fill_2 FILLER_14_2510 ();
 sg13g2_decap_4 FILLER_14_2534 ();
 sg13g2_decap_4 FILLER_14_2550 ();
 sg13g2_decap_8 FILLER_14_2559 ();
 sg13g2_fill_2 FILLER_14_2566 ();
 sg13g2_fill_1 FILLER_14_2568 ();
 sg13g2_decap_8 FILLER_14_2579 ();
 sg13g2_decap_4 FILLER_14_2586 ();
 sg13g2_fill_1 FILLER_14_2624 ();
 sg13g2_fill_2 FILLER_14_2645 ();
 sg13g2_fill_1 FILLER_14_2647 ();
 sg13g2_decap_4 FILLER_14_2661 ();
 sg13g2_fill_1 FILLER_14_2665 ();
 sg13g2_fill_1 FILLER_14_2687 ();
 sg13g2_decap_8 FILLER_14_2717 ();
 sg13g2_decap_4 FILLER_14_2724 ();
 sg13g2_decap_4 FILLER_14_2732 ();
 sg13g2_fill_1 FILLER_14_2736 ();
 sg13g2_fill_1 FILLER_14_2751 ();
 sg13g2_fill_2 FILLER_14_2845 ();
 sg13g2_fill_1 FILLER_14_2847 ();
 sg13g2_decap_8 FILLER_14_2861 ();
 sg13g2_decap_4 FILLER_14_2868 ();
 sg13g2_decap_4 FILLER_14_2879 ();
 sg13g2_fill_1 FILLER_14_2883 ();
 sg13g2_decap_8 FILLER_14_2895 ();
 sg13g2_decap_4 FILLER_14_2902 ();
 sg13g2_fill_1 FILLER_14_2916 ();
 sg13g2_fill_2 FILLER_14_2937 ();
 sg13g2_decap_8 FILLER_14_2964 ();
 sg13g2_decap_4 FILLER_14_2971 ();
 sg13g2_decap_8 FILLER_14_2993 ();
 sg13g2_decap_4 FILLER_14_3000 ();
 sg13g2_fill_1 FILLER_14_3004 ();
 sg13g2_decap_8 FILLER_14_3079 ();
 sg13g2_decap_8 FILLER_14_3086 ();
 sg13g2_decap_8 FILLER_14_3093 ();
 sg13g2_fill_2 FILLER_14_3115 ();
 sg13g2_fill_1 FILLER_14_3135 ();
 sg13g2_fill_2 FILLER_14_3187 ();
 sg13g2_fill_1 FILLER_14_3189 ();
 sg13g2_decap_8 FILLER_14_3225 ();
 sg13g2_decap_8 FILLER_14_3232 ();
 sg13g2_decap_8 FILLER_14_3239 ();
 sg13g2_decap_8 FILLER_14_3246 ();
 sg13g2_decap_8 FILLER_14_3253 ();
 sg13g2_decap_8 FILLER_14_3260 ();
 sg13g2_decap_8 FILLER_14_3267 ();
 sg13g2_decap_8 FILLER_14_3274 ();
 sg13g2_decap_8 FILLER_14_3281 ();
 sg13g2_decap_8 FILLER_14_3288 ();
 sg13g2_decap_8 FILLER_14_3295 ();
 sg13g2_decap_8 FILLER_14_3302 ();
 sg13g2_decap_8 FILLER_14_3309 ();
 sg13g2_decap_8 FILLER_14_3316 ();
 sg13g2_decap_8 FILLER_14_3323 ();
 sg13g2_decap_8 FILLER_14_3330 ();
 sg13g2_decap_8 FILLER_14_3337 ();
 sg13g2_decap_8 FILLER_14_3344 ();
 sg13g2_decap_8 FILLER_14_3351 ();
 sg13g2_decap_8 FILLER_14_3358 ();
 sg13g2_decap_8 FILLER_14_3365 ();
 sg13g2_decap_8 FILLER_14_3372 ();
 sg13g2_decap_8 FILLER_14_3379 ();
 sg13g2_decap_8 FILLER_14_3386 ();
 sg13g2_decap_8 FILLER_14_3393 ();
 sg13g2_decap_8 FILLER_14_3400 ();
 sg13g2_decap_8 FILLER_14_3407 ();
 sg13g2_decap_8 FILLER_14_3414 ();
 sg13g2_decap_8 FILLER_14_3421 ();
 sg13g2_decap_8 FILLER_14_3428 ();
 sg13g2_decap_8 FILLER_14_3435 ();
 sg13g2_decap_8 FILLER_14_3442 ();
 sg13g2_decap_8 FILLER_14_3449 ();
 sg13g2_decap_8 FILLER_14_3456 ();
 sg13g2_decap_8 FILLER_14_3463 ();
 sg13g2_decap_8 FILLER_14_3470 ();
 sg13g2_decap_8 FILLER_14_3477 ();
 sg13g2_decap_8 FILLER_14_3484 ();
 sg13g2_decap_8 FILLER_14_3491 ();
 sg13g2_decap_8 FILLER_14_3498 ();
 sg13g2_decap_8 FILLER_14_3505 ();
 sg13g2_decap_8 FILLER_14_3512 ();
 sg13g2_decap_8 FILLER_14_3519 ();
 sg13g2_decap_8 FILLER_14_3526 ();
 sg13g2_decap_8 FILLER_14_3533 ();
 sg13g2_decap_8 FILLER_14_3540 ();
 sg13g2_decap_8 FILLER_14_3547 ();
 sg13g2_decap_8 FILLER_14_3554 ();
 sg13g2_decap_8 FILLER_14_3561 ();
 sg13g2_decap_8 FILLER_14_3568 ();
 sg13g2_decap_4 FILLER_14_3575 ();
 sg13g2_fill_1 FILLER_14_3579 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_4 FILLER_15_294 ();
 sg13g2_decap_4 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_339 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_fill_1 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_513 ();
 sg13g2_decap_4 FILLER_15_520 ();
 sg13g2_decap_8 FILLER_15_552 ();
 sg13g2_decap_4 FILLER_15_559 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_fill_1 FILLER_15_603 ();
 sg13g2_decap_4 FILLER_15_622 ();
 sg13g2_fill_2 FILLER_15_626 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_decap_4 FILLER_15_639 ();
 sg13g2_fill_1 FILLER_15_643 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_fill_1 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_681 ();
 sg13g2_decap_4 FILLER_15_688 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_fill_2 FILLER_15_759 ();
 sg13g2_fill_1 FILLER_15_761 ();
 sg13g2_fill_2 FILLER_15_781 ();
 sg13g2_decap_4 FILLER_15_792 ();
 sg13g2_fill_1 FILLER_15_825 ();
 sg13g2_fill_1 FILLER_15_837 ();
 sg13g2_decap_4 FILLER_15_860 ();
 sg13g2_fill_1 FILLER_15_864 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_fill_1 FILLER_15_883 ();
 sg13g2_decap_8 FILLER_15_896 ();
 sg13g2_decap_8 FILLER_15_903 ();
 sg13g2_fill_1 FILLER_15_910 ();
 sg13g2_fill_2 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_933 ();
 sg13g2_fill_2 FILLER_15_944 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_fill_2 FILLER_15_973 ();
 sg13g2_fill_1 FILLER_15_975 ();
 sg13g2_decap_4 FILLER_15_988 ();
 sg13g2_fill_1 FILLER_15_1051 ();
 sg13g2_fill_2 FILLER_15_1065 ();
 sg13g2_fill_2 FILLER_15_1072 ();
 sg13g2_fill_2 FILLER_15_1087 ();
 sg13g2_decap_8 FILLER_15_1093 ();
 sg13g2_fill_2 FILLER_15_1100 ();
 sg13g2_fill_1 FILLER_15_1102 ();
 sg13g2_fill_1 FILLER_15_1106 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_fill_1 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1168 ();
 sg13g2_fill_2 FILLER_15_1175 ();
 sg13g2_fill_1 FILLER_15_1177 ();
 sg13g2_fill_1 FILLER_15_1189 ();
 sg13g2_fill_2 FILLER_15_1196 ();
 sg13g2_fill_2 FILLER_15_1205 ();
 sg13g2_fill_1 FILLER_15_1221 ();
 sg13g2_decap_8 FILLER_15_1235 ();
 sg13g2_decap_4 FILLER_15_1242 ();
 sg13g2_fill_2 FILLER_15_1274 ();
 sg13g2_fill_2 FILLER_15_1285 ();
 sg13g2_fill_1 FILLER_15_1287 ();
 sg13g2_fill_2 FILLER_15_1309 ();
 sg13g2_fill_2 FILLER_15_1338 ();
 sg13g2_fill_1 FILLER_15_1348 ();
 sg13g2_decap_8 FILLER_15_1354 ();
 sg13g2_fill_2 FILLER_15_1382 ();
 sg13g2_fill_2 FILLER_15_1391 ();
 sg13g2_decap_8 FILLER_15_1418 ();
 sg13g2_fill_2 FILLER_15_1425 ();
 sg13g2_fill_1 FILLER_15_1427 ();
 sg13g2_fill_2 FILLER_15_1459 ();
 sg13g2_decap_4 FILLER_15_1482 ();
 sg13g2_decap_4 FILLER_15_1514 ();
 sg13g2_fill_2 FILLER_15_1518 ();
 sg13g2_fill_2 FILLER_15_1537 ();
 sg13g2_fill_1 FILLER_15_1539 ();
 sg13g2_fill_2 FILLER_15_1548 ();
 sg13g2_decap_4 FILLER_15_1561 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_fill_1 FILLER_15_1582 ();
 sg13g2_decap_8 FILLER_15_1587 ();
 sg13g2_decap_8 FILLER_15_1594 ();
 sg13g2_fill_2 FILLER_15_1601 ();
 sg13g2_fill_1 FILLER_15_1603 ();
 sg13g2_fill_2 FILLER_15_1617 ();
 sg13g2_fill_1 FILLER_15_1619 ();
 sg13g2_fill_2 FILLER_15_1627 ();
 sg13g2_fill_1 FILLER_15_1629 ();
 sg13g2_fill_2 FILLER_15_1643 ();
 sg13g2_decap_8 FILLER_15_1660 ();
 sg13g2_fill_2 FILLER_15_1667 ();
 sg13g2_fill_1 FILLER_15_1669 ();
 sg13g2_decap_8 FILLER_15_1690 ();
 sg13g2_fill_1 FILLER_15_1697 ();
 sg13g2_fill_1 FILLER_15_1703 ();
 sg13g2_fill_2 FILLER_15_1715 ();
 sg13g2_fill_1 FILLER_15_1717 ();
 sg13g2_decap_4 FILLER_15_1721 ();
 sg13g2_fill_2 FILLER_15_1725 ();
 sg13g2_decap_8 FILLER_15_1732 ();
 sg13g2_fill_2 FILLER_15_1739 ();
 sg13g2_decap_8 FILLER_15_1797 ();
 sg13g2_decap_4 FILLER_15_1804 ();
 sg13g2_fill_2 FILLER_15_1808 ();
 sg13g2_fill_2 FILLER_15_1836 ();
 sg13g2_fill_2 FILLER_15_1861 ();
 sg13g2_decap_8 FILLER_15_1867 ();
 sg13g2_fill_1 FILLER_15_1874 ();
 sg13g2_fill_1 FILLER_15_1912 ();
 sg13g2_decap_8 FILLER_15_1918 ();
 sg13g2_fill_2 FILLER_15_1925 ();
 sg13g2_fill_1 FILLER_15_1927 ();
 sg13g2_fill_2 FILLER_15_1933 ();
 sg13g2_decap_8 FILLER_15_1944 ();
 sg13g2_decap_4 FILLER_15_1951 ();
 sg13g2_fill_2 FILLER_15_1955 ();
 sg13g2_fill_2 FILLER_15_1962 ();
 sg13g2_fill_1 FILLER_15_1964 ();
 sg13g2_fill_1 FILLER_15_1970 ();
 sg13g2_decap_8 FILLER_15_1977 ();
 sg13g2_fill_1 FILLER_15_1984 ();
 sg13g2_decap_4 FILLER_15_1993 ();
 sg13g2_fill_1 FILLER_15_1997 ();
 sg13g2_fill_2 FILLER_15_2013 ();
 sg13g2_fill_1 FILLER_15_2015 ();
 sg13g2_decap_8 FILLER_15_2042 ();
 sg13g2_decap_8 FILLER_15_2049 ();
 sg13g2_decap_8 FILLER_15_2056 ();
 sg13g2_fill_2 FILLER_15_2063 ();
 sg13g2_fill_1 FILLER_15_2065 ();
 sg13g2_fill_2 FILLER_15_2163 ();
 sg13g2_decap_8 FILLER_15_2191 ();
 sg13g2_fill_2 FILLER_15_2202 ();
 sg13g2_fill_2 FILLER_15_2217 ();
 sg13g2_fill_1 FILLER_15_2219 ();
 sg13g2_fill_1 FILLER_15_2237 ();
 sg13g2_fill_2 FILLER_15_2251 ();
 sg13g2_decap_4 FILLER_15_2265 ();
 sg13g2_decap_8 FILLER_15_2274 ();
 sg13g2_decap_8 FILLER_15_2281 ();
 sg13g2_decap_4 FILLER_15_2288 ();
 sg13g2_fill_2 FILLER_15_2302 ();
 sg13g2_decap_8 FILLER_15_2309 ();
 sg13g2_decap_4 FILLER_15_2316 ();
 sg13g2_fill_2 FILLER_15_2320 ();
 sg13g2_decap_8 FILLER_15_2344 ();
 sg13g2_fill_1 FILLER_15_2351 ();
 sg13g2_decap_4 FILLER_15_2367 ();
 sg13g2_decap_8 FILLER_15_2379 ();
 sg13g2_decap_8 FILLER_15_2386 ();
 sg13g2_decap_4 FILLER_15_2428 ();
 sg13g2_fill_2 FILLER_15_2432 ();
 sg13g2_decap_8 FILLER_15_2467 ();
 sg13g2_fill_2 FILLER_15_2474 ();
 sg13g2_decap_8 FILLER_15_2489 ();
 sg13g2_decap_8 FILLER_15_2496 ();
 sg13g2_decap_4 FILLER_15_2503 ();
 sg13g2_fill_1 FILLER_15_2507 ();
 sg13g2_fill_2 FILLER_15_2521 ();
 sg13g2_decap_4 FILLER_15_2532 ();
 sg13g2_fill_1 FILLER_15_2541 ();
 sg13g2_decap_4 FILLER_15_2550 ();
 sg13g2_fill_1 FILLER_15_2554 ();
 sg13g2_fill_2 FILLER_15_2560 ();
 sg13g2_decap_4 FILLER_15_2573 ();
 sg13g2_fill_2 FILLER_15_2577 ();
 sg13g2_decap_8 FILLER_15_2583 ();
 sg13g2_fill_2 FILLER_15_2590 ();
 sg13g2_decap_8 FILLER_15_2608 ();
 sg13g2_fill_2 FILLER_15_2615 ();
 sg13g2_fill_1 FILLER_15_2617 ();
 sg13g2_decap_4 FILLER_15_2639 ();
 sg13g2_decap_8 FILLER_15_2659 ();
 sg13g2_decap_4 FILLER_15_2666 ();
 sg13g2_decap_8 FILLER_15_2688 ();
 sg13g2_decap_8 FILLER_15_2695 ();
 sg13g2_fill_1 FILLER_15_2702 ();
 sg13g2_decap_8 FILLER_15_2706 ();
 sg13g2_decap_4 FILLER_15_2713 ();
 sg13g2_fill_1 FILLER_15_2717 ();
 sg13g2_decap_4 FILLER_15_2734 ();
 sg13g2_fill_2 FILLER_15_2743 ();
 sg13g2_fill_2 FILLER_15_2780 ();
 sg13g2_fill_1 FILLER_15_2786 ();
 sg13g2_decap_4 FILLER_15_2796 ();
 sg13g2_fill_1 FILLER_15_2800 ();
 sg13g2_decap_4 FILLER_15_2804 ();
 sg13g2_decap_8 FILLER_15_2812 ();
 sg13g2_fill_1 FILLER_15_2819 ();
 sg13g2_decap_8 FILLER_15_2836 ();
 sg13g2_fill_2 FILLER_15_2843 ();
 sg13g2_decap_4 FILLER_15_2873 ();
 sg13g2_fill_2 FILLER_15_2877 ();
 sg13g2_fill_1 FILLER_15_2907 ();
 sg13g2_fill_1 FILLER_15_2913 ();
 sg13g2_decap_4 FILLER_15_2922 ();
 sg13g2_fill_1 FILLER_15_2926 ();
 sg13g2_decap_4 FILLER_15_2946 ();
 sg13g2_fill_1 FILLER_15_2957 ();
 sg13g2_decap_8 FILLER_15_2970 ();
 sg13g2_fill_1 FILLER_15_2977 ();
 sg13g2_fill_1 FILLER_15_2983 ();
 sg13g2_decap_4 FILLER_15_3016 ();
 sg13g2_fill_2 FILLER_15_3039 ();
 sg13g2_decap_8 FILLER_15_3050 ();
 sg13g2_decap_4 FILLER_15_3057 ();
 sg13g2_decap_4 FILLER_15_3066 ();
 sg13g2_fill_2 FILLER_15_3070 ();
 sg13g2_fill_2 FILLER_15_3076 ();
 sg13g2_decap_4 FILLER_15_3099 ();
 sg13g2_fill_2 FILLER_15_3110 ();
 sg13g2_fill_1 FILLER_15_3112 ();
 sg13g2_fill_1 FILLER_15_3129 ();
 sg13g2_fill_2 FILLER_15_3146 ();
 sg13g2_decap_4 FILLER_15_3163 ();
 sg13g2_fill_2 FILLER_15_3167 ();
 sg13g2_fill_1 FILLER_15_3187 ();
 sg13g2_decap_8 FILLER_15_3209 ();
 sg13g2_decap_8 FILLER_15_3216 ();
 sg13g2_decap_8 FILLER_15_3223 ();
 sg13g2_decap_8 FILLER_15_3230 ();
 sg13g2_fill_2 FILLER_15_3237 ();
 sg13g2_decap_8 FILLER_15_3246 ();
 sg13g2_decap_8 FILLER_15_3253 ();
 sg13g2_decap_8 FILLER_15_3260 ();
 sg13g2_decap_8 FILLER_15_3267 ();
 sg13g2_decap_8 FILLER_15_3274 ();
 sg13g2_decap_8 FILLER_15_3281 ();
 sg13g2_decap_8 FILLER_15_3288 ();
 sg13g2_decap_8 FILLER_15_3295 ();
 sg13g2_decap_8 FILLER_15_3302 ();
 sg13g2_decap_8 FILLER_15_3309 ();
 sg13g2_decap_8 FILLER_15_3316 ();
 sg13g2_decap_8 FILLER_15_3323 ();
 sg13g2_decap_8 FILLER_15_3330 ();
 sg13g2_decap_8 FILLER_15_3337 ();
 sg13g2_decap_8 FILLER_15_3344 ();
 sg13g2_decap_8 FILLER_15_3351 ();
 sg13g2_decap_8 FILLER_15_3358 ();
 sg13g2_decap_8 FILLER_15_3365 ();
 sg13g2_decap_8 FILLER_15_3372 ();
 sg13g2_decap_8 FILLER_15_3379 ();
 sg13g2_decap_8 FILLER_15_3386 ();
 sg13g2_decap_8 FILLER_15_3393 ();
 sg13g2_decap_8 FILLER_15_3400 ();
 sg13g2_decap_8 FILLER_15_3407 ();
 sg13g2_decap_8 FILLER_15_3414 ();
 sg13g2_decap_8 FILLER_15_3421 ();
 sg13g2_decap_8 FILLER_15_3428 ();
 sg13g2_decap_8 FILLER_15_3435 ();
 sg13g2_decap_8 FILLER_15_3442 ();
 sg13g2_decap_8 FILLER_15_3449 ();
 sg13g2_decap_8 FILLER_15_3456 ();
 sg13g2_decap_8 FILLER_15_3463 ();
 sg13g2_decap_8 FILLER_15_3470 ();
 sg13g2_decap_8 FILLER_15_3477 ();
 sg13g2_decap_8 FILLER_15_3484 ();
 sg13g2_decap_8 FILLER_15_3491 ();
 sg13g2_decap_8 FILLER_15_3498 ();
 sg13g2_decap_8 FILLER_15_3505 ();
 sg13g2_decap_8 FILLER_15_3512 ();
 sg13g2_decap_8 FILLER_15_3519 ();
 sg13g2_decap_8 FILLER_15_3526 ();
 sg13g2_decap_8 FILLER_15_3533 ();
 sg13g2_decap_8 FILLER_15_3540 ();
 sg13g2_decap_8 FILLER_15_3547 ();
 sg13g2_decap_8 FILLER_15_3554 ();
 sg13g2_decap_8 FILLER_15_3561 ();
 sg13g2_decap_8 FILLER_15_3568 ();
 sg13g2_decap_4 FILLER_15_3575 ();
 sg13g2_fill_1 FILLER_15_3579 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_338 ();
 sg13g2_fill_1 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_fill_2 FILLER_16_375 ();
 sg13g2_fill_1 FILLER_16_377 ();
 sg13g2_fill_1 FILLER_16_392 ();
 sg13g2_decap_4 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_16_415 ();
 sg13g2_decap_4 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_16_432 ();
 sg13g2_fill_2 FILLER_16_443 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_8 FILLER_16_464 ();
 sg13g2_decap_4 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_495 ();
 sg13g2_decap_8 FILLER_16_502 ();
 sg13g2_fill_1 FILLER_16_509 ();
 sg13g2_fill_1 FILLER_16_514 ();
 sg13g2_decap_4 FILLER_16_533 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_fill_2 FILLER_16_567 ();
 sg13g2_fill_1 FILLER_16_569 ();
 sg13g2_decap_4 FILLER_16_598 ();
 sg13g2_fill_1 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_635 ();
 sg13g2_decap_4 FILLER_16_670 ();
 sg13g2_fill_2 FILLER_16_674 ();
 sg13g2_fill_1 FILLER_16_718 ();
 sg13g2_fill_2 FILLER_16_728 ();
 sg13g2_decap_4 FILLER_16_743 ();
 sg13g2_fill_1 FILLER_16_747 ();
 sg13g2_fill_2 FILLER_16_756 ();
 sg13g2_fill_1 FILLER_16_758 ();
 sg13g2_decap_4 FILLER_16_792 ();
 sg13g2_fill_1 FILLER_16_796 ();
 sg13g2_fill_2 FILLER_16_816 ();
 sg13g2_fill_1 FILLER_16_826 ();
 sg13g2_fill_2 FILLER_16_870 ();
 sg13g2_fill_1 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_880 ();
 sg13g2_fill_2 FILLER_16_887 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_4 FILLER_16_899 ();
 sg13g2_fill_1 FILLER_16_903 ();
 sg13g2_fill_2 FILLER_16_935 ();
 sg13g2_fill_1 FILLER_16_937 ();
 sg13g2_fill_2 FILLER_16_951 ();
 sg13g2_fill_2 FILLER_16_971 ();
 sg13g2_fill_1 FILLER_16_973 ();
 sg13g2_fill_1 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_993 ();
 sg13g2_decap_8 FILLER_16_1000 ();
 sg13g2_fill_1 FILLER_16_1007 ();
 sg13g2_decap_4 FILLER_16_1017 ();
 sg13g2_fill_2 FILLER_16_1021 ();
 sg13g2_fill_2 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_decap_4 FILLER_16_1036 ();
 sg13g2_fill_2 FILLER_16_1040 ();
 sg13g2_decap_8 FILLER_16_1053 ();
 sg13g2_fill_2 FILLER_16_1060 ();
 sg13g2_fill_1 FILLER_16_1062 ();
 sg13g2_fill_1 FILLER_16_1067 ();
 sg13g2_decap_8 FILLER_16_1089 ();
 sg13g2_fill_2 FILLER_16_1096 ();
 sg13g2_fill_1 FILLER_16_1098 ();
 sg13g2_fill_2 FILLER_16_1120 ();
 sg13g2_fill_1 FILLER_16_1122 ();
 sg13g2_fill_2 FILLER_16_1136 ();
 sg13g2_decap_8 FILLER_16_1159 ();
 sg13g2_decap_4 FILLER_16_1166 ();
 sg13g2_fill_1 FILLER_16_1170 ();
 sg13g2_decap_4 FILLER_16_1176 ();
 sg13g2_fill_2 FILLER_16_1180 ();
 sg13g2_fill_2 FILLER_16_1200 ();
 sg13g2_decap_4 FILLER_16_1209 ();
 sg13g2_fill_1 FILLER_16_1213 ();
 sg13g2_decap_8 FILLER_16_1244 ();
 sg13g2_decap_8 FILLER_16_1255 ();
 sg13g2_fill_1 FILLER_16_1262 ();
 sg13g2_fill_2 FILLER_16_1293 ();
 sg13g2_decap_8 FILLER_16_1353 ();
 sg13g2_decap_8 FILLER_16_1360 ();
 sg13g2_fill_2 FILLER_16_1367 ();
 sg13g2_fill_1 FILLER_16_1369 ();
 sg13g2_decap_8 FILLER_16_1388 ();
 sg13g2_fill_1 FILLER_16_1395 ();
 sg13g2_decap_8 FILLER_16_1424 ();
 sg13g2_fill_2 FILLER_16_1459 ();
 sg13g2_fill_1 FILLER_16_1461 ();
 sg13g2_decap_8 FILLER_16_1478 ();
 sg13g2_fill_1 FILLER_16_1485 ();
 sg13g2_decap_8 FILLER_16_1507 ();
 sg13g2_decap_4 FILLER_16_1514 ();
 sg13g2_fill_2 FILLER_16_1518 ();
 sg13g2_decap_8 FILLER_16_1535 ();
 sg13g2_fill_1 FILLER_16_1542 ();
 sg13g2_fill_1 FILLER_16_1591 ();
 sg13g2_decap_8 FILLER_16_1643 ();
 sg13g2_fill_1 FILLER_16_1650 ();
 sg13g2_fill_1 FILLER_16_1674 ();
 sg13g2_decap_8 FILLER_16_1685 ();
 sg13g2_decap_4 FILLER_16_1692 ();
 sg13g2_fill_2 FILLER_16_1696 ();
 sg13g2_fill_2 FILLER_16_1706 ();
 sg13g2_fill_1 FILLER_16_1708 ();
 sg13g2_decap_4 FILLER_16_1752 ();
 sg13g2_fill_2 FILLER_16_1756 ();
 sg13g2_decap_8 FILLER_16_1800 ();
 sg13g2_decap_8 FILLER_16_1807 ();
 sg13g2_fill_2 FILLER_16_1814 ();
 sg13g2_fill_1 FILLER_16_1829 ();
 sg13g2_fill_1 FILLER_16_1868 ();
 sg13g2_decap_4 FILLER_16_1884 ();
 sg13g2_fill_1 FILLER_16_1888 ();
 sg13g2_decap_8 FILLER_16_1893 ();
 sg13g2_fill_2 FILLER_16_1904 ();
 sg13g2_fill_1 FILLER_16_1906 ();
 sg13g2_fill_2 FILLER_16_1916 ();
 sg13g2_fill_2 FILLER_16_1930 ();
 sg13g2_fill_1 FILLER_16_1932 ();
 sg13g2_decap_4 FILLER_16_1953 ();
 sg13g2_fill_1 FILLER_16_1981 ();
 sg13g2_decap_8 FILLER_16_1991 ();
 sg13g2_decap_4 FILLER_16_1998 ();
 sg13g2_fill_1 FILLER_16_2033 ();
 sg13g2_decap_4 FILLER_16_2069 ();
 sg13g2_fill_1 FILLER_16_2073 ();
 sg13g2_decap_8 FILLER_16_2100 ();
 sg13g2_decap_4 FILLER_16_2107 ();
 sg13g2_decap_8 FILLER_16_2115 ();
 sg13g2_decap_4 FILLER_16_2122 ();
 sg13g2_fill_2 FILLER_16_2126 ();
 sg13g2_fill_2 FILLER_16_2132 ();
 sg13g2_fill_2 FILLER_16_2152 ();
 sg13g2_fill_2 FILLER_16_2176 ();
 sg13g2_fill_2 FILLER_16_2194 ();
 sg13g2_decap_8 FILLER_16_2200 ();
 sg13g2_fill_2 FILLER_16_2240 ();
 sg13g2_fill_1 FILLER_16_2242 ();
 sg13g2_fill_2 FILLER_16_2262 ();
 sg13g2_fill_2 FILLER_16_2282 ();
 sg13g2_decap_8 FILLER_16_2312 ();
 sg13g2_decap_4 FILLER_16_2319 ();
 sg13g2_fill_1 FILLER_16_2323 ();
 sg13g2_decap_8 FILLER_16_2336 ();
 sg13g2_decap_8 FILLER_16_2343 ();
 sg13g2_decap_8 FILLER_16_2350 ();
 sg13g2_decap_8 FILLER_16_2357 ();
 sg13g2_fill_1 FILLER_16_2364 ();
 sg13g2_decap_8 FILLER_16_2393 ();
 sg13g2_decap_4 FILLER_16_2417 ();
 sg13g2_decap_4 FILLER_16_2425 ();
 sg13g2_decap_8 FILLER_16_2442 ();
 sg13g2_decap_4 FILLER_16_2449 ();
 sg13g2_fill_2 FILLER_16_2459 ();
 sg13g2_fill_2 FILLER_16_2470 ();
 sg13g2_fill_1 FILLER_16_2472 ();
 sg13g2_decap_4 FILLER_16_2491 ();
 sg13g2_fill_2 FILLER_16_2495 ();
 sg13g2_fill_2 FILLER_16_2502 ();
 sg13g2_fill_2 FILLER_16_2517 ();
 sg13g2_fill_1 FILLER_16_2519 ();
 sg13g2_decap_8 FILLER_16_2537 ();
 sg13g2_decap_4 FILLER_16_2544 ();
 sg13g2_fill_2 FILLER_16_2548 ();
 sg13g2_fill_2 FILLER_16_2572 ();
 sg13g2_fill_2 FILLER_16_2602 ();
 sg13g2_decap_4 FILLER_16_2617 ();
 sg13g2_fill_1 FILLER_16_2621 ();
 sg13g2_fill_1 FILLER_16_2663 ();
 sg13g2_decap_4 FILLER_16_2668 ();
 sg13g2_fill_1 FILLER_16_2672 ();
 sg13g2_fill_1 FILLER_16_2686 ();
 sg13g2_fill_2 FILLER_16_2709 ();
 sg13g2_decap_4 FILLER_16_2747 ();
 sg13g2_fill_1 FILLER_16_2751 ();
 sg13g2_fill_2 FILLER_16_2802 ();
 sg13g2_decap_8 FILLER_16_2814 ();
 sg13g2_fill_2 FILLER_16_2821 ();
 sg13g2_fill_2 FILLER_16_2855 ();
 sg13g2_decap_8 FILLER_16_2870 ();
 sg13g2_fill_2 FILLER_16_2877 ();
 sg13g2_decap_8 FILLER_16_2892 ();
 sg13g2_decap_4 FILLER_16_2899 ();
 sg13g2_decap_8 FILLER_16_2921 ();
 sg13g2_decap_4 FILLER_16_2928 ();
 sg13g2_fill_1 FILLER_16_2932 ();
 sg13g2_fill_2 FILLER_16_2951 ();
 sg13g2_fill_1 FILLER_16_2953 ();
 sg13g2_fill_1 FILLER_16_2959 ();
 sg13g2_decap_8 FILLER_16_2983 ();
 sg13g2_decap_4 FILLER_16_2990 ();
 sg13g2_fill_1 FILLER_16_2994 ();
 sg13g2_decap_8 FILLER_16_2999 ();
 sg13g2_decap_8 FILLER_16_3006 ();
 sg13g2_fill_2 FILLER_16_3013 ();
 sg13g2_fill_1 FILLER_16_3015 ();
 sg13g2_decap_8 FILLER_16_3022 ();
 sg13g2_decap_8 FILLER_16_3029 ();
 sg13g2_fill_1 FILLER_16_3036 ();
 sg13g2_fill_2 FILLER_16_3055 ();
 sg13g2_decap_8 FILLER_16_3070 ();
 sg13g2_decap_4 FILLER_16_3077 ();
 sg13g2_fill_2 FILLER_16_3081 ();
 sg13g2_decap_8 FILLER_16_3099 ();
 sg13g2_fill_1 FILLER_16_3106 ();
 sg13g2_decap_4 FILLER_16_3112 ();
 sg13g2_decap_8 FILLER_16_3131 ();
 sg13g2_fill_1 FILLER_16_3138 ();
 sg13g2_decap_8 FILLER_16_3144 ();
 sg13g2_decap_4 FILLER_16_3151 ();
 sg13g2_decap_8 FILLER_16_3160 ();
 sg13g2_fill_2 FILLER_16_3167 ();
 sg13g2_fill_1 FILLER_16_3169 ();
 sg13g2_fill_2 FILLER_16_3219 ();
 sg13g2_fill_1 FILLER_16_3225 ();
 sg13g2_decap_8 FILLER_16_3254 ();
 sg13g2_decap_8 FILLER_16_3261 ();
 sg13g2_decap_8 FILLER_16_3268 ();
 sg13g2_decap_8 FILLER_16_3275 ();
 sg13g2_decap_8 FILLER_16_3282 ();
 sg13g2_decap_8 FILLER_16_3289 ();
 sg13g2_decap_8 FILLER_16_3296 ();
 sg13g2_decap_8 FILLER_16_3303 ();
 sg13g2_decap_8 FILLER_16_3310 ();
 sg13g2_decap_8 FILLER_16_3317 ();
 sg13g2_decap_8 FILLER_16_3324 ();
 sg13g2_decap_8 FILLER_16_3331 ();
 sg13g2_decap_8 FILLER_16_3338 ();
 sg13g2_decap_8 FILLER_16_3345 ();
 sg13g2_decap_8 FILLER_16_3352 ();
 sg13g2_decap_8 FILLER_16_3359 ();
 sg13g2_decap_8 FILLER_16_3366 ();
 sg13g2_decap_8 FILLER_16_3373 ();
 sg13g2_decap_8 FILLER_16_3380 ();
 sg13g2_decap_8 FILLER_16_3387 ();
 sg13g2_decap_8 FILLER_16_3394 ();
 sg13g2_decap_8 FILLER_16_3401 ();
 sg13g2_decap_8 FILLER_16_3408 ();
 sg13g2_decap_8 FILLER_16_3415 ();
 sg13g2_decap_8 FILLER_16_3422 ();
 sg13g2_decap_8 FILLER_16_3429 ();
 sg13g2_decap_8 FILLER_16_3436 ();
 sg13g2_decap_8 FILLER_16_3443 ();
 sg13g2_decap_8 FILLER_16_3450 ();
 sg13g2_decap_8 FILLER_16_3457 ();
 sg13g2_decap_8 FILLER_16_3464 ();
 sg13g2_decap_8 FILLER_16_3471 ();
 sg13g2_decap_8 FILLER_16_3478 ();
 sg13g2_decap_8 FILLER_16_3485 ();
 sg13g2_decap_8 FILLER_16_3492 ();
 sg13g2_decap_8 FILLER_16_3499 ();
 sg13g2_decap_8 FILLER_16_3506 ();
 sg13g2_decap_8 FILLER_16_3513 ();
 sg13g2_decap_8 FILLER_16_3520 ();
 sg13g2_decap_8 FILLER_16_3527 ();
 sg13g2_decap_8 FILLER_16_3534 ();
 sg13g2_decap_8 FILLER_16_3541 ();
 sg13g2_decap_8 FILLER_16_3548 ();
 sg13g2_decap_8 FILLER_16_3555 ();
 sg13g2_decap_8 FILLER_16_3562 ();
 sg13g2_decap_8 FILLER_16_3569 ();
 sg13g2_decap_4 FILLER_16_3576 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_447 ();
 sg13g2_decap_8 FILLER_17_463 ();
 sg13g2_fill_2 FILLER_17_470 ();
 sg13g2_fill_2 FILLER_17_487 ();
 sg13g2_fill_1 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_555 ();
 sg13g2_fill_1 FILLER_17_562 ();
 sg13g2_fill_2 FILLER_17_572 ();
 sg13g2_fill_1 FILLER_17_574 ();
 sg13g2_fill_1 FILLER_17_579 ();
 sg13g2_decap_8 FILLER_17_587 ();
 sg13g2_decap_8 FILLER_17_594 ();
 sg13g2_fill_2 FILLER_17_614 ();
 sg13g2_fill_1 FILLER_17_616 ();
 sg13g2_decap_4 FILLER_17_642 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_fill_2 FILLER_17_663 ();
 sg13g2_fill_2 FILLER_17_678 ();
 sg13g2_fill_1 FILLER_17_680 ();
 sg13g2_decap_4 FILLER_17_692 ();
 sg13g2_fill_1 FILLER_17_696 ();
 sg13g2_fill_2 FILLER_17_709 ();
 sg13g2_fill_1 FILLER_17_732 ();
 sg13g2_decap_4 FILLER_17_737 ();
 sg13g2_decap_8 FILLER_17_754 ();
 sg13g2_decap_4 FILLER_17_761 ();
 sg13g2_fill_2 FILLER_17_765 ();
 sg13g2_decap_8 FILLER_17_789 ();
 sg13g2_decap_8 FILLER_17_811 ();
 sg13g2_decap_4 FILLER_17_825 ();
 sg13g2_decap_8 FILLER_17_919 ();
 sg13g2_decap_8 FILLER_17_926 ();
 sg13g2_decap_8 FILLER_17_933 ();
 sg13g2_decap_4 FILLER_17_952 ();
 sg13g2_fill_2 FILLER_17_956 ();
 sg13g2_fill_1 FILLER_17_976 ();
 sg13g2_decap_4 FILLER_17_999 ();
 sg13g2_fill_1 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1026 ();
 sg13g2_decap_4 FILLER_17_1033 ();
 sg13g2_decap_4 FILLER_17_1059 ();
 sg13g2_fill_2 FILLER_17_1078 ();
 sg13g2_fill_1 FILLER_17_1080 ();
 sg13g2_decap_8 FILLER_17_1091 ();
 sg13g2_fill_1 FILLER_17_1175 ();
 sg13g2_fill_2 FILLER_17_1198 ();
 sg13g2_fill_2 FILLER_17_1209 ();
 sg13g2_fill_1 FILLER_17_1229 ();
 sg13g2_fill_2 FILLER_17_1263 ();
 sg13g2_fill_2 FILLER_17_1290 ();
 sg13g2_fill_2 FILLER_17_1321 ();
 sg13g2_fill_1 FILLER_17_1336 ();
 sg13g2_fill_2 FILLER_17_1346 ();
 sg13g2_fill_2 FILLER_17_1386 ();
 sg13g2_fill_1 FILLER_17_1388 ();
 sg13g2_fill_1 FILLER_17_1405 ();
 sg13g2_fill_2 FILLER_17_1446 ();
 sg13g2_fill_1 FILLER_17_1448 ();
 sg13g2_fill_2 FILLER_17_1462 ();
 sg13g2_decap_4 FILLER_17_1474 ();
 sg13g2_fill_1 FILLER_17_1478 ();
 sg13g2_decap_8 FILLER_17_1507 ();
 sg13g2_decap_8 FILLER_17_1514 ();
 sg13g2_decap_4 FILLER_17_1574 ();
 sg13g2_fill_1 FILLER_17_1578 ();
 sg13g2_decap_4 FILLER_17_1633 ();
 sg13g2_fill_2 FILLER_17_1637 ();
 sg13g2_decap_8 FILLER_17_1696 ();
 sg13g2_decap_8 FILLER_17_1703 ();
 sg13g2_decap_4 FILLER_17_1710 ();
 sg13g2_fill_2 FILLER_17_1714 ();
 sg13g2_fill_1 FILLER_17_1728 ();
 sg13g2_decap_8 FILLER_17_1733 ();
 sg13g2_decap_8 FILLER_17_1740 ();
 sg13g2_decap_8 FILLER_17_1747 ();
 sg13g2_fill_1 FILLER_17_1754 ();
 sg13g2_fill_1 FILLER_17_1763 ();
 sg13g2_decap_4 FILLER_17_1769 ();
 sg13g2_fill_2 FILLER_17_1773 ();
 sg13g2_fill_2 FILLER_17_1788 ();
 sg13g2_fill_2 FILLER_17_1803 ();
 sg13g2_fill_1 FILLER_17_1805 ();
 sg13g2_fill_1 FILLER_17_1832 ();
 sg13g2_decap_4 FILLER_17_1871 ();
 sg13g2_fill_2 FILLER_17_1875 ();
 sg13g2_fill_2 FILLER_17_1882 ();
 sg13g2_decap_8 FILLER_17_1888 ();
 sg13g2_fill_2 FILLER_17_1895 ();
 sg13g2_decap_8 FILLER_17_1914 ();
 sg13g2_fill_2 FILLER_17_1921 ();
 sg13g2_fill_1 FILLER_17_1935 ();
 sg13g2_fill_2 FILLER_17_1944 ();
 sg13g2_fill_2 FILLER_17_1951 ();
 sg13g2_fill_1 FILLER_17_1962 ();
 sg13g2_fill_2 FILLER_17_1969 ();
 sg13g2_fill_1 FILLER_17_1971 ();
 sg13g2_decap_4 FILLER_17_1986 ();
 sg13g2_fill_2 FILLER_17_1990 ();
 sg13g2_decap_8 FILLER_17_2016 ();
 sg13g2_fill_1 FILLER_17_2023 ();
 sg13g2_fill_1 FILLER_17_2029 ();
 sg13g2_decap_4 FILLER_17_2043 ();
 sg13g2_decap_8 FILLER_17_2051 ();
 sg13g2_decap_8 FILLER_17_2058 ();
 sg13g2_decap_4 FILLER_17_2065 ();
 sg13g2_fill_2 FILLER_17_2069 ();
 sg13g2_fill_2 FILLER_17_2103 ();
 sg13g2_fill_1 FILLER_17_2105 ();
 sg13g2_fill_2 FILLER_17_2147 ();
 sg13g2_fill_1 FILLER_17_2149 ();
 sg13g2_decap_8 FILLER_17_2170 ();
 sg13g2_decap_4 FILLER_17_2177 ();
 sg13g2_fill_1 FILLER_17_2181 ();
 sg13g2_fill_2 FILLER_17_2186 ();
 sg13g2_decap_8 FILLER_17_2204 ();
 sg13g2_fill_1 FILLER_17_2211 ();
 sg13g2_decap_8 FILLER_17_2217 ();
 sg13g2_decap_8 FILLER_17_2224 ();
 sg13g2_decap_8 FILLER_17_2231 ();
 sg13g2_decap_8 FILLER_17_2238 ();
 sg13g2_fill_2 FILLER_17_2245 ();
 sg13g2_decap_4 FILLER_17_2261 ();
 sg13g2_fill_1 FILLER_17_2265 ();
 sg13g2_decap_8 FILLER_17_2287 ();
 sg13g2_fill_2 FILLER_17_2294 ();
 sg13g2_fill_1 FILLER_17_2311 ();
 sg13g2_fill_1 FILLER_17_2326 ();
 sg13g2_fill_2 FILLER_17_2355 ();
 sg13g2_decap_4 FILLER_17_2411 ();
 sg13g2_fill_1 FILLER_17_2415 ();
 sg13g2_decap_4 FILLER_17_2444 ();
 sg13g2_fill_2 FILLER_17_2448 ();
 sg13g2_fill_2 FILLER_17_2472 ();
 sg13g2_fill_1 FILLER_17_2474 ();
 sg13g2_fill_1 FILLER_17_2488 ();
 sg13g2_fill_2 FILLER_17_2519 ();
 sg13g2_fill_1 FILLER_17_2521 ();
 sg13g2_fill_2 FILLER_17_2527 ();
 sg13g2_fill_1 FILLER_17_2529 ();
 sg13g2_decap_4 FILLER_17_2538 ();
 sg13g2_fill_1 FILLER_17_2542 ();
 sg13g2_fill_2 FILLER_17_2554 ();
 sg13g2_fill_1 FILLER_17_2561 ();
 sg13g2_decap_4 FILLER_17_2590 ();
 sg13g2_decap_4 FILLER_17_2617 ();
 sg13g2_fill_1 FILLER_17_2621 ();
 sg13g2_decap_4 FILLER_17_2635 ();
 sg13g2_fill_2 FILLER_17_2639 ();
 sg13g2_fill_1 FILLER_17_2645 ();
 sg13g2_fill_2 FILLER_17_2708 ();
 sg13g2_fill_2 FILLER_17_2726 ();
 sg13g2_fill_1 FILLER_17_2728 ();
 sg13g2_fill_1 FILLER_17_2738 ();
 sg13g2_fill_2 FILLER_17_2765 ();
 sg13g2_decap_8 FILLER_17_2789 ();
 sg13g2_fill_1 FILLER_17_2815 ();
 sg13g2_decap_8 FILLER_17_2827 ();
 sg13g2_decap_8 FILLER_17_2834 ();
 sg13g2_decap_8 FILLER_17_2841 ();
 sg13g2_decap_8 FILLER_17_2865 ();
 sg13g2_decap_4 FILLER_17_2872 ();
 sg13g2_fill_1 FILLER_17_2876 ();
 sg13g2_decap_4 FILLER_17_2910 ();
 sg13g2_decap_8 FILLER_17_2937 ();
 sg13g2_decap_8 FILLER_17_2944 ();
 sg13g2_decap_8 FILLER_17_2951 ();
 sg13g2_decap_4 FILLER_17_2958 ();
 sg13g2_fill_1 FILLER_17_2962 ();
 sg13g2_fill_1 FILLER_17_2968 ();
 sg13g2_fill_2 FILLER_17_2979 ();
 sg13g2_decap_4 FILLER_17_3018 ();
 sg13g2_fill_2 FILLER_17_3022 ();
 sg13g2_decap_4 FILLER_17_3054 ();
 sg13g2_fill_2 FILLER_17_3076 ();
 sg13g2_fill_1 FILLER_17_3078 ();
 sg13g2_decap_8 FILLER_17_3105 ();
 sg13g2_fill_2 FILLER_17_3112 ();
 sg13g2_fill_1 FILLER_17_3114 ();
 sg13g2_decap_8 FILLER_17_3128 ();
 sg13g2_fill_1 FILLER_17_3135 ();
 sg13g2_fill_2 FILLER_17_3144 ();
 sg13g2_decap_4 FILLER_17_3172 ();
 sg13g2_fill_1 FILLER_17_3181 ();
 sg13g2_decap_4 FILLER_17_3187 ();
 sg13g2_fill_2 FILLER_17_3191 ();
 sg13g2_fill_1 FILLER_17_3211 ();
 sg13g2_fill_2 FILLER_17_3235 ();
 sg13g2_decap_8 FILLER_17_3257 ();
 sg13g2_decap_8 FILLER_17_3264 ();
 sg13g2_decap_8 FILLER_17_3271 ();
 sg13g2_decap_8 FILLER_17_3278 ();
 sg13g2_decap_8 FILLER_17_3285 ();
 sg13g2_decap_8 FILLER_17_3292 ();
 sg13g2_decap_8 FILLER_17_3299 ();
 sg13g2_decap_8 FILLER_17_3306 ();
 sg13g2_decap_8 FILLER_17_3313 ();
 sg13g2_decap_8 FILLER_17_3320 ();
 sg13g2_decap_8 FILLER_17_3327 ();
 sg13g2_decap_8 FILLER_17_3334 ();
 sg13g2_decap_8 FILLER_17_3341 ();
 sg13g2_decap_8 FILLER_17_3348 ();
 sg13g2_decap_8 FILLER_17_3355 ();
 sg13g2_decap_8 FILLER_17_3362 ();
 sg13g2_decap_8 FILLER_17_3369 ();
 sg13g2_decap_8 FILLER_17_3376 ();
 sg13g2_decap_8 FILLER_17_3383 ();
 sg13g2_decap_8 FILLER_17_3390 ();
 sg13g2_decap_8 FILLER_17_3397 ();
 sg13g2_decap_8 FILLER_17_3404 ();
 sg13g2_decap_8 FILLER_17_3411 ();
 sg13g2_decap_8 FILLER_17_3418 ();
 sg13g2_decap_8 FILLER_17_3425 ();
 sg13g2_decap_8 FILLER_17_3432 ();
 sg13g2_decap_8 FILLER_17_3439 ();
 sg13g2_decap_8 FILLER_17_3446 ();
 sg13g2_decap_8 FILLER_17_3453 ();
 sg13g2_decap_8 FILLER_17_3460 ();
 sg13g2_decap_8 FILLER_17_3467 ();
 sg13g2_decap_8 FILLER_17_3474 ();
 sg13g2_decap_8 FILLER_17_3481 ();
 sg13g2_decap_8 FILLER_17_3488 ();
 sg13g2_decap_8 FILLER_17_3495 ();
 sg13g2_decap_8 FILLER_17_3502 ();
 sg13g2_decap_8 FILLER_17_3509 ();
 sg13g2_decap_8 FILLER_17_3516 ();
 sg13g2_decap_8 FILLER_17_3523 ();
 sg13g2_decap_8 FILLER_17_3530 ();
 sg13g2_decap_8 FILLER_17_3537 ();
 sg13g2_decap_8 FILLER_17_3544 ();
 sg13g2_decap_8 FILLER_17_3551 ();
 sg13g2_decap_8 FILLER_17_3558 ();
 sg13g2_decap_8 FILLER_17_3565 ();
 sg13g2_decap_8 FILLER_17_3572 ();
 sg13g2_fill_1 FILLER_17_3579 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_decap_4 FILLER_18_376 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_decap_4 FILLER_18_390 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_fill_1 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_fill_2 FILLER_18_416 ();
 sg13g2_fill_1 FILLER_18_418 ();
 sg13g2_fill_2 FILLER_18_422 ();
 sg13g2_decap_8 FILLER_18_428 ();
 sg13g2_decap_4 FILLER_18_435 ();
 sg13g2_fill_2 FILLER_18_452 ();
 sg13g2_fill_1 FILLER_18_470 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_4 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_4 FILLER_18_513 ();
 sg13g2_fill_2 FILLER_18_517 ();
 sg13g2_fill_1 FILLER_18_528 ();
 sg13g2_decap_8 FILLER_18_538 ();
 sg13g2_decap_8 FILLER_18_545 ();
 sg13g2_decap_4 FILLER_18_552 ();
 sg13g2_fill_2 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_579 ();
 sg13g2_decap_4 FILLER_18_586 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_fill_1 FILLER_18_620 ();
 sg13g2_fill_2 FILLER_18_656 ();
 sg13g2_decap_8 FILLER_18_671 ();
 sg13g2_decap_4 FILLER_18_678 ();
 sg13g2_fill_1 FILLER_18_682 ();
 sg13g2_fill_2 FILLER_18_711 ();
 sg13g2_fill_1 FILLER_18_741 ();
 sg13g2_decap_4 FILLER_18_747 ();
 sg13g2_decap_4 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_4 FILLER_18_784 ();
 sg13g2_fill_2 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_4 FILLER_18_812 ();
 sg13g2_fill_1 FILLER_18_853 ();
 sg13g2_decap_8 FILLER_18_867 ();
 sg13g2_decap_8 FILLER_18_874 ();
 sg13g2_fill_2 FILLER_18_881 ();
 sg13g2_fill_1 FILLER_18_883 ();
 sg13g2_decap_8 FILLER_18_903 ();
 sg13g2_decap_4 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_927 ();
 sg13g2_decap_4 FILLER_18_941 ();
 sg13g2_fill_2 FILLER_18_945 ();
 sg13g2_fill_2 FILLER_18_960 ();
 sg13g2_fill_1 FILLER_18_962 ();
 sg13g2_decap_4 FILLER_18_976 ();
 sg13g2_decap_4 FILLER_18_1004 ();
 sg13g2_fill_1 FILLER_18_1008 ();
 sg13g2_fill_1 FILLER_18_1036 ();
 sg13g2_fill_2 FILLER_18_1050 ();
 sg13g2_decap_8 FILLER_18_1080 ();
 sg13g2_decap_8 FILLER_18_1087 ();
 sg13g2_decap_8 FILLER_18_1094 ();
 sg13g2_fill_2 FILLER_18_1101 ();
 sg13g2_decap_4 FILLER_18_1116 ();
 sg13g2_fill_1 FILLER_18_1120 ();
 sg13g2_decap_8 FILLER_18_1132 ();
 sg13g2_fill_2 FILLER_18_1139 ();
 sg13g2_fill_1 FILLER_18_1141 ();
 sg13g2_decap_4 FILLER_18_1149 ();
 sg13g2_decap_4 FILLER_18_1157 ();
 sg13g2_fill_2 FILLER_18_1161 ();
 sg13g2_fill_1 FILLER_18_1189 ();
 sg13g2_fill_1 FILLER_18_1196 ();
 sg13g2_fill_2 FILLER_18_1233 ();
 sg13g2_fill_1 FILLER_18_1235 ();
 sg13g2_decap_4 FILLER_18_1256 ();
 sg13g2_fill_2 FILLER_18_1348 ();
 sg13g2_decap_8 FILLER_18_1376 ();
 sg13g2_decap_8 FILLER_18_1383 ();
 sg13g2_decap_8 FILLER_18_1390 ();
 sg13g2_decap_8 FILLER_18_1429 ();
 sg13g2_decap_4 FILLER_18_1436 ();
 sg13g2_fill_1 FILLER_18_1440 ();
 sg13g2_decap_8 FILLER_18_1458 ();
 sg13g2_decap_4 FILLER_18_1465 ();
 sg13g2_fill_1 FILLER_18_1469 ();
 sg13g2_fill_1 FILLER_18_1489 ();
 sg13g2_decap_8 FILLER_18_1522 ();
 sg13g2_decap_8 FILLER_18_1533 ();
 sg13g2_fill_2 FILLER_18_1540 ();
 sg13g2_fill_1 FILLER_18_1542 ();
 sg13g2_fill_2 FILLER_18_1575 ();
 sg13g2_fill_1 FILLER_18_1577 ();
 sg13g2_decap_4 FILLER_18_1591 ();
 sg13g2_fill_1 FILLER_18_1595 ();
 sg13g2_fill_1 FILLER_18_1609 ();
 sg13g2_fill_1 FILLER_18_1614 ();
 sg13g2_decap_8 FILLER_18_1628 ();
 sg13g2_fill_2 FILLER_18_1663 ();
 sg13g2_decap_4 FILLER_18_1668 ();
 sg13g2_fill_1 FILLER_18_1672 ();
 sg13g2_decap_8 FILLER_18_1677 ();
 sg13g2_fill_1 FILLER_18_1710 ();
 sg13g2_decap_4 FILLER_18_1733 ();
 sg13g2_fill_1 FILLER_18_1737 ();
 sg13g2_decap_4 FILLER_18_1745 ();
 sg13g2_fill_2 FILLER_18_1768 ();
 sg13g2_fill_1 FILLER_18_1770 ();
 sg13g2_fill_2 FILLER_18_1797 ();
 sg13g2_fill_2 FILLER_18_1807 ();
 sg13g2_fill_1 FILLER_18_1809 ();
 sg13g2_decap_8 FILLER_18_1820 ();
 sg13g2_decap_4 FILLER_18_1827 ();
 sg13g2_fill_2 FILLER_18_1831 ();
 sg13g2_decap_8 FILLER_18_1850 ();
 sg13g2_decap_8 FILLER_18_1869 ();
 sg13g2_fill_2 FILLER_18_1876 ();
 sg13g2_fill_1 FILLER_18_1878 ();
 sg13g2_fill_2 FILLER_18_1920 ();
 sg13g2_fill_1 FILLER_18_1931 ();
 sg13g2_decap_8 FILLER_18_1942 ();
 sg13g2_fill_2 FILLER_18_1949 ();
 sg13g2_fill_2 FILLER_18_1980 ();
 sg13g2_decap_8 FILLER_18_1995 ();
 sg13g2_decap_8 FILLER_18_2002 ();
 sg13g2_fill_2 FILLER_18_2014 ();
 sg13g2_fill_1 FILLER_18_2016 ();
 sg13g2_decap_4 FILLER_18_2022 ();
 sg13g2_fill_1 FILLER_18_2044 ();
 sg13g2_fill_1 FILLER_18_2070 ();
 sg13g2_fill_1 FILLER_18_2085 ();
 sg13g2_decap_8 FILLER_18_2090 ();
 sg13g2_decap_4 FILLER_18_2097 ();
 sg13g2_fill_2 FILLER_18_2101 ();
 sg13g2_decap_8 FILLER_18_2116 ();
 sg13g2_decap_8 FILLER_18_2123 ();
 sg13g2_decap_8 FILLER_18_2130 ();
 sg13g2_fill_2 FILLER_18_2137 ();
 sg13g2_fill_2 FILLER_18_2152 ();
 sg13g2_decap_4 FILLER_18_2185 ();
 sg13g2_fill_2 FILLER_18_2189 ();
 sg13g2_fill_2 FILLER_18_2212 ();
 sg13g2_decap_8 FILLER_18_2247 ();
 sg13g2_decap_4 FILLER_18_2254 ();
 sg13g2_fill_2 FILLER_18_2263 ();
 sg13g2_fill_1 FILLER_18_2265 ();
 sg13g2_fill_2 FILLER_18_2283 ();
 sg13g2_decap_4 FILLER_18_2290 ();
 sg13g2_decap_8 FILLER_18_2309 ();
 sg13g2_decap_4 FILLER_18_2316 ();
 sg13g2_fill_1 FILLER_18_2328 ();
 sg13g2_decap_8 FILLER_18_2342 ();
 sg13g2_fill_2 FILLER_18_2366 ();
 sg13g2_fill_1 FILLER_18_2368 ();
 sg13g2_decap_8 FILLER_18_2381 ();
 sg13g2_decap_8 FILLER_18_2388 ();
 sg13g2_decap_8 FILLER_18_2434 ();
 sg13g2_decap_8 FILLER_18_2441 ();
 sg13g2_fill_1 FILLER_18_2448 ();
 sg13g2_decap_4 FILLER_18_2470 ();
 sg13g2_fill_2 FILLER_18_2474 ();
 sg13g2_decap_8 FILLER_18_2485 ();
 sg13g2_decap_4 FILLER_18_2492 ();
 sg13g2_fill_1 FILLER_18_2496 ();
 sg13g2_decap_8 FILLER_18_2501 ();
 sg13g2_decap_8 FILLER_18_2508 ();
 sg13g2_decap_8 FILLER_18_2533 ();
 sg13g2_fill_2 FILLER_18_2540 ();
 sg13g2_decap_8 FILLER_18_2579 ();
 sg13g2_fill_2 FILLER_18_2586 ();
 sg13g2_fill_1 FILLER_18_2588 ();
 sg13g2_fill_2 FILLER_18_2602 ();
 sg13g2_decap_4 FILLER_18_2632 ();
 sg13g2_fill_2 FILLER_18_2636 ();
 sg13g2_decap_4 FILLER_18_2659 ();
 sg13g2_fill_1 FILLER_18_2663 ();
 sg13g2_decap_8 FILLER_18_2676 ();
 sg13g2_fill_2 FILLER_18_2683 ();
 sg13g2_fill_1 FILLER_18_2685 ();
 sg13g2_decap_8 FILLER_18_2700 ();
 sg13g2_decap_4 FILLER_18_2707 ();
 sg13g2_fill_1 FILLER_18_2711 ();
 sg13g2_decap_8 FILLER_18_2724 ();
 sg13g2_fill_1 FILLER_18_2731 ();
 sg13g2_fill_2 FILLER_18_2743 ();
 sg13g2_fill_1 FILLER_18_2745 ();
 sg13g2_decap_4 FILLER_18_2756 ();
 sg13g2_fill_2 FILLER_18_2785 ();
 sg13g2_fill_2 FILLER_18_2795 ();
 sg13g2_fill_1 FILLER_18_2818 ();
 sg13g2_fill_2 FILLER_18_2848 ();
 sg13g2_fill_1 FILLER_18_2850 ();
 sg13g2_decap_4 FILLER_18_2877 ();
 sg13g2_fill_1 FILLER_18_2881 ();
 sg13g2_decap_8 FILLER_18_2886 ();
 sg13g2_fill_2 FILLER_18_2893 ();
 sg13g2_fill_2 FILLER_18_2914 ();
 sg13g2_decap_4 FILLER_18_2921 ();
 sg13g2_decap_8 FILLER_18_2944 ();
 sg13g2_decap_8 FILLER_18_2951 ();
 sg13g2_fill_2 FILLER_18_2969 ();
 sg13g2_decap_8 FILLER_18_2987 ();
 sg13g2_decap_8 FILLER_18_2994 ();
 sg13g2_fill_1 FILLER_18_3001 ();
 sg13g2_fill_1 FILLER_18_3011 ();
 sg13g2_fill_2 FILLER_18_3040 ();
 sg13g2_fill_1 FILLER_18_3042 ();
 sg13g2_fill_1 FILLER_18_3048 ();
 sg13g2_fill_2 FILLER_18_3079 ();
 sg13g2_fill_1 FILLER_18_3081 ();
 sg13g2_decap_8 FILLER_18_3096 ();
 sg13g2_fill_2 FILLER_18_3103 ();
 sg13g2_fill_2 FILLER_18_3121 ();
 sg13g2_fill_1 FILLER_18_3123 ();
 sg13g2_decap_8 FILLER_18_3142 ();
 sg13g2_decap_8 FILLER_18_3149 ();
 sg13g2_fill_1 FILLER_18_3156 ();
 sg13g2_fill_2 FILLER_18_3183 ();
 sg13g2_decap_4 FILLER_18_3190 ();
 sg13g2_fill_2 FILLER_18_3202 ();
 sg13g2_fill_1 FILLER_18_3208 ();
 sg13g2_fill_2 FILLER_18_3228 ();
 sg13g2_fill_1 FILLER_18_3230 ();
 sg13g2_decap_8 FILLER_18_3250 ();
 sg13g2_decap_8 FILLER_18_3257 ();
 sg13g2_decap_8 FILLER_18_3264 ();
 sg13g2_decap_8 FILLER_18_3271 ();
 sg13g2_decap_8 FILLER_18_3278 ();
 sg13g2_decap_8 FILLER_18_3285 ();
 sg13g2_decap_8 FILLER_18_3292 ();
 sg13g2_decap_8 FILLER_18_3299 ();
 sg13g2_decap_8 FILLER_18_3306 ();
 sg13g2_decap_8 FILLER_18_3313 ();
 sg13g2_decap_8 FILLER_18_3320 ();
 sg13g2_decap_8 FILLER_18_3327 ();
 sg13g2_decap_8 FILLER_18_3334 ();
 sg13g2_decap_8 FILLER_18_3341 ();
 sg13g2_decap_8 FILLER_18_3348 ();
 sg13g2_decap_8 FILLER_18_3355 ();
 sg13g2_decap_8 FILLER_18_3362 ();
 sg13g2_decap_8 FILLER_18_3369 ();
 sg13g2_decap_8 FILLER_18_3376 ();
 sg13g2_decap_8 FILLER_18_3383 ();
 sg13g2_decap_8 FILLER_18_3390 ();
 sg13g2_decap_8 FILLER_18_3397 ();
 sg13g2_decap_8 FILLER_18_3404 ();
 sg13g2_decap_8 FILLER_18_3411 ();
 sg13g2_decap_8 FILLER_18_3418 ();
 sg13g2_decap_8 FILLER_18_3425 ();
 sg13g2_decap_8 FILLER_18_3432 ();
 sg13g2_decap_8 FILLER_18_3439 ();
 sg13g2_decap_8 FILLER_18_3446 ();
 sg13g2_decap_8 FILLER_18_3453 ();
 sg13g2_decap_8 FILLER_18_3460 ();
 sg13g2_decap_8 FILLER_18_3467 ();
 sg13g2_decap_8 FILLER_18_3474 ();
 sg13g2_decap_8 FILLER_18_3481 ();
 sg13g2_decap_8 FILLER_18_3488 ();
 sg13g2_decap_8 FILLER_18_3495 ();
 sg13g2_decap_8 FILLER_18_3502 ();
 sg13g2_decap_8 FILLER_18_3509 ();
 sg13g2_decap_8 FILLER_18_3516 ();
 sg13g2_decap_8 FILLER_18_3523 ();
 sg13g2_decap_8 FILLER_18_3530 ();
 sg13g2_decap_8 FILLER_18_3537 ();
 sg13g2_decap_8 FILLER_18_3544 ();
 sg13g2_decap_8 FILLER_18_3551 ();
 sg13g2_decap_8 FILLER_18_3558 ();
 sg13g2_decap_8 FILLER_18_3565 ();
 sg13g2_decap_8 FILLER_18_3572 ();
 sg13g2_fill_1 FILLER_18_3579 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_254 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_decap_4 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_399 ();
 sg13g2_decap_4 FILLER_19_423 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_2 FILLER_19_442 ();
 sg13g2_fill_1 FILLER_19_456 ();
 sg13g2_decap_8 FILLER_19_467 ();
 sg13g2_decap_4 FILLER_19_474 ();
 sg13g2_fill_2 FILLER_19_478 ();
 sg13g2_decap_8 FILLER_19_485 ();
 sg13g2_fill_2 FILLER_19_492 ();
 sg13g2_fill_1 FILLER_19_494 ();
 sg13g2_fill_2 FILLER_19_511 ();
 sg13g2_fill_1 FILLER_19_513 ();
 sg13g2_fill_2 FILLER_19_522 ();
 sg13g2_fill_1 FILLER_19_524 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_decap_4 FILLER_19_590 ();
 sg13g2_fill_1 FILLER_19_594 ();
 sg13g2_fill_2 FILLER_19_605 ();
 sg13g2_fill_2 FILLER_19_614 ();
 sg13g2_fill_2 FILLER_19_627 ();
 sg13g2_fill_2 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_645 ();
 sg13g2_fill_2 FILLER_19_652 ();
 sg13g2_fill_1 FILLER_19_654 ();
 sg13g2_fill_2 FILLER_19_665 ();
 sg13g2_decap_4 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_fill_2 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_723 ();
 sg13g2_decap_8 FILLER_19_730 ();
 sg13g2_fill_2 FILLER_19_755 ();
 sg13g2_fill_1 FILLER_19_757 ();
 sg13g2_fill_2 FILLER_19_780 ();
 sg13g2_fill_1 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_804 ();
 sg13g2_decap_4 FILLER_19_811 ();
 sg13g2_fill_1 FILLER_19_819 ();
 sg13g2_fill_1 FILLER_19_833 ();
 sg13g2_decap_4 FILLER_19_878 ();
 sg13g2_fill_2 FILLER_19_882 ();
 sg13g2_fill_1 FILLER_19_944 ();
 sg13g2_decap_4 FILLER_19_960 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_fill_2 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_995 ();
 sg13g2_decap_8 FILLER_19_1002 ();
 sg13g2_fill_2 FILLER_19_1009 ();
 sg13g2_fill_1 FILLER_19_1011 ();
 sg13g2_fill_2 FILLER_19_1021 ();
 sg13g2_decap_8 FILLER_19_1028 ();
 sg13g2_fill_2 FILLER_19_1035 ();
 sg13g2_fill_1 FILLER_19_1037 ();
 sg13g2_decap_4 FILLER_19_1061 ();
 sg13g2_decap_8 FILLER_19_1082 ();
 sg13g2_decap_8 FILLER_19_1089 ();
 sg13g2_fill_1 FILLER_19_1096 ();
 sg13g2_decap_4 FILLER_19_1122 ();
 sg13g2_fill_2 FILLER_19_1131 ();
 sg13g2_fill_1 FILLER_19_1133 ();
 sg13g2_decap_4 FILLER_19_1162 ();
 sg13g2_fill_2 FILLER_19_1166 ();
 sg13g2_decap_8 FILLER_19_1207 ();
 sg13g2_decap_8 FILLER_19_1214 ();
 sg13g2_fill_2 FILLER_19_1221 ();
 sg13g2_decap_4 FILLER_19_1227 ();
 sg13g2_fill_2 FILLER_19_1231 ();
 sg13g2_decap_8 FILLER_19_1250 ();
 sg13g2_fill_2 FILLER_19_1257 ();
 sg13g2_fill_1 FILLER_19_1259 ();
 sg13g2_fill_2 FILLER_19_1291 ();
 sg13g2_fill_2 FILLER_19_1319 ();
 sg13g2_decap_8 FILLER_19_1338 ();
 sg13g2_decap_8 FILLER_19_1379 ();
 sg13g2_fill_1 FILLER_19_1386 ();
 sg13g2_fill_2 FILLER_19_1400 ();
 sg13g2_fill_2 FILLER_19_1415 ();
 sg13g2_fill_1 FILLER_19_1417 ();
 sg13g2_decap_4 FILLER_19_1423 ();
 sg13g2_fill_2 FILLER_19_1427 ();
 sg13g2_fill_2 FILLER_19_1434 ();
 sg13g2_fill_1 FILLER_19_1436 ();
 sg13g2_fill_1 FILLER_19_1472 ();
 sg13g2_fill_1 FILLER_19_1513 ();
 sg13g2_decap_8 FILLER_19_1518 ();
 sg13g2_fill_2 FILLER_19_1525 ();
 sg13g2_fill_1 FILLER_19_1527 ();
 sg13g2_decap_8 FILLER_19_1545 ();
 sg13g2_fill_2 FILLER_19_1552 ();
 sg13g2_decap_8 FILLER_19_1584 ();
 sg13g2_decap_8 FILLER_19_1591 ();
 sg13g2_fill_2 FILLER_19_1598 ();
 sg13g2_fill_1 FILLER_19_1600 ();
 sg13g2_fill_2 FILLER_19_1633 ();
 sg13g2_fill_1 FILLER_19_1635 ();
 sg13g2_fill_2 FILLER_19_1641 ();
 sg13g2_decap_8 FILLER_19_1652 ();
 sg13g2_decap_8 FILLER_19_1659 ();
 sg13g2_decap_8 FILLER_19_1666 ();
 sg13g2_fill_2 FILLER_19_1673 ();
 sg13g2_decap_8 FILLER_19_1682 ();
 sg13g2_decap_4 FILLER_19_1689 ();
 sg13g2_fill_1 FILLER_19_1693 ();
 sg13g2_decap_8 FILLER_19_1704 ();
 sg13g2_decap_4 FILLER_19_1711 ();
 sg13g2_fill_2 FILLER_19_1729 ();
 sg13g2_fill_1 FILLER_19_1731 ();
 sg13g2_decap_8 FILLER_19_1751 ();
 sg13g2_decap_8 FILLER_19_1758 ();
 sg13g2_decap_8 FILLER_19_1765 ();
 sg13g2_fill_2 FILLER_19_1772 ();
 sg13g2_fill_1 FILLER_19_1774 ();
 sg13g2_decap_4 FILLER_19_1792 ();
 sg13g2_fill_1 FILLER_19_1796 ();
 sg13g2_decap_8 FILLER_19_1829 ();
 sg13g2_fill_1 FILLER_19_1849 ();
 sg13g2_fill_1 FILLER_19_1863 ();
 sg13g2_decap_4 FILLER_19_1877 ();
 sg13g2_decap_8 FILLER_19_1895 ();
 sg13g2_fill_1 FILLER_19_1902 ();
 sg13g2_decap_4 FILLER_19_1917 ();
 sg13g2_decap_4 FILLER_19_1958 ();
 sg13g2_fill_1 FILLER_19_1965 ();
 sg13g2_fill_1 FILLER_19_1969 ();
 sg13g2_decap_4 FILLER_19_1998 ();
 sg13g2_fill_1 FILLER_19_2002 ();
 sg13g2_fill_2 FILLER_19_2017 ();
 sg13g2_fill_1 FILLER_19_2019 ();
 sg13g2_fill_2 FILLER_19_2049 ();
 sg13g2_fill_1 FILLER_19_2051 ();
 sg13g2_fill_2 FILLER_19_2065 ();
 sg13g2_fill_1 FILLER_19_2067 ();
 sg13g2_decap_4 FILLER_19_2109 ();
 sg13g2_fill_1 FILLER_19_2141 ();
 sg13g2_fill_2 FILLER_19_2173 ();
 sg13g2_decap_8 FILLER_19_2218 ();
 sg13g2_decap_8 FILLER_19_2225 ();
 sg13g2_decap_4 FILLER_19_2232 ();
 sg13g2_fill_1 FILLER_19_2236 ();
 sg13g2_fill_2 FILLER_19_2245 ();
 sg13g2_fill_1 FILLER_19_2247 ();
 sg13g2_decap_4 FILLER_19_2253 ();
 sg13g2_fill_1 FILLER_19_2278 ();
 sg13g2_decap_8 FILLER_19_2307 ();
 sg13g2_fill_2 FILLER_19_2314 ();
 sg13g2_fill_1 FILLER_19_2333 ();
 sg13g2_decap_8 FILLER_19_2384 ();
 sg13g2_decap_4 FILLER_19_2391 ();
 sg13g2_fill_2 FILLER_19_2430 ();
 sg13g2_fill_1 FILLER_19_2432 ();
 sg13g2_fill_1 FILLER_19_2506 ();
 sg13g2_fill_2 FILLER_19_2521 ();
 sg13g2_fill_1 FILLER_19_2550 ();
 sg13g2_decap_4 FILLER_19_2556 ();
 sg13g2_fill_1 FILLER_19_2560 ();
 sg13g2_fill_2 FILLER_19_2578 ();
 sg13g2_decap_8 FILLER_19_2622 ();
 sg13g2_decap_4 FILLER_19_2629 ();
 sg13g2_fill_1 FILLER_19_2633 ();
 sg13g2_fill_1 FILLER_19_2646 ();
 sg13g2_fill_2 FILLER_19_2652 ();
 sg13g2_decap_8 FILLER_19_2666 ();
 sg13g2_decap_4 FILLER_19_2673 ();
 sg13g2_fill_1 FILLER_19_2677 ();
 sg13g2_decap_8 FILLER_19_2686 ();
 sg13g2_decap_8 FILLER_19_2693 ();
 sg13g2_decap_4 FILLER_19_2700 ();
 sg13g2_fill_1 FILLER_19_2704 ();
 sg13g2_decap_8 FILLER_19_2716 ();
 sg13g2_fill_2 FILLER_19_2723 ();
 sg13g2_decap_4 FILLER_19_2746 ();
 sg13g2_fill_1 FILLER_19_2755 ();
 sg13g2_decap_4 FILLER_19_2761 ();
 sg13g2_decap_4 FILLER_19_2777 ();
 sg13g2_fill_2 FILLER_19_2781 ();
 sg13g2_decap_4 FILLER_19_2787 ();
 sg13g2_fill_1 FILLER_19_2791 ();
 sg13g2_decap_8 FILLER_19_2814 ();
 sg13g2_fill_1 FILLER_19_2821 ();
 sg13g2_decap_8 FILLER_19_2836 ();
 sg13g2_decap_4 FILLER_19_2843 ();
 sg13g2_decap_4 FILLER_19_2891 ();
 sg13g2_fill_2 FILLER_19_2900 ();
 sg13g2_fill_1 FILLER_19_2902 ();
 sg13g2_decap_4 FILLER_19_2921 ();
 sg13g2_decap_4 FILLER_19_2940 ();
 sg13g2_fill_2 FILLER_19_2948 ();
 sg13g2_decap_8 FILLER_19_2962 ();
 sg13g2_decap_8 FILLER_19_2985 ();
 sg13g2_decap_4 FILLER_19_2992 ();
 sg13g2_fill_2 FILLER_19_3004 ();
 sg13g2_fill_1 FILLER_19_3006 ();
 sg13g2_decap_8 FILLER_19_3027 ();
 sg13g2_decap_8 FILLER_19_3034 ();
 sg13g2_fill_1 FILLER_19_3041 ();
 sg13g2_fill_2 FILLER_19_3057 ();
 sg13g2_decap_8 FILLER_19_3069 ();
 sg13g2_decap_4 FILLER_19_3076 ();
 sg13g2_fill_1 FILLER_19_3080 ();
 sg13g2_fill_2 FILLER_19_3128 ();
 sg13g2_fill_1 FILLER_19_3134 ();
 sg13g2_fill_1 FILLER_19_3139 ();
 sg13g2_decap_8 FILLER_19_3151 ();
 sg13g2_decap_4 FILLER_19_3158 ();
 sg13g2_decap_8 FILLER_19_3177 ();
 sg13g2_decap_4 FILLER_19_3184 ();
 sg13g2_fill_2 FILLER_19_3200 ();
 sg13g2_decap_8 FILLER_19_3206 ();
 sg13g2_decap_8 FILLER_19_3213 ();
 sg13g2_fill_2 FILLER_19_3220 ();
 sg13g2_fill_1 FILLER_19_3232 ();
 sg13g2_decap_8 FILLER_19_3258 ();
 sg13g2_decap_8 FILLER_19_3265 ();
 sg13g2_decap_8 FILLER_19_3272 ();
 sg13g2_fill_2 FILLER_19_3279 ();
 sg13g2_fill_1 FILLER_19_3281 ();
 sg13g2_decap_8 FILLER_19_3313 ();
 sg13g2_fill_2 FILLER_19_3320 ();
 sg13g2_decap_8 FILLER_19_3330 ();
 sg13g2_decap_8 FILLER_19_3337 ();
 sg13g2_decap_8 FILLER_19_3344 ();
 sg13g2_decap_8 FILLER_19_3351 ();
 sg13g2_decap_8 FILLER_19_3358 ();
 sg13g2_decap_8 FILLER_19_3365 ();
 sg13g2_decap_8 FILLER_19_3372 ();
 sg13g2_decap_8 FILLER_19_3379 ();
 sg13g2_decap_8 FILLER_19_3386 ();
 sg13g2_decap_8 FILLER_19_3393 ();
 sg13g2_decap_8 FILLER_19_3400 ();
 sg13g2_decap_8 FILLER_19_3407 ();
 sg13g2_decap_8 FILLER_19_3414 ();
 sg13g2_decap_8 FILLER_19_3421 ();
 sg13g2_decap_8 FILLER_19_3428 ();
 sg13g2_decap_8 FILLER_19_3435 ();
 sg13g2_decap_8 FILLER_19_3442 ();
 sg13g2_decap_8 FILLER_19_3449 ();
 sg13g2_decap_8 FILLER_19_3456 ();
 sg13g2_decap_8 FILLER_19_3463 ();
 sg13g2_decap_8 FILLER_19_3470 ();
 sg13g2_decap_8 FILLER_19_3477 ();
 sg13g2_decap_8 FILLER_19_3484 ();
 sg13g2_decap_8 FILLER_19_3491 ();
 sg13g2_decap_8 FILLER_19_3498 ();
 sg13g2_decap_8 FILLER_19_3505 ();
 sg13g2_decap_8 FILLER_19_3512 ();
 sg13g2_decap_8 FILLER_19_3519 ();
 sg13g2_decap_8 FILLER_19_3526 ();
 sg13g2_decap_8 FILLER_19_3533 ();
 sg13g2_decap_8 FILLER_19_3540 ();
 sg13g2_decap_8 FILLER_19_3547 ();
 sg13g2_decap_8 FILLER_19_3554 ();
 sg13g2_decap_8 FILLER_19_3561 ();
 sg13g2_decap_8 FILLER_19_3568 ();
 sg13g2_decap_4 FILLER_19_3575 ();
 sg13g2_fill_1 FILLER_19_3579 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_decap_4 FILLER_20_446 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_2 FILLER_20_462 ();
 sg13g2_fill_1 FILLER_20_475 ();
 sg13g2_fill_1 FILLER_20_492 ();
 sg13g2_fill_2 FILLER_20_512 ();
 sg13g2_fill_2 FILLER_20_519 ();
 sg13g2_fill_1 FILLER_20_521 ();
 sg13g2_fill_2 FILLER_20_548 ();
 sg13g2_decap_4 FILLER_20_588 ();
 sg13g2_fill_1 FILLER_20_592 ();
 sg13g2_fill_1 FILLER_20_607 ();
 sg13g2_decap_4 FILLER_20_617 ();
 sg13g2_fill_2 FILLER_20_626 ();
 sg13g2_fill_1 FILLER_20_628 ();
 sg13g2_decap_4 FILLER_20_646 ();
 sg13g2_fill_1 FILLER_20_650 ();
 sg13g2_fill_2 FILLER_20_660 ();
 sg13g2_fill_1 FILLER_20_662 ();
 sg13g2_fill_2 FILLER_20_677 ();
 sg13g2_fill_1 FILLER_20_724 ();
 sg13g2_fill_1 FILLER_20_731 ();
 sg13g2_decap_4 FILLER_20_748 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_766 ();
 sg13g2_fill_1 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_fill_2 FILLER_20_785 ();
 sg13g2_fill_1 FILLER_20_787 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_4 FILLER_20_805 ();
 sg13g2_fill_1 FILLER_20_809 ();
 sg13g2_decap_4 FILLER_20_838 ();
 sg13g2_fill_2 FILLER_20_842 ();
 sg13g2_decap_4 FILLER_20_870 ();
 sg13g2_fill_2 FILLER_20_874 ();
 sg13g2_fill_2 FILLER_20_910 ();
 sg13g2_fill_1 FILLER_20_922 ();
 sg13g2_decap_4 FILLER_20_931 ();
 sg13g2_fill_1 FILLER_20_935 ();
 sg13g2_fill_2 FILLER_20_960 ();
 sg13g2_fill_1 FILLER_20_962 ();
 sg13g2_decap_8 FILLER_20_973 ();
 sg13g2_fill_2 FILLER_20_980 ();
 sg13g2_fill_1 FILLER_20_982 ();
 sg13g2_fill_1 FILLER_20_988 ();
 sg13g2_fill_2 FILLER_20_993 ();
 sg13g2_decap_8 FILLER_20_1000 ();
 sg13g2_fill_1 FILLER_20_1007 ();
 sg13g2_decap_8 FILLER_20_1029 ();
 sg13g2_fill_2 FILLER_20_1036 ();
 sg13g2_decap_8 FILLER_20_1057 ();
 sg13g2_decap_8 FILLER_20_1064 ();
 sg13g2_decap_4 FILLER_20_1076 ();
 sg13g2_fill_2 FILLER_20_1080 ();
 sg13g2_fill_2 FILLER_20_1123 ();
 sg13g2_fill_2 FILLER_20_1138 ();
 sg13g2_decap_8 FILLER_20_1144 ();
 sg13g2_fill_1 FILLER_20_1151 ();
 sg13g2_decap_8 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1169 ();
 sg13g2_fill_2 FILLER_20_1176 ();
 sg13g2_fill_1 FILLER_20_1178 ();
 sg13g2_fill_2 FILLER_20_1220 ();
 sg13g2_fill_1 FILLER_20_1222 ();
 sg13g2_decap_4 FILLER_20_1249 ();
 sg13g2_fill_2 FILLER_20_1266 ();
 sg13g2_decap_4 FILLER_20_1277 ();
 sg13g2_fill_2 FILLER_20_1281 ();
 sg13g2_decap_4 FILLER_20_1311 ();
 sg13g2_decap_8 FILLER_20_1334 ();
 sg13g2_decap_8 FILLER_20_1341 ();
 sg13g2_fill_2 FILLER_20_1400 ();
 sg13g2_decap_4 FILLER_20_1406 ();
 sg13g2_fill_2 FILLER_20_1410 ();
 sg13g2_fill_2 FILLER_20_1420 ();
 sg13g2_fill_1 FILLER_20_1434 ();
 sg13g2_decap_8 FILLER_20_1445 ();
 sg13g2_fill_1 FILLER_20_1452 ();
 sg13g2_decap_4 FILLER_20_1458 ();
 sg13g2_fill_1 FILLER_20_1462 ();
 sg13g2_decap_8 FILLER_20_1467 ();
 sg13g2_decap_8 FILLER_20_1474 ();
 sg13g2_fill_2 FILLER_20_1485 ();
 sg13g2_fill_1 FILLER_20_1487 ();
 sg13g2_decap_8 FILLER_20_1501 ();
 sg13g2_fill_1 FILLER_20_1508 ();
 sg13g2_decap_8 FILLER_20_1537 ();
 sg13g2_fill_1 FILLER_20_1576 ();
 sg13g2_decap_4 FILLER_20_1587 ();
 sg13g2_fill_1 FILLER_20_1599 ();
 sg13g2_fill_1 FILLER_20_1628 ();
 sg13g2_decap_8 FILLER_20_1661 ();
 sg13g2_decap_8 FILLER_20_1696 ();
 sg13g2_decap_8 FILLER_20_1703 ();
 sg13g2_decap_4 FILLER_20_1710 ();
 sg13g2_fill_1 FILLER_20_1714 ();
 sg13g2_decap_8 FILLER_20_1753 ();
 sg13g2_decap_4 FILLER_20_1760 ();
 sg13g2_fill_1 FILLER_20_1764 ();
 sg13g2_fill_1 FILLER_20_1799 ();
 sg13g2_fill_2 FILLER_20_1813 ();
 sg13g2_decap_8 FILLER_20_1825 ();
 sg13g2_decap_8 FILLER_20_1832 ();
 sg13g2_decap_4 FILLER_20_1839 ();
 sg13g2_fill_2 FILLER_20_1843 ();
 sg13g2_decap_8 FILLER_20_1862 ();
 sg13g2_decap_4 FILLER_20_1869 ();
 sg13g2_fill_2 FILLER_20_1910 ();
 sg13g2_fill_1 FILLER_20_1917 ();
 sg13g2_decap_4 FILLER_20_1926 ();
 sg13g2_fill_2 FILLER_20_1930 ();
 sg13g2_decap_8 FILLER_20_1978 ();
 sg13g2_decap_8 FILLER_20_1985 ();
 sg13g2_decap_4 FILLER_20_1992 ();
 sg13g2_fill_2 FILLER_20_1996 ();
 sg13g2_fill_1 FILLER_20_2006 ();
 sg13g2_decap_8 FILLER_20_2011 ();
 sg13g2_fill_1 FILLER_20_2025 ();
 sg13g2_fill_1 FILLER_20_2033 ();
 sg13g2_decap_8 FILLER_20_2039 ();
 sg13g2_decap_8 FILLER_20_2046 ();
 sg13g2_fill_2 FILLER_20_2053 ();
 sg13g2_decap_8 FILLER_20_2068 ();
 sg13g2_decap_8 FILLER_20_2075 ();
 sg13g2_decap_8 FILLER_20_2088 ();
 sg13g2_fill_2 FILLER_20_2095 ();
 sg13g2_fill_1 FILLER_20_2097 ();
 sg13g2_fill_2 FILLER_20_2115 ();
 sg13g2_fill_1 FILLER_20_2117 ();
 sg13g2_decap_4 FILLER_20_2122 ();
 sg13g2_decap_4 FILLER_20_2139 ();
 sg13g2_fill_2 FILLER_20_2161 ();
 sg13g2_decap_8 FILLER_20_2171 ();
 sg13g2_fill_1 FILLER_20_2188 ();
 sg13g2_fill_2 FILLER_20_2201 ();
 sg13g2_fill_1 FILLER_20_2208 ();
 sg13g2_fill_2 FILLER_20_2219 ();
 sg13g2_fill_1 FILLER_20_2221 ();
 sg13g2_fill_1 FILLER_20_2227 ();
 sg13g2_fill_2 FILLER_20_2237 ();
 sg13g2_fill_1 FILLER_20_2239 ();
 sg13g2_fill_1 FILLER_20_2248 ();
 sg13g2_decap_8 FILLER_20_2310 ();
 sg13g2_fill_1 FILLER_20_2317 ();
 sg13g2_fill_2 FILLER_20_2339 ();
 sg13g2_decap_4 FILLER_20_2360 ();
 sg13g2_fill_1 FILLER_20_2364 ();
 sg13g2_fill_1 FILLER_20_2402 ();
 sg13g2_fill_1 FILLER_20_2418 ();
 sg13g2_decap_8 FILLER_20_2428 ();
 sg13g2_fill_2 FILLER_20_2448 ();
 sg13g2_decap_8 FILLER_20_2476 ();
 sg13g2_fill_2 FILLER_20_2487 ();
 sg13g2_fill_2 FILLER_20_2503 ();
 sg13g2_fill_1 FILLER_20_2505 ();
 sg13g2_fill_2 FILLER_20_2526 ();
 sg13g2_fill_2 FILLER_20_2547 ();
 sg13g2_fill_1 FILLER_20_2549 ();
 sg13g2_decap_8 FILLER_20_2582 ();
 sg13g2_fill_2 FILLER_20_2589 ();
 sg13g2_fill_1 FILLER_20_2591 ();
 sg13g2_fill_2 FILLER_20_2605 ();
 sg13g2_fill_1 FILLER_20_2607 ();
 sg13g2_fill_2 FILLER_20_2630 ();
 sg13g2_fill_1 FILLER_20_2632 ();
 sg13g2_decap_8 FILLER_20_2656 ();
 sg13g2_fill_2 FILLER_20_2663 ();
 sg13g2_fill_1 FILLER_20_2665 ();
 sg13g2_decap_4 FILLER_20_2757 ();
 sg13g2_decap_4 FILLER_20_2769 ();
 sg13g2_fill_2 FILLER_20_2786 ();
 sg13g2_fill_1 FILLER_20_2788 ();
 sg13g2_decap_8 FILLER_20_2812 ();
 sg13g2_fill_2 FILLER_20_2819 ();
 sg13g2_decap_8 FILLER_20_2838 ();
 sg13g2_fill_2 FILLER_20_2845 ();
 sg13g2_decap_4 FILLER_20_2857 ();
 sg13g2_fill_2 FILLER_20_2861 ();
 sg13g2_decap_8 FILLER_20_2872 ();
 sg13g2_decap_8 FILLER_20_2879 ();
 sg13g2_decap_4 FILLER_20_2886 ();
 sg13g2_fill_2 FILLER_20_2890 ();
 sg13g2_decap_4 FILLER_20_2900 ();
 sg13g2_fill_2 FILLER_20_2913 ();
 sg13g2_decap_4 FILLER_20_2926 ();
 sg13g2_fill_2 FILLER_20_2940 ();
 sg13g2_fill_1 FILLER_20_2952 ();
 sg13g2_fill_2 FILLER_20_2963 ();
 sg13g2_fill_1 FILLER_20_2965 ();
 sg13g2_decap_8 FILLER_20_2991 ();
 sg13g2_fill_1 FILLER_20_2998 ();
 sg13g2_fill_1 FILLER_20_3004 ();
 sg13g2_decap_8 FILLER_20_3008 ();
 sg13g2_fill_1 FILLER_20_3015 ();
 sg13g2_fill_1 FILLER_20_3028 ();
 sg13g2_fill_1 FILLER_20_3037 ();
 sg13g2_decap_4 FILLER_20_3056 ();
 sg13g2_fill_1 FILLER_20_3060 ();
 sg13g2_decap_8 FILLER_20_3068 ();
 sg13g2_fill_1 FILLER_20_3075 ();
 sg13g2_decap_8 FILLER_20_3081 ();
 sg13g2_fill_2 FILLER_20_3088 ();
 sg13g2_fill_2 FILLER_20_3094 ();
 sg13g2_decap_8 FILLER_20_3101 ();
 sg13g2_fill_1 FILLER_20_3108 ();
 sg13g2_decap_4 FILLER_20_3122 ();
 sg13g2_fill_2 FILLER_20_3188 ();
 sg13g2_fill_1 FILLER_20_3190 ();
 sg13g2_fill_1 FILLER_20_3196 ();
 sg13g2_decap_8 FILLER_20_3225 ();
 sg13g2_decap_4 FILLER_20_3241 ();
 sg13g2_fill_1 FILLER_20_3245 ();
 sg13g2_fill_2 FILLER_20_3306 ();
 sg13g2_fill_1 FILLER_20_3308 ();
 sg13g2_fill_1 FILLER_20_3347 ();
 sg13g2_decap_8 FILLER_20_3352 ();
 sg13g2_decap_8 FILLER_20_3359 ();
 sg13g2_decap_8 FILLER_20_3366 ();
 sg13g2_decap_8 FILLER_20_3373 ();
 sg13g2_decap_8 FILLER_20_3380 ();
 sg13g2_decap_8 FILLER_20_3387 ();
 sg13g2_decap_8 FILLER_20_3394 ();
 sg13g2_decap_8 FILLER_20_3401 ();
 sg13g2_decap_8 FILLER_20_3408 ();
 sg13g2_decap_8 FILLER_20_3415 ();
 sg13g2_decap_8 FILLER_20_3422 ();
 sg13g2_decap_8 FILLER_20_3429 ();
 sg13g2_decap_8 FILLER_20_3436 ();
 sg13g2_decap_8 FILLER_20_3443 ();
 sg13g2_decap_8 FILLER_20_3450 ();
 sg13g2_decap_8 FILLER_20_3457 ();
 sg13g2_decap_8 FILLER_20_3464 ();
 sg13g2_decap_8 FILLER_20_3471 ();
 sg13g2_decap_8 FILLER_20_3478 ();
 sg13g2_decap_8 FILLER_20_3485 ();
 sg13g2_decap_8 FILLER_20_3492 ();
 sg13g2_decap_8 FILLER_20_3499 ();
 sg13g2_decap_8 FILLER_20_3506 ();
 sg13g2_decap_8 FILLER_20_3513 ();
 sg13g2_decap_8 FILLER_20_3520 ();
 sg13g2_decap_8 FILLER_20_3527 ();
 sg13g2_decap_8 FILLER_20_3534 ();
 sg13g2_decap_8 FILLER_20_3541 ();
 sg13g2_decap_8 FILLER_20_3548 ();
 sg13g2_decap_8 FILLER_20_3555 ();
 sg13g2_decap_8 FILLER_20_3562 ();
 sg13g2_decap_8 FILLER_20_3569 ();
 sg13g2_decap_4 FILLER_20_3576 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_4 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_4 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_363 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_decap_4 FILLER_21_379 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_4 FILLER_21_440 ();
 sg13g2_decap_4 FILLER_21_465 ();
 sg13g2_fill_2 FILLER_21_469 ();
 sg13g2_fill_1 FILLER_21_485 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_4 FILLER_21_521 ();
 sg13g2_fill_2 FILLER_21_566 ();
 sg13g2_fill_1 FILLER_21_568 ();
 sg13g2_fill_2 FILLER_21_583 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_fill_2 FILLER_21_619 ();
 sg13g2_fill_1 FILLER_21_639 ();
 sg13g2_fill_2 FILLER_21_645 ();
 sg13g2_decap_4 FILLER_21_655 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_fill_1 FILLER_21_700 ();
 sg13g2_fill_1 FILLER_21_707 ();
 sg13g2_fill_2 FILLER_21_717 ();
 sg13g2_fill_1 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_748 ();
 sg13g2_decap_4 FILLER_21_776 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_4 FILLER_21_807 ();
 sg13g2_fill_2 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_837 ();
 sg13g2_fill_2 FILLER_21_844 ();
 sg13g2_fill_1 FILLER_21_846 ();
 sg13g2_fill_2 FILLER_21_864 ();
 sg13g2_decap_8 FILLER_21_891 ();
 sg13g2_decap_4 FILLER_21_898 ();
 sg13g2_fill_1 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_928 ();
 sg13g2_decap_4 FILLER_21_935 ();
 sg13g2_fill_1 FILLER_21_939 ();
 sg13g2_fill_2 FILLER_21_953 ();
 sg13g2_fill_1 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_962 ();
 sg13g2_fill_2 FILLER_21_969 ();
 sg13g2_fill_1 FILLER_21_971 ();
 sg13g2_fill_1 FILLER_21_981 ();
 sg13g2_decap_4 FILLER_21_997 ();
 sg13g2_fill_2 FILLER_21_1001 ();
 sg13g2_decap_4 FILLER_21_1031 ();
 sg13g2_fill_1 FILLER_21_1035 ();
 sg13g2_decap_8 FILLER_21_1061 ();
 sg13g2_decap_4 FILLER_21_1068 ();
 sg13g2_decap_4 FILLER_21_1096 ();
 sg13g2_decap_8 FILLER_21_1104 ();
 sg13g2_decap_4 FILLER_21_1111 ();
 sg13g2_fill_1 FILLER_21_1115 ();
 sg13g2_decap_8 FILLER_21_1133 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_4 FILLER_21_1147 ();
 sg13g2_decap_8 FILLER_21_1167 ();
 sg13g2_decap_8 FILLER_21_1193 ();
 sg13g2_fill_2 FILLER_21_1200 ();
 sg13g2_fill_1 FILLER_21_1202 ();
 sg13g2_fill_2 FILLER_21_1213 ();
 sg13g2_fill_1 FILLER_21_1215 ();
 sg13g2_decap_4 FILLER_21_1249 ();
 sg13g2_fill_2 FILLER_21_1266 ();
 sg13g2_decap_8 FILLER_21_1276 ();
 sg13g2_decap_4 FILLER_21_1283 ();
 sg13g2_fill_1 FILLER_21_1287 ();
 sg13g2_decap_8 FILLER_21_1292 ();
 sg13g2_fill_2 FILLER_21_1299 ();
 sg13g2_fill_2 FILLER_21_1322 ();
 sg13g2_fill_1 FILLER_21_1324 ();
 sg13g2_decap_8 FILLER_21_1338 ();
 sg13g2_decap_4 FILLER_21_1350 ();
 sg13g2_fill_2 FILLER_21_1354 ();
 sg13g2_fill_2 FILLER_21_1377 ();
 sg13g2_fill_1 FILLER_21_1379 ();
 sg13g2_decap_4 FILLER_21_1385 ();
 sg13g2_fill_1 FILLER_21_1389 ();
 sg13g2_decap_4 FILLER_21_1398 ();
 sg13g2_fill_2 FILLER_21_1406 ();
 sg13g2_fill_1 FILLER_21_1408 ();
 sg13g2_fill_2 FILLER_21_1442 ();
 sg13g2_fill_1 FILLER_21_1444 ();
 sg13g2_fill_1 FILLER_21_1458 ();
 sg13g2_decap_4 FILLER_21_1475 ();
 sg13g2_fill_1 FILLER_21_1479 ();
 sg13g2_decap_8 FILLER_21_1498 ();
 sg13g2_decap_4 FILLER_21_1505 ();
 sg13g2_fill_1 FILLER_21_1517 ();
 sg13g2_fill_2 FILLER_21_1523 ();
 sg13g2_fill_1 FILLER_21_1525 ();
 sg13g2_decap_8 FILLER_21_1529 ();
 sg13g2_fill_2 FILLER_21_1536 ();
 sg13g2_fill_2 FILLER_21_1553 ();
 sg13g2_fill_1 FILLER_21_1555 ();
 sg13g2_decap_8 FILLER_21_1580 ();
 sg13g2_decap_4 FILLER_21_1587 ();
 sg13g2_fill_1 FILLER_21_1591 ();
 sg13g2_fill_2 FILLER_21_1611 ();
 sg13g2_fill_1 FILLER_21_1613 ();
 sg13g2_decap_8 FILLER_21_1619 ();
 sg13g2_decap_8 FILLER_21_1626 ();
 sg13g2_fill_2 FILLER_21_1633 ();
 sg13g2_fill_1 FILLER_21_1654 ();
 sg13g2_fill_1 FILLER_21_1659 ();
 sg13g2_fill_2 FILLER_21_1682 ();
 sg13g2_fill_1 FILLER_21_1684 ();
 sg13g2_decap_8 FILLER_21_1713 ();
 sg13g2_decap_4 FILLER_21_1725 ();
 sg13g2_fill_2 FILLER_21_1729 ();
 sg13g2_fill_1 FILLER_21_1735 ();
 sg13g2_decap_4 FILLER_21_1748 ();
 sg13g2_fill_1 FILLER_21_1752 ();
 sg13g2_decap_8 FILLER_21_1766 ();
 sg13g2_decap_8 FILLER_21_1790 ();
 sg13g2_decap_4 FILLER_21_1797 ();
 sg13g2_decap_4 FILLER_21_1805 ();
 sg13g2_fill_1 FILLER_21_1809 ();
 sg13g2_decap_8 FILLER_21_1828 ();
 sg13g2_fill_1 FILLER_21_1835 ();
 sg13g2_fill_2 FILLER_21_1868 ();
 sg13g2_fill_1 FILLER_21_1877 ();
 sg13g2_fill_1 FILLER_21_1888 ();
 sg13g2_decap_8 FILLER_21_1899 ();
 sg13g2_decap_4 FILLER_21_1906 ();
 sg13g2_fill_2 FILLER_21_1910 ();
 sg13g2_fill_1 FILLER_21_1916 ();
 sg13g2_decap_4 FILLER_21_1922 ();
 sg13g2_fill_2 FILLER_21_1935 ();
 sg13g2_fill_2 FILLER_21_1953 ();
 sg13g2_fill_1 FILLER_21_1955 ();
 sg13g2_decap_8 FILLER_21_1986 ();
 sg13g2_fill_1 FILLER_21_1993 ();
 sg13g2_fill_1 FILLER_21_2053 ();
 sg13g2_fill_1 FILLER_21_2105 ();
 sg13g2_fill_2 FILLER_21_2127 ();
 sg13g2_fill_1 FILLER_21_2129 ();
 sg13g2_fill_1 FILLER_21_2172 ();
 sg13g2_fill_2 FILLER_21_2201 ();
 sg13g2_fill_2 FILLER_21_2224 ();
 sg13g2_fill_1 FILLER_21_2226 ();
 sg13g2_fill_2 FILLER_21_2243 ();
 sg13g2_fill_1 FILLER_21_2245 ();
 sg13g2_decap_8 FILLER_21_2254 ();
 sg13g2_fill_1 FILLER_21_2261 ();
 sg13g2_fill_1 FILLER_21_2267 ();
 sg13g2_decap_8 FILLER_21_2272 ();
 sg13g2_decap_8 FILLER_21_2279 ();
 sg13g2_decap_8 FILLER_21_2286 ();
 sg13g2_fill_2 FILLER_21_2293 ();
 sg13g2_fill_1 FILLER_21_2295 ();
 sg13g2_decap_4 FILLER_21_2300 ();
 sg13g2_fill_1 FILLER_21_2304 ();
 sg13g2_fill_2 FILLER_21_2318 ();
 sg13g2_fill_1 FILLER_21_2320 ();
 sg13g2_fill_1 FILLER_21_2326 ();
 sg13g2_decap_8 FILLER_21_2340 ();
 sg13g2_fill_1 FILLER_21_2347 ();
 sg13g2_decap_8 FILLER_21_2364 ();
 sg13g2_fill_2 FILLER_21_2376 ();
 sg13g2_fill_1 FILLER_21_2378 ();
 sg13g2_fill_1 FILLER_21_2383 ();
 sg13g2_decap_8 FILLER_21_2387 ();
 sg13g2_fill_2 FILLER_21_2394 ();
 sg13g2_fill_1 FILLER_21_2396 ();
 sg13g2_decap_4 FILLER_21_2423 ();
 sg13g2_fill_2 FILLER_21_2455 ();
 sg13g2_fill_1 FILLER_21_2457 ();
 sg13g2_decap_4 FILLER_21_2476 ();
 sg13g2_fill_2 FILLER_21_2480 ();
 sg13g2_decap_8 FILLER_21_2486 ();
 sg13g2_fill_2 FILLER_21_2493 ();
 sg13g2_decap_8 FILLER_21_2500 ();
 sg13g2_fill_2 FILLER_21_2507 ();
 sg13g2_fill_1 FILLER_21_2509 ();
 sg13g2_fill_2 FILLER_21_2544 ();
 sg13g2_decap_8 FILLER_21_2549 ();
 sg13g2_decap_4 FILLER_21_2556 ();
 sg13g2_fill_1 FILLER_21_2560 ();
 sg13g2_decap_8 FILLER_21_2569 ();
 sg13g2_decap_8 FILLER_21_2576 ();
 sg13g2_decap_8 FILLER_21_2583 ();
 sg13g2_fill_2 FILLER_21_2590 ();
 sg13g2_decap_8 FILLER_21_2596 ();
 sg13g2_fill_2 FILLER_21_2603 ();
 sg13g2_decap_8 FILLER_21_2609 ();
 sg13g2_fill_2 FILLER_21_2616 ();
 sg13g2_fill_1 FILLER_21_2618 ();
 sg13g2_decap_8 FILLER_21_2647 ();
 sg13g2_fill_2 FILLER_21_2654 ();
 sg13g2_fill_1 FILLER_21_2656 ();
 sg13g2_fill_2 FILLER_21_2675 ();
 sg13g2_fill_1 FILLER_21_2677 ();
 sg13g2_decap_8 FILLER_21_2689 ();
 sg13g2_decap_8 FILLER_21_2696 ();
 sg13g2_decap_4 FILLER_21_2703 ();
 sg13g2_fill_1 FILLER_21_2707 ();
 sg13g2_fill_1 FILLER_21_2721 ();
 sg13g2_decap_8 FILLER_21_2753 ();
 sg13g2_fill_2 FILLER_21_2760 ();
 sg13g2_fill_1 FILLER_21_2782 ();
 sg13g2_decap_4 FILLER_21_2801 ();
 sg13g2_fill_1 FILLER_21_2805 ();
 sg13g2_decap_8 FILLER_21_2812 ();
 sg13g2_decap_8 FILLER_21_2819 ();
 sg13g2_fill_2 FILLER_21_2826 ();
 sg13g2_fill_1 FILLER_21_2828 ();
 sg13g2_decap_4 FILLER_21_2833 ();
 sg13g2_fill_1 FILLER_21_2837 ();
 sg13g2_fill_1 FILLER_21_2875 ();
 sg13g2_fill_1 FILLER_21_2885 ();
 sg13g2_decap_4 FILLER_21_2892 ();
 sg13g2_fill_2 FILLER_21_2896 ();
 sg13g2_fill_2 FILLER_21_2909 ();
 sg13g2_fill_1 FILLER_21_2911 ();
 sg13g2_fill_1 FILLER_21_2920 ();
 sg13g2_fill_2 FILLER_21_2926 ();
 sg13g2_fill_1 FILLER_21_2928 ();
 sg13g2_decap_8 FILLER_21_2941 ();
 sg13g2_decap_4 FILLER_21_2948 ();
 sg13g2_fill_1 FILLER_21_2952 ();
 sg13g2_decap_4 FILLER_21_2966 ();
 sg13g2_decap_8 FILLER_21_2984 ();
 sg13g2_decap_4 FILLER_21_2991 ();
 sg13g2_fill_1 FILLER_21_2995 ();
 sg13g2_fill_2 FILLER_21_3018 ();
 sg13g2_fill_1 FILLER_21_3020 ();
 sg13g2_fill_1 FILLER_21_3029 ();
 sg13g2_decap_4 FILLER_21_3060 ();
 sg13g2_fill_1 FILLER_21_3064 ();
 sg13g2_decap_8 FILLER_21_3105 ();
 sg13g2_fill_1 FILLER_21_3112 ();
 sg13g2_fill_1 FILLER_21_3118 ();
 sg13g2_fill_2 FILLER_21_3137 ();
 sg13g2_decap_8 FILLER_21_3144 ();
 sg13g2_decap_4 FILLER_21_3151 ();
 sg13g2_fill_2 FILLER_21_3155 ();
 sg13g2_decap_4 FILLER_21_3183 ();
 sg13g2_decap_4 FILLER_21_3192 ();
 sg13g2_decap_8 FILLER_21_3201 ();
 sg13g2_decap_8 FILLER_21_3213 ();
 sg13g2_fill_1 FILLER_21_3220 ();
 sg13g2_fill_2 FILLER_21_3249 ();
 sg13g2_decap_8 FILLER_21_3255 ();
 sg13g2_decap_4 FILLER_21_3262 ();
 sg13g2_fill_1 FILLER_21_3266 ();
 sg13g2_fill_1 FILLER_21_3285 ();
 sg13g2_fill_2 FILLER_21_3320 ();
 sg13g2_fill_2 FILLER_21_3328 ();
 sg13g2_fill_2 FILLER_21_3348 ();
 sg13g2_decap_8 FILLER_21_3359 ();
 sg13g2_decap_8 FILLER_21_3366 ();
 sg13g2_decap_8 FILLER_21_3373 ();
 sg13g2_decap_8 FILLER_21_3380 ();
 sg13g2_decap_8 FILLER_21_3387 ();
 sg13g2_decap_8 FILLER_21_3394 ();
 sg13g2_decap_8 FILLER_21_3401 ();
 sg13g2_decap_8 FILLER_21_3408 ();
 sg13g2_decap_8 FILLER_21_3415 ();
 sg13g2_decap_8 FILLER_21_3422 ();
 sg13g2_decap_8 FILLER_21_3429 ();
 sg13g2_decap_8 FILLER_21_3436 ();
 sg13g2_decap_8 FILLER_21_3443 ();
 sg13g2_decap_8 FILLER_21_3450 ();
 sg13g2_decap_8 FILLER_21_3457 ();
 sg13g2_decap_8 FILLER_21_3464 ();
 sg13g2_decap_8 FILLER_21_3471 ();
 sg13g2_decap_8 FILLER_21_3478 ();
 sg13g2_decap_8 FILLER_21_3485 ();
 sg13g2_decap_8 FILLER_21_3492 ();
 sg13g2_decap_8 FILLER_21_3499 ();
 sg13g2_decap_8 FILLER_21_3506 ();
 sg13g2_decap_8 FILLER_21_3513 ();
 sg13g2_decap_8 FILLER_21_3520 ();
 sg13g2_decap_8 FILLER_21_3527 ();
 sg13g2_decap_8 FILLER_21_3534 ();
 sg13g2_decap_8 FILLER_21_3541 ();
 sg13g2_decap_8 FILLER_21_3548 ();
 sg13g2_decap_8 FILLER_21_3555 ();
 sg13g2_decap_8 FILLER_21_3562 ();
 sg13g2_decap_8 FILLER_21_3569 ();
 sg13g2_decap_4 FILLER_21_3576 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_217 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_438 ();
 sg13g2_decap_4 FILLER_22_448 ();
 sg13g2_fill_2 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_463 ();
 sg13g2_decap_4 FILLER_22_470 ();
 sg13g2_fill_2 FILLER_22_474 ();
 sg13g2_fill_2 FILLER_22_493 ();
 sg13g2_fill_2 FILLER_22_522 ();
 sg13g2_fill_1 FILLER_22_524 ();
 sg13g2_fill_2 FILLER_22_564 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_628 ();
 sg13g2_decap_4 FILLER_22_635 ();
 sg13g2_decap_4 FILLER_22_657 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_4 FILLER_22_691 ();
 sg13g2_fill_2 FILLER_22_722 ();
 sg13g2_decap_4 FILLER_22_740 ();
 sg13g2_fill_2 FILLER_22_744 ();
 sg13g2_fill_2 FILLER_22_777 ();
 sg13g2_decap_4 FILLER_22_806 ();
 sg13g2_fill_1 FILLER_22_810 ();
 sg13g2_fill_2 FILLER_22_889 ();
 sg13g2_decap_4 FILLER_22_898 ();
 sg13g2_decap_8 FILLER_22_906 ();
 sg13g2_decap_4 FILLER_22_913 ();
 sg13g2_decap_4 FILLER_22_925 ();
 sg13g2_fill_2 FILLER_22_929 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_fill_1 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_955 ();
 sg13g2_decap_4 FILLER_22_962 ();
 sg13g2_fill_2 FILLER_22_980 ();
 sg13g2_decap_8 FILLER_22_993 ();
 sg13g2_fill_2 FILLER_22_1000 ();
 sg13g2_fill_1 FILLER_22_1002 ();
 sg13g2_decap_4 FILLER_22_1008 ();
 sg13g2_fill_2 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1031 ();
 sg13g2_fill_2 FILLER_22_1038 ();
 sg13g2_fill_1 FILLER_22_1040 ();
 sg13g2_decap_8 FILLER_22_1051 ();
 sg13g2_decap_4 FILLER_22_1058 ();
 sg13g2_fill_2 FILLER_22_1062 ();
 sg13g2_fill_1 FILLER_22_1067 ();
 sg13g2_decap_8 FILLER_22_1092 ();
 sg13g2_fill_2 FILLER_22_1099 ();
 sg13g2_fill_1 FILLER_22_1112 ();
 sg13g2_fill_2 FILLER_22_1132 ();
 sg13g2_fill_2 FILLER_22_1155 ();
 sg13g2_fill_1 FILLER_22_1157 ();
 sg13g2_decap_8 FILLER_22_1187 ();
 sg13g2_fill_2 FILLER_22_1194 ();
 sg13g2_fill_1 FILLER_22_1196 ();
 sg13g2_fill_2 FILLER_22_1214 ();
 sg13g2_fill_2 FILLER_22_1231 ();
 sg13g2_decap_4 FILLER_22_1258 ();
 sg13g2_fill_2 FILLER_22_1262 ();
 sg13g2_decap_4 FILLER_22_1288 ();
 sg13g2_fill_2 FILLER_22_1292 ();
 sg13g2_fill_2 FILLER_22_1343 ();
 sg13g2_fill_1 FILLER_22_1345 ();
 sg13g2_decap_4 FILLER_22_1370 ();
 sg13g2_fill_2 FILLER_22_1374 ();
 sg13g2_decap_8 FILLER_22_1381 ();
 sg13g2_fill_1 FILLER_22_1388 ();
 sg13g2_fill_2 FILLER_22_1410 ();
 sg13g2_fill_1 FILLER_22_1412 ();
 sg13g2_fill_1 FILLER_22_1418 ();
 sg13g2_decap_8 FILLER_22_1443 ();
 sg13g2_decap_8 FILLER_22_1450 ();
 sg13g2_decap_4 FILLER_22_1457 ();
 sg13g2_fill_2 FILLER_22_1461 ();
 sg13g2_decap_4 FILLER_22_1466 ();
 sg13g2_fill_2 FILLER_22_1470 ();
 sg13g2_decap_8 FILLER_22_1479 ();
 sg13g2_fill_2 FILLER_22_1507 ();
 sg13g2_fill_1 FILLER_22_1509 ();
 sg13g2_fill_2 FILLER_22_1527 ();
 sg13g2_fill_2 FILLER_22_1541 ();
 sg13g2_decap_4 FILLER_22_1563 ();
 sg13g2_fill_1 FILLER_22_1567 ();
 sg13g2_fill_1 FILLER_22_1573 ();
 sg13g2_fill_1 FILLER_22_1584 ();
 sg13g2_fill_2 FILLER_22_1644 ();
 sg13g2_fill_2 FILLER_22_1684 ();
 sg13g2_fill_2 FILLER_22_1702 ();
 sg13g2_decap_8 FILLER_22_1750 ();
 sg13g2_decap_4 FILLER_22_1757 ();
 sg13g2_fill_2 FILLER_22_1761 ();
 sg13g2_fill_2 FILLER_22_1772 ();
 sg13g2_decap_8 FILLER_22_1789 ();
 sg13g2_fill_1 FILLER_22_1796 ();
 sg13g2_decap_4 FILLER_22_1810 ();
 sg13g2_decap_4 FILLER_22_1858 ();
 sg13g2_decap_8 FILLER_22_1890 ();
 sg13g2_decap_4 FILLER_22_1897 ();
 sg13g2_fill_2 FILLER_22_1901 ();
 sg13g2_decap_8 FILLER_22_1940 ();
 sg13g2_fill_2 FILLER_22_1947 ();
 sg13g2_decap_4 FILLER_22_1962 ();
 sg13g2_fill_2 FILLER_22_1966 ();
 sg13g2_decap_8 FILLER_22_2008 ();
 sg13g2_decap_8 FILLER_22_2015 ();
 sg13g2_fill_2 FILLER_22_2022 ();
 sg13g2_decap_4 FILLER_22_2029 ();
 sg13g2_decap_4 FILLER_22_2044 ();
 sg13g2_fill_1 FILLER_22_2048 ();
 sg13g2_fill_2 FILLER_22_2063 ();
 sg13g2_fill_1 FILLER_22_2065 ();
 sg13g2_fill_2 FILLER_22_2075 ();
 sg13g2_fill_1 FILLER_22_2077 ();
 sg13g2_fill_1 FILLER_22_2087 ();
 sg13g2_fill_2 FILLER_22_2102 ();
 sg13g2_fill_1 FILLER_22_2104 ();
 sg13g2_decap_8 FILLER_22_2113 ();
 sg13g2_decap_8 FILLER_22_2120 ();
 sg13g2_fill_2 FILLER_22_2127 ();
 sg13g2_fill_1 FILLER_22_2129 ();
 sg13g2_decap_8 FILLER_22_2151 ();
 sg13g2_decap_8 FILLER_22_2158 ();
 sg13g2_fill_1 FILLER_22_2168 ();
 sg13g2_fill_2 FILLER_22_2175 ();
 sg13g2_fill_1 FILLER_22_2177 ();
 sg13g2_decap_4 FILLER_22_2182 ();
 sg13g2_fill_1 FILLER_22_2186 ();
 sg13g2_decap_8 FILLER_22_2190 ();
 sg13g2_decap_4 FILLER_22_2203 ();
 sg13g2_fill_1 FILLER_22_2207 ();
 sg13g2_decap_8 FILLER_22_2236 ();
 sg13g2_fill_1 FILLER_22_2243 ();
 sg13g2_fill_1 FILLER_22_2257 ();
 sg13g2_decap_8 FILLER_22_2274 ();
 sg13g2_decap_8 FILLER_22_2281 ();
 sg13g2_fill_2 FILLER_22_2288 ();
 sg13g2_fill_1 FILLER_22_2290 ();
 sg13g2_decap_4 FILLER_22_2323 ();
 sg13g2_fill_2 FILLER_22_2340 ();
 sg13g2_fill_1 FILLER_22_2346 ();
 sg13g2_decap_4 FILLER_22_2363 ();
 sg13g2_decap_8 FILLER_22_2388 ();
 sg13g2_fill_1 FILLER_22_2400 ();
 sg13g2_decap_4 FILLER_22_2422 ();
 sg13g2_fill_1 FILLER_22_2426 ();
 sg13g2_decap_8 FILLER_22_2440 ();
 sg13g2_decap_4 FILLER_22_2447 ();
 sg13g2_fill_2 FILLER_22_2451 ();
 sg13g2_decap_4 FILLER_22_2467 ();
 sg13g2_fill_2 FILLER_22_2471 ();
 sg13g2_decap_8 FILLER_22_2477 ();
 sg13g2_decap_8 FILLER_22_2484 ();
 sg13g2_fill_2 FILLER_22_2491 ();
 sg13g2_fill_2 FILLER_22_2501 ();
 sg13g2_fill_1 FILLER_22_2520 ();
 sg13g2_decap_4 FILLER_22_2531 ();
 sg13g2_fill_2 FILLER_22_2557 ();
 sg13g2_fill_1 FILLER_22_2559 ();
 sg13g2_fill_2 FILLER_22_2616 ();
 sg13g2_fill_1 FILLER_22_2626 ();
 sg13g2_fill_1 FILLER_22_2636 ();
 sg13g2_fill_2 FILLER_22_2651 ();
 sg13g2_fill_1 FILLER_22_2670 ();
 sg13g2_decap_4 FILLER_22_2684 ();
 sg13g2_fill_1 FILLER_22_2688 ();
 sg13g2_decap_8 FILLER_22_2717 ();
 sg13g2_fill_2 FILLER_22_2724 ();
 sg13g2_fill_2 FILLER_22_2745 ();
 sg13g2_decap_8 FILLER_22_2779 ();
 sg13g2_decap_4 FILLER_22_2791 ();
 sg13g2_fill_2 FILLER_22_2795 ();
 sg13g2_fill_2 FILLER_22_2846 ();
 sg13g2_decap_8 FILLER_22_2861 ();
 sg13g2_fill_2 FILLER_22_2934 ();
 sg13g2_fill_1 FILLER_22_2936 ();
 sg13g2_decap_8 FILLER_22_2941 ();
 sg13g2_decap_4 FILLER_22_2948 ();
 sg13g2_fill_1 FILLER_22_2952 ();
 sg13g2_fill_1 FILLER_22_2968 ();
 sg13g2_fill_2 FILLER_22_2983 ();
 sg13g2_fill_1 FILLER_22_2985 ();
 sg13g2_decap_8 FILLER_22_2999 ();
 sg13g2_decap_4 FILLER_22_3006 ();
 sg13g2_decap_4 FILLER_22_3029 ();
 sg13g2_fill_1 FILLER_22_3033 ();
 sg13g2_decap_8 FILLER_22_3048 ();
 sg13g2_decap_4 FILLER_22_3055 ();
 sg13g2_fill_1 FILLER_22_3059 ();
 sg13g2_decap_4 FILLER_22_3063 ();
 sg13g2_fill_1 FILLER_22_3072 ();
 sg13g2_decap_8 FILLER_22_3086 ();
 sg13g2_decap_4 FILLER_22_3093 ();
 sg13g2_fill_2 FILLER_22_3110 ();
 sg13g2_decap_8 FILLER_22_3130 ();
 sg13g2_decap_4 FILLER_22_3137 ();
 sg13g2_fill_2 FILLER_22_3145 ();
 sg13g2_fill_2 FILLER_22_3184 ();
 sg13g2_fill_1 FILLER_22_3197 ();
 sg13g2_fill_1 FILLER_22_3208 ();
 sg13g2_fill_1 FILLER_22_3218 ();
 sg13g2_fill_1 FILLER_22_3230 ();
 sg13g2_decap_8 FILLER_22_3243 ();
 sg13g2_fill_2 FILLER_22_3277 ();
 sg13g2_decap_8 FILLER_22_3371 ();
 sg13g2_decap_8 FILLER_22_3378 ();
 sg13g2_decap_8 FILLER_22_3385 ();
 sg13g2_decap_8 FILLER_22_3392 ();
 sg13g2_decap_8 FILLER_22_3399 ();
 sg13g2_decap_8 FILLER_22_3406 ();
 sg13g2_decap_8 FILLER_22_3413 ();
 sg13g2_decap_8 FILLER_22_3420 ();
 sg13g2_decap_8 FILLER_22_3427 ();
 sg13g2_decap_8 FILLER_22_3434 ();
 sg13g2_decap_8 FILLER_22_3441 ();
 sg13g2_decap_8 FILLER_22_3448 ();
 sg13g2_decap_8 FILLER_22_3455 ();
 sg13g2_decap_8 FILLER_22_3462 ();
 sg13g2_decap_8 FILLER_22_3469 ();
 sg13g2_decap_8 FILLER_22_3476 ();
 sg13g2_decap_8 FILLER_22_3483 ();
 sg13g2_decap_8 FILLER_22_3490 ();
 sg13g2_decap_8 FILLER_22_3497 ();
 sg13g2_decap_8 FILLER_22_3504 ();
 sg13g2_decap_8 FILLER_22_3511 ();
 sg13g2_decap_8 FILLER_22_3518 ();
 sg13g2_decap_8 FILLER_22_3525 ();
 sg13g2_decap_8 FILLER_22_3532 ();
 sg13g2_decap_8 FILLER_22_3539 ();
 sg13g2_decap_8 FILLER_22_3546 ();
 sg13g2_decap_8 FILLER_22_3553 ();
 sg13g2_decap_8 FILLER_22_3560 ();
 sg13g2_decap_8 FILLER_22_3567 ();
 sg13g2_decap_4 FILLER_22_3574 ();
 sg13g2_fill_2 FILLER_22_3578 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_201 ();
 sg13g2_decap_8 FILLER_23_208 ();
 sg13g2_decap_4 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_240 ();
 sg13g2_decap_4 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_4 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_4 FILLER_23_386 ();
 sg13g2_fill_1 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_4 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_463 ();
 sg13g2_fill_2 FILLER_23_470 ();
 sg13g2_fill_1 FILLER_23_541 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_fill_2 FILLER_23_785 ();
 sg13g2_fill_2 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_832 ();
 sg13g2_fill_2 FILLER_23_839 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_1 FILLER_23_860 ();
 sg13g2_decap_4 FILLER_23_866 ();
 sg13g2_fill_2 FILLER_23_895 ();
 sg13g2_decap_4 FILLER_23_925 ();
 sg13g2_fill_2 FILLER_23_957 ();
 sg13g2_fill_1 FILLER_23_959 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_4 FILLER_23_992 ();
 sg13g2_fill_1 FILLER_23_996 ();
 sg13g2_fill_1 FILLER_23_1015 ();
 sg13g2_decap_4 FILLER_23_1033 ();
 sg13g2_fill_1 FILLER_23_1037 ();
 sg13g2_fill_2 FILLER_23_1056 ();
 sg13g2_fill_1 FILLER_23_1058 ();
 sg13g2_fill_2 FILLER_23_1064 ();
 sg13g2_decap_8 FILLER_23_1092 ();
 sg13g2_decap_8 FILLER_23_1099 ();
 sg13g2_fill_1 FILLER_23_1106 ();
 sg13g2_decap_4 FILLER_23_1112 ();
 sg13g2_fill_1 FILLER_23_1116 ();
 sg13g2_decap_8 FILLER_23_1135 ();
 sg13g2_decap_8 FILLER_23_1142 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_fill_1 FILLER_23_1161 ();
 sg13g2_fill_2 FILLER_23_1175 ();
 sg13g2_fill_1 FILLER_23_1177 ();
 sg13g2_decap_4 FILLER_23_1183 ();
 sg13g2_fill_1 FILLER_23_1187 ();
 sg13g2_fill_2 FILLER_23_1209 ();
 sg13g2_fill_1 FILLER_23_1211 ();
 sg13g2_fill_2 FILLER_23_1224 ();
 sg13g2_fill_2 FILLER_23_1231 ();
 sg13g2_decap_8 FILLER_23_1253 ();
 sg13g2_decap_4 FILLER_23_1260 ();
 sg13g2_fill_1 FILLER_23_1264 ();
 sg13g2_decap_8 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_fill_1 FILLER_23_1306 ();
 sg13g2_decap_4 FILLER_23_1320 ();
 sg13g2_fill_1 FILLER_23_1324 ();
 sg13g2_decap_4 FILLER_23_1341 ();
 sg13g2_fill_1 FILLER_23_1362 ();
 sg13g2_decap_4 FILLER_23_1376 ();
 sg13g2_fill_1 FILLER_23_1398 ();
 sg13g2_decap_4 FILLER_23_1407 ();
 sg13g2_fill_2 FILLER_23_1421 ();
 sg13g2_decap_8 FILLER_23_1436 ();
 sg13g2_decap_4 FILLER_23_1443 ();
 sg13g2_decap_8 FILLER_23_1454 ();
 sg13g2_decap_4 FILLER_23_1461 ();
 sg13g2_fill_2 FILLER_23_1465 ();
 sg13g2_decap_8 FILLER_23_1500 ();
 sg13g2_fill_1 FILLER_23_1507 ();
 sg13g2_decap_8 FILLER_23_1523 ();
 sg13g2_decap_8 FILLER_23_1530 ();
 sg13g2_fill_2 FILLER_23_1549 ();
 sg13g2_fill_2 FILLER_23_1564 ();
 sg13g2_fill_1 FILLER_23_1566 ();
 sg13g2_fill_2 FILLER_23_1611 ();
 sg13g2_fill_1 FILLER_23_1613 ();
 sg13g2_decap_8 FILLER_23_1626 ();
 sg13g2_decap_4 FILLER_23_1633 ();
 sg13g2_decap_4 FILLER_23_1642 ();
 sg13g2_fill_2 FILLER_23_1646 ();
 sg13g2_decap_8 FILLER_23_1665 ();
 sg13g2_fill_2 FILLER_23_1672 ();
 sg13g2_fill_1 FILLER_23_1674 ();
 sg13g2_fill_2 FILLER_23_1695 ();
 sg13g2_fill_1 FILLER_23_1697 ();
 sg13g2_fill_2 FILLER_23_1706 ();
 sg13g2_fill_1 FILLER_23_1708 ();
 sg13g2_decap_8 FILLER_23_1713 ();
 sg13g2_decap_8 FILLER_23_1720 ();
 sg13g2_decap_8 FILLER_23_1727 ();
 sg13g2_fill_1 FILLER_23_1734 ();
 sg13g2_decap_8 FILLER_23_1782 ();
 sg13g2_decap_8 FILLER_23_1789 ();
 sg13g2_decap_8 FILLER_23_1801 ();
 sg13g2_decap_8 FILLER_23_1808 ();
 sg13g2_decap_4 FILLER_23_1815 ();
 sg13g2_decap_8 FILLER_23_1823 ();
 sg13g2_decap_4 FILLER_23_1830 ();
 sg13g2_decap_4 FILLER_23_1862 ();
 sg13g2_fill_1 FILLER_23_1866 ();
 sg13g2_decap_8 FILLER_23_1871 ();
 sg13g2_decap_4 FILLER_23_1878 ();
 sg13g2_fill_1 FILLER_23_1882 ();
 sg13g2_fill_2 FILLER_23_1910 ();
 sg13g2_fill_1 FILLER_23_1912 ();
 sg13g2_decap_4 FILLER_23_1921 ();
 sg13g2_decap_8 FILLER_23_1936 ();
 sg13g2_decap_8 FILLER_23_1943 ();
 sg13g2_decap_8 FILLER_23_1950 ();
 sg13g2_fill_1 FILLER_23_1957 ();
 sg13g2_decap_8 FILLER_23_1964 ();
 sg13g2_fill_1 FILLER_23_1971 ();
 sg13g2_fill_2 FILLER_23_1985 ();
 sg13g2_decap_4 FILLER_23_1992 ();
 sg13g2_fill_1 FILLER_23_1996 ();
 sg13g2_decap_4 FILLER_23_2001 ();
 sg13g2_fill_2 FILLER_23_2005 ();
 sg13g2_fill_2 FILLER_23_2010 ();
 sg13g2_decap_8 FILLER_23_2017 ();
 sg13g2_fill_2 FILLER_23_2024 ();
 sg13g2_fill_1 FILLER_23_2045 ();
 sg13g2_fill_2 FILLER_23_2067 ();
 sg13g2_fill_1 FILLER_23_2095 ();
 sg13g2_decap_8 FILLER_23_2113 ();
 sg13g2_decap_8 FILLER_23_2120 ();
 sg13g2_fill_2 FILLER_23_2127 ();
 sg13g2_fill_1 FILLER_23_2129 ();
 sg13g2_fill_2 FILLER_23_2158 ();
 sg13g2_decap_4 FILLER_23_2176 ();
 sg13g2_fill_1 FILLER_23_2180 ();
 sg13g2_decap_4 FILLER_23_2255 ();
 sg13g2_fill_2 FILLER_23_2291 ();
 sg13g2_fill_1 FILLER_23_2293 ();
 sg13g2_fill_2 FILLER_23_2333 ();
 sg13g2_fill_1 FILLER_23_2343 ();
 sg13g2_decap_8 FILLER_23_2356 ();
 sg13g2_decap_4 FILLER_23_2363 ();
 sg13g2_fill_2 FILLER_23_2367 ();
 sg13g2_decap_8 FILLER_23_2387 ();
 sg13g2_decap_4 FILLER_23_2394 ();
 sg13g2_decap_8 FILLER_23_2413 ();
 sg13g2_decap_8 FILLER_23_2420 ();
 sg13g2_fill_2 FILLER_23_2427 ();
 sg13g2_decap_8 FILLER_23_2437 ();
 sg13g2_fill_2 FILLER_23_2457 ();
 sg13g2_fill_1 FILLER_23_2459 ();
 sg13g2_fill_2 FILLER_23_2464 ();
 sg13g2_fill_1 FILLER_23_2466 ();
 sg13g2_fill_2 FILLER_23_2524 ();
 sg13g2_fill_1 FILLER_23_2526 ();
 sg13g2_fill_2 FILLER_23_2548 ();
 sg13g2_fill_1 FILLER_23_2550 ();
 sg13g2_decap_4 FILLER_23_2567 ();
 sg13g2_fill_1 FILLER_23_2571 ();
 sg13g2_decap_4 FILLER_23_2581 ();
 sg13g2_fill_1 FILLER_23_2585 ();
 sg13g2_fill_1 FILLER_23_2604 ();
 sg13g2_fill_2 FILLER_23_2617 ();
 sg13g2_fill_1 FILLER_23_2619 ();
 sg13g2_decap_4 FILLER_23_2625 ();
 sg13g2_fill_1 FILLER_23_2629 ();
 sg13g2_fill_2 FILLER_23_2648 ();
 sg13g2_fill_1 FILLER_23_2650 ();
 sg13g2_fill_2 FILLER_23_2659 ();
 sg13g2_fill_1 FILLER_23_2666 ();
 sg13g2_decap_8 FILLER_23_2677 ();
 sg13g2_decap_4 FILLER_23_2684 ();
 sg13g2_decap_8 FILLER_23_2699 ();
 sg13g2_decap_8 FILLER_23_2706 ();
 sg13g2_fill_1 FILLER_23_2713 ();
 sg13g2_decap_8 FILLER_23_2718 ();
 sg13g2_fill_1 FILLER_23_2725 ();
 sg13g2_decap_8 FILLER_23_2746 ();
 sg13g2_decap_8 FILLER_23_2753 ();
 sg13g2_decap_8 FILLER_23_2770 ();
 sg13g2_decap_4 FILLER_23_2777 ();
 sg13g2_decap_8 FILLER_23_2797 ();
 sg13g2_decap_4 FILLER_23_2804 ();
 sg13g2_fill_1 FILLER_23_2808 ();
 sg13g2_fill_2 FILLER_23_2827 ();
 sg13g2_fill_1 FILLER_23_2829 ();
 sg13g2_decap_8 FILLER_23_2833 ();
 sg13g2_fill_2 FILLER_23_2840 ();
 sg13g2_fill_2 FILLER_23_2930 ();
 sg13g2_fill_2 FILLER_23_2995 ();
 sg13g2_fill_2 FILLER_23_3016 ();
 sg13g2_fill_2 FILLER_23_3029 ();
 sg13g2_fill_1 FILLER_23_3031 ();
 sg13g2_fill_2 FILLER_23_3055 ();
 sg13g2_fill_1 FILLER_23_3057 ();
 sg13g2_fill_2 FILLER_23_3071 ();
 sg13g2_fill_2 FILLER_23_3086 ();
 sg13g2_fill_2 FILLER_23_3091 ();
 sg13g2_fill_1 FILLER_23_3093 ();
 sg13g2_fill_2 FILLER_23_3102 ();
 sg13g2_fill_1 FILLER_23_3104 ();
 sg13g2_fill_2 FILLER_23_3119 ();
 sg13g2_decap_8 FILLER_23_3126 ();
 sg13g2_fill_2 FILLER_23_3133 ();
 sg13g2_fill_1 FILLER_23_3135 ();
 sg13g2_decap_4 FILLER_23_3159 ();
 sg13g2_fill_1 FILLER_23_3163 ();
 sg13g2_decap_8 FILLER_23_3181 ();
 sg13g2_fill_2 FILLER_23_3188 ();
 sg13g2_decap_8 FILLER_23_3213 ();
 sg13g2_decap_4 FILLER_23_3220 ();
 sg13g2_fill_1 FILLER_23_3224 ();
 sg13g2_fill_2 FILLER_23_3253 ();
 sg13g2_decap_8 FILLER_23_3262 ();
 sg13g2_fill_2 FILLER_23_3298 ();
 sg13g2_fill_2 FILLER_23_3313 ();
 sg13g2_decap_8 FILLER_23_3349 ();
 sg13g2_decap_8 FILLER_23_3365 ();
 sg13g2_decap_8 FILLER_23_3372 ();
 sg13g2_decap_8 FILLER_23_3379 ();
 sg13g2_decap_8 FILLER_23_3386 ();
 sg13g2_decap_8 FILLER_23_3393 ();
 sg13g2_decap_8 FILLER_23_3400 ();
 sg13g2_decap_8 FILLER_23_3407 ();
 sg13g2_decap_8 FILLER_23_3414 ();
 sg13g2_decap_8 FILLER_23_3421 ();
 sg13g2_decap_8 FILLER_23_3428 ();
 sg13g2_decap_8 FILLER_23_3435 ();
 sg13g2_decap_8 FILLER_23_3442 ();
 sg13g2_decap_8 FILLER_23_3449 ();
 sg13g2_decap_8 FILLER_23_3456 ();
 sg13g2_decap_8 FILLER_23_3463 ();
 sg13g2_decap_8 FILLER_23_3470 ();
 sg13g2_decap_8 FILLER_23_3477 ();
 sg13g2_decap_8 FILLER_23_3484 ();
 sg13g2_decap_8 FILLER_23_3491 ();
 sg13g2_decap_8 FILLER_23_3498 ();
 sg13g2_decap_8 FILLER_23_3505 ();
 sg13g2_decap_8 FILLER_23_3512 ();
 sg13g2_decap_8 FILLER_23_3519 ();
 sg13g2_decap_8 FILLER_23_3526 ();
 sg13g2_decap_8 FILLER_23_3533 ();
 sg13g2_decap_8 FILLER_23_3540 ();
 sg13g2_decap_8 FILLER_23_3547 ();
 sg13g2_decap_8 FILLER_23_3554 ();
 sg13g2_decap_8 FILLER_23_3561 ();
 sg13g2_decap_8 FILLER_23_3568 ();
 sg13g2_decap_4 FILLER_23_3575 ();
 sg13g2_fill_1 FILLER_23_3579 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_24_415 ();
 sg13g2_fill_1 FILLER_24_419 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_442 ();
 sg13g2_fill_1 FILLER_24_471 ();
 sg13g2_decap_8 FILLER_24_481 ();
 sg13g2_decap_8 FILLER_24_488 ();
 sg13g2_decap_8 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_fill_2 FILLER_24_516 ();
 sg13g2_fill_1 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_4 FILLER_24_571 ();
 sg13g2_fill_2 FILLER_24_575 ();
 sg13g2_fill_1 FILLER_24_590 ();
 sg13g2_fill_1 FILLER_24_595 ();
 sg13g2_fill_1 FILLER_24_605 ();
 sg13g2_fill_1 FILLER_24_610 ();
 sg13g2_decap_8 FILLER_24_624 ();
 sg13g2_fill_2 FILLER_24_631 ();
 sg13g2_fill_2 FILLER_24_680 ();
 sg13g2_decap_4 FILLER_24_691 ();
 sg13g2_fill_2 FILLER_24_695 ();
 sg13g2_fill_1 FILLER_24_734 ();
 sg13g2_decap_4 FILLER_24_771 ();
 sg13g2_fill_1 FILLER_24_775 ();
 sg13g2_fill_1 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_fill_1 FILLER_24_803 ();
 sg13g2_fill_2 FILLER_24_816 ();
 sg13g2_fill_2 FILLER_24_842 ();
 sg13g2_fill_1 FILLER_24_844 ();
 sg13g2_fill_2 FILLER_24_850 ();
 sg13g2_decap_4 FILLER_24_870 ();
 sg13g2_fill_1 FILLER_24_892 ();
 sg13g2_decap_8 FILLER_24_898 ();
 sg13g2_decap_8 FILLER_24_905 ();
 sg13g2_fill_2 FILLER_24_912 ();
 sg13g2_decap_8 FILLER_24_933 ();
 sg13g2_decap_8 FILLER_24_940 ();
 sg13g2_decap_8 FILLER_24_947 ();
 sg13g2_decap_4 FILLER_24_954 ();
 sg13g2_fill_1 FILLER_24_958 ();
 sg13g2_decap_8 FILLER_24_985 ();
 sg13g2_decap_8 FILLER_24_1010 ();
 sg13g2_decap_4 FILLER_24_1017 ();
 sg13g2_fill_2 FILLER_24_1021 ();
 sg13g2_decap_8 FILLER_24_1033 ();
 sg13g2_fill_1 FILLER_24_1040 ();
 sg13g2_decap_8 FILLER_24_1058 ();
 sg13g2_decap_4 FILLER_24_1065 ();
 sg13g2_fill_2 FILLER_24_1097 ();
 sg13g2_fill_1 FILLER_24_1099 ();
 sg13g2_fill_2 FILLER_24_1118 ();
 sg13g2_fill_1 FILLER_24_1120 ();
 sg13g2_decap_8 FILLER_24_1142 ();
 sg13g2_decap_4 FILLER_24_1149 ();
 sg13g2_decap_8 FILLER_24_1168 ();
 sg13g2_decap_8 FILLER_24_1182 ();
 sg13g2_fill_1 FILLER_24_1189 ();
 sg13g2_fill_2 FILLER_24_1204 ();
 sg13g2_decap_8 FILLER_24_1238 ();
 sg13g2_decap_8 FILLER_24_1245 ();
 sg13g2_decap_8 FILLER_24_1252 ();
 sg13g2_decap_8 FILLER_24_1259 ();
 sg13g2_decap_4 FILLER_24_1266 ();
 sg13g2_decap_4 FILLER_24_1301 ();
 sg13g2_decap_4 FILLER_24_1310 ();
 sg13g2_fill_2 FILLER_24_1336 ();
 sg13g2_decap_8 FILLER_24_1350 ();
 sg13g2_decap_4 FILLER_24_1357 ();
 sg13g2_fill_1 FILLER_24_1361 ();
 sg13g2_decap_4 FILLER_24_1376 ();
 sg13g2_fill_2 FILLER_24_1380 ();
 sg13g2_fill_2 FILLER_24_1391 ();
 sg13g2_fill_1 FILLER_24_1393 ();
 sg13g2_decap_4 FILLER_24_1407 ();
 sg13g2_fill_1 FILLER_24_1411 ();
 sg13g2_decap_8 FILLER_24_1430 ();
 sg13g2_decap_8 FILLER_24_1437 ();
 sg13g2_fill_1 FILLER_24_1472 ();
 sg13g2_decap_8 FILLER_24_1477 ();
 sg13g2_decap_4 FILLER_24_1493 ();
 sg13g2_fill_2 FILLER_24_1497 ();
 sg13g2_decap_4 FILLER_24_1512 ();
 sg13g2_decap_4 FILLER_24_1525 ();
 sg13g2_fill_2 FILLER_24_1529 ();
 sg13g2_decap_4 FILLER_24_1540 ();
 sg13g2_fill_1 FILLER_24_1544 ();
 sg13g2_decap_8 FILLER_24_1559 ();
 sg13g2_decap_8 FILLER_24_1566 ();
 sg13g2_decap_4 FILLER_24_1573 ();
 sg13g2_fill_1 FILLER_24_1577 ();
 sg13g2_decap_8 FILLER_24_1583 ();
 sg13g2_decap_4 FILLER_24_1590 ();
 sg13g2_fill_1 FILLER_24_1594 ();
 sg13g2_fill_1 FILLER_24_1603 ();
 sg13g2_fill_1 FILLER_24_1614 ();
 sg13g2_fill_1 FILLER_24_1624 ();
 sg13g2_fill_2 FILLER_24_1630 ();
 sg13g2_fill_1 FILLER_24_1632 ();
 sg13g2_decap_8 FILLER_24_1664 ();
 sg13g2_decap_4 FILLER_24_1671 ();
 sg13g2_decap_8 FILLER_24_1715 ();
 sg13g2_fill_2 FILLER_24_1722 ();
 sg13g2_fill_1 FILLER_24_1724 ();
 sg13g2_decap_8 FILLER_24_1754 ();
 sg13g2_decap_4 FILLER_24_1761 ();
 sg13g2_fill_1 FILLER_24_1765 ();
 sg13g2_fill_2 FILLER_24_1776 ();
 sg13g2_decap_8 FILLER_24_1811 ();
 sg13g2_decap_4 FILLER_24_1818 ();
 sg13g2_fill_1 FILLER_24_1822 ();
 sg13g2_decap_8 FILLER_24_1847 ();
 sg13g2_fill_1 FILLER_24_1854 ();
 sg13g2_fill_2 FILLER_24_1861 ();
 sg13g2_decap_8 FILLER_24_1873 ();
 sg13g2_decap_8 FILLER_24_1880 ();
 sg13g2_fill_2 FILLER_24_1893 ();
 sg13g2_fill_2 FILLER_24_1899 ();
 sg13g2_fill_1 FILLER_24_1901 ();
 sg13g2_fill_2 FILLER_24_1914 ();
 sg13g2_fill_2 FILLER_24_1929 ();
 sg13g2_fill_2 FILLER_24_1950 ();
 sg13g2_fill_1 FILLER_24_1972 ();
 sg13g2_fill_2 FILLER_24_1978 ();
 sg13g2_fill_1 FILLER_24_1980 ();
 sg13g2_decap_8 FILLER_24_1989 ();
 sg13g2_fill_2 FILLER_24_1996 ();
 sg13g2_fill_2 FILLER_24_2028 ();
 sg13g2_fill_2 FILLER_24_2038 ();
 sg13g2_fill_2 FILLER_24_2053 ();
 sg13g2_fill_2 FILLER_24_2063 ();
 sg13g2_decap_4 FILLER_24_2074 ();
 sg13g2_fill_1 FILLER_24_2078 ();
 sg13g2_decap_8 FILLER_24_2117 ();
 sg13g2_decap_8 FILLER_24_2124 ();
 sg13g2_decap_8 FILLER_24_2134 ();
 sg13g2_fill_1 FILLER_24_2141 ();
 sg13g2_decap_8 FILLER_24_2155 ();
 sg13g2_fill_1 FILLER_24_2194 ();
 sg13g2_decap_8 FILLER_24_2199 ();
 sg13g2_decap_8 FILLER_24_2206 ();
 sg13g2_fill_2 FILLER_24_2213 ();
 sg13g2_decap_4 FILLER_24_2254 ();
 sg13g2_fill_1 FILLER_24_2258 ();
 sg13g2_decap_8 FILLER_24_2276 ();
 sg13g2_fill_2 FILLER_24_2283 ();
 sg13g2_decap_8 FILLER_24_2300 ();
 sg13g2_decap_4 FILLER_24_2307 ();
 sg13g2_fill_1 FILLER_24_2311 ();
 sg13g2_fill_1 FILLER_24_2329 ();
 sg13g2_fill_2 FILLER_24_2353 ();
 sg13g2_fill_2 FILLER_24_2371 ();
 sg13g2_fill_1 FILLER_24_2373 ();
 sg13g2_fill_2 FILLER_24_2384 ();
 sg13g2_decap_8 FILLER_24_2391 ();
 sg13g2_fill_2 FILLER_24_2398 ();
 sg13g2_fill_2 FILLER_24_2417 ();
 sg13g2_fill_1 FILLER_24_2419 ();
 sg13g2_fill_1 FILLER_24_2441 ();
 sg13g2_decap_8 FILLER_24_2483 ();
 sg13g2_fill_1 FILLER_24_2490 ();
 sg13g2_decap_4 FILLER_24_2522 ();
 sg13g2_fill_1 FILLER_24_2554 ();
 sg13g2_fill_2 FILLER_24_2638 ();
 sg13g2_fill_1 FILLER_24_2640 ();
 sg13g2_fill_2 FILLER_24_2654 ();
 sg13g2_decap_8 FILLER_24_2669 ();
 sg13g2_fill_2 FILLER_24_2676 ();
 sg13g2_decap_8 FILLER_24_2685 ();
 sg13g2_decap_8 FILLER_24_2692 ();
 sg13g2_decap_4 FILLER_24_2699 ();
 sg13g2_fill_2 FILLER_24_2703 ();
 sg13g2_fill_2 FILLER_24_2720 ();
 sg13g2_fill_2 FILLER_24_2752 ();
 sg13g2_fill_2 FILLER_24_2776 ();
 sg13g2_fill_1 FILLER_24_2778 ();
 sg13g2_fill_1 FILLER_24_2784 ();
 sg13g2_decap_8 FILLER_24_2801 ();
 sg13g2_fill_1 FILLER_24_2825 ();
 sg13g2_decap_4 FILLER_24_2867 ();
 sg13g2_decap_8 FILLER_24_2935 ();
 sg13g2_decap_8 FILLER_24_2942 ();
 sg13g2_decap_4 FILLER_24_2949 ();
 sg13g2_decap_8 FILLER_24_2969 ();
 sg13g2_decap_8 FILLER_24_2976 ();
 sg13g2_decap_8 FILLER_24_2992 ();
 sg13g2_fill_1 FILLER_24_2999 ();
 sg13g2_decap_4 FILLER_24_3009 ();
 sg13g2_decap_4 FILLER_24_3030 ();
 sg13g2_fill_1 FILLER_24_3034 ();
 sg13g2_decap_8 FILLER_24_3043 ();
 sg13g2_fill_2 FILLER_24_3050 ();
 sg13g2_fill_2 FILLER_24_3064 ();
 sg13g2_fill_1 FILLER_24_3066 ();
 sg13g2_decap_4 FILLER_24_3083 ();
 sg13g2_decap_4 FILLER_24_3095 ();
 sg13g2_fill_2 FILLER_24_3099 ();
 sg13g2_decap_8 FILLER_24_3106 ();
 sg13g2_fill_2 FILLER_24_3113 ();
 sg13g2_decap_8 FILLER_24_3127 ();
 sg13g2_decap_4 FILLER_24_3134 ();
 sg13g2_fill_1 FILLER_24_3138 ();
 sg13g2_fill_2 FILLER_24_3143 ();
 sg13g2_fill_1 FILLER_24_3145 ();
 sg13g2_decap_8 FILLER_24_3164 ();
 sg13g2_decap_8 FILLER_24_3171 ();
 sg13g2_decap_8 FILLER_24_3178 ();
 sg13g2_decap_8 FILLER_24_3204 ();
 sg13g2_decap_4 FILLER_24_3211 ();
 sg13g2_fill_1 FILLER_24_3215 ();
 sg13g2_decap_8 FILLER_24_3243 ();
 sg13g2_decap_8 FILLER_24_3250 ();
 sg13g2_decap_4 FILLER_24_3257 ();
 sg13g2_fill_2 FILLER_24_3308 ();
 sg13g2_fill_1 FILLER_24_3310 ();
 sg13g2_fill_2 FILLER_24_3324 ();
 sg13g2_fill_1 FILLER_24_3326 ();
 sg13g2_fill_2 FILLER_24_3344 ();
 sg13g2_decap_8 FILLER_24_3374 ();
 sg13g2_decap_8 FILLER_24_3381 ();
 sg13g2_decap_8 FILLER_24_3388 ();
 sg13g2_decap_8 FILLER_24_3395 ();
 sg13g2_decap_8 FILLER_24_3402 ();
 sg13g2_decap_8 FILLER_24_3409 ();
 sg13g2_decap_8 FILLER_24_3416 ();
 sg13g2_decap_8 FILLER_24_3423 ();
 sg13g2_decap_8 FILLER_24_3430 ();
 sg13g2_decap_8 FILLER_24_3437 ();
 sg13g2_decap_8 FILLER_24_3444 ();
 sg13g2_decap_8 FILLER_24_3451 ();
 sg13g2_decap_8 FILLER_24_3458 ();
 sg13g2_decap_8 FILLER_24_3465 ();
 sg13g2_decap_8 FILLER_24_3472 ();
 sg13g2_decap_8 FILLER_24_3479 ();
 sg13g2_decap_8 FILLER_24_3486 ();
 sg13g2_decap_8 FILLER_24_3493 ();
 sg13g2_decap_8 FILLER_24_3500 ();
 sg13g2_decap_8 FILLER_24_3507 ();
 sg13g2_decap_8 FILLER_24_3514 ();
 sg13g2_decap_8 FILLER_24_3521 ();
 sg13g2_decap_8 FILLER_24_3528 ();
 sg13g2_decap_8 FILLER_24_3535 ();
 sg13g2_decap_8 FILLER_24_3542 ();
 sg13g2_decap_8 FILLER_24_3549 ();
 sg13g2_decap_8 FILLER_24_3556 ();
 sg13g2_decap_8 FILLER_24_3563 ();
 sg13g2_decap_8 FILLER_24_3570 ();
 sg13g2_fill_2 FILLER_24_3577 ();
 sg13g2_fill_1 FILLER_24_3579 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_4 FILLER_25_349 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_decap_4 FILLER_25_390 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_25_432 ();
 sg13g2_decap_4 FILLER_25_439 ();
 sg13g2_fill_2 FILLER_25_443 ();
 sg13g2_fill_2 FILLER_25_452 ();
 sg13g2_fill_1 FILLER_25_454 ();
 sg13g2_decap_4 FILLER_25_461 ();
 sg13g2_fill_2 FILLER_25_478 ();
 sg13g2_fill_1 FILLER_25_480 ();
 sg13g2_fill_2 FILLER_25_489 ();
 sg13g2_decap_8 FILLER_25_503 ();
 sg13g2_decap_8 FILLER_25_528 ();
 sg13g2_decap_4 FILLER_25_535 ();
 sg13g2_fill_2 FILLER_25_539 ();
 sg13g2_fill_1 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_558 ();
 sg13g2_decap_8 FILLER_25_565 ();
 sg13g2_fill_1 FILLER_25_572 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_fill_1 FILLER_25_613 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_4 FILLER_25_672 ();
 sg13g2_fill_2 FILLER_25_708 ();
 sg13g2_fill_2 FILLER_25_723 ();
 sg13g2_fill_2 FILLER_25_734 ();
 sg13g2_fill_2 FILLER_25_744 ();
 sg13g2_fill_1 FILLER_25_746 ();
 sg13g2_fill_2 FILLER_25_762 ();
 sg13g2_fill_1 FILLER_25_769 ();
 sg13g2_decap_4 FILLER_25_774 ();
 sg13g2_fill_2 FILLER_25_778 ();
 sg13g2_decap_4 FILLER_25_824 ();
 sg13g2_fill_1 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_fill_1 FILLER_25_854 ();
 sg13g2_fill_2 FILLER_25_859 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_1 FILLER_25_889 ();
 sg13g2_decap_8 FILLER_25_903 ();
 sg13g2_fill_1 FILLER_25_910 ();
 sg13g2_decap_8 FILLER_25_936 ();
 sg13g2_fill_2 FILLER_25_943 ();
 sg13g2_fill_1 FILLER_25_945 ();
 sg13g2_decap_4 FILLER_25_951 ();
 sg13g2_fill_1 FILLER_25_955 ();
 sg13g2_decap_4 FILLER_25_960 ();
 sg13g2_decap_8 FILLER_25_983 ();
 sg13g2_fill_2 FILLER_25_990 ();
 sg13g2_fill_1 FILLER_25_992 ();
 sg13g2_fill_2 FILLER_25_1013 ();
 sg13g2_fill_1 FILLER_25_1015 ();
 sg13g2_decap_4 FILLER_25_1032 ();
 sg13g2_decap_8 FILLER_25_1041 ();
 sg13g2_fill_1 FILLER_25_1048 ();
 sg13g2_decap_8 FILLER_25_1057 ();
 sg13g2_fill_2 FILLER_25_1064 ();
 sg13g2_fill_2 FILLER_25_1092 ();
 sg13g2_fill_1 FILLER_25_1094 ();
 sg13g2_fill_2 FILLER_25_1116 ();
 sg13g2_fill_2 FILLER_25_1138 ();
 sg13g2_fill_1 FILLER_25_1140 ();
 sg13g2_fill_2 FILLER_25_1159 ();
 sg13g2_fill_1 FILLER_25_1161 ();
 sg13g2_decap_4 FILLER_25_1167 ();
 sg13g2_fill_2 FILLER_25_1171 ();
 sg13g2_fill_2 FILLER_25_1201 ();
 sg13g2_fill_1 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1210 ();
 sg13g2_fill_2 FILLER_25_1217 ();
 sg13g2_fill_1 FILLER_25_1219 ();
 sg13g2_decap_8 FILLER_25_1225 ();
 sg13g2_decap_4 FILLER_25_1232 ();
 sg13g2_fill_2 FILLER_25_1271 ();
 sg13g2_fill_1 FILLER_25_1273 ();
 sg13g2_decap_8 FILLER_25_1287 ();
 sg13g2_fill_1 FILLER_25_1294 ();
 sg13g2_decap_8 FILLER_25_1314 ();
 sg13g2_decap_8 FILLER_25_1321 ();
 sg13g2_decap_4 FILLER_25_1328 ();
 sg13g2_fill_2 FILLER_25_1332 ();
 sg13g2_fill_1 FILLER_25_1343 ();
 sg13g2_decap_8 FILLER_25_1349 ();
 sg13g2_decap_4 FILLER_25_1356 ();
 sg13g2_fill_1 FILLER_25_1360 ();
 sg13g2_fill_1 FILLER_25_1393 ();
 sg13g2_fill_2 FILLER_25_1399 ();
 sg13g2_decap_4 FILLER_25_1409 ();
 sg13g2_fill_2 FILLER_25_1413 ();
 sg13g2_fill_2 FILLER_25_1448 ();
 sg13g2_fill_1 FILLER_25_1454 ();
 sg13g2_decap_8 FILLER_25_1465 ();
 sg13g2_decap_8 FILLER_25_1472 ();
 sg13g2_decap_4 FILLER_25_1479 ();
 sg13g2_fill_2 FILLER_25_1483 ();
 sg13g2_fill_2 FILLER_25_1507 ();
 sg13g2_fill_1 FILLER_25_1509 ();
 sg13g2_decap_8 FILLER_25_1542 ();
 sg13g2_fill_2 FILLER_25_1549 ();
 sg13g2_fill_1 FILLER_25_1551 ();
 sg13g2_fill_1 FILLER_25_1559 ();
 sg13g2_decap_4 FILLER_25_1591 ();
 sg13g2_fill_1 FILLER_25_1595 ();
 sg13g2_fill_2 FILLER_25_1609 ();
 sg13g2_fill_2 FILLER_25_1619 ();
 sg13g2_decap_8 FILLER_25_1637 ();
 sg13g2_decap_8 FILLER_25_1644 ();
 sg13g2_decap_4 FILLER_25_1651 ();
 sg13g2_fill_1 FILLER_25_1655 ();
 sg13g2_decap_8 FILLER_25_1661 ();
 sg13g2_decap_8 FILLER_25_1668 ();
 sg13g2_decap_8 FILLER_25_1675 ();
 sg13g2_fill_2 FILLER_25_1691 ();
 sg13g2_fill_2 FILLER_25_1717 ();
 sg13g2_fill_1 FILLER_25_1719 ();
 sg13g2_fill_1 FILLER_25_1730 ();
 sg13g2_fill_2 FILLER_25_1735 ();
 sg13g2_decap_4 FILLER_25_1747 ();
 sg13g2_fill_1 FILLER_25_1751 ();
 sg13g2_decap_4 FILLER_25_1758 ();
 sg13g2_fill_1 FILLER_25_1762 ();
 sg13g2_fill_2 FILLER_25_1776 ();
 sg13g2_decap_8 FILLER_25_1801 ();
 sg13g2_fill_1 FILLER_25_1812 ();
 sg13g2_fill_2 FILLER_25_1822 ();
 sg13g2_decap_8 FILLER_25_1837 ();
 sg13g2_decap_4 FILLER_25_1844 ();
 sg13g2_fill_2 FILLER_25_1848 ();
 sg13g2_fill_1 FILLER_25_1858 ();
 sg13g2_fill_2 FILLER_25_1881 ();
 sg13g2_fill_1 FILLER_25_1883 ();
 sg13g2_decap_8 FILLER_25_1910 ();
 sg13g2_fill_2 FILLER_25_1917 ();
 sg13g2_fill_1 FILLER_25_1919 ();
 sg13g2_fill_2 FILLER_25_1942 ();
 sg13g2_fill_2 FILLER_25_1957 ();
 sg13g2_fill_1 FILLER_25_1959 ();
 sg13g2_decap_8 FILLER_25_1999 ();
 sg13g2_fill_2 FILLER_25_2006 ();
 sg13g2_fill_1 FILLER_25_2011 ();
 sg13g2_decap_8 FILLER_25_2016 ();
 sg13g2_decap_8 FILLER_25_2023 ();
 sg13g2_decap_4 FILLER_25_2030 ();
 sg13g2_fill_2 FILLER_25_2034 ();
 sg13g2_decap_4 FILLER_25_2044 ();
 sg13g2_fill_2 FILLER_25_2048 ();
 sg13g2_fill_2 FILLER_25_2055 ();
 sg13g2_fill_2 FILLER_25_2062 ();
 sg13g2_fill_1 FILLER_25_2072 ();
 sg13g2_fill_1 FILLER_25_2091 ();
 sg13g2_fill_2 FILLER_25_2101 ();
 sg13g2_decap_8 FILLER_25_2114 ();
 sg13g2_decap_4 FILLER_25_2121 ();
 sg13g2_fill_2 FILLER_25_2125 ();
 sg13g2_fill_2 FILLER_25_2154 ();
 sg13g2_fill_2 FILLER_25_2166 ();
 sg13g2_decap_8 FILLER_25_2175 ();
 sg13g2_decap_4 FILLER_25_2182 ();
 sg13g2_decap_8 FILLER_25_2200 ();
 sg13g2_decap_4 FILLER_25_2207 ();
 sg13g2_fill_1 FILLER_25_2211 ();
 sg13g2_fill_2 FILLER_25_2229 ();
 sg13g2_fill_2 FILLER_25_2329 ();
 sg13g2_decap_8 FILLER_25_2343 ();
 sg13g2_decap_4 FILLER_25_2350 ();
 sg13g2_decap_8 FILLER_25_2367 ();
 sg13g2_decap_8 FILLER_25_2391 ();
 sg13g2_decap_8 FILLER_25_2398 ();
 sg13g2_decap_8 FILLER_25_2420 ();
 sg13g2_fill_1 FILLER_25_2427 ();
 sg13g2_decap_4 FILLER_25_2437 ();
 sg13g2_fill_1 FILLER_25_2456 ();
 sg13g2_fill_2 FILLER_25_2460 ();
 sg13g2_decap_8 FILLER_25_2490 ();
 sg13g2_fill_2 FILLER_25_2497 ();
 sg13g2_decap_8 FILLER_25_2503 ();
 sg13g2_decap_8 FILLER_25_2510 ();
 sg13g2_decap_8 FILLER_25_2517 ();
 sg13g2_decap_4 FILLER_25_2524 ();
 sg13g2_decap_8 FILLER_25_2540 ();
 sg13g2_decap_8 FILLER_25_2547 ();
 sg13g2_decap_8 FILLER_25_2554 ();
 sg13g2_fill_1 FILLER_25_2574 ();
 sg13g2_decap_4 FILLER_25_2580 ();
 sg13g2_decap_8 FILLER_25_2612 ();
 sg13g2_decap_8 FILLER_25_2619 ();
 sg13g2_decap_4 FILLER_25_2642 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_decap_4 FILLER_25_2669 ();
 sg13g2_fill_2 FILLER_25_2673 ();
 sg13g2_fill_2 FILLER_25_2703 ();
 sg13g2_fill_1 FILLER_25_2705 ();
 sg13g2_decap_8 FILLER_25_2724 ();
 sg13g2_fill_2 FILLER_25_2748 ();
 sg13g2_fill_1 FILLER_25_2750 ();
 sg13g2_fill_2 FILLER_25_2784 ();
 sg13g2_fill_1 FILLER_25_2786 ();
 sg13g2_fill_2 FILLER_25_2792 ();
 sg13g2_fill_1 FILLER_25_2794 ();
 sg13g2_decap_4 FILLER_25_2803 ();
 sg13g2_decap_8 FILLER_25_2827 ();
 sg13g2_decap_4 FILLER_25_2834 ();
 sg13g2_fill_2 FILLER_25_2838 ();
 sg13g2_decap_8 FILLER_25_2844 ();
 sg13g2_fill_1 FILLER_25_2866 ();
 sg13g2_decap_4 FILLER_25_2871 ();
 sg13g2_fill_2 FILLER_25_2875 ();
 sg13g2_decap_4 FILLER_25_2884 ();
 sg13g2_decap_8 FILLER_25_2893 ();
 sg13g2_decap_8 FILLER_25_2900 ();
 sg13g2_fill_2 FILLER_25_2907 ();
 sg13g2_decap_8 FILLER_25_2918 ();
 sg13g2_decap_4 FILLER_25_2925 ();
 sg13g2_fill_1 FILLER_25_2929 ();
 sg13g2_decap_4 FILLER_25_2933 ();
 sg13g2_fill_1 FILLER_25_2937 ();
 sg13g2_decap_4 FILLER_25_2949 ();
 sg13g2_fill_1 FILLER_25_2984 ();
 sg13g2_decap_4 FILLER_25_3013 ();
 sg13g2_decap_8 FILLER_25_3045 ();
 sg13g2_fill_2 FILLER_25_3052 ();
 sg13g2_fill_1 FILLER_25_3054 ();
 sg13g2_fill_2 FILLER_25_3090 ();
 sg13g2_decap_8 FILLER_25_3120 ();
 sg13g2_decap_8 FILLER_25_3127 ();
 sg13g2_fill_2 FILLER_25_3134 ();
 sg13g2_fill_1 FILLER_25_3136 ();
 sg13g2_fill_2 FILLER_25_3142 ();
 sg13g2_fill_2 FILLER_25_3169 ();
 sg13g2_fill_2 FILLER_25_3192 ();
 sg13g2_fill_1 FILLER_25_3194 ();
 sg13g2_fill_1 FILLER_25_3213 ();
 sg13g2_fill_1 FILLER_25_3231 ();
 sg13g2_fill_1 FILLER_25_3248 ();
 sg13g2_fill_2 FILLER_25_3277 ();
 sg13g2_fill_2 FILLER_25_3299 ();
 sg13g2_decap_4 FILLER_25_3342 ();
 sg13g2_decap_8 FILLER_25_3359 ();
 sg13g2_decap_8 FILLER_25_3366 ();
 sg13g2_decap_8 FILLER_25_3373 ();
 sg13g2_decap_8 FILLER_25_3380 ();
 sg13g2_decap_8 FILLER_25_3387 ();
 sg13g2_decap_8 FILLER_25_3394 ();
 sg13g2_decap_8 FILLER_25_3401 ();
 sg13g2_decap_8 FILLER_25_3408 ();
 sg13g2_decap_8 FILLER_25_3415 ();
 sg13g2_decap_8 FILLER_25_3422 ();
 sg13g2_decap_8 FILLER_25_3429 ();
 sg13g2_decap_8 FILLER_25_3436 ();
 sg13g2_decap_8 FILLER_25_3443 ();
 sg13g2_decap_8 FILLER_25_3450 ();
 sg13g2_decap_8 FILLER_25_3457 ();
 sg13g2_decap_8 FILLER_25_3464 ();
 sg13g2_decap_8 FILLER_25_3471 ();
 sg13g2_decap_8 FILLER_25_3478 ();
 sg13g2_decap_8 FILLER_25_3485 ();
 sg13g2_decap_8 FILLER_25_3492 ();
 sg13g2_decap_8 FILLER_25_3499 ();
 sg13g2_decap_8 FILLER_25_3506 ();
 sg13g2_decap_8 FILLER_25_3513 ();
 sg13g2_decap_8 FILLER_25_3520 ();
 sg13g2_decap_8 FILLER_25_3527 ();
 sg13g2_decap_8 FILLER_25_3534 ();
 sg13g2_decap_8 FILLER_25_3541 ();
 sg13g2_decap_8 FILLER_25_3548 ();
 sg13g2_decap_8 FILLER_25_3555 ();
 sg13g2_decap_8 FILLER_25_3562 ();
 sg13g2_decap_8 FILLER_25_3569 ();
 sg13g2_decap_4 FILLER_25_3576 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_4 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_4 FILLER_26_418 ();
 sg13g2_fill_2 FILLER_26_422 ();
 sg13g2_decap_4 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_26_433 ();
 sg13g2_decap_4 FILLER_26_439 ();
 sg13g2_fill_2 FILLER_26_476 ();
 sg13g2_fill_1 FILLER_26_478 ();
 sg13g2_fill_2 FILLER_26_487 ();
 sg13g2_fill_2 FILLER_26_495 ();
 sg13g2_fill_1 FILLER_26_497 ();
 sg13g2_fill_1 FILLER_26_511 ();
 sg13g2_fill_1 FILLER_26_520 ();
 sg13g2_fill_1 FILLER_26_539 ();
 sg13g2_fill_2 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_578 ();
 sg13g2_fill_2 FILLER_26_597 ();
 sg13g2_decap_4 FILLER_26_632 ();
 sg13g2_fill_2 FILLER_26_636 ();
 sg13g2_fill_2 FILLER_26_651 ();
 sg13g2_fill_1 FILLER_26_675 ();
 sg13g2_decap_4 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_751 ();
 sg13g2_decap_4 FILLER_26_794 ();
 sg13g2_decap_4 FILLER_26_811 ();
 sg13g2_fill_1 FILLER_26_815 ();
 sg13g2_fill_1 FILLER_26_829 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_fill_2 FILLER_26_858 ();
 sg13g2_fill_1 FILLER_26_860 ();
 sg13g2_fill_2 FILLER_26_874 ();
 sg13g2_fill_2 FILLER_26_888 ();
 sg13g2_fill_1 FILLER_26_890 ();
 sg13g2_fill_2 FILLER_26_901 ();
 sg13g2_fill_1 FILLER_26_903 ();
 sg13g2_fill_1 FILLER_26_920 ();
 sg13g2_decap_8 FILLER_26_988 ();
 sg13g2_fill_1 FILLER_26_995 ();
 sg13g2_decap_8 FILLER_26_1009 ();
 sg13g2_decap_8 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1023 ();
 sg13g2_fill_1 FILLER_26_1025 ();
 sg13g2_decap_4 FILLER_26_1031 ();
 sg13g2_fill_1 FILLER_26_1035 ();
 sg13g2_fill_2 FILLER_26_1048 ();
 sg13g2_decap_8 FILLER_26_1063 ();
 sg13g2_decap_8 FILLER_26_1070 ();
 sg13g2_decap_4 FILLER_26_1077 ();
 sg13g2_fill_2 FILLER_26_1081 ();
 sg13g2_decap_4 FILLER_26_1096 ();
 sg13g2_decap_4 FILLER_26_1116 ();
 sg13g2_fill_2 FILLER_26_1134 ();
 sg13g2_fill_1 FILLER_26_1136 ();
 sg13g2_decap_4 FILLER_26_1146 ();
 sg13g2_decap_8 FILLER_26_1166 ();
 sg13g2_decap_4 FILLER_26_1173 ();
 sg13g2_fill_1 FILLER_26_1177 ();
 sg13g2_decap_8 FILLER_26_1182 ();
 sg13g2_decap_8 FILLER_26_1189 ();
 sg13g2_fill_2 FILLER_26_1196 ();
 sg13g2_fill_1 FILLER_26_1198 ();
 sg13g2_decap_8 FILLER_26_1217 ();
 sg13g2_decap_8 FILLER_26_1224 ();
 sg13g2_fill_1 FILLER_26_1231 ();
 sg13g2_decap_8 FILLER_26_1256 ();
 sg13g2_fill_2 FILLER_26_1263 ();
 sg13g2_fill_1 FILLER_26_1265 ();
 sg13g2_fill_2 FILLER_26_1319 ();
 sg13g2_fill_2 FILLER_26_1338 ();
 sg13g2_fill_1 FILLER_26_1340 ();
 sg13g2_decap_4 FILLER_26_1362 ();
 sg13g2_decap_8 FILLER_26_1384 ();
 sg13g2_decap_4 FILLER_26_1391 ();
 sg13g2_fill_2 FILLER_26_1395 ();
 sg13g2_decap_8 FILLER_26_1410 ();
 sg13g2_decap_4 FILLER_26_1417 ();
 sg13g2_fill_1 FILLER_26_1421 ();
 sg13g2_fill_1 FILLER_26_1430 ();
 sg13g2_fill_2 FILLER_26_1445 ();
 sg13g2_fill_1 FILLER_26_1447 ();
 sg13g2_decap_8 FILLER_26_1501 ();
 sg13g2_decap_4 FILLER_26_1523 ();
 sg13g2_fill_1 FILLER_26_1527 ();
 sg13g2_fill_2 FILLER_26_1538 ();
 sg13g2_decap_4 FILLER_26_1545 ();
 sg13g2_fill_1 FILLER_26_1549 ();
 sg13g2_fill_2 FILLER_26_1566 ();
 sg13g2_fill_1 FILLER_26_1568 ();
 sg13g2_decap_4 FILLER_26_1573 ();
 sg13g2_decap_4 FILLER_26_1581 ();
 sg13g2_fill_1 FILLER_26_1585 ();
 sg13g2_fill_2 FILLER_26_1590 ();
 sg13g2_fill_1 FILLER_26_1592 ();
 sg13g2_fill_1 FILLER_26_1606 ();
 sg13g2_fill_2 FILLER_26_1646 ();
 sg13g2_fill_1 FILLER_26_1648 ();
 sg13g2_decap_4 FILLER_26_1666 ();
 sg13g2_fill_2 FILLER_26_1670 ();
 sg13g2_fill_2 FILLER_26_1698 ();
 sg13g2_fill_1 FILLER_26_1700 ();
 sg13g2_fill_1 FILLER_26_1710 ();
 sg13g2_fill_2 FILLER_26_1715 ();
 sg13g2_decap_4 FILLER_26_1748 ();
 sg13g2_fill_1 FILLER_26_1752 ();
 sg13g2_fill_2 FILLER_26_1761 ();
 sg13g2_decap_8 FILLER_26_1767 ();
 sg13g2_decap_8 FILLER_26_1774 ();
 sg13g2_fill_1 FILLER_26_1781 ();
 sg13g2_fill_1 FILLER_26_1790 ();
 sg13g2_fill_2 FILLER_26_1796 ();
 sg13g2_decap_4 FILLER_26_1817 ();
 sg13g2_fill_1 FILLER_26_1821 ();
 sg13g2_decap_8 FILLER_26_1826 ();
 sg13g2_fill_1 FILLER_26_1833 ();
 sg13g2_decap_8 FILLER_26_1849 ();
 sg13g2_fill_2 FILLER_26_1856 ();
 sg13g2_fill_2 FILLER_26_1871 ();
 sg13g2_fill_2 FILLER_26_1913 ();
 sg13g2_decap_8 FILLER_26_1941 ();
 sg13g2_fill_1 FILLER_26_1948 ();
 sg13g2_fill_2 FILLER_26_1999 ();
 sg13g2_fill_1 FILLER_26_2001 ();
 sg13g2_fill_2 FILLER_26_2005 ();
 sg13g2_fill_2 FILLER_26_2035 ();
 sg13g2_fill_1 FILLER_26_2037 ();
 sg13g2_fill_2 FILLER_26_2046 ();
 sg13g2_fill_1 FILLER_26_2048 ();
 sg13g2_decap_8 FILLER_26_2066 ();
 sg13g2_decap_4 FILLER_26_2073 ();
 sg13g2_fill_1 FILLER_26_2077 ();
 sg13g2_fill_1 FILLER_26_2093 ();
 sg13g2_fill_1 FILLER_26_2103 ();
 sg13g2_decap_8 FILLER_26_2136 ();
 sg13g2_decap_4 FILLER_26_2143 ();
 sg13g2_fill_1 FILLER_26_2147 ();
 sg13g2_fill_2 FILLER_26_2194 ();
 sg13g2_decap_4 FILLER_26_2209 ();
 sg13g2_fill_1 FILLER_26_2213 ();
 sg13g2_decap_4 FILLER_26_2242 ();
 sg13g2_fill_1 FILLER_26_2246 ();
 sg13g2_decap_8 FILLER_26_2276 ();
 sg13g2_fill_2 FILLER_26_2283 ();
 sg13g2_fill_2 FILLER_26_2293 ();
 sg13g2_fill_2 FILLER_26_2300 ();
 sg13g2_fill_2 FILLER_26_2310 ();
 sg13g2_decap_8 FILLER_26_2320 ();
 sg13g2_fill_1 FILLER_26_2327 ();
 sg13g2_decap_8 FILLER_26_2338 ();
 sg13g2_decap_8 FILLER_26_2345 ();
 sg13g2_decap_8 FILLER_26_2352 ();
 sg13g2_fill_1 FILLER_26_2359 ();
 sg13g2_decap_8 FILLER_26_2370 ();
 sg13g2_decap_4 FILLER_26_2377 ();
 sg13g2_fill_2 FILLER_26_2399 ();
 sg13g2_decap_4 FILLER_26_2416 ();
 sg13g2_fill_2 FILLER_26_2420 ();
 sg13g2_fill_1 FILLER_26_2442 ();
 sg13g2_decap_8 FILLER_26_2449 ();
 sg13g2_decap_8 FILLER_26_2456 ();
 sg13g2_decap_4 FILLER_26_2463 ();
 sg13g2_fill_1 FILLER_26_2485 ();
 sg13g2_decap_8 FILLER_26_2496 ();
 sg13g2_decap_4 FILLER_26_2503 ();
 sg13g2_decap_8 FILLER_26_2517 ();
 sg13g2_fill_2 FILLER_26_2524 ();
 sg13g2_fill_1 FILLER_26_2526 ();
 sg13g2_decap_8 FILLER_26_2548 ();
 sg13g2_decap_8 FILLER_26_2555 ();
 sg13g2_decap_4 FILLER_26_2562 ();
 sg13g2_fill_2 FILLER_26_2588 ();
 sg13g2_decap_4 FILLER_26_2594 ();
 sg13g2_fill_2 FILLER_26_2598 ();
 sg13g2_fill_1 FILLER_26_2662 ();
 sg13g2_decap_8 FILLER_26_2673 ();
 sg13g2_decap_8 FILLER_26_2704 ();
 sg13g2_decap_4 FILLER_26_2711 ();
 sg13g2_fill_1 FILLER_26_2715 ();
 sg13g2_fill_1 FILLER_26_2721 ();
 sg13g2_fill_2 FILLER_26_2727 ();
 sg13g2_fill_2 FILLER_26_2734 ();
 sg13g2_fill_1 FILLER_26_2736 ();
 sg13g2_fill_2 FILLER_26_2746 ();
 sg13g2_fill_1 FILLER_26_2748 ();
 sg13g2_fill_2 FILLER_26_2777 ();
 sg13g2_fill_1 FILLER_26_2779 ();
 sg13g2_fill_2 FILLER_26_2804 ();
 sg13g2_decap_4 FILLER_26_2810 ();
 sg13g2_fill_1 FILLER_26_2819 ();
 sg13g2_decap_8 FILLER_26_2835 ();
 sg13g2_fill_2 FILLER_26_2842 ();
 sg13g2_fill_2 FILLER_26_2853 ();
 sg13g2_fill_1 FILLER_26_2855 ();
 sg13g2_fill_2 FILLER_26_2878 ();
 sg13g2_fill_1 FILLER_26_2880 ();
 sg13g2_fill_2 FILLER_26_2901 ();
 sg13g2_fill_1 FILLER_26_2903 ();
 sg13g2_fill_1 FILLER_26_2909 ();
 sg13g2_fill_2 FILLER_26_2926 ();
 sg13g2_decap_8 FILLER_26_2961 ();
 sg13g2_decap_8 FILLER_26_2968 ();
 sg13g2_decap_8 FILLER_26_2975 ();
 sg13g2_decap_8 FILLER_26_2995 ();
 sg13g2_decap_4 FILLER_26_3006 ();
 sg13g2_fill_2 FILLER_26_3010 ();
 sg13g2_decap_4 FILLER_26_3026 ();
 sg13g2_fill_2 FILLER_26_3030 ();
 sg13g2_decap_8 FILLER_26_3037 ();
 sg13g2_fill_2 FILLER_26_3051 ();
 sg13g2_fill_1 FILLER_26_3053 ();
 sg13g2_fill_1 FILLER_26_3082 ();
 sg13g2_fill_2 FILLER_26_3096 ();
 sg13g2_decap_4 FILLER_26_3102 ();
 sg13g2_fill_1 FILLER_26_3113 ();
 sg13g2_decap_8 FILLER_26_3124 ();
 sg13g2_decap_4 FILLER_26_3131 ();
 sg13g2_decap_8 FILLER_26_3143 ();
 sg13g2_decap_4 FILLER_26_3162 ();
 sg13g2_fill_2 FILLER_26_3177 ();
 sg13g2_fill_1 FILLER_26_3188 ();
 sg13g2_fill_2 FILLER_26_3229 ();
 sg13g2_fill_2 FILLER_26_3250 ();
 sg13g2_fill_1 FILLER_26_3252 ();
 sg13g2_fill_2 FILLER_26_3294 ();
 sg13g2_fill_1 FILLER_26_3296 ();
 sg13g2_decap_8 FILLER_26_3301 ();
 sg13g2_fill_2 FILLER_26_3308 ();
 sg13g2_fill_1 FILLER_26_3310 ();
 sg13g2_fill_1 FILLER_26_3315 ();
 sg13g2_decap_8 FILLER_26_3366 ();
 sg13g2_decap_8 FILLER_26_3373 ();
 sg13g2_decap_8 FILLER_26_3380 ();
 sg13g2_decap_8 FILLER_26_3387 ();
 sg13g2_decap_8 FILLER_26_3394 ();
 sg13g2_decap_8 FILLER_26_3401 ();
 sg13g2_decap_8 FILLER_26_3408 ();
 sg13g2_decap_8 FILLER_26_3415 ();
 sg13g2_decap_8 FILLER_26_3422 ();
 sg13g2_decap_8 FILLER_26_3429 ();
 sg13g2_decap_8 FILLER_26_3436 ();
 sg13g2_decap_8 FILLER_26_3443 ();
 sg13g2_decap_8 FILLER_26_3450 ();
 sg13g2_decap_8 FILLER_26_3457 ();
 sg13g2_decap_8 FILLER_26_3464 ();
 sg13g2_decap_8 FILLER_26_3471 ();
 sg13g2_decap_8 FILLER_26_3478 ();
 sg13g2_decap_8 FILLER_26_3485 ();
 sg13g2_decap_8 FILLER_26_3492 ();
 sg13g2_decap_8 FILLER_26_3499 ();
 sg13g2_decap_8 FILLER_26_3506 ();
 sg13g2_decap_8 FILLER_26_3513 ();
 sg13g2_decap_8 FILLER_26_3520 ();
 sg13g2_decap_8 FILLER_26_3527 ();
 sg13g2_decap_8 FILLER_26_3534 ();
 sg13g2_decap_8 FILLER_26_3541 ();
 sg13g2_decap_8 FILLER_26_3548 ();
 sg13g2_decap_8 FILLER_26_3555 ();
 sg13g2_decap_8 FILLER_26_3562 ();
 sg13g2_decap_8 FILLER_26_3569 ();
 sg13g2_decap_4 FILLER_26_3576 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_4 FILLER_27_397 ();
 sg13g2_fill_2 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_27_417 ();
 sg13g2_fill_1 FILLER_27_419 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_27_437 ();
 sg13g2_fill_2 FILLER_27_444 ();
 sg13g2_fill_1 FILLER_27_446 ();
 sg13g2_fill_1 FILLER_27_457 ();
 sg13g2_fill_1 FILLER_27_467 ();
 sg13g2_fill_2 FILLER_27_473 ();
 sg13g2_fill_1 FILLER_27_475 ();
 sg13g2_decap_4 FILLER_27_494 ();
 sg13g2_fill_1 FILLER_27_498 ();
 sg13g2_decap_4 FILLER_27_516 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_fill_1 FILLER_27_532 ();
 sg13g2_fill_1 FILLER_27_544 ();
 sg13g2_decap_8 FILLER_27_558 ();
 sg13g2_decap_8 FILLER_27_565 ();
 sg13g2_fill_2 FILLER_27_577 ();
 sg13g2_fill_1 FILLER_27_579 ();
 sg13g2_fill_1 FILLER_27_585 ();
 sg13g2_decap_4 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_4 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_670 ();
 sg13g2_fill_2 FILLER_27_677 ();
 sg13g2_fill_1 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_710 ();
 sg13g2_fill_2 FILLER_27_717 ();
 sg13g2_fill_2 FILLER_27_741 ();
 sg13g2_decap_4 FILLER_27_755 ();
 sg13g2_fill_1 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_780 ();
 sg13g2_fill_2 FILLER_27_787 ();
 sg13g2_fill_1 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_794 ();
 sg13g2_fill_2 FILLER_27_801 ();
 sg13g2_fill_1 FILLER_27_803 ();
 sg13g2_fill_2 FILLER_27_858 ();
 sg13g2_fill_1 FILLER_27_860 ();
 sg13g2_fill_1 FILLER_27_874 ();
 sg13g2_fill_2 FILLER_27_896 ();
 sg13g2_fill_2 FILLER_27_914 ();
 sg13g2_fill_1 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_956 ();
 sg13g2_fill_2 FILLER_27_963 ();
 sg13g2_fill_1 FILLER_27_969 ();
 sg13g2_decap_4 FILLER_27_982 ();
 sg13g2_fill_2 FILLER_27_986 ();
 sg13g2_fill_2 FILLER_27_1001 ();
 sg13g2_fill_1 FILLER_27_1008 ();
 sg13g2_fill_2 FILLER_27_1014 ();
 sg13g2_decap_4 FILLER_27_1031 ();
 sg13g2_fill_1 FILLER_27_1035 ();
 sg13g2_decap_8 FILLER_27_1054 ();
 sg13g2_decap_4 FILLER_27_1061 ();
 sg13g2_fill_1 FILLER_27_1065 ();
 sg13g2_fill_1 FILLER_27_1076 ();
 sg13g2_decap_4 FILLER_27_1082 ();
 sg13g2_fill_2 FILLER_27_1086 ();
 sg13g2_fill_2 FILLER_27_1101 ();
 sg13g2_fill_1 FILLER_27_1103 ();
 sg13g2_fill_2 FILLER_27_1112 ();
 sg13g2_fill_1 FILLER_27_1114 ();
 sg13g2_fill_2 FILLER_27_1132 ();
 sg13g2_decap_4 FILLER_27_1142 ();
 sg13g2_fill_2 FILLER_27_1156 ();
 sg13g2_fill_2 FILLER_27_1171 ();
 sg13g2_fill_1 FILLER_27_1173 ();
 sg13g2_fill_1 FILLER_27_1184 ();
 sg13g2_fill_2 FILLER_27_1194 ();
 sg13g2_fill_1 FILLER_27_1196 ();
 sg13g2_decap_8 FILLER_27_1210 ();
 sg13g2_fill_2 FILLER_27_1217 ();
 sg13g2_fill_1 FILLER_27_1219 ();
 sg13g2_decap_4 FILLER_27_1235 ();
 sg13g2_fill_2 FILLER_27_1239 ();
 sg13g2_fill_2 FILLER_27_1269 ();
 sg13g2_fill_1 FILLER_27_1271 ();
 sg13g2_fill_1 FILLER_27_1309 ();
 sg13g2_fill_2 FILLER_27_1315 ();
 sg13g2_fill_1 FILLER_27_1317 ();
 sg13g2_decap_8 FILLER_27_1339 ();
 sg13g2_fill_1 FILLER_27_1346 ();
 sg13g2_fill_2 FILLER_27_1360 ();
 sg13g2_decap_8 FILLER_27_1381 ();
 sg13g2_decap_4 FILLER_27_1417 ();
 sg13g2_fill_2 FILLER_27_1445 ();
 sg13g2_fill_1 FILLER_27_1472 ();
 sg13g2_decap_8 FILLER_27_1491 ();
 sg13g2_fill_2 FILLER_27_1498 ();
 sg13g2_fill_2 FILLER_27_1523 ();
 sg13g2_fill_1 FILLER_27_1525 ();
 sg13g2_fill_1 FILLER_27_1531 ();
 sg13g2_fill_2 FILLER_27_1536 ();
 sg13g2_fill_2 FILLER_27_1555 ();
 sg13g2_fill_2 FILLER_27_1572 ();
 sg13g2_decap_8 FILLER_27_1586 ();
 sg13g2_decap_4 FILLER_27_1593 ();
 sg13g2_decap_4 FILLER_27_1612 ();
 sg13g2_fill_2 FILLER_27_1616 ();
 sg13g2_fill_2 FILLER_27_1630 ();
 sg13g2_fill_2 FILLER_27_1646 ();
 sg13g2_fill_1 FILLER_27_1648 ();
 sg13g2_decap_8 FILLER_27_1670 ();
 sg13g2_decap_8 FILLER_27_1677 ();
 sg13g2_decap_8 FILLER_27_1711 ();
 sg13g2_fill_2 FILLER_27_1718 ();
 sg13g2_fill_1 FILLER_27_1720 ();
 sg13g2_decap_4 FILLER_27_1729 ();
 sg13g2_fill_2 FILLER_27_1737 ();
 sg13g2_fill_1 FILLER_27_1739 ();
 sg13g2_decap_8 FILLER_27_1774 ();
 sg13g2_decap_4 FILLER_27_1781 ();
 sg13g2_fill_2 FILLER_27_1785 ();
 sg13g2_fill_2 FILLER_27_1807 ();
 sg13g2_decap_8 FILLER_27_1821 ();
 sg13g2_fill_2 FILLER_27_1828 ();
 sg13g2_fill_2 FILLER_27_1847 ();
 sg13g2_fill_2 FILLER_27_1857 ();
 sg13g2_decap_8 FILLER_27_1869 ();
 sg13g2_fill_2 FILLER_27_1876 ();
 sg13g2_fill_2 FILLER_27_1898 ();
 sg13g2_fill_1 FILLER_27_1900 ();
 sg13g2_fill_2 FILLER_27_1917 ();
 sg13g2_fill_2 FILLER_27_1925 ();
 sg13g2_fill_1 FILLER_27_1927 ();
 sg13g2_fill_2 FILLER_27_1934 ();
 sg13g2_fill_1 FILLER_27_1936 ();
 sg13g2_decap_8 FILLER_27_1946 ();
 sg13g2_fill_2 FILLER_27_1953 ();
 sg13g2_decap_8 FILLER_27_1967 ();
 sg13g2_decap_4 FILLER_27_1974 ();
 sg13g2_fill_1 FILLER_27_1978 ();
 sg13g2_decap_8 FILLER_27_1990 ();
 sg13g2_fill_2 FILLER_27_1997 ();
 sg13g2_fill_1 FILLER_27_1999 ();
 sg13g2_fill_2 FILLER_27_2031 ();
 sg13g2_fill_1 FILLER_27_2033 ();
 sg13g2_decap_8 FILLER_27_2056 ();
 sg13g2_decap_4 FILLER_27_2063 ();
 sg13g2_fill_1 FILLER_27_2067 ();
 sg13g2_decap_8 FILLER_27_2117 ();
 sg13g2_decap_8 FILLER_27_2124 ();
 sg13g2_fill_2 FILLER_27_2131 ();
 sg13g2_decap_8 FILLER_27_2146 ();
 sg13g2_decap_8 FILLER_27_2179 ();
 sg13g2_fill_2 FILLER_27_2186 ();
 sg13g2_decap_8 FILLER_27_2209 ();
 sg13g2_decap_4 FILLER_27_2216 ();
 sg13g2_decap_4 FILLER_27_2224 ();
 sg13g2_fill_1 FILLER_27_2228 ();
 sg13g2_decap_8 FILLER_27_2249 ();
 sg13g2_fill_1 FILLER_27_2256 ();
 sg13g2_decap_8 FILLER_27_2276 ();
 sg13g2_decap_8 FILLER_27_2283 ();
 sg13g2_decap_4 FILLER_27_2290 ();
 sg13g2_fill_2 FILLER_27_2309 ();
 sg13g2_fill_1 FILLER_27_2311 ();
 sg13g2_decap_8 FILLER_27_2332 ();
 sg13g2_fill_2 FILLER_27_2383 ();
 sg13g2_fill_2 FILLER_27_2402 ();
 sg13g2_fill_1 FILLER_27_2404 ();
 sg13g2_decap_8 FILLER_27_2410 ();
 sg13g2_decap_8 FILLER_27_2417 ();
 sg13g2_decap_8 FILLER_27_2424 ();
 sg13g2_fill_2 FILLER_27_2431 ();
 sg13g2_fill_1 FILLER_27_2442 ();
 sg13g2_decap_8 FILLER_27_2452 ();
 sg13g2_decap_8 FILLER_27_2459 ();
 sg13g2_fill_2 FILLER_27_2466 ();
 sg13g2_fill_1 FILLER_27_2468 ();
 sg13g2_decap_4 FILLER_27_2479 ();
 sg13g2_fill_2 FILLER_27_2516 ();
 sg13g2_decap_8 FILLER_27_2526 ();
 sg13g2_decap_8 FILLER_27_2542 ();
 sg13g2_fill_2 FILLER_27_2549 ();
 sg13g2_fill_1 FILLER_27_2551 ();
 sg13g2_fill_2 FILLER_27_2565 ();
 sg13g2_decap_8 FILLER_27_2593 ();
 sg13g2_decap_8 FILLER_27_2600 ();
 sg13g2_decap_4 FILLER_27_2607 ();
 sg13g2_decap_4 FILLER_27_2624 ();
 sg13g2_decap_8 FILLER_27_2641 ();
 sg13g2_decap_4 FILLER_27_2648 ();
 sg13g2_fill_2 FILLER_27_2657 ();
 sg13g2_fill_1 FILLER_27_2659 ();
 sg13g2_fill_2 FILLER_27_2665 ();
 sg13g2_fill_1 FILLER_27_2667 ();
 sg13g2_fill_2 FILLER_27_2691 ();
 sg13g2_fill_1 FILLER_27_2706 ();
 sg13g2_decap_8 FILLER_27_2731 ();
 sg13g2_decap_8 FILLER_27_2738 ();
 sg13g2_fill_1 FILLER_27_2771 ();
 sg13g2_fill_2 FILLER_27_2785 ();
 sg13g2_decap_4 FILLER_27_2815 ();
 sg13g2_fill_2 FILLER_27_2819 ();
 sg13g2_decap_8 FILLER_27_2852 ();
 sg13g2_decap_8 FILLER_27_2868 ();
 sg13g2_fill_1 FILLER_27_2875 ();
 sg13g2_fill_2 FILLER_27_2888 ();
 sg13g2_fill_1 FILLER_27_2890 ();
 sg13g2_decap_4 FILLER_27_2904 ();
 sg13g2_decap_8 FILLER_27_2922 ();
 sg13g2_decap_4 FILLER_27_2929 ();
 sg13g2_fill_2 FILLER_27_2933 ();
 sg13g2_fill_2 FILLER_27_2940 ();
 sg13g2_fill_1 FILLER_27_2942 ();
 sg13g2_fill_2 FILLER_27_2961 ();
 sg13g2_fill_1 FILLER_27_2963 ();
 sg13g2_decap_4 FILLER_27_2969 ();
 sg13g2_fill_2 FILLER_27_2983 ();
 sg13g2_fill_2 FILLER_27_2991 ();
 sg13g2_fill_1 FILLER_27_2993 ();
 sg13g2_fill_2 FILLER_27_3010 ();
 sg13g2_fill_2 FILLER_27_3025 ();
 sg13g2_fill_2 FILLER_27_3040 ();
 sg13g2_decap_4 FILLER_27_3095 ();
 sg13g2_fill_2 FILLER_27_3132 ();
 sg13g2_decap_4 FILLER_27_3157 ();
 sg13g2_fill_2 FILLER_27_3161 ();
 sg13g2_fill_1 FILLER_27_3187 ();
 sg13g2_fill_2 FILLER_27_3193 ();
 sg13g2_decap_8 FILLER_27_3240 ();
 sg13g2_decap_4 FILLER_27_3247 ();
 sg13g2_fill_2 FILLER_27_3251 ();
 sg13g2_fill_2 FILLER_27_3279 ();
 sg13g2_fill_2 FILLER_27_3286 ();
 sg13g2_decap_4 FILLER_27_3337 ();
 sg13g2_fill_2 FILLER_27_3341 ();
 sg13g2_decap_8 FILLER_27_3347 ();
 sg13g2_decap_8 FILLER_27_3354 ();
 sg13g2_decap_8 FILLER_27_3361 ();
 sg13g2_decap_8 FILLER_27_3368 ();
 sg13g2_decap_8 FILLER_27_3375 ();
 sg13g2_decap_8 FILLER_27_3382 ();
 sg13g2_decap_8 FILLER_27_3389 ();
 sg13g2_decap_8 FILLER_27_3396 ();
 sg13g2_decap_8 FILLER_27_3403 ();
 sg13g2_decap_8 FILLER_27_3410 ();
 sg13g2_decap_8 FILLER_27_3417 ();
 sg13g2_decap_8 FILLER_27_3424 ();
 sg13g2_decap_8 FILLER_27_3431 ();
 sg13g2_decap_8 FILLER_27_3438 ();
 sg13g2_decap_8 FILLER_27_3445 ();
 sg13g2_decap_8 FILLER_27_3452 ();
 sg13g2_decap_8 FILLER_27_3459 ();
 sg13g2_decap_8 FILLER_27_3466 ();
 sg13g2_decap_8 FILLER_27_3473 ();
 sg13g2_decap_8 FILLER_27_3480 ();
 sg13g2_decap_8 FILLER_27_3487 ();
 sg13g2_decap_8 FILLER_27_3494 ();
 sg13g2_decap_8 FILLER_27_3501 ();
 sg13g2_decap_8 FILLER_27_3508 ();
 sg13g2_decap_8 FILLER_27_3515 ();
 sg13g2_decap_8 FILLER_27_3522 ();
 sg13g2_decap_8 FILLER_27_3529 ();
 sg13g2_decap_8 FILLER_27_3536 ();
 sg13g2_decap_8 FILLER_27_3543 ();
 sg13g2_decap_8 FILLER_27_3550 ();
 sg13g2_decap_8 FILLER_27_3557 ();
 sg13g2_decap_8 FILLER_27_3564 ();
 sg13g2_decap_8 FILLER_27_3571 ();
 sg13g2_fill_2 FILLER_27_3578 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_4 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_4 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_396 ();
 sg13g2_fill_2 FILLER_28_462 ();
 sg13g2_fill_1 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_530 ();
 sg13g2_fill_2 FILLER_28_568 ();
 sg13g2_fill_1 FILLER_28_570 ();
 sg13g2_fill_2 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_fill_1 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_fill_2 FILLER_28_634 ();
 sg13g2_fill_2 FILLER_28_640 ();
 sg13g2_fill_1 FILLER_28_651 ();
 sg13g2_fill_2 FILLER_28_665 ();
 sg13g2_fill_1 FILLER_28_667 ();
 sg13g2_decap_8 FILLER_28_688 ();
 sg13g2_decap_4 FILLER_28_695 ();
 sg13g2_fill_2 FILLER_28_709 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_fill_2 FILLER_28_722 ();
 sg13g2_decap_4 FILLER_28_756 ();
 sg13g2_fill_2 FILLER_28_760 ();
 sg13g2_fill_2 FILLER_28_775 ();
 sg13g2_fill_1 FILLER_28_777 ();
 sg13g2_fill_2 FILLER_28_783 ();
 sg13g2_fill_1 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_fill_2 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_fill_2 FILLER_28_876 ();
 sg13g2_fill_2 FILLER_28_883 ();
 sg13g2_decap_8 FILLER_28_896 ();
 sg13g2_decap_8 FILLER_28_903 ();
 sg13g2_fill_2 FILLER_28_910 ();
 sg13g2_fill_1 FILLER_28_912 ();
 sg13g2_decap_4 FILLER_28_922 ();
 sg13g2_decap_8 FILLER_28_931 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_949 ();
 sg13g2_decap_4 FILLER_28_956 ();
 sg13g2_fill_2 FILLER_28_988 ();
 sg13g2_fill_1 FILLER_28_990 ();
 sg13g2_fill_2 FILLER_28_996 ();
 sg13g2_fill_1 FILLER_28_998 ();
 sg13g2_decap_4 FILLER_28_1012 ();
 sg13g2_fill_2 FILLER_28_1029 ();
 sg13g2_fill_2 FILLER_28_1039 ();
 sg13g2_decap_8 FILLER_28_1050 ();
 sg13g2_decap_4 FILLER_28_1057 ();
 sg13g2_fill_2 FILLER_28_1061 ();
 sg13g2_decap_8 FILLER_28_1083 ();
 sg13g2_fill_1 FILLER_28_1090 ();
 sg13g2_decap_4 FILLER_28_1112 ();
 sg13g2_fill_1 FILLER_28_1116 ();
 sg13g2_decap_4 FILLER_28_1135 ();
 sg13g2_fill_1 FILLER_28_1139 ();
 sg13g2_decap_4 FILLER_28_1160 ();
 sg13g2_fill_1 FILLER_28_1164 ();
 sg13g2_fill_2 FILLER_28_1170 ();
 sg13g2_fill_2 FILLER_28_1177 ();
 sg13g2_decap_8 FILLER_28_1191 ();
 sg13g2_fill_2 FILLER_28_1198 ();
 sg13g2_fill_1 FILLER_28_1200 ();
 sg13g2_decap_8 FILLER_28_1234 ();
 sg13g2_decap_8 FILLER_28_1252 ();
 sg13g2_decap_8 FILLER_28_1268 ();
 sg13g2_fill_2 FILLER_28_1275 ();
 sg13g2_fill_1 FILLER_28_1277 ();
 sg13g2_decap_8 FILLER_28_1282 ();
 sg13g2_decap_8 FILLER_28_1289 ();
 sg13g2_fill_1 FILLER_28_1296 ();
 sg13g2_fill_1 FILLER_28_1305 ();
 sg13g2_decap_8 FILLER_28_1311 ();
 sg13g2_fill_2 FILLER_28_1318 ();
 sg13g2_fill_1 FILLER_28_1320 ();
 sg13g2_decap_8 FILLER_28_1335 ();
 sg13g2_decap_8 FILLER_28_1342 ();
 sg13g2_fill_1 FILLER_28_1349 ();
 sg13g2_fill_2 FILLER_28_1355 ();
 sg13g2_fill_1 FILLER_28_1357 ();
 sg13g2_fill_1 FILLER_28_1368 ();
 sg13g2_decap_8 FILLER_28_1377 ();
 sg13g2_decap_4 FILLER_28_1384 ();
 sg13g2_fill_1 FILLER_28_1388 ();
 sg13g2_decap_8 FILLER_28_1413 ();
 sg13g2_decap_8 FILLER_28_1420 ();
 sg13g2_fill_2 FILLER_28_1427 ();
 sg13g2_fill_1 FILLER_28_1429 ();
 sg13g2_decap_4 FILLER_28_1440 ();
 sg13g2_fill_1 FILLER_28_1444 ();
 sg13g2_decap_4 FILLER_28_1462 ();
 sg13g2_decap_4 FILLER_28_1505 ();
 sg13g2_fill_2 FILLER_28_1509 ();
 sg13g2_fill_2 FILLER_28_1521 ();
 sg13g2_fill_2 FILLER_28_1531 ();
 sg13g2_fill_1 FILLER_28_1533 ();
 sg13g2_fill_2 FILLER_28_1544 ();
 sg13g2_fill_1 FILLER_28_1546 ();
 sg13g2_decap_8 FILLER_28_1555 ();
 sg13g2_fill_2 FILLER_28_1562 ();
 sg13g2_fill_1 FILLER_28_1564 ();
 sg13g2_decap_4 FILLER_28_1577 ();
 sg13g2_fill_2 FILLER_28_1589 ();
 sg13g2_decap_8 FILLER_28_1612 ();
 sg13g2_fill_2 FILLER_28_1619 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_4 FILLER_28_1638 ();
 sg13g2_fill_2 FILLER_28_1642 ();
 sg13g2_decap_8 FILLER_28_1669 ();
 sg13g2_fill_1 FILLER_28_1676 ();
 sg13g2_fill_2 FILLER_28_1701 ();
 sg13g2_fill_1 FILLER_28_1703 ();
 sg13g2_fill_1 FILLER_28_1712 ();
 sg13g2_fill_2 FILLER_28_1721 ();
 sg13g2_fill_1 FILLER_28_1723 ();
 sg13g2_fill_1 FILLER_28_1743 ();
 sg13g2_fill_1 FILLER_28_1759 ();
 sg13g2_decap_8 FILLER_28_1764 ();
 sg13g2_fill_2 FILLER_28_1807 ();
 sg13g2_fill_1 FILLER_28_1809 ();
 sg13g2_fill_1 FILLER_28_1816 ();
 sg13g2_fill_2 FILLER_28_1821 ();
 sg13g2_fill_2 FILLER_28_1843 ();
 sg13g2_decap_4 FILLER_28_1868 ();
 sg13g2_decap_8 FILLER_28_1875 ();
 sg13g2_fill_2 FILLER_28_1882 ();
 sg13g2_fill_1 FILLER_28_1884 ();
 sg13g2_decap_8 FILLER_28_1892 ();
 sg13g2_decap_8 FILLER_28_1899 ();
 sg13g2_fill_2 FILLER_28_1913 ();
 sg13g2_fill_1 FILLER_28_1933 ();
 sg13g2_decap_8 FILLER_28_1965 ();
 sg13g2_decap_8 FILLER_28_1972 ();
 sg13g2_decap_8 FILLER_28_1979 ();
 sg13g2_decap_4 FILLER_28_1986 ();
 sg13g2_fill_2 FILLER_28_1990 ();
 sg13g2_decap_8 FILLER_28_1997 ();
 sg13g2_decap_4 FILLER_28_2004 ();
 sg13g2_fill_1 FILLER_28_2008 ();
 sg13g2_decap_4 FILLER_28_2013 ();
 sg13g2_fill_1 FILLER_28_2017 ();
 sg13g2_decap_4 FILLER_28_2027 ();
 sg13g2_fill_2 FILLER_28_2047 ();
 sg13g2_decap_4 FILLER_28_2076 ();
 sg13g2_fill_1 FILLER_28_2092 ();
 sg13g2_fill_2 FILLER_28_2106 ();
 sg13g2_fill_1 FILLER_28_2108 ();
 sg13g2_decap_4 FILLER_28_2113 ();
 sg13g2_fill_1 FILLER_28_2126 ();
 sg13g2_decap_4 FILLER_28_2140 ();
 sg13g2_fill_2 FILLER_28_2165 ();
 sg13g2_fill_1 FILLER_28_2167 ();
 sg13g2_decap_4 FILLER_28_2173 ();
 sg13g2_fill_1 FILLER_28_2177 ();
 sg13g2_fill_2 FILLER_28_2182 ();
 sg13g2_fill_2 FILLER_28_2203 ();
 sg13g2_decap_8 FILLER_28_2214 ();
 sg13g2_fill_2 FILLER_28_2221 ();
 sg13g2_decap_8 FILLER_28_2227 ();
 sg13g2_decap_8 FILLER_28_2250 ();
 sg13g2_decap_8 FILLER_28_2257 ();
 sg13g2_decap_4 FILLER_28_2264 ();
 sg13g2_fill_1 FILLER_28_2268 ();
 sg13g2_decap_8 FILLER_28_2274 ();
 sg13g2_decap_8 FILLER_28_2281 ();
 sg13g2_decap_8 FILLER_28_2292 ();
 sg13g2_decap_8 FILLER_28_2304 ();
 sg13g2_fill_1 FILLER_28_2311 ();
 sg13g2_decap_8 FILLER_28_2317 ();
 sg13g2_fill_1 FILLER_28_2324 ();
 sg13g2_decap_8 FILLER_28_2330 ();
 sg13g2_decap_4 FILLER_28_2337 ();
 sg13g2_decap_4 FILLER_28_2349 ();
 sg13g2_fill_1 FILLER_28_2353 ();
 sg13g2_decap_4 FILLER_28_2364 ();
 sg13g2_decap_4 FILLER_28_2383 ();
 sg13g2_fill_2 FILLER_28_2387 ();
 sg13g2_fill_1 FILLER_28_2408 ();
 sg13g2_fill_1 FILLER_28_2421 ();
 sg13g2_decap_4 FILLER_28_2426 ();
 sg13g2_fill_1 FILLER_28_2435 ();
 sg13g2_decap_8 FILLER_28_2446 ();
 sg13g2_fill_2 FILLER_28_2453 ();
 sg13g2_fill_1 FILLER_28_2455 ();
 sg13g2_fill_2 FILLER_28_2469 ();
 sg13g2_fill_1 FILLER_28_2471 ();
 sg13g2_decap_4 FILLER_28_2488 ();
 sg13g2_decap_4 FILLER_28_2500 ();
 sg13g2_fill_2 FILLER_28_2504 ();
 sg13g2_decap_4 FILLER_28_2544 ();
 sg13g2_fill_2 FILLER_28_2565 ();
 sg13g2_decap_8 FILLER_28_2588 ();
 sg13g2_decap_8 FILLER_28_2595 ();
 sg13g2_fill_2 FILLER_28_2602 ();
 sg13g2_fill_1 FILLER_28_2604 ();
 sg13g2_decap_8 FILLER_28_2622 ();
 sg13g2_fill_2 FILLER_28_2629 ();
 sg13g2_fill_1 FILLER_28_2652 ();
 sg13g2_decap_4 FILLER_28_2700 ();
 sg13g2_fill_1 FILLER_28_2704 ();
 sg13g2_fill_1 FILLER_28_2709 ();
 sg13g2_decap_8 FILLER_28_2734 ();
 sg13g2_decap_4 FILLER_28_2741 ();
 sg13g2_fill_2 FILLER_28_2745 ();
 sg13g2_decap_8 FILLER_28_2760 ();
 sg13g2_fill_2 FILLER_28_2767 ();
 sg13g2_fill_1 FILLER_28_2800 ();
 sg13g2_decap_8 FILLER_28_2833 ();
 sg13g2_decap_4 FILLER_28_2840 ();
 sg13g2_fill_1 FILLER_28_2844 ();
 sg13g2_decap_4 FILLER_28_2849 ();
 sg13g2_fill_1 FILLER_28_2853 ();
 sg13g2_decap_4 FILLER_28_2867 ();
 sg13g2_decap_8 FILLER_28_2897 ();
 sg13g2_fill_2 FILLER_28_2904 ();
 sg13g2_decap_8 FILLER_28_2922 ();
 sg13g2_fill_2 FILLER_28_2929 ();
 sg13g2_fill_1 FILLER_28_2931 ();
 sg13g2_decap_8 FILLER_28_2950 ();
 sg13g2_fill_2 FILLER_28_2977 ();
 sg13g2_fill_1 FILLER_28_2979 ();
 sg13g2_decap_8 FILLER_28_2990 ();
 sg13g2_decap_4 FILLER_28_2997 ();
 sg13g2_fill_1 FILLER_28_3009 ();
 sg13g2_decap_4 FILLER_28_3027 ();
 sg13g2_fill_1 FILLER_28_3031 ();
 sg13g2_decap_8 FILLER_28_3050 ();
 sg13g2_decap_8 FILLER_28_3057 ();
 sg13g2_decap_4 FILLER_28_3064 ();
 sg13g2_fill_2 FILLER_28_3096 ();
 sg13g2_decap_8 FILLER_28_3129 ();
 sg13g2_decap_8 FILLER_28_3136 ();
 sg13g2_fill_2 FILLER_28_3154 ();
 sg13g2_fill_1 FILLER_28_3156 ();
 sg13g2_fill_2 FILLER_28_3192 ();
 sg13g2_decap_4 FILLER_28_3198 ();
 sg13g2_fill_1 FILLER_28_3202 ();
 sg13g2_decap_4 FILLER_28_3212 ();
 sg13g2_fill_1 FILLER_28_3216 ();
 sg13g2_fill_2 FILLER_28_3231 ();
 sg13g2_fill_2 FILLER_28_3237 ();
 sg13g2_fill_2 FILLER_28_3261 ();
 sg13g2_fill_1 FILLER_28_3263 ();
 sg13g2_fill_1 FILLER_28_3317 ();
 sg13g2_fill_2 FILLER_28_3331 ();
 sg13g2_decap_8 FILLER_28_3346 ();
 sg13g2_decap_8 FILLER_28_3353 ();
 sg13g2_decap_8 FILLER_28_3360 ();
 sg13g2_decap_8 FILLER_28_3367 ();
 sg13g2_decap_8 FILLER_28_3374 ();
 sg13g2_decap_8 FILLER_28_3381 ();
 sg13g2_decap_8 FILLER_28_3388 ();
 sg13g2_decap_8 FILLER_28_3395 ();
 sg13g2_decap_8 FILLER_28_3402 ();
 sg13g2_decap_8 FILLER_28_3409 ();
 sg13g2_decap_8 FILLER_28_3416 ();
 sg13g2_decap_8 FILLER_28_3423 ();
 sg13g2_decap_8 FILLER_28_3430 ();
 sg13g2_decap_8 FILLER_28_3437 ();
 sg13g2_decap_8 FILLER_28_3444 ();
 sg13g2_decap_8 FILLER_28_3451 ();
 sg13g2_decap_8 FILLER_28_3458 ();
 sg13g2_decap_8 FILLER_28_3465 ();
 sg13g2_decap_8 FILLER_28_3472 ();
 sg13g2_decap_8 FILLER_28_3479 ();
 sg13g2_decap_8 FILLER_28_3486 ();
 sg13g2_decap_8 FILLER_28_3493 ();
 sg13g2_decap_8 FILLER_28_3500 ();
 sg13g2_decap_8 FILLER_28_3507 ();
 sg13g2_decap_8 FILLER_28_3514 ();
 sg13g2_decap_8 FILLER_28_3521 ();
 sg13g2_decap_8 FILLER_28_3528 ();
 sg13g2_decap_8 FILLER_28_3535 ();
 sg13g2_decap_8 FILLER_28_3542 ();
 sg13g2_decap_8 FILLER_28_3549 ();
 sg13g2_decap_8 FILLER_28_3556 ();
 sg13g2_decap_8 FILLER_28_3563 ();
 sg13g2_decap_8 FILLER_28_3570 ();
 sg13g2_fill_2 FILLER_28_3577 ();
 sg13g2_fill_1 FILLER_28_3579 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_2 FILLER_29_421 ();
 sg13g2_decap_4 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_29_437 ();
 sg13g2_decap_4 FILLER_29_444 ();
 sg13g2_fill_1 FILLER_29_467 ();
 sg13g2_fill_1 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_fill_2 FILLER_29_504 ();
 sg13g2_fill_1 FILLER_29_506 ();
 sg13g2_decap_4 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_526 ();
 sg13g2_fill_2 FILLER_29_533 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_fill_2 FILLER_29_546 ();
 sg13g2_decap_4 FILLER_29_552 ();
 sg13g2_fill_1 FILLER_29_556 ();
 sg13g2_decap_4 FILLER_29_598 ();
 sg13g2_fill_1 FILLER_29_602 ();
 sg13g2_fill_2 FILLER_29_659 ();
 sg13g2_fill_2 FILLER_29_685 ();
 sg13g2_decap_4 FILLER_29_700 ();
 sg13g2_fill_2 FILLER_29_704 ();
 sg13g2_fill_1 FILLER_29_734 ();
 sg13g2_decap_4 FILLER_29_739 ();
 sg13g2_fill_2 FILLER_29_756 ();
 sg13g2_fill_1 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_2 FILLER_29_861 ();
 sg13g2_fill_1 FILLER_29_863 ();
 sg13g2_fill_2 FILLER_29_876 ();
 sg13g2_fill_1 FILLER_29_878 ();
 sg13g2_decap_4 FILLER_29_908 ();
 sg13g2_fill_1 FILLER_29_912 ();
 sg13g2_decap_4 FILLER_29_917 ();
 sg13g2_fill_1 FILLER_29_921 ();
 sg13g2_fill_1 FILLER_29_926 ();
 sg13g2_decap_4 FILLER_29_961 ();
 sg13g2_fill_2 FILLER_29_965 ();
 sg13g2_decap_4 FILLER_29_974 ();
 sg13g2_fill_1 FILLER_29_978 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_fill_1 FILLER_29_1011 ();
 sg13g2_fill_2 FILLER_29_1017 ();
 sg13g2_fill_1 FILLER_29_1019 ();
 sg13g2_decap_8 FILLER_29_1029 ();
 sg13g2_fill_2 FILLER_29_1044 ();
 sg13g2_decap_8 FILLER_29_1056 ();
 sg13g2_decap_8 FILLER_29_1063 ();
 sg13g2_decap_8 FILLER_29_1075 ();
 sg13g2_decap_4 FILLER_29_1082 ();
 sg13g2_fill_1 FILLER_29_1086 ();
 sg13g2_decap_4 FILLER_29_1114 ();
 sg13g2_fill_1 FILLER_29_1118 ();
 sg13g2_decap_4 FILLER_29_1137 ();
 sg13g2_fill_1 FILLER_29_1141 ();
 sg13g2_decap_8 FILLER_29_1166 ();
 sg13g2_fill_2 FILLER_29_1173 ();
 sg13g2_fill_1 FILLER_29_1175 ();
 sg13g2_fill_2 FILLER_29_1184 ();
 sg13g2_fill_1 FILLER_29_1186 ();
 sg13g2_decap_4 FILLER_29_1192 ();
 sg13g2_fill_1 FILLER_29_1196 ();
 sg13g2_decap_4 FILLER_29_1212 ();
 sg13g2_fill_1 FILLER_29_1216 ();
 sg13g2_decap_4 FILLER_29_1247 ();
 sg13g2_decap_8 FILLER_29_1272 ();
 sg13g2_decap_8 FILLER_29_1279 ();
 sg13g2_decap_4 FILLER_29_1286 ();
 sg13g2_fill_2 FILLER_29_1290 ();
 sg13g2_fill_2 FILLER_29_1319 ();
 sg13g2_decap_4 FILLER_29_1341 ();
 sg13g2_fill_2 FILLER_29_1345 ();
 sg13g2_fill_1 FILLER_29_1354 ();
 sg13g2_decap_8 FILLER_29_1376 ();
 sg13g2_fill_2 FILLER_29_1383 ();
 sg13g2_fill_1 FILLER_29_1385 ();
 sg13g2_fill_2 FILLER_29_1400 ();
 sg13g2_fill_1 FILLER_29_1402 ();
 sg13g2_decap_4 FILLER_29_1419 ();
 sg13g2_fill_1 FILLER_29_1423 ();
 sg13g2_decap_8 FILLER_29_1467 ();
 sg13g2_decap_8 FILLER_29_1489 ();
 sg13g2_decap_8 FILLER_29_1496 ();
 sg13g2_fill_2 FILLER_29_1503 ();
 sg13g2_fill_2 FILLER_29_1529 ();
 sg13g2_decap_8 FILLER_29_1539 ();
 sg13g2_fill_1 FILLER_29_1546 ();
 sg13g2_decap_8 FILLER_29_1575 ();
 sg13g2_decap_4 FILLER_29_1582 ();
 sg13g2_fill_2 FILLER_29_1586 ();
 sg13g2_fill_1 FILLER_29_1601 ();
 sg13g2_decap_4 FILLER_29_1610 ();
 sg13g2_fill_2 FILLER_29_1623 ();
 sg13g2_decap_8 FILLER_29_1640 ();
 sg13g2_fill_2 FILLER_29_1647 ();
 sg13g2_decap_8 FILLER_29_1663 ();
 sg13g2_fill_2 FILLER_29_1683 ();
 sg13g2_fill_1 FILLER_29_1716 ();
 sg13g2_fill_2 FILLER_29_1732 ();
 sg13g2_fill_1 FILLER_29_1734 ();
 sg13g2_decap_4 FILLER_29_1765 ();
 sg13g2_fill_2 FILLER_29_1769 ();
 sg13g2_fill_2 FILLER_29_1803 ();
 sg13g2_fill_2 FILLER_29_1818 ();
 sg13g2_fill_1 FILLER_29_1824 ();
 sg13g2_decap_4 FILLER_29_1838 ();
 sg13g2_fill_2 FILLER_29_1842 ();
 sg13g2_fill_2 FILLER_29_1853 ();
 sg13g2_decap_4 FILLER_29_1861 ();
 sg13g2_fill_2 FILLER_29_1865 ();
 sg13g2_fill_2 FILLER_29_1901 ();
 sg13g2_fill_1 FILLER_29_1903 ();
 sg13g2_fill_1 FILLER_29_1941 ();
 sg13g2_fill_2 FILLER_29_1949 ();
 sg13g2_fill_1 FILLER_29_1951 ();
 sg13g2_fill_1 FILLER_29_1962 ();
 sg13g2_decap_8 FILLER_29_1972 ();
 sg13g2_fill_2 FILLER_29_1979 ();
 sg13g2_fill_1 FILLER_29_1981 ();
 sg13g2_fill_1 FILLER_29_2005 ();
 sg13g2_decap_8 FILLER_29_2017 ();
 sg13g2_fill_2 FILLER_29_2024 ();
 sg13g2_fill_2 FILLER_29_2052 ();
 sg13g2_decap_4 FILLER_29_2058 ();
 sg13g2_fill_1 FILLER_29_2062 ();
 sg13g2_fill_2 FILLER_29_2103 ();
 sg13g2_fill_1 FILLER_29_2105 ();
 sg13g2_fill_1 FILLER_29_2119 ();
 sg13g2_fill_1 FILLER_29_2133 ();
 sg13g2_decap_4 FILLER_29_2139 ();
 sg13g2_decap_8 FILLER_29_2147 ();
 sg13g2_fill_1 FILLER_29_2154 ();
 sg13g2_decap_8 FILLER_29_2176 ();
 sg13g2_decap_8 FILLER_29_2183 ();
 sg13g2_fill_1 FILLER_29_2190 ();
 sg13g2_fill_1 FILLER_29_2200 ();
 sg13g2_decap_4 FILLER_29_2225 ();
 sg13g2_fill_1 FILLER_29_2229 ();
 sg13g2_fill_2 FILLER_29_2247 ();
 sg13g2_fill_1 FILLER_29_2249 ();
 sg13g2_decap_4 FILLER_29_2278 ();
 sg13g2_fill_1 FILLER_29_2282 ();
 sg13g2_decap_4 FILLER_29_2288 ();
 sg13g2_fill_2 FILLER_29_2296 ();
 sg13g2_fill_1 FILLER_29_2298 ();
 sg13g2_fill_1 FILLER_29_2308 ();
 sg13g2_decap_4 FILLER_29_2314 ();
 sg13g2_fill_2 FILLER_29_2324 ();
 sg13g2_fill_1 FILLER_29_2326 ();
 sg13g2_fill_1 FILLER_29_2340 ();
 sg13g2_decap_8 FILLER_29_2350 ();
 sg13g2_decap_8 FILLER_29_2357 ();
 sg13g2_decap_8 FILLER_29_2364 ();
 sg13g2_decap_8 FILLER_29_2371 ();
 sg13g2_fill_2 FILLER_29_2378 ();
 sg13g2_fill_1 FILLER_29_2380 ();
 sg13g2_decap_4 FILLER_29_2389 ();
 sg13g2_fill_1 FILLER_29_2393 ();
 sg13g2_fill_2 FILLER_29_2416 ();
 sg13g2_decap_4 FILLER_29_2432 ();
 sg13g2_fill_2 FILLER_29_2439 ();
 sg13g2_fill_1 FILLER_29_2441 ();
 sg13g2_decap_4 FILLER_29_2455 ();
 sg13g2_decap_4 FILLER_29_2464 ();
 sg13g2_fill_1 FILLER_29_2468 ();
 sg13g2_fill_2 FILLER_29_2473 ();
 sg13g2_fill_2 FILLER_29_2479 ();
 sg13g2_fill_1 FILLER_29_2481 ();
 sg13g2_fill_2 FILLER_29_2486 ();
 sg13g2_fill_1 FILLER_29_2488 ();
 sg13g2_decap_8 FILLER_29_2494 ();
 sg13g2_decap_8 FILLER_29_2501 ();
 sg13g2_fill_2 FILLER_29_2508 ();
 sg13g2_decap_4 FILLER_29_2526 ();
 sg13g2_fill_2 FILLER_29_2546 ();
 sg13g2_fill_1 FILLER_29_2548 ();
 sg13g2_decap_8 FILLER_29_2561 ();
 sg13g2_decap_8 FILLER_29_2568 ();
 sg13g2_decap_8 FILLER_29_2583 ();
 sg13g2_decap_8 FILLER_29_2590 ();
 sg13g2_decap_8 FILLER_29_2597 ();
 sg13g2_fill_1 FILLER_29_2604 ();
 sg13g2_fill_1 FILLER_29_2631 ();
 sg13g2_decap_4 FILLER_29_2645 ();
 sg13g2_decap_8 FILLER_29_2659 ();
 sg13g2_decap_8 FILLER_29_2666 ();
 sg13g2_decap_8 FILLER_29_2673 ();
 sg13g2_decap_8 FILLER_29_2680 ();
 sg13g2_fill_2 FILLER_29_2687 ();
 sg13g2_fill_2 FILLER_29_2705 ();
 sg13g2_fill_1 FILLER_29_2707 ();
 sg13g2_decap_4 FILLER_29_2712 ();
 sg13g2_fill_1 FILLER_29_2733 ();
 sg13g2_decap_4 FILLER_29_2779 ();
 sg13g2_decap_4 FILLER_29_2787 ();
 sg13g2_decap_8 FILLER_29_2800 ();
 sg13g2_decap_4 FILLER_29_2835 ();
 sg13g2_fill_2 FILLER_29_2839 ();
 sg13g2_fill_2 FILLER_29_2847 ();
 sg13g2_fill_1 FILLER_29_2853 ();
 sg13g2_fill_2 FILLER_29_2874 ();
 sg13g2_fill_1 FILLER_29_2876 ();
 sg13g2_decap_8 FILLER_29_2889 ();
 sg13g2_decap_4 FILLER_29_2896 ();
 sg13g2_fill_1 FILLER_29_2900 ();
 sg13g2_decap_8 FILLER_29_2907 ();
 sg13g2_decap_8 FILLER_29_2914 ();
 sg13g2_fill_2 FILLER_29_2921 ();
 sg13g2_decap_4 FILLER_29_2931 ();
 sg13g2_decap_8 FILLER_29_2943 ();
 sg13g2_decap_8 FILLER_29_2950 ();
 sg13g2_fill_2 FILLER_29_2957 ();
 sg13g2_fill_1 FILLER_29_2959 ();
 sg13g2_fill_1 FILLER_29_2976 ();
 sg13g2_fill_2 FILLER_29_2997 ();
 sg13g2_decap_8 FILLER_29_3020 ();
 sg13g2_decap_4 FILLER_29_3027 ();
 sg13g2_fill_2 FILLER_29_3031 ();
 sg13g2_decap_8 FILLER_29_3050 ();
 sg13g2_decap_8 FILLER_29_3057 ();
 sg13g2_fill_1 FILLER_29_3064 ();
 sg13g2_fill_2 FILLER_29_3070 ();
 sg13g2_fill_2 FILLER_29_3094 ();
 sg13g2_fill_1 FILLER_29_3109 ();
 sg13g2_fill_2 FILLER_29_3174 ();
 sg13g2_fill_1 FILLER_29_3204 ();
 sg13g2_decap_8 FILLER_29_3218 ();
 sg13g2_fill_2 FILLER_29_3225 ();
 sg13g2_fill_1 FILLER_29_3227 ();
 sg13g2_fill_1 FILLER_29_3256 ();
 sg13g2_decap_8 FILLER_29_3261 ();
 sg13g2_fill_1 FILLER_29_3268 ();
 sg13g2_decap_8 FILLER_29_3294 ();
 sg13g2_decap_4 FILLER_29_3301 ();
 sg13g2_fill_2 FILLER_29_3305 ();
 sg13g2_fill_2 FILLER_29_3340 ();
 sg13g2_decap_4 FILLER_29_3345 ();
 sg13g2_fill_2 FILLER_29_3349 ();
 sg13g2_decap_8 FILLER_29_3379 ();
 sg13g2_decap_8 FILLER_29_3386 ();
 sg13g2_decap_8 FILLER_29_3393 ();
 sg13g2_decap_8 FILLER_29_3400 ();
 sg13g2_decap_8 FILLER_29_3407 ();
 sg13g2_decap_8 FILLER_29_3414 ();
 sg13g2_decap_8 FILLER_29_3421 ();
 sg13g2_decap_8 FILLER_29_3428 ();
 sg13g2_decap_8 FILLER_29_3435 ();
 sg13g2_decap_8 FILLER_29_3442 ();
 sg13g2_decap_8 FILLER_29_3449 ();
 sg13g2_decap_8 FILLER_29_3456 ();
 sg13g2_decap_8 FILLER_29_3463 ();
 sg13g2_decap_8 FILLER_29_3470 ();
 sg13g2_decap_8 FILLER_29_3477 ();
 sg13g2_decap_8 FILLER_29_3484 ();
 sg13g2_decap_8 FILLER_29_3491 ();
 sg13g2_decap_8 FILLER_29_3498 ();
 sg13g2_decap_8 FILLER_29_3505 ();
 sg13g2_decap_8 FILLER_29_3512 ();
 sg13g2_decap_8 FILLER_29_3519 ();
 sg13g2_decap_8 FILLER_29_3526 ();
 sg13g2_decap_8 FILLER_29_3533 ();
 sg13g2_decap_8 FILLER_29_3540 ();
 sg13g2_decap_8 FILLER_29_3547 ();
 sg13g2_decap_8 FILLER_29_3554 ();
 sg13g2_decap_8 FILLER_29_3561 ();
 sg13g2_decap_8 FILLER_29_3568 ();
 sg13g2_decap_4 FILLER_29_3575 ();
 sg13g2_fill_1 FILLER_29_3579 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_decap_8 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_fill_2 FILLER_30_419 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_4 FILLER_30_441 ();
 sg13g2_fill_1 FILLER_30_445 ();
 sg13g2_fill_1 FILLER_30_451 ();
 sg13g2_decap_8 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_472 ();
 sg13g2_fill_1 FILLER_30_488 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_fill_2 FILLER_30_508 ();
 sg13g2_fill_1 FILLER_30_525 ();
 sg13g2_fill_2 FILLER_30_551 ();
 sg13g2_fill_1 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_fill_1 FILLER_30_574 ();
 sg13g2_fill_1 FILLER_30_579 ();
 sg13g2_decap_8 FILLER_30_591 ();
 sg13g2_decap_8 FILLER_30_598 ();
 sg13g2_decap_4 FILLER_30_605 ();
 sg13g2_decap_8 FILLER_30_613 ();
 sg13g2_fill_2 FILLER_30_620 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_634 ();
 sg13g2_decap_4 FILLER_30_641 ();
 sg13g2_fill_1 FILLER_30_645 ();
 sg13g2_decap_8 FILLER_30_659 ();
 sg13g2_decap_4 FILLER_30_666 ();
 sg13g2_fill_2 FILLER_30_670 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_4 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_754 ();
 sg13g2_fill_1 FILLER_30_761 ();
 sg13g2_fill_1 FILLER_30_779 ();
 sg13g2_fill_1 FILLER_30_784 ();
 sg13g2_fill_2 FILLER_30_803 ();
 sg13g2_fill_1 FILLER_30_805 ();
 sg13g2_fill_2 FILLER_30_815 ();
 sg13g2_fill_1 FILLER_30_850 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_4 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_886 ();
 sg13g2_fill_1 FILLER_30_893 ();
 sg13g2_fill_2 FILLER_30_899 ();
 sg13g2_fill_1 FILLER_30_901 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_4 FILLER_30_945 ();
 sg13g2_fill_1 FILLER_30_949 ();
 sg13g2_fill_1 FILLER_30_993 ();
 sg13g2_fill_2 FILLER_30_1006 ();
 sg13g2_fill_1 FILLER_30_1008 ();
 sg13g2_fill_2 FILLER_30_1032 ();
 sg13g2_decap_4 FILLER_30_1052 ();
 sg13g2_fill_1 FILLER_30_1056 ();
 sg13g2_decap_8 FILLER_30_1086 ();
 sg13g2_decap_8 FILLER_30_1093 ();
 sg13g2_fill_1 FILLER_30_1100 ();
 sg13g2_decap_8 FILLER_30_1127 ();
 sg13g2_decap_4 FILLER_30_1134 ();
 sg13g2_decap_8 FILLER_30_1158 ();
 sg13g2_fill_2 FILLER_30_1165 ();
 sg13g2_fill_1 FILLER_30_1167 ();
 sg13g2_fill_2 FILLER_30_1214 ();
 sg13g2_fill_1 FILLER_30_1216 ();
 sg13g2_decap_4 FILLER_30_1247 ();
 sg13g2_fill_1 FILLER_30_1251 ();
 sg13g2_decap_4 FILLER_30_1276 ();
 sg13g2_fill_2 FILLER_30_1280 ();
 sg13g2_decap_8 FILLER_30_1295 ();
 sg13g2_fill_2 FILLER_30_1316 ();
 sg13g2_decap_8 FILLER_30_1346 ();
 sg13g2_decap_8 FILLER_30_1353 ();
 sg13g2_fill_1 FILLER_30_1360 ();
 sg13g2_fill_2 FILLER_30_1377 ();
 sg13g2_fill_2 FILLER_30_1384 ();
 sg13g2_fill_2 FILLER_30_1390 ();
 sg13g2_decap_8 FILLER_30_1413 ();
 sg13g2_decap_8 FILLER_30_1420 ();
 sg13g2_fill_2 FILLER_30_1427 ();
 sg13g2_fill_1 FILLER_30_1429 ();
 sg13g2_decap_8 FILLER_30_1444 ();
 sg13g2_fill_2 FILLER_30_1456 ();
 sg13g2_decap_8 FILLER_30_1462 ();
 sg13g2_decap_4 FILLER_30_1469 ();
 sg13g2_fill_2 FILLER_30_1473 ();
 sg13g2_decap_8 FILLER_30_1492 ();
 sg13g2_decap_8 FILLER_30_1499 ();
 sg13g2_fill_2 FILLER_30_1506 ();
 sg13g2_fill_2 FILLER_30_1526 ();
 sg13g2_fill_1 FILLER_30_1528 ();
 sg13g2_decap_8 FILLER_30_1546 ();
 sg13g2_fill_1 FILLER_30_1553 ();
 sg13g2_decap_4 FILLER_30_1559 ();
 sg13g2_fill_1 FILLER_30_1563 ();
 sg13g2_decap_8 FILLER_30_1567 ();
 sg13g2_decap_8 FILLER_30_1574 ();
 sg13g2_fill_2 FILLER_30_1593 ();
 sg13g2_fill_2 FILLER_30_1600 ();
 sg13g2_decap_8 FILLER_30_1615 ();
 sg13g2_decap_4 FILLER_30_1622 ();
 sg13g2_fill_2 FILLER_30_1626 ();
 sg13g2_fill_1 FILLER_30_1659 ();
 sg13g2_decap_8 FILLER_30_1667 ();
 sg13g2_fill_2 FILLER_30_1674 ();
 sg13g2_fill_1 FILLER_30_1682 ();
 sg13g2_decap_4 FILLER_30_1686 ();
 sg13g2_fill_1 FILLER_30_1690 ();
 sg13g2_decap_8 FILLER_30_1695 ();
 sg13g2_fill_2 FILLER_30_1702 ();
 sg13g2_fill_1 FILLER_30_1704 ();
 sg13g2_decap_8 FILLER_30_1761 ();
 sg13g2_decap_4 FILLER_30_1768 ();
 sg13g2_decap_4 FILLER_30_1776 ();
 sg13g2_decap_8 FILLER_30_1804 ();
 sg13g2_decap_8 FILLER_30_1811 ();
 sg13g2_fill_1 FILLER_30_1818 ();
 sg13g2_fill_2 FILLER_30_1823 ();
 sg13g2_fill_2 FILLER_30_1853 ();
 sg13g2_fill_2 FILLER_30_1877 ();
 sg13g2_decap_8 FILLER_30_1886 ();
 sg13g2_decap_4 FILLER_30_1893 ();
 sg13g2_fill_1 FILLER_30_1934 ();
 sg13g2_fill_1 FILLER_30_1944 ();
 sg13g2_fill_1 FILLER_30_1981 ();
 sg13g2_decap_8 FILLER_30_1994 ();
 sg13g2_fill_2 FILLER_30_2001 ();
 sg13g2_decap_8 FILLER_30_2025 ();
 sg13g2_fill_2 FILLER_30_2032 ();
 sg13g2_fill_1 FILLER_30_2034 ();
 sg13g2_decap_8 FILLER_30_2040 ();
 sg13g2_decap_4 FILLER_30_2047 ();
 sg13g2_fill_1 FILLER_30_2055 ();
 sg13g2_decap_8 FILLER_30_2064 ();
 sg13g2_decap_8 FILLER_30_2093 ();
 sg13g2_decap_8 FILLER_30_2100 ();
 sg13g2_fill_1 FILLER_30_2107 ();
 sg13g2_decap_8 FILLER_30_2129 ();
 sg13g2_decap_4 FILLER_30_2157 ();
 sg13g2_decap_8 FILLER_30_2169 ();
 sg13g2_decap_8 FILLER_30_2179 ();
 sg13g2_decap_4 FILLER_30_2192 ();
 sg13g2_fill_1 FILLER_30_2196 ();
 sg13g2_decap_8 FILLER_30_2213 ();
 sg13g2_decap_4 FILLER_30_2220 ();
 sg13g2_fill_1 FILLER_30_2245 ();
 sg13g2_fill_2 FILLER_30_2263 ();
 sg13g2_decap_4 FILLER_30_2271 ();
 sg13g2_fill_2 FILLER_30_2275 ();
 sg13g2_decap_4 FILLER_30_2285 ();
 sg13g2_decap_8 FILLER_30_2311 ();
 sg13g2_fill_2 FILLER_30_2318 ();
 sg13g2_fill_1 FILLER_30_2325 ();
 sg13g2_fill_1 FILLER_30_2339 ();
 sg13g2_decap_8 FILLER_30_2344 ();
 sg13g2_decap_4 FILLER_30_2351 ();
 sg13g2_decap_4 FILLER_30_2374 ();
 sg13g2_decap_8 FILLER_30_2391 ();
 sg13g2_fill_2 FILLER_30_2398 ();
 sg13g2_fill_1 FILLER_30_2400 ();
 sg13g2_decap_8 FILLER_30_2414 ();
 sg13g2_fill_1 FILLER_30_2421 ();
 sg13g2_decap_8 FILLER_30_2440 ();
 sg13g2_decap_8 FILLER_30_2455 ();
 sg13g2_decap_8 FILLER_30_2462 ();
 sg13g2_decap_8 FILLER_30_2469 ();
 sg13g2_fill_1 FILLER_30_2476 ();
 sg13g2_fill_2 FILLER_30_2490 ();
 sg13g2_fill_1 FILLER_30_2492 ();
 sg13g2_fill_2 FILLER_30_2498 ();
 sg13g2_fill_1 FILLER_30_2500 ();
 sg13g2_decap_8 FILLER_30_2514 ();
 sg13g2_decap_8 FILLER_30_2521 ();
 sg13g2_decap_8 FILLER_30_2528 ();
 sg13g2_fill_2 FILLER_30_2535 ();
 sg13g2_fill_1 FILLER_30_2537 ();
 sg13g2_decap_8 FILLER_30_2560 ();
 sg13g2_fill_1 FILLER_30_2580 ();
 sg13g2_decap_8 FILLER_30_2597 ();
 sg13g2_decap_8 FILLER_30_2604 ();
 sg13g2_fill_1 FILLER_30_2637 ();
 sg13g2_decap_4 FILLER_30_2645 ();
 sg13g2_decap_4 FILLER_30_2670 ();
 sg13g2_decap_4 FILLER_30_2679 ();
 sg13g2_decap_8 FILLER_30_2688 ();
 sg13g2_decap_8 FILLER_30_2699 ();
 sg13g2_decap_8 FILLER_30_2706 ();
 sg13g2_fill_2 FILLER_30_2719 ();
 sg13g2_decap_8 FILLER_30_2733 ();
 sg13g2_decap_4 FILLER_30_2740 ();
 sg13g2_fill_1 FILLER_30_2744 ();
 sg13g2_fill_1 FILLER_30_2777 ();
 sg13g2_decap_4 FILLER_30_2806 ();
 sg13g2_fill_2 FILLER_30_2818 ();
 sg13g2_fill_2 FILLER_30_2847 ();
 sg13g2_decap_8 FILLER_30_2865 ();
 sg13g2_decap_8 FILLER_30_2889 ();
 sg13g2_decap_8 FILLER_30_2906 ();
 sg13g2_fill_2 FILLER_30_2913 ();
 sg13g2_fill_1 FILLER_30_2915 ();
 sg13g2_decap_8 FILLER_30_2936 ();
 sg13g2_fill_2 FILLER_30_2948 ();
 sg13g2_decap_8 FILLER_30_2964 ();
 sg13g2_decap_8 FILLER_30_2971 ();
 sg13g2_fill_2 FILLER_30_2978 ();
 sg13g2_fill_1 FILLER_30_2980 ();
 sg13g2_decap_8 FILLER_30_2994 ();
 sg13g2_decap_4 FILLER_30_3001 ();
 sg13g2_decap_8 FILLER_30_3011 ();
 sg13g2_fill_2 FILLER_30_3018 ();
 sg13g2_fill_2 FILLER_30_3024 ();
 sg13g2_fill_2 FILLER_30_3042 ();
 sg13g2_decap_8 FILLER_30_3052 ();
 sg13g2_fill_2 FILLER_30_3059 ();
 sg13g2_fill_1 FILLER_30_3061 ();
 sg13g2_fill_2 FILLER_30_3089 ();
 sg13g2_fill_2 FILLER_30_3131 ();
 sg13g2_fill_2 FILLER_30_3169 ();
 sg13g2_fill_2 FILLER_30_3194 ();
 sg13g2_decap_8 FILLER_30_3233 ();
 sg13g2_decap_4 FILLER_30_3240 ();
 sg13g2_fill_1 FILLER_30_3244 ();
 sg13g2_decap_4 FILLER_30_3295 ();
 sg13g2_fill_1 FILLER_30_3299 ();
 sg13g2_fill_2 FILLER_30_3310 ();
 sg13g2_fill_1 FILLER_30_3312 ();
 sg13g2_fill_2 FILLER_30_3345 ();
 sg13g2_decap_4 FILLER_30_3360 ();
 sg13g2_fill_2 FILLER_30_3364 ();
 sg13g2_decap_8 FILLER_30_3375 ();
 sg13g2_decap_8 FILLER_30_3382 ();
 sg13g2_decap_8 FILLER_30_3389 ();
 sg13g2_decap_8 FILLER_30_3396 ();
 sg13g2_decap_8 FILLER_30_3403 ();
 sg13g2_decap_8 FILLER_30_3410 ();
 sg13g2_decap_8 FILLER_30_3417 ();
 sg13g2_decap_8 FILLER_30_3424 ();
 sg13g2_decap_8 FILLER_30_3431 ();
 sg13g2_decap_8 FILLER_30_3438 ();
 sg13g2_decap_8 FILLER_30_3445 ();
 sg13g2_decap_8 FILLER_30_3452 ();
 sg13g2_decap_8 FILLER_30_3459 ();
 sg13g2_decap_8 FILLER_30_3466 ();
 sg13g2_decap_8 FILLER_30_3473 ();
 sg13g2_decap_8 FILLER_30_3480 ();
 sg13g2_decap_8 FILLER_30_3487 ();
 sg13g2_decap_8 FILLER_30_3494 ();
 sg13g2_decap_8 FILLER_30_3501 ();
 sg13g2_decap_8 FILLER_30_3508 ();
 sg13g2_decap_8 FILLER_30_3515 ();
 sg13g2_decap_8 FILLER_30_3522 ();
 sg13g2_decap_8 FILLER_30_3529 ();
 sg13g2_decap_8 FILLER_30_3536 ();
 sg13g2_decap_8 FILLER_30_3543 ();
 sg13g2_decap_8 FILLER_30_3550 ();
 sg13g2_decap_8 FILLER_30_3557 ();
 sg13g2_decap_8 FILLER_30_3564 ();
 sg13g2_decap_8 FILLER_30_3571 ();
 sg13g2_fill_2 FILLER_30_3578 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_205 ();
 sg13g2_decap_4 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_fill_2 FILLER_31_385 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_404 ();
 sg13g2_fill_2 FILLER_31_411 ();
 sg13g2_fill_2 FILLER_31_418 ();
 sg13g2_fill_1 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_431 ();
 sg13g2_decap_8 FILLER_31_461 ();
 sg13g2_decap_8 FILLER_31_468 ();
 sg13g2_fill_2 FILLER_31_475 ();
 sg13g2_decap_8 FILLER_31_486 ();
 sg13g2_fill_2 FILLER_31_493 ();
 sg13g2_fill_1 FILLER_31_495 ();
 sg13g2_fill_2 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_decap_8 FILLER_31_559 ();
 sg13g2_decap_8 FILLER_31_566 ();
 sg13g2_fill_2 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_599 ();
 sg13g2_decap_8 FILLER_31_606 ();
 sg13g2_fill_2 FILLER_31_613 ();
 sg13g2_decap_4 FILLER_31_632 ();
 sg13g2_fill_1 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_decap_4 FILLER_31_666 ();
 sg13g2_fill_1 FILLER_31_670 ();
 sg13g2_decap_4 FILLER_31_676 ();
 sg13g2_fill_1 FILLER_31_680 ();
 sg13g2_fill_2 FILLER_31_685 ();
 sg13g2_decap_4 FILLER_31_705 ();
 sg13g2_fill_1 FILLER_31_709 ();
 sg13g2_fill_1 FILLER_31_728 ();
 sg13g2_decap_4 FILLER_31_781 ();
 sg13g2_fill_2 FILLER_31_785 ();
 sg13g2_decap_4 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_4 FILLER_31_821 ();
 sg13g2_fill_2 FILLER_31_825 ();
 sg13g2_decap_4 FILLER_31_832 ();
 sg13g2_fill_1 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_4 FILLER_31_861 ();
 sg13g2_decap_4 FILLER_31_880 ();
 sg13g2_fill_1 FILLER_31_904 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_4 FILLER_31_917 ();
 sg13g2_decap_4 FILLER_31_936 ();
 sg13g2_fill_1 FILLER_31_940 ();
 sg13g2_fill_2 FILLER_31_957 ();
 sg13g2_fill_1 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_fill_1 FILLER_31_980 ();
 sg13g2_fill_1 FILLER_31_985 ();
 sg13g2_decap_8 FILLER_31_995 ();
 sg13g2_fill_1 FILLER_31_1017 ();
 sg13g2_fill_2 FILLER_31_1024 ();
 sg13g2_fill_1 FILLER_31_1026 ();
 sg13g2_decap_8 FILLER_31_1075 ();
 sg13g2_fill_2 FILLER_31_1082 ();
 sg13g2_decap_8 FILLER_31_1088 ();
 sg13g2_decap_8 FILLER_31_1095 ();
 sg13g2_decap_4 FILLER_31_1102 ();
 sg13g2_fill_1 FILLER_31_1106 ();
 sg13g2_fill_1 FILLER_31_1123 ();
 sg13g2_decap_8 FILLER_31_1156 ();
 sg13g2_decap_8 FILLER_31_1163 ();
 sg13g2_fill_1 FILLER_31_1170 ();
 sg13g2_decap_4 FILLER_31_1179 ();
 sg13g2_fill_2 FILLER_31_1183 ();
 sg13g2_fill_2 FILLER_31_1210 ();
 sg13g2_fill_2 FILLER_31_1237 ();
 sg13g2_fill_1 FILLER_31_1239 ();
 sg13g2_decap_4 FILLER_31_1265 ();
 sg13g2_fill_2 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1280 ();
 sg13g2_decap_4 FILLER_31_1287 ();
 sg13g2_decap_8 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1302 ();
 sg13g2_fill_2 FILLER_31_1309 ();
 sg13g2_decap_8 FILLER_31_1347 ();
 sg13g2_decap_4 FILLER_31_1354 ();
 sg13g2_fill_1 FILLER_31_1358 ();
 sg13g2_fill_1 FILLER_31_1377 ();
 sg13g2_fill_1 FILLER_31_1386 ();
 sg13g2_fill_2 FILLER_31_1392 ();
 sg13g2_fill_1 FILLER_31_1399 ();
 sg13g2_decap_4 FILLER_31_1417 ();
 sg13g2_fill_2 FILLER_31_1421 ();
 sg13g2_fill_2 FILLER_31_1453 ();
 sg13g2_fill_1 FILLER_31_1455 ();
 sg13g2_decap_8 FILLER_31_1468 ();
 sg13g2_decap_8 FILLER_31_1485 ();
 sg13g2_fill_2 FILLER_31_1492 ();
 sg13g2_fill_1 FILLER_31_1494 ();
 sg13g2_decap_4 FILLER_31_1504 ();
 sg13g2_fill_1 FILLER_31_1508 ();
 sg13g2_fill_1 FILLER_31_1513 ();
 sg13g2_decap_8 FILLER_31_1527 ();
 sg13g2_fill_1 FILLER_31_1534 ();
 sg13g2_decap_8 FILLER_31_1546 ();
 sg13g2_decap_4 FILLER_31_1553 ();
 sg13g2_fill_1 FILLER_31_1557 ();
 sg13g2_decap_8 FILLER_31_1573 ();
 sg13g2_fill_1 FILLER_31_1589 ();
 sg13g2_fill_2 FILLER_31_1603 ();
 sg13g2_fill_1 FILLER_31_1605 ();
 sg13g2_fill_2 FILLER_31_1634 ();
 sg13g2_fill_1 FILLER_31_1636 ();
 sg13g2_fill_1 FILLER_31_1654 ();
 sg13g2_decap_8 FILLER_31_1692 ();
 sg13g2_decap_4 FILLER_31_1699 ();
 sg13g2_decap_8 FILLER_31_1721 ();
 sg13g2_decap_8 FILLER_31_1728 ();
 sg13g2_fill_2 FILLER_31_1735 ();
 sg13g2_fill_1 FILLER_31_1737 ();
 sg13g2_decap_8 FILLER_31_1742 ();
 sg13g2_decap_4 FILLER_31_1749 ();
 sg13g2_fill_2 FILLER_31_1765 ();
 sg13g2_decap_4 FILLER_31_1835 ();
 sg13g2_fill_2 FILLER_31_1839 ();
 sg13g2_fill_2 FILLER_31_1851 ();
 sg13g2_fill_1 FILLER_31_1853 ();
 sg13g2_decap_4 FILLER_31_1904 ();
 sg13g2_fill_2 FILLER_31_1929 ();
 sg13g2_fill_1 FILLER_31_1931 ();
 sg13g2_decap_8 FILLER_31_1952 ();
 sg13g2_fill_1 FILLER_31_1959 ();
 sg13g2_decap_8 FILLER_31_1985 ();
 sg13g2_decap_8 FILLER_31_1992 ();
 sg13g2_fill_2 FILLER_31_1999 ();
 sg13g2_fill_1 FILLER_31_2001 ();
 sg13g2_fill_1 FILLER_31_2027 ();
 sg13g2_decap_8 FILLER_31_2048 ();
 sg13g2_fill_2 FILLER_31_2055 ();
 sg13g2_decap_4 FILLER_31_2099 ();
 sg13g2_fill_2 FILLER_31_2124 ();
 sg13g2_fill_2 FILLER_31_2134 ();
 sg13g2_fill_1 FILLER_31_2136 ();
 sg13g2_decap_8 FILLER_31_2152 ();
 sg13g2_decap_8 FILLER_31_2159 ();
 sg13g2_decap_4 FILLER_31_2166 ();
 sg13g2_fill_1 FILLER_31_2170 ();
 sg13g2_fill_2 FILLER_31_2196 ();
 sg13g2_decap_8 FILLER_31_2211 ();
 sg13g2_decap_4 FILLER_31_2218 ();
 sg13g2_decap_4 FILLER_31_2244 ();
 sg13g2_fill_1 FILLER_31_2265 ();
 sg13g2_decap_4 FILLER_31_2275 ();
 sg13g2_decap_4 FILLER_31_2284 ();
 sg13g2_fill_2 FILLER_31_2288 ();
 sg13g2_decap_4 FILLER_31_2307 ();
 sg13g2_fill_1 FILLER_31_2311 ();
 sg13g2_decap_8 FILLER_31_2325 ();
 sg13g2_decap_8 FILLER_31_2332 ();
 sg13g2_decap_8 FILLER_31_2339 ();
 sg13g2_decap_4 FILLER_31_2346 ();
 sg13g2_fill_2 FILLER_31_2372 ();
 sg13g2_decap_8 FILLER_31_2395 ();
 sg13g2_decap_4 FILLER_31_2411 ();
 sg13g2_fill_2 FILLER_31_2440 ();
 sg13g2_fill_1 FILLER_31_2442 ();
 sg13g2_fill_1 FILLER_31_2469 ();
 sg13g2_fill_2 FILLER_31_2495 ();
 sg13g2_decap_4 FILLER_31_2522 ();
 sg13g2_fill_2 FILLER_31_2526 ();
 sg13g2_decap_4 FILLER_31_2533 ();
 sg13g2_fill_2 FILLER_31_2537 ();
 sg13g2_fill_2 FILLER_31_2546 ();
 sg13g2_decap_4 FILLER_31_2561 ();
 sg13g2_fill_1 FILLER_31_2571 ();
 sg13g2_fill_2 FILLER_31_2580 ();
 sg13g2_fill_1 FILLER_31_2582 ();
 sg13g2_fill_2 FILLER_31_2605 ();
 sg13g2_fill_1 FILLER_31_2607 ();
 sg13g2_decap_8 FILLER_31_2629 ();
 sg13g2_decap_8 FILLER_31_2636 ();
 sg13g2_decap_8 FILLER_31_2643 ();
 sg13g2_fill_2 FILLER_31_2655 ();
 sg13g2_fill_1 FILLER_31_2662 ();
 sg13g2_fill_1 FILLER_31_2671 ();
 sg13g2_fill_2 FILLER_31_2676 ();
 sg13g2_decap_4 FILLER_31_2683 ();
 sg13g2_decap_8 FILLER_31_2703 ();
 sg13g2_decap_4 FILLER_31_2710 ();
 sg13g2_fill_1 FILLER_31_2714 ();
 sg13g2_fill_2 FILLER_31_2736 ();
 sg13g2_decap_4 FILLER_31_2747 ();
 sg13g2_fill_1 FILLER_31_2751 ();
 sg13g2_decap_8 FILLER_31_2790 ();
 sg13g2_decap_8 FILLER_31_2797 ();
 sg13g2_fill_2 FILLER_31_2804 ();
 sg13g2_fill_2 FILLER_31_2811 ();
 sg13g2_fill_1 FILLER_31_2813 ();
 sg13g2_fill_2 FILLER_31_2819 ();
 sg13g2_fill_1 FILLER_31_2821 ();
 sg13g2_fill_1 FILLER_31_2826 ();
 sg13g2_decap_4 FILLER_31_2840 ();
 sg13g2_decap_8 FILLER_31_2849 ();
 sg13g2_decap_8 FILLER_31_2856 ();
 sg13g2_fill_1 FILLER_31_2863 ();
 sg13g2_fill_1 FILLER_31_2889 ();
 sg13g2_fill_2 FILLER_31_2895 ();
 sg13g2_fill_1 FILLER_31_2897 ();
 sg13g2_fill_1 FILLER_31_2911 ();
 sg13g2_fill_1 FILLER_31_2924 ();
 sg13g2_decap_8 FILLER_31_2930 ();
 sg13g2_decap_8 FILLER_31_2937 ();
 sg13g2_decap_4 FILLER_31_2950 ();
 sg13g2_decap_4 FILLER_31_2962 ();
 sg13g2_fill_2 FILLER_31_2966 ();
 sg13g2_fill_2 FILLER_31_2981 ();
 sg13g2_fill_1 FILLER_31_2983 ();
 sg13g2_decap_4 FILLER_31_3000 ();
 sg13g2_fill_1 FILLER_31_3009 ();
 sg13g2_fill_1 FILLER_31_3018 ();
 sg13g2_decap_8 FILLER_31_3035 ();
 sg13g2_decap_8 FILLER_31_3042 ();
 sg13g2_fill_2 FILLER_31_3049 ();
 sg13g2_fill_1 FILLER_31_3051 ();
 sg13g2_fill_2 FILLER_31_3057 ();
 sg13g2_fill_1 FILLER_31_3059 ();
 sg13g2_fill_2 FILLER_31_3081 ();
 sg13g2_fill_1 FILLER_31_3088 ();
 sg13g2_fill_1 FILLER_31_3129 ();
 sg13g2_fill_1 FILLER_31_3135 ();
 sg13g2_fill_2 FILLER_31_3172 ();
 sg13g2_fill_2 FILLER_31_3187 ();
 sg13g2_fill_1 FILLER_31_3189 ();
 sg13g2_decap_8 FILLER_31_3217 ();
 sg13g2_decap_4 FILLER_31_3224 ();
 sg13g2_fill_2 FILLER_31_3246 ();
 sg13g2_decap_8 FILLER_31_3266 ();
 sg13g2_decap_4 FILLER_31_3273 ();
 sg13g2_fill_1 FILLER_31_3277 ();
 sg13g2_decap_4 FILLER_31_3291 ();
 sg13g2_fill_1 FILLER_31_3295 ();
 sg13g2_fill_2 FILLER_31_3321 ();
 sg13g2_fill_2 FILLER_31_3339 ();
 sg13g2_fill_2 FILLER_31_3355 ();
 sg13g2_decap_8 FILLER_31_3360 ();
 sg13g2_fill_1 FILLER_31_3367 ();
 sg13g2_fill_2 FILLER_31_3372 ();
 sg13g2_decap_8 FILLER_31_3383 ();
 sg13g2_decap_8 FILLER_31_3390 ();
 sg13g2_decap_8 FILLER_31_3397 ();
 sg13g2_decap_8 FILLER_31_3404 ();
 sg13g2_decap_8 FILLER_31_3411 ();
 sg13g2_decap_8 FILLER_31_3418 ();
 sg13g2_decap_8 FILLER_31_3425 ();
 sg13g2_decap_8 FILLER_31_3432 ();
 sg13g2_decap_8 FILLER_31_3439 ();
 sg13g2_decap_8 FILLER_31_3446 ();
 sg13g2_decap_8 FILLER_31_3453 ();
 sg13g2_decap_8 FILLER_31_3460 ();
 sg13g2_decap_8 FILLER_31_3467 ();
 sg13g2_decap_8 FILLER_31_3474 ();
 sg13g2_decap_8 FILLER_31_3481 ();
 sg13g2_decap_8 FILLER_31_3488 ();
 sg13g2_decap_8 FILLER_31_3495 ();
 sg13g2_decap_8 FILLER_31_3502 ();
 sg13g2_decap_8 FILLER_31_3509 ();
 sg13g2_decap_8 FILLER_31_3516 ();
 sg13g2_decap_8 FILLER_31_3523 ();
 sg13g2_decap_8 FILLER_31_3530 ();
 sg13g2_decap_8 FILLER_31_3537 ();
 sg13g2_decap_8 FILLER_31_3544 ();
 sg13g2_decap_8 FILLER_31_3551 ();
 sg13g2_decap_8 FILLER_31_3558 ();
 sg13g2_decap_8 FILLER_31_3565 ();
 sg13g2_decap_8 FILLER_31_3572 ();
 sg13g2_fill_1 FILLER_31_3579 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_fill_2 FILLER_32_435 ();
 sg13g2_fill_2 FILLER_32_455 ();
 sg13g2_fill_1 FILLER_32_462 ();
 sg13g2_decap_4 FILLER_32_504 ();
 sg13g2_fill_2 FILLER_32_508 ();
 sg13g2_fill_2 FILLER_32_533 ();
 sg13g2_fill_2 FILLER_32_545 ();
 sg13g2_decap_8 FILLER_32_563 ();
 sg13g2_decap_4 FILLER_32_570 ();
 sg13g2_fill_2 FILLER_32_574 ();
 sg13g2_fill_2 FILLER_32_589 ();
 sg13g2_fill_2 FILLER_32_605 ();
 sg13g2_fill_2 FILLER_32_612 ();
 sg13g2_decap_4 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_656 ();
 sg13g2_decap_4 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_4 FILLER_32_707 ();
 sg13g2_fill_2 FILLER_32_732 ();
 sg13g2_fill_1 FILLER_32_734 ();
 sg13g2_fill_1 FILLER_32_752 ();
 sg13g2_fill_2 FILLER_32_763 ();
 sg13g2_decap_4 FILLER_32_773 ();
 sg13g2_fill_2 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_fill_2 FILLER_32_822 ();
 sg13g2_fill_1 FILLER_32_824 ();
 sg13g2_fill_1 FILLER_32_838 ();
 sg13g2_fill_2 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_fill_2 FILLER_32_864 ();
 sg13g2_decap_4 FILLER_32_870 ();
 sg13g2_fill_2 FILLER_32_874 ();
 sg13g2_decap_8 FILLER_32_881 ();
 sg13g2_fill_2 FILLER_32_888 ();
 sg13g2_fill_1 FILLER_32_890 ();
 sg13g2_fill_2 FILLER_32_897 ();
 sg13g2_fill_1 FILLER_32_899 ();
 sg13g2_decap_8 FILLER_32_905 ();
 sg13g2_fill_1 FILLER_32_912 ();
 sg13g2_fill_2 FILLER_32_930 ();
 sg13g2_fill_1 FILLER_32_932 ();
 sg13g2_fill_1 FILLER_32_938 ();
 sg13g2_fill_1 FILLER_32_951 ();
 sg13g2_fill_2 FILLER_32_955 ();
 sg13g2_fill_2 FILLER_32_969 ();
 sg13g2_fill_2 FILLER_32_983 ();
 sg13g2_fill_1 FILLER_32_1040 ();
 sg13g2_decap_8 FILLER_32_1048 ();
 sg13g2_decap_4 FILLER_32_1055 ();
 sg13g2_fill_1 FILLER_32_1059 ();
 sg13g2_fill_1 FILLER_32_1077 ();
 sg13g2_fill_1 FILLER_32_1106 ();
 sg13g2_fill_1 FILLER_32_1135 ();
 sg13g2_fill_2 FILLER_32_1154 ();
 sg13g2_fill_1 FILLER_32_1171 ();
 sg13g2_fill_2 FILLER_32_1180 ();
 sg13g2_fill_1 FILLER_32_1182 ();
 sg13g2_fill_2 FILLER_32_1196 ();
 sg13g2_fill_1 FILLER_32_1198 ();
 sg13g2_fill_2 FILLER_32_1210 ();
 sg13g2_fill_1 FILLER_32_1212 ();
 sg13g2_fill_2 FILLER_32_1230 ();
 sg13g2_fill_1 FILLER_32_1232 ();
 sg13g2_decap_4 FILLER_32_1241 ();
 sg13g2_fill_1 FILLER_32_1245 ();
 sg13g2_decap_4 FILLER_32_1255 ();
 sg13g2_decap_4 FILLER_32_1267 ();
 sg13g2_fill_2 FILLER_32_1284 ();
 sg13g2_decap_4 FILLER_32_1314 ();
 sg13g2_fill_1 FILLER_32_1318 ();
 sg13g2_fill_2 FILLER_32_1328 ();
 sg13g2_decap_8 FILLER_32_1341 ();
 sg13g2_decap_8 FILLER_32_1348 ();
 sg13g2_fill_2 FILLER_32_1355 ();
 sg13g2_decap_4 FILLER_32_1363 ();
 sg13g2_fill_1 FILLER_32_1367 ();
 sg13g2_fill_2 FILLER_32_1377 ();
 sg13g2_fill_1 FILLER_32_1391 ();
 sg13g2_decap_8 FILLER_32_1402 ();
 sg13g2_decap_8 FILLER_32_1409 ();
 sg13g2_decap_8 FILLER_32_1416 ();
 sg13g2_fill_2 FILLER_32_1423 ();
 sg13g2_decap_4 FILLER_32_1460 ();
 sg13g2_decap_4 FILLER_32_1469 ();
 sg13g2_fill_2 FILLER_32_1473 ();
 sg13g2_decap_4 FILLER_32_1490 ();
 sg13g2_decap_4 FILLER_32_1531 ();
 sg13g2_fill_2 FILLER_32_1535 ();
 sg13g2_fill_2 FILLER_32_1540 ();
 sg13g2_decap_4 FILLER_32_1546 ();
 sg13g2_fill_1 FILLER_32_1550 ();
 sg13g2_fill_1 FILLER_32_1560 ();
 sg13g2_decap_8 FILLER_32_1643 ();
 sg13g2_fill_2 FILLER_32_1650 ();
 sg13g2_fill_1 FILLER_32_1652 ();
 sg13g2_decap_8 FILLER_32_1665 ();
 sg13g2_fill_2 FILLER_32_1672 ();
 sg13g2_fill_1 FILLER_32_1674 ();
 sg13g2_fill_1 FILLER_32_1715 ();
 sg13g2_fill_2 FILLER_32_1721 ();
 sg13g2_fill_2 FILLER_32_1741 ();
 sg13g2_decap_8 FILLER_32_1746 ();
 sg13g2_fill_2 FILLER_32_1753 ();
 sg13g2_decap_4 FILLER_32_1783 ();
 sg13g2_fill_1 FILLER_32_1787 ();
 sg13g2_decap_8 FILLER_32_1807 ();
 sg13g2_fill_2 FILLER_32_1814 ();
 sg13g2_decap_8 FILLER_32_1830 ();
 sg13g2_fill_1 FILLER_32_1861 ();
 sg13g2_decap_8 FILLER_32_1866 ();
 sg13g2_decap_8 FILLER_32_1873 ();
 sg13g2_decap_4 FILLER_32_1880 ();
 sg13g2_fill_2 FILLER_32_1884 ();
 sg13g2_decap_8 FILLER_32_1906 ();
 sg13g2_decap_8 FILLER_32_1913 ();
 sg13g2_fill_1 FILLER_32_1920 ();
 sg13g2_fill_2 FILLER_32_1925 ();
 sg13g2_decap_8 FILLER_32_1932 ();
 sg13g2_decap_8 FILLER_32_1939 ();
 sg13g2_decap_8 FILLER_32_1993 ();
 sg13g2_decap_4 FILLER_32_2000 ();
 sg13g2_fill_2 FILLER_32_2004 ();
 sg13g2_decap_8 FILLER_32_2019 ();
 sg13g2_decap_8 FILLER_32_2026 ();
 sg13g2_decap_8 FILLER_32_2038 ();
 sg13g2_decap_8 FILLER_32_2094 ();
 sg13g2_decap_8 FILLER_32_2101 ();
 sg13g2_decap_8 FILLER_32_2108 ();
 sg13g2_decap_8 FILLER_32_2115 ();
 sg13g2_fill_2 FILLER_32_2122 ();
 sg13g2_fill_1 FILLER_32_2124 ();
 sg13g2_decap_4 FILLER_32_2131 ();
 sg13g2_fill_2 FILLER_32_2135 ();
 sg13g2_fill_1 FILLER_32_2160 ();
 sg13g2_fill_1 FILLER_32_2165 ();
 sg13g2_decap_8 FILLER_32_2184 ();
 sg13g2_decap_4 FILLER_32_2191 ();
 sg13g2_fill_2 FILLER_32_2195 ();
 sg13g2_fill_1 FILLER_32_2207 ();
 sg13g2_decap_8 FILLER_32_2213 ();
 sg13g2_decap_4 FILLER_32_2220 ();
 sg13g2_decap_8 FILLER_32_2232 ();
 sg13g2_fill_2 FILLER_32_2239 ();
 sg13g2_fill_1 FILLER_32_2241 ();
 sg13g2_fill_1 FILLER_32_2259 ();
 sg13g2_decap_8 FILLER_32_2264 ();
 sg13g2_fill_2 FILLER_32_2276 ();
 sg13g2_decap_8 FILLER_32_2286 ();
 sg13g2_fill_2 FILLER_32_2293 ();
 sg13g2_decap_8 FILLER_32_2334 ();
 sg13g2_decap_8 FILLER_32_2341 ();
 sg13g2_decap_8 FILLER_32_2348 ();
 sg13g2_fill_1 FILLER_32_2355 ();
 sg13g2_decap_8 FILLER_32_2369 ();
 sg13g2_fill_2 FILLER_32_2376 ();
 sg13g2_fill_2 FILLER_32_2396 ();
 sg13g2_fill_1 FILLER_32_2398 ();
 sg13g2_decap_4 FILLER_32_2414 ();
 sg13g2_fill_2 FILLER_32_2418 ();
 sg13g2_fill_2 FILLER_32_2440 ();
 sg13g2_fill_1 FILLER_32_2442 ();
 sg13g2_fill_1 FILLER_32_2448 ();
 sg13g2_fill_1 FILLER_32_2457 ();
 sg13g2_decap_8 FILLER_32_2463 ();
 sg13g2_decap_4 FILLER_32_2470 ();
 sg13g2_decap_8 FILLER_32_2489 ();
 sg13g2_decap_8 FILLER_32_2496 ();
 sg13g2_fill_1 FILLER_32_2503 ();
 sg13g2_fill_1 FILLER_32_2509 ();
 sg13g2_decap_4 FILLER_32_2515 ();
 sg13g2_decap_4 FILLER_32_2539 ();
 sg13g2_decap_4 FILLER_32_2547 ();
 sg13g2_decap_4 FILLER_32_2566 ();
 sg13g2_fill_1 FILLER_32_2570 ();
 sg13g2_decap_8 FILLER_32_2592 ();
 sg13g2_decap_8 FILLER_32_2599 ();
 sg13g2_decap_4 FILLER_32_2606 ();
 sg13g2_fill_1 FILLER_32_2610 ();
 sg13g2_decap_4 FILLER_32_2633 ();
 sg13g2_fill_2 FILLER_32_2637 ();
 sg13g2_fill_1 FILLER_32_2643 ();
 sg13g2_fill_1 FILLER_32_2652 ();
 sg13g2_fill_2 FILLER_32_2658 ();
 sg13g2_fill_1 FILLER_32_2660 ();
 sg13g2_fill_2 FILLER_32_2665 ();
 sg13g2_fill_2 FILLER_32_2682 ();
 sg13g2_fill_1 FILLER_32_2684 ();
 sg13g2_fill_1 FILLER_32_2690 ();
 sg13g2_decap_8 FILLER_32_2712 ();
 sg13g2_decap_4 FILLER_32_2719 ();
 sg13g2_fill_2 FILLER_32_2723 ();
 sg13g2_decap_8 FILLER_32_2782 ();
 sg13g2_decap_4 FILLER_32_2799 ();
 sg13g2_fill_1 FILLER_32_2814 ();
 sg13g2_decap_8 FILLER_32_2826 ();
 sg13g2_decap_8 FILLER_32_2833 ();
 sg13g2_fill_2 FILLER_32_2840 ();
 sg13g2_fill_1 FILLER_32_2842 ();
 sg13g2_decap_8 FILLER_32_2862 ();
 sg13g2_decap_4 FILLER_32_2869 ();
 sg13g2_fill_2 FILLER_32_2877 ();
 sg13g2_decap_4 FILLER_32_2883 ();
 sg13g2_fill_1 FILLER_32_2887 ();
 sg13g2_fill_2 FILLER_32_2892 ();
 sg13g2_decap_8 FILLER_32_2903 ();
 sg13g2_fill_2 FILLER_32_2910 ();
 sg13g2_decap_8 FILLER_32_2937 ();
 sg13g2_decap_8 FILLER_32_2967 ();
 sg13g2_fill_2 FILLER_32_2974 ();
 sg13g2_fill_1 FILLER_32_2976 ();
 sg13g2_decap_8 FILLER_32_2993 ();
 sg13g2_decap_4 FILLER_32_3000 ();
 sg13g2_fill_1 FILLER_32_3004 ();
 sg13g2_decap_8 FILLER_32_3014 ();
 sg13g2_decap_8 FILLER_32_3021 ();
 sg13g2_fill_2 FILLER_32_3091 ();
 sg13g2_fill_2 FILLER_32_3098 ();
 sg13g2_fill_2 FILLER_32_3113 ();
 sg13g2_fill_1 FILLER_32_3129 ();
 sg13g2_fill_2 FILLER_32_3148 ();
 sg13g2_fill_2 FILLER_32_3177 ();
 sg13g2_fill_2 FILLER_32_3189 ();
 sg13g2_decap_8 FILLER_32_3218 ();
 sg13g2_fill_1 FILLER_32_3225 ();
 sg13g2_decap_4 FILLER_32_3298 ();
 sg13g2_fill_2 FILLER_32_3302 ();
 sg13g2_decap_8 FILLER_32_3314 ();
 sg13g2_fill_2 FILLER_32_3321 ();
 sg13g2_fill_1 FILLER_32_3331 ();
 sg13g2_decap_4 FILLER_32_3345 ();
 sg13g2_fill_1 FILLER_32_3349 ();
 sg13g2_fill_2 FILLER_32_3360 ();
 sg13g2_fill_1 FILLER_32_3362 ();
 sg13g2_decap_8 FILLER_32_3391 ();
 sg13g2_decap_8 FILLER_32_3398 ();
 sg13g2_decap_8 FILLER_32_3405 ();
 sg13g2_decap_8 FILLER_32_3412 ();
 sg13g2_decap_8 FILLER_32_3419 ();
 sg13g2_decap_8 FILLER_32_3426 ();
 sg13g2_decap_8 FILLER_32_3433 ();
 sg13g2_decap_8 FILLER_32_3440 ();
 sg13g2_decap_8 FILLER_32_3447 ();
 sg13g2_decap_8 FILLER_32_3454 ();
 sg13g2_decap_8 FILLER_32_3461 ();
 sg13g2_decap_8 FILLER_32_3468 ();
 sg13g2_decap_8 FILLER_32_3475 ();
 sg13g2_decap_8 FILLER_32_3482 ();
 sg13g2_decap_8 FILLER_32_3489 ();
 sg13g2_decap_8 FILLER_32_3496 ();
 sg13g2_decap_8 FILLER_32_3503 ();
 sg13g2_decap_8 FILLER_32_3510 ();
 sg13g2_decap_8 FILLER_32_3517 ();
 sg13g2_decap_8 FILLER_32_3524 ();
 sg13g2_decap_8 FILLER_32_3531 ();
 sg13g2_decap_8 FILLER_32_3538 ();
 sg13g2_decap_8 FILLER_32_3545 ();
 sg13g2_decap_8 FILLER_32_3552 ();
 sg13g2_decap_8 FILLER_32_3559 ();
 sg13g2_decap_8 FILLER_32_3566 ();
 sg13g2_decap_8 FILLER_32_3573 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_4 FILLER_33_369 ();
 sg13g2_decap_4 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_fill_2 FILLER_33_417 ();
 sg13g2_fill_2 FILLER_33_430 ();
 sg13g2_fill_2 FILLER_33_445 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_fill_2 FILLER_33_487 ();
 sg13g2_decap_4 FILLER_33_502 ();
 sg13g2_fill_2 FILLER_33_506 ();
 sg13g2_fill_1 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_524 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_decap_4 FILLER_33_545 ();
 sg13g2_decap_8 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_562 ();
 sg13g2_decap_4 FILLER_33_572 ();
 sg13g2_fill_1 FILLER_33_576 ();
 sg13g2_decap_8 FILLER_33_593 ();
 sg13g2_decap_8 FILLER_33_600 ();
 sg13g2_fill_2 FILLER_33_615 ();
 sg13g2_decap_4 FILLER_33_636 ();
 sg13g2_fill_1 FILLER_33_640 ();
 sg13g2_decap_8 FILLER_33_652 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_decap_4 FILLER_33_682 ();
 sg13g2_fill_1 FILLER_33_686 ();
 sg13g2_decap_4 FILLER_33_701 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_738 ();
 sg13g2_decap_4 FILLER_33_745 ();
 sg13g2_fill_2 FILLER_33_749 ();
 sg13g2_fill_2 FILLER_33_756 ();
 sg13g2_decap_4 FILLER_33_780 ();
 sg13g2_fill_1 FILLER_33_784 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_801 ();
 sg13g2_fill_2 FILLER_33_808 ();
 sg13g2_decap_8 FILLER_33_815 ();
 sg13g2_decap_4 FILLER_33_827 ();
 sg13g2_fill_1 FILLER_33_831 ();
 sg13g2_fill_1 FILLER_33_857 ();
 sg13g2_decap_4 FILLER_33_881 ();
 sg13g2_fill_2 FILLER_33_903 ();
 sg13g2_decap_4 FILLER_33_918 ();
 sg13g2_fill_1 FILLER_33_922 ();
 sg13g2_fill_1 FILLER_33_961 ();
 sg13g2_decap_8 FILLER_33_1003 ();
 sg13g2_fill_1 FILLER_33_1010 ();
 sg13g2_fill_1 FILLER_33_1020 ();
 sg13g2_fill_2 FILLER_33_1034 ();
 sg13g2_fill_1 FILLER_33_1064 ();
 sg13g2_fill_1 FILLER_33_1093 ();
 sg13g2_decap_8 FILLER_33_1097 ();
 sg13g2_fill_1 FILLER_33_1104 ();
 sg13g2_fill_2 FILLER_33_1124 ();
 sg13g2_fill_2 FILLER_33_1129 ();
 sg13g2_fill_2 FILLER_33_1179 ();
 sg13g2_decap_4 FILLER_33_1190 ();
 sg13g2_fill_2 FILLER_33_1200 ();
 sg13g2_fill_1 FILLER_33_1202 ();
 sg13g2_decap_4 FILLER_33_1215 ();
 sg13g2_fill_1 FILLER_33_1219 ();
 sg13g2_fill_2 FILLER_33_1248 ();
 sg13g2_fill_1 FILLER_33_1250 ();
 sg13g2_fill_1 FILLER_33_1272 ();
 sg13g2_decap_8 FILLER_33_1289 ();
 sg13g2_fill_2 FILLER_33_1296 ();
 sg13g2_fill_1 FILLER_33_1397 ();
 sg13g2_decap_8 FILLER_33_1401 ();
 sg13g2_decap_8 FILLER_33_1408 ();
 sg13g2_fill_1 FILLER_33_1415 ();
 sg13g2_decap_4 FILLER_33_1423 ();
 sg13g2_fill_2 FILLER_33_1427 ();
 sg13g2_fill_1 FILLER_33_1449 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_4 FILLER_33_1519 ();
 sg13g2_decap_4 FILLER_33_1532 ();
 sg13g2_fill_1 FILLER_33_1536 ();
 sg13g2_fill_1 FILLER_33_1565 ();
 sg13g2_fill_1 FILLER_33_1570 ();
 sg13g2_fill_2 FILLER_33_1595 ();
 sg13g2_fill_2 FILLER_33_1625 ();
 sg13g2_decap_8 FILLER_33_1635 ();
 sg13g2_decap_4 FILLER_33_1642 ();
 sg13g2_fill_2 FILLER_33_1646 ();
 sg13g2_fill_1 FILLER_33_1666 ();
 sg13g2_decap_4 FILLER_33_1675 ();
 sg13g2_fill_1 FILLER_33_1679 ();
 sg13g2_decap_8 FILLER_33_1684 ();
 sg13g2_fill_2 FILLER_33_1691 ();
 sg13g2_fill_1 FILLER_33_1693 ();
 sg13g2_fill_2 FILLER_33_1719 ();
 sg13g2_fill_1 FILLER_33_1721 ();
 sg13g2_fill_1 FILLER_33_1735 ();
 sg13g2_decap_8 FILLER_33_1739 ();
 sg13g2_decap_8 FILLER_33_1746 ();
 sg13g2_fill_2 FILLER_33_1753 ();
 sg13g2_decap_8 FILLER_33_1769 ();
 sg13g2_decap_8 FILLER_33_1776 ();
 sg13g2_decap_4 FILLER_33_1783 ();
 sg13g2_fill_1 FILLER_33_1787 ();
 sg13g2_fill_2 FILLER_33_1816 ();
 sg13g2_decap_8 FILLER_33_1834 ();
 sg13g2_fill_1 FILLER_33_1841 ();
 sg13g2_decap_4 FILLER_33_1847 ();
 sg13g2_decap_8 FILLER_33_1859 ();
 sg13g2_decap_4 FILLER_33_1866 ();
 sg13g2_fill_1 FILLER_33_1870 ();
 sg13g2_decap_8 FILLER_33_1887 ();
 sg13g2_fill_2 FILLER_33_1894 ();
 sg13g2_fill_1 FILLER_33_1896 ();
 sg13g2_decap_4 FILLER_33_1906 ();
 sg13g2_fill_1 FILLER_33_1910 ();
 sg13g2_fill_2 FILLER_33_1924 ();
 sg13g2_decap_8 FILLER_33_1938 ();
 sg13g2_decap_8 FILLER_33_1961 ();
 sg13g2_fill_1 FILLER_33_1968 ();
 sg13g2_fill_2 FILLER_33_1977 ();
 sg13g2_fill_1 FILLER_33_1979 ();
 sg13g2_decap_8 FILLER_33_1986 ();
 sg13g2_fill_2 FILLER_33_1993 ();
 sg13g2_fill_1 FILLER_33_2008 ();
 sg13g2_decap_4 FILLER_33_2021 ();
 sg13g2_fill_1 FILLER_33_2037 ();
 sg13g2_decap_4 FILLER_33_2059 ();
 sg13g2_decap_4 FILLER_33_2111 ();
 sg13g2_fill_1 FILLER_33_2115 ();
 sg13g2_decap_4 FILLER_33_2120 ();
 sg13g2_fill_2 FILLER_33_2124 ();
 sg13g2_decap_4 FILLER_33_2131 ();
 sg13g2_fill_1 FILLER_33_2135 ();
 sg13g2_decap_4 FILLER_33_2157 ();
 sg13g2_fill_2 FILLER_33_2166 ();
 sg13g2_fill_1 FILLER_33_2168 ();
 sg13g2_decap_8 FILLER_33_2188 ();
 sg13g2_fill_2 FILLER_33_2195 ();
 sg13g2_fill_1 FILLER_33_2197 ();
 sg13g2_fill_1 FILLER_33_2211 ();
 sg13g2_fill_2 FILLER_33_2224 ();
 sg13g2_fill_1 FILLER_33_2226 ();
 sg13g2_decap_8 FILLER_33_2239 ();
 sg13g2_fill_2 FILLER_33_2246 ();
 sg13g2_fill_1 FILLER_33_2248 ();
 sg13g2_decap_8 FILLER_33_2253 ();
 sg13g2_fill_2 FILLER_33_2270 ();
 sg13g2_fill_1 FILLER_33_2272 ();
 sg13g2_decap_4 FILLER_33_2301 ();
 sg13g2_fill_1 FILLER_33_2309 ();
 sg13g2_decap_4 FILLER_33_2315 ();
 sg13g2_fill_1 FILLER_33_2319 ();
 sg13g2_fill_2 FILLER_33_2352 ();
 sg13g2_decap_8 FILLER_33_2364 ();
 sg13g2_fill_2 FILLER_33_2371 ();
 sg13g2_fill_1 FILLER_33_2373 ();
 sg13g2_fill_2 FILLER_33_2392 ();
 sg13g2_fill_1 FILLER_33_2394 ();
 sg13g2_decap_8 FILLER_33_2405 ();
 sg13g2_decap_8 FILLER_33_2412 ();
 sg13g2_decap_4 FILLER_33_2419 ();
 sg13g2_fill_2 FILLER_33_2448 ();
 sg13g2_decap_4 FILLER_33_2468 ();
 sg13g2_fill_2 FILLER_33_2472 ();
 sg13g2_decap_4 FILLER_33_2496 ();
 sg13g2_fill_1 FILLER_33_2500 ();
 sg13g2_decap_4 FILLER_33_2543 ();
 sg13g2_fill_2 FILLER_33_2547 ();
 sg13g2_decap_8 FILLER_33_2567 ();
 sg13g2_decap_4 FILLER_33_2574 ();
 sg13g2_fill_2 FILLER_33_2578 ();
 sg13g2_decap_4 FILLER_33_2588 ();
 sg13g2_fill_2 FILLER_33_2592 ();
 sg13g2_decap_4 FILLER_33_2600 ();
 sg13g2_fill_1 FILLER_33_2604 ();
 sg13g2_decap_4 FILLER_33_2629 ();
 sg13g2_fill_1 FILLER_33_2633 ();
 sg13g2_decap_4 FILLER_33_2659 ();
 sg13g2_fill_2 FILLER_33_2663 ();
 sg13g2_fill_2 FILLER_33_2670 ();
 sg13g2_fill_2 FILLER_33_2684 ();
 sg13g2_fill_2 FILLER_33_2692 ();
 sg13g2_decap_8 FILLER_33_2711 ();
 sg13g2_decap_8 FILLER_33_2718 ();
 sg13g2_decap_4 FILLER_33_2725 ();
 sg13g2_fill_2 FILLER_33_2729 ();
 sg13g2_fill_2 FILLER_33_2736 ();
 sg13g2_fill_1 FILLER_33_2738 ();
 sg13g2_decap_8 FILLER_33_2744 ();
 sg13g2_fill_2 FILLER_33_2751 ();
 sg13g2_decap_8 FILLER_33_2778 ();
 sg13g2_decap_4 FILLER_33_2801 ();
 sg13g2_fill_1 FILLER_33_2805 ();
 sg13g2_decap_4 FILLER_33_2831 ();
 sg13g2_fill_1 FILLER_33_2835 ();
 sg13g2_fill_1 FILLER_33_2844 ();
 sg13g2_decap_4 FILLER_33_2867 ();
 sg13g2_fill_2 FILLER_33_2884 ();
 sg13g2_decap_8 FILLER_33_2902 ();
 sg13g2_decap_4 FILLER_33_2909 ();
 sg13g2_fill_1 FILLER_33_2925 ();
 sg13g2_decap_8 FILLER_33_2934 ();
 sg13g2_fill_2 FILLER_33_2941 ();
 sg13g2_decap_8 FILLER_33_2970 ();
 sg13g2_fill_2 FILLER_33_2977 ();
 sg13g2_fill_1 FILLER_33_2984 ();
 sg13g2_fill_2 FILLER_33_2997 ();
 sg13g2_fill_1 FILLER_33_2999 ();
 sg13g2_fill_1 FILLER_33_3023 ();
 sg13g2_decap_8 FILLER_33_3029 ();
 sg13g2_decap_8 FILLER_33_3036 ();
 sg13g2_decap_4 FILLER_33_3043 ();
 sg13g2_fill_1 FILLER_33_3047 ();
 sg13g2_decap_8 FILLER_33_3063 ();
 sg13g2_decap_8 FILLER_33_3070 ();
 sg13g2_fill_1 FILLER_33_3118 ();
 sg13g2_fill_1 FILLER_33_3134 ();
 sg13g2_fill_2 FILLER_33_3162 ();
 sg13g2_fill_1 FILLER_33_3164 ();
 sg13g2_fill_1 FILLER_33_3192 ();
 sg13g2_fill_2 FILLER_33_3212 ();
 sg13g2_decap_4 FILLER_33_3223 ();
 sg13g2_fill_1 FILLER_33_3227 ();
 sg13g2_fill_2 FILLER_33_3251 ();
 sg13g2_decap_4 FILLER_33_3262 ();
 sg13g2_fill_1 FILLER_33_3285 ();
 sg13g2_decap_8 FILLER_33_3307 ();
 sg13g2_decap_4 FILLER_33_3314 ();
 sg13g2_decap_8 FILLER_33_3338 ();
 sg13g2_decap_8 FILLER_33_3376 ();
 sg13g2_decap_8 FILLER_33_3383 ();
 sg13g2_decap_8 FILLER_33_3390 ();
 sg13g2_decap_8 FILLER_33_3397 ();
 sg13g2_decap_8 FILLER_33_3404 ();
 sg13g2_decap_8 FILLER_33_3411 ();
 sg13g2_decap_8 FILLER_33_3418 ();
 sg13g2_decap_8 FILLER_33_3425 ();
 sg13g2_decap_8 FILLER_33_3432 ();
 sg13g2_decap_8 FILLER_33_3439 ();
 sg13g2_decap_8 FILLER_33_3446 ();
 sg13g2_decap_8 FILLER_33_3453 ();
 sg13g2_decap_8 FILLER_33_3460 ();
 sg13g2_decap_8 FILLER_33_3467 ();
 sg13g2_decap_8 FILLER_33_3474 ();
 sg13g2_decap_8 FILLER_33_3481 ();
 sg13g2_decap_8 FILLER_33_3488 ();
 sg13g2_decap_8 FILLER_33_3495 ();
 sg13g2_decap_8 FILLER_33_3502 ();
 sg13g2_decap_8 FILLER_33_3509 ();
 sg13g2_decap_8 FILLER_33_3516 ();
 sg13g2_decap_8 FILLER_33_3523 ();
 sg13g2_decap_8 FILLER_33_3530 ();
 sg13g2_decap_8 FILLER_33_3537 ();
 sg13g2_decap_8 FILLER_33_3544 ();
 sg13g2_decap_8 FILLER_33_3551 ();
 sg13g2_decap_8 FILLER_33_3558 ();
 sg13g2_decap_8 FILLER_33_3565 ();
 sg13g2_decap_8 FILLER_33_3572 ();
 sg13g2_fill_1 FILLER_33_3579 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_4 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_262 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_34_445 ();
 sg13g2_decap_8 FILLER_34_452 ();
 sg13g2_fill_2 FILLER_34_459 ();
 sg13g2_fill_2 FILLER_34_474 ();
 sg13g2_fill_1 FILLER_34_488 ();
 sg13g2_fill_2 FILLER_34_507 ();
 sg13g2_fill_1 FILLER_34_509 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_527 ();
 sg13g2_fill_2 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_536 ();
 sg13g2_decap_4 FILLER_34_541 ();
 sg13g2_fill_1 FILLER_34_545 ();
 sg13g2_fill_1 FILLER_34_593 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_decap_4 FILLER_34_625 ();
 sg13g2_fill_1 FILLER_34_629 ();
 sg13g2_decap_4 FILLER_34_644 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_decap_4 FILLER_34_661 ();
 sg13g2_fill_1 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_decap_4 FILLER_34_676 ();
 sg13g2_fill_2 FILLER_34_698 ();
 sg13g2_fill_1 FILLER_34_700 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_731 ();
 sg13g2_decap_8 FILLER_34_738 ();
 sg13g2_fill_1 FILLER_34_758 ();
 sg13g2_fill_2 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_4 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_fill_2 FILLER_34_813 ();
 sg13g2_decap_4 FILLER_34_835 ();
 sg13g2_decap_8 FILLER_34_869 ();
 sg13g2_decap_8 FILLER_34_876 ();
 sg13g2_decap_8 FILLER_34_883 ();
 sg13g2_fill_2 FILLER_34_890 ();
 sg13g2_fill_1 FILLER_34_892 ();
 sg13g2_fill_2 FILLER_34_898 ();
 sg13g2_fill_1 FILLER_34_900 ();
 sg13g2_decap_4 FILLER_34_917 ();
 sg13g2_fill_1 FILLER_34_921 ();
 sg13g2_decap_8 FILLER_34_934 ();
 sg13g2_fill_2 FILLER_34_941 ();
 sg13g2_fill_1 FILLER_34_943 ();
 sg13g2_decap_8 FILLER_34_957 ();
 sg13g2_decap_4 FILLER_34_964 ();
 sg13g2_fill_1 FILLER_34_968 ();
 sg13g2_decap_4 FILLER_34_975 ();
 sg13g2_fill_1 FILLER_34_979 ();
 sg13g2_fill_2 FILLER_34_984 ();
 sg13g2_decap_4 FILLER_34_1011 ();
 sg13g2_fill_1 FILLER_34_1015 ();
 sg13g2_decap_4 FILLER_34_1065 ();
 sg13g2_fill_1 FILLER_34_1069 ();
 sg13g2_decap_4 FILLER_34_1083 ();
 sg13g2_fill_1 FILLER_34_1087 ();
 sg13g2_decap_4 FILLER_34_1116 ();
 sg13g2_decap_4 FILLER_34_1146 ();
 sg13g2_decap_8 FILLER_34_1178 ();
 sg13g2_fill_2 FILLER_34_1185 ();
 sg13g2_decap_8 FILLER_34_1203 ();
 sg13g2_fill_1 FILLER_34_1210 ();
 sg13g2_decap_8 FILLER_34_1221 ();
 sg13g2_fill_2 FILLER_34_1228 ();
 sg13g2_decap_4 FILLER_34_1267 ();
 sg13g2_decap_4 FILLER_34_1287 ();
 sg13g2_fill_1 FILLER_34_1291 ();
 sg13g2_decap_4 FILLER_34_1317 ();
 sg13g2_fill_2 FILLER_34_1334 ();
 sg13g2_fill_1 FILLER_34_1336 ();
 sg13g2_fill_2 FILLER_34_1365 ();
 sg13g2_fill_1 FILLER_34_1367 ();
 sg13g2_decap_4 FILLER_34_1372 ();
 sg13g2_fill_2 FILLER_34_1376 ();
 sg13g2_fill_2 FILLER_34_1383 ();
 sg13g2_fill_1 FILLER_34_1453 ();
 sg13g2_decap_8 FILLER_34_1473 ();
 sg13g2_fill_1 FILLER_34_1488 ();
 sg13g2_decap_8 FILLER_34_1493 ();
 sg13g2_fill_2 FILLER_34_1500 ();
 sg13g2_fill_1 FILLER_34_1502 ();
 sg13g2_decap_4 FILLER_34_1513 ();
 sg13g2_fill_2 FILLER_34_1517 ();
 sg13g2_fill_1 FILLER_34_1535 ();
 sg13g2_decap_4 FILLER_34_1542 ();
 sg13g2_fill_1 FILLER_34_1546 ();
 sg13g2_fill_2 FILLER_34_1552 ();
 sg13g2_fill_2 FILLER_34_1561 ();
 sg13g2_fill_1 FILLER_34_1563 ();
 sg13g2_fill_2 FILLER_34_1568 ();
 sg13g2_fill_2 FILLER_34_1620 ();
 sg13g2_decap_8 FILLER_34_1640 ();
 sg13g2_decap_4 FILLER_34_1647 ();
 sg13g2_fill_2 FILLER_34_1651 ();
 sg13g2_fill_2 FILLER_34_1665 ();
 sg13g2_fill_1 FILLER_34_1667 ();
 sg13g2_decap_8 FILLER_34_1680 ();
 sg13g2_fill_2 FILLER_34_1687 ();
 sg13g2_fill_1 FILLER_34_1689 ();
 sg13g2_decap_8 FILLER_34_1695 ();
 sg13g2_fill_1 FILLER_34_1702 ();
 sg13g2_decap_8 FILLER_34_1713 ();
 sg13g2_decap_4 FILLER_34_1720 ();
 sg13g2_fill_2 FILLER_34_1747 ();
 sg13g2_fill_1 FILLER_34_1749 ();
 sg13g2_decap_4 FILLER_34_1761 ();
 sg13g2_fill_2 FILLER_34_1773 ();
 sg13g2_decap_8 FILLER_34_1783 ();
 sg13g2_decap_8 FILLER_34_1807 ();
 sg13g2_decap_4 FILLER_34_1814 ();
 sg13g2_fill_1 FILLER_34_1827 ();
 sg13g2_decap_8 FILLER_34_1832 ();
 sg13g2_fill_2 FILLER_34_1839 ();
 sg13g2_fill_1 FILLER_34_1841 ();
 sg13g2_fill_1 FILLER_34_1847 ();
 sg13g2_decap_8 FILLER_34_1867 ();
 sg13g2_fill_2 FILLER_34_1874 ();
 sg13g2_fill_1 FILLER_34_1876 ();
 sg13g2_decap_4 FILLER_34_1898 ();
 sg13g2_fill_2 FILLER_34_1902 ();
 sg13g2_decap_4 FILLER_34_1912 ();
 sg13g2_fill_2 FILLER_34_1916 ();
 sg13g2_fill_2 FILLER_34_1921 ();
 sg13g2_decap_4 FILLER_34_1927 ();
 sg13g2_fill_2 FILLER_34_1931 ();
 sg13g2_decap_4 FILLER_34_1945 ();
 sg13g2_fill_2 FILLER_34_1949 ();
 sg13g2_decap_8 FILLER_34_1957 ();
 sg13g2_decap_8 FILLER_34_1964 ();
 sg13g2_fill_2 FILLER_34_1990 ();
 sg13g2_fill_1 FILLER_34_1992 ();
 sg13g2_fill_1 FILLER_34_2008 ();
 sg13g2_decap_4 FILLER_34_2014 ();
 sg13g2_fill_2 FILLER_34_2022 ();
 sg13g2_decap_4 FILLER_34_2036 ();
 sg13g2_fill_2 FILLER_34_2040 ();
 sg13g2_fill_1 FILLER_34_2046 ();
 sg13g2_fill_2 FILLER_34_2052 ();
 sg13g2_fill_1 FILLER_34_2054 ();
 sg13g2_decap_8 FILLER_34_2060 ();
 sg13g2_decap_4 FILLER_34_2067 ();
 sg13g2_fill_2 FILLER_34_2071 ();
 sg13g2_fill_1 FILLER_34_2077 ();
 sg13g2_fill_1 FILLER_34_2091 ();
 sg13g2_fill_2 FILLER_34_2105 ();
 sg13g2_fill_1 FILLER_34_2113 ();
 sg13g2_decap_8 FILLER_34_2155 ();
 sg13g2_decap_8 FILLER_34_2162 ();
 sg13g2_fill_1 FILLER_34_2174 ();
 sg13g2_decap_8 FILLER_34_2184 ();
 sg13g2_decap_4 FILLER_34_2191 ();
 sg13g2_fill_1 FILLER_34_2195 ();
 sg13g2_decap_8 FILLER_34_2212 ();
 sg13g2_decap_4 FILLER_34_2219 ();
 sg13g2_fill_2 FILLER_34_2223 ();
 sg13g2_decap_8 FILLER_34_2230 ();
 sg13g2_fill_1 FILLER_34_2237 ();
 sg13g2_fill_1 FILLER_34_2246 ();
 sg13g2_decap_8 FILLER_34_2282 ();
 sg13g2_decap_8 FILLER_34_2289 ();
 sg13g2_decap_8 FILLER_34_2296 ();
 sg13g2_fill_2 FILLER_34_2303 ();
 sg13g2_fill_2 FILLER_34_2310 ();
 sg13g2_fill_1 FILLER_34_2312 ();
 sg13g2_fill_1 FILLER_34_2330 ();
 sg13g2_decap_4 FILLER_34_2341 ();
 sg13g2_fill_1 FILLER_34_2353 ();
 sg13g2_decap_8 FILLER_34_2364 ();
 sg13g2_decap_8 FILLER_34_2371 ();
 sg13g2_fill_2 FILLER_34_2378 ();
 sg13g2_decap_8 FILLER_34_2389 ();
 sg13g2_fill_2 FILLER_34_2396 ();
 sg13g2_fill_1 FILLER_34_2398 ();
 sg13g2_decap_8 FILLER_34_2413 ();
 sg13g2_decap_8 FILLER_34_2420 ();
 sg13g2_decap_8 FILLER_34_2427 ();
 sg13g2_fill_1 FILLER_34_2434 ();
 sg13g2_fill_1 FILLER_34_2440 ();
 sg13g2_fill_2 FILLER_34_2451 ();
 sg13g2_fill_1 FILLER_34_2453 ();
 sg13g2_decap_8 FILLER_34_2468 ();
 sg13g2_fill_2 FILLER_34_2475 ();
 sg13g2_fill_2 FILLER_34_2483 ();
 sg13g2_fill_1 FILLER_34_2485 ();
 sg13g2_fill_2 FILLER_34_2491 ();
 sg13g2_decap_4 FILLER_34_2501 ();
 sg13g2_fill_1 FILLER_34_2505 ();
 sg13g2_decap_8 FILLER_34_2510 ();
 sg13g2_decap_8 FILLER_34_2517 ();
 sg13g2_decap_8 FILLER_34_2524 ();
 sg13g2_decap_8 FILLER_34_2531 ();
 sg13g2_fill_1 FILLER_34_2538 ();
 sg13g2_decap_8 FILLER_34_2566 ();
 sg13g2_fill_2 FILLER_34_2573 ();
 sg13g2_decap_8 FILLER_34_2593 ();
 sg13g2_decap_8 FILLER_34_2600 ();
 sg13g2_decap_4 FILLER_34_2607 ();
 sg13g2_fill_1 FILLER_34_2611 ();
 sg13g2_decap_4 FILLER_34_2624 ();
 sg13g2_fill_2 FILLER_34_2628 ();
 sg13g2_fill_1 FILLER_34_2642 ();
 sg13g2_decap_8 FILLER_34_2648 ();
 sg13g2_fill_2 FILLER_34_2655 ();
 sg13g2_fill_1 FILLER_34_2657 ();
 sg13g2_fill_1 FILLER_34_2663 ();
 sg13g2_decap_8 FILLER_34_2677 ();
 sg13g2_decap_8 FILLER_34_2684 ();
 sg13g2_fill_2 FILLER_34_2691 ();
 sg13g2_fill_2 FILLER_34_2701 ();
 sg13g2_fill_1 FILLER_34_2703 ();
 sg13g2_decap_8 FILLER_34_2717 ();
 sg13g2_decap_4 FILLER_34_2724 ();
 sg13g2_fill_1 FILLER_34_2728 ();
 sg13g2_decap_4 FILLER_34_2742 ();
 sg13g2_fill_1 FILLER_34_2763 ();
 sg13g2_decap_8 FILLER_34_2768 ();
 sg13g2_decap_8 FILLER_34_2775 ();
 sg13g2_decap_4 FILLER_34_2782 ();
 sg13g2_fill_1 FILLER_34_2786 ();
 sg13g2_decap_4 FILLER_34_2798 ();
 sg13g2_fill_2 FILLER_34_2802 ();
 sg13g2_fill_2 FILLER_34_2808 ();
 sg13g2_decap_8 FILLER_34_2826 ();
 sg13g2_fill_2 FILLER_34_2833 ();
 sg13g2_fill_1 FILLER_34_2835 ();
 sg13g2_decap_4 FILLER_34_2871 ();
 sg13g2_fill_2 FILLER_34_2875 ();
 sg13g2_fill_1 FILLER_34_2885 ();
 sg13g2_fill_2 FILLER_34_2902 ();
 sg13g2_fill_1 FILLER_34_2904 ();
 sg13g2_decap_8 FILLER_34_2931 ();
 sg13g2_fill_1 FILLER_34_2938 ();
 sg13g2_decap_8 FILLER_34_2964 ();
 sg13g2_fill_2 FILLER_34_2971 ();
 sg13g2_fill_1 FILLER_34_3009 ();
 sg13g2_fill_2 FILLER_34_3016 ();
 sg13g2_fill_1 FILLER_34_3018 ();
 sg13g2_fill_2 FILLER_34_3060 ();
 sg13g2_fill_1 FILLER_34_3062 ();
 sg13g2_fill_1 FILLER_34_3090 ();
 sg13g2_fill_2 FILLER_34_3104 ();
 sg13g2_fill_1 FILLER_34_3106 ();
 sg13g2_fill_1 FILLER_34_3112 ();
 sg13g2_fill_2 FILLER_34_3123 ();
 sg13g2_fill_1 FILLER_34_3125 ();
 sg13g2_fill_1 FILLER_34_3148 ();
 sg13g2_decap_8 FILLER_34_3185 ();
 sg13g2_fill_2 FILLER_34_3202 ();
 sg13g2_fill_1 FILLER_34_3204 ();
 sg13g2_decap_8 FILLER_34_3232 ();
 sg13g2_decap_4 FILLER_34_3287 ();
 sg13g2_decap_4 FILLER_34_3314 ();
 sg13g2_fill_1 FILLER_34_3318 ();
 sg13g2_fill_1 FILLER_34_3344 ();
 sg13g2_fill_2 FILLER_34_3357 ();
 sg13g2_decap_4 FILLER_34_3372 ();
 sg13g2_fill_2 FILLER_34_3376 ();
 sg13g2_decap_8 FILLER_34_3384 ();
 sg13g2_decap_8 FILLER_34_3391 ();
 sg13g2_decap_8 FILLER_34_3398 ();
 sg13g2_fill_1 FILLER_34_3405 ();
 sg13g2_decap_8 FILLER_34_3410 ();
 sg13g2_decap_8 FILLER_34_3417 ();
 sg13g2_decap_8 FILLER_34_3424 ();
 sg13g2_decap_8 FILLER_34_3431 ();
 sg13g2_decap_8 FILLER_34_3438 ();
 sg13g2_decap_8 FILLER_34_3445 ();
 sg13g2_decap_8 FILLER_34_3452 ();
 sg13g2_decap_8 FILLER_34_3459 ();
 sg13g2_decap_8 FILLER_34_3466 ();
 sg13g2_decap_8 FILLER_34_3473 ();
 sg13g2_decap_8 FILLER_34_3480 ();
 sg13g2_decap_8 FILLER_34_3487 ();
 sg13g2_decap_8 FILLER_34_3494 ();
 sg13g2_decap_8 FILLER_34_3501 ();
 sg13g2_decap_8 FILLER_34_3508 ();
 sg13g2_decap_8 FILLER_34_3515 ();
 sg13g2_decap_8 FILLER_34_3522 ();
 sg13g2_decap_8 FILLER_34_3529 ();
 sg13g2_decap_8 FILLER_34_3536 ();
 sg13g2_decap_8 FILLER_34_3543 ();
 sg13g2_decap_8 FILLER_34_3550 ();
 sg13g2_decap_8 FILLER_34_3557 ();
 sg13g2_decap_8 FILLER_34_3564 ();
 sg13g2_decap_8 FILLER_34_3571 ();
 sg13g2_fill_2 FILLER_34_3578 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_430 ();
 sg13g2_fill_1 FILLER_35_461 ();
 sg13g2_decap_8 FILLER_35_550 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_8 FILLER_35_568 ();
 sg13g2_decap_8 FILLER_35_575 ();
 sg13g2_decap_8 FILLER_35_589 ();
 sg13g2_fill_2 FILLER_35_596 ();
 sg13g2_fill_1 FILLER_35_598 ();
 sg13g2_decap_4 FILLER_35_629 ();
 sg13g2_fill_2 FILLER_35_656 ();
 sg13g2_decap_4 FILLER_35_668 ();
 sg13g2_fill_2 FILLER_35_685 ();
 sg13g2_fill_2 FILLER_35_702 ();
 sg13g2_fill_2 FILLER_35_717 ();
 sg13g2_fill_2 FILLER_35_727 ();
 sg13g2_decap_8 FILLER_35_737 ();
 sg13g2_fill_2 FILLER_35_744 ();
 sg13g2_fill_1 FILLER_35_746 ();
 sg13g2_fill_1 FILLER_35_755 ();
 sg13g2_decap_4 FILLER_35_768 ();
 sg13g2_decap_8 FILLER_35_775 ();
 sg13g2_fill_2 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_fill_1 FILLER_35_826 ();
 sg13g2_decap_4 FILLER_35_840 ();
 sg13g2_fill_1 FILLER_35_844 ();
 sg13g2_fill_2 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_35_874 ();
 sg13g2_fill_2 FILLER_35_881 ();
 sg13g2_decap_8 FILLER_35_915 ();
 sg13g2_decap_4 FILLER_35_922 ();
 sg13g2_fill_2 FILLER_35_935 ();
 sg13g2_fill_1 FILLER_35_937 ();
 sg13g2_fill_2 FILLER_35_959 ();
 sg13g2_decap_4 FILLER_35_992 ();
 sg13g2_fill_1 FILLER_35_1041 ();
 sg13g2_fill_1 FILLER_35_1046 ();
 sg13g2_decap_8 FILLER_35_1060 ();
 sg13g2_fill_2 FILLER_35_1072 ();
 sg13g2_fill_1 FILLER_35_1074 ();
 sg13g2_fill_2 FILLER_35_1088 ();
 sg13g2_fill_2 FILLER_35_1107 ();
 sg13g2_fill_1 FILLER_35_1109 ();
 sg13g2_fill_2 FILLER_35_1114 ();
 sg13g2_fill_1 FILLER_35_1116 ();
 sg13g2_fill_1 FILLER_35_1144 ();
 sg13g2_decap_4 FILLER_35_1150 ();
 sg13g2_fill_1 FILLER_35_1154 ();
 sg13g2_decap_4 FILLER_35_1159 ();
 sg13g2_fill_2 FILLER_35_1163 ();
 sg13g2_decap_8 FILLER_35_1170 ();
 sg13g2_decap_4 FILLER_35_1177 ();
 sg13g2_fill_2 FILLER_35_1181 ();
 sg13g2_fill_2 FILLER_35_1223 ();
 sg13g2_decap_8 FILLER_35_1229 ();
 sg13g2_decap_8 FILLER_35_1236 ();
 sg13g2_fill_1 FILLER_35_1243 ();
 sg13g2_decap_8 FILLER_35_1248 ();
 sg13g2_decap_8 FILLER_35_1255 ();
 sg13g2_decap_4 FILLER_35_1262 ();
 sg13g2_decap_8 FILLER_35_1279 ();
 sg13g2_fill_2 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1322 ();
 sg13g2_fill_1 FILLER_35_1329 ();
 sg13g2_decap_8 FILLER_35_1335 ();
 sg13g2_decap_4 FILLER_35_1346 ();
 sg13g2_fill_1 FILLER_35_1350 ();
 sg13g2_decap_8 FILLER_35_1368 ();
 sg13g2_decap_4 FILLER_35_1380 ();
 sg13g2_fill_1 FILLER_35_1384 ();
 sg13g2_decap_8 FILLER_35_1401 ();
 sg13g2_decap_8 FILLER_35_1408 ();
 sg13g2_decap_8 FILLER_35_1415 ();
 sg13g2_decap_4 FILLER_35_1422 ();
 sg13g2_decap_4 FILLER_35_1442 ();
 sg13g2_decap_8 FILLER_35_1464 ();
 sg13g2_decap_4 FILLER_35_1471 ();
 sg13g2_decap_4 FILLER_35_1492 ();
 sg13g2_fill_2 FILLER_35_1523 ();
 sg13g2_decap_8 FILLER_35_1534 ();
 sg13g2_decap_4 FILLER_35_1541 ();
 sg13g2_fill_2 FILLER_35_1549 ();
 sg13g2_fill_2 FILLER_35_1577 ();
 sg13g2_decap_4 FILLER_35_1608 ();
 sg13g2_fill_2 FILLER_35_1620 ();
 sg13g2_decap_8 FILLER_35_1639 ();
 sg13g2_fill_1 FILLER_35_1646 ();
 sg13g2_fill_1 FILLER_35_1681 ();
 sg13g2_decap_4 FILLER_35_1702 ();
 sg13g2_decap_8 FILLER_35_1719 ();
 sg13g2_decap_8 FILLER_35_1787 ();
 sg13g2_decap_8 FILLER_35_1794 ();
 sg13g2_decap_4 FILLER_35_1801 ();
 sg13g2_fill_1 FILLER_35_1805 ();
 sg13g2_fill_2 FILLER_35_1811 ();
 sg13g2_fill_2 FILLER_35_1821 ();
 sg13g2_fill_1 FILLER_35_1823 ();
 sg13g2_fill_1 FILLER_35_1836 ();
 sg13g2_decap_4 FILLER_35_1857 ();
 sg13g2_fill_2 FILLER_35_1861 ();
 sg13g2_decap_4 FILLER_35_1882 ();
 sg13g2_fill_1 FILLER_35_1892 ();
 sg13g2_fill_2 FILLER_35_1898 ();
 sg13g2_fill_1 FILLER_35_1900 ();
 sg13g2_decap_4 FILLER_35_1921 ();
 sg13g2_fill_1 FILLER_35_1925 ();
 sg13g2_decap_8 FILLER_35_1931 ();
 sg13g2_fill_2 FILLER_35_1944 ();
 sg13g2_decap_8 FILLER_35_1966 ();
 sg13g2_fill_2 FILLER_35_1973 ();
 sg13g2_fill_1 FILLER_35_1987 ();
 sg13g2_fill_2 FILLER_35_1998 ();
 sg13g2_decap_8 FILLER_35_2006 ();
 sg13g2_decap_4 FILLER_35_2013 ();
 sg13g2_fill_1 FILLER_35_2017 ();
 sg13g2_decap_4 FILLER_35_2032 ();
 sg13g2_fill_2 FILLER_35_2036 ();
 sg13g2_fill_2 FILLER_35_2055 ();
 sg13g2_fill_1 FILLER_35_2057 ();
 sg13g2_fill_2 FILLER_35_2063 ();
 sg13g2_fill_1 FILLER_35_2078 ();
 sg13g2_fill_1 FILLER_35_2117 ();
 sg13g2_fill_2 FILLER_35_2131 ();
 sg13g2_fill_1 FILLER_35_2133 ();
 sg13g2_decap_4 FILLER_35_2140 ();
 sg13g2_decap_8 FILLER_35_2152 ();
 sg13g2_fill_2 FILLER_35_2159 ();
 sg13g2_fill_1 FILLER_35_2161 ();
 sg13g2_fill_1 FILLER_35_2199 ();
 sg13g2_fill_2 FILLER_35_2218 ();
 sg13g2_fill_1 FILLER_35_2220 ();
 sg13g2_decap_4 FILLER_35_2242 ();
 sg13g2_fill_2 FILLER_35_2246 ();
 sg13g2_decap_8 FILLER_35_2254 ();
 sg13g2_fill_2 FILLER_35_2261 ();
 sg13g2_fill_1 FILLER_35_2263 ();
 sg13g2_fill_1 FILLER_35_2280 ();
 sg13g2_decap_4 FILLER_35_2301 ();
 sg13g2_decap_4 FILLER_35_2313 ();
 sg13g2_fill_1 FILLER_35_2317 ();
 sg13g2_decap_8 FILLER_35_2339 ();
 sg13g2_decap_8 FILLER_35_2346 ();
 sg13g2_fill_2 FILLER_35_2353 ();
 sg13g2_decap_4 FILLER_35_2397 ();
 sg13g2_decap_4 FILLER_35_2422 ();
 sg13g2_fill_2 FILLER_35_2426 ();
 sg13g2_decap_8 FILLER_35_2446 ();
 sg13g2_decap_4 FILLER_35_2453 ();
 sg13g2_fill_2 FILLER_35_2467 ();
 sg13g2_decap_8 FILLER_35_2477 ();
 sg13g2_fill_1 FILLER_35_2484 ();
 sg13g2_fill_2 FILLER_35_2523 ();
 sg13g2_fill_2 FILLER_35_2543 ();
 sg13g2_fill_1 FILLER_35_2557 ();
 sg13g2_fill_1 FILLER_35_2563 ();
 sg13g2_decap_8 FILLER_35_2570 ();
 sg13g2_fill_1 FILLER_35_2577 ();
 sg13g2_decap_8 FILLER_35_2600 ();
 sg13g2_decap_8 FILLER_35_2622 ();
 sg13g2_decap_8 FILLER_35_2629 ();
 sg13g2_fill_2 FILLER_35_2636 ();
 sg13g2_fill_1 FILLER_35_2638 ();
 sg13g2_decap_8 FILLER_35_2654 ();
 sg13g2_decap_4 FILLER_35_2661 ();
 sg13g2_fill_2 FILLER_35_2687 ();
 sg13g2_fill_1 FILLER_35_2707 ();
 sg13g2_decap_8 FILLER_35_2717 ();
 sg13g2_decap_4 FILLER_35_2740 ();
 sg13g2_fill_1 FILLER_35_2744 ();
 sg13g2_fill_2 FILLER_35_2749 ();
 sg13g2_decap_8 FILLER_35_2769 ();
 sg13g2_decap_4 FILLER_35_2776 ();
 sg13g2_fill_2 FILLER_35_2780 ();
 sg13g2_fill_2 FILLER_35_2795 ();
 sg13g2_decap_4 FILLER_35_2813 ();
 sg13g2_fill_2 FILLER_35_2817 ();
 sg13g2_fill_2 FILLER_35_2827 ();
 sg13g2_decap_8 FILLER_35_2835 ();
 sg13g2_fill_2 FILLER_35_2842 ();
 sg13g2_decap_8 FILLER_35_2853 ();
 sg13g2_fill_2 FILLER_35_2860 ();
 sg13g2_fill_1 FILLER_35_2862 ();
 sg13g2_fill_1 FILLER_35_2872 ();
 sg13g2_fill_1 FILLER_35_2899 ();
 sg13g2_fill_2 FILLER_35_2913 ();
 sg13g2_decap_8 FILLER_35_2938 ();
 sg13g2_fill_1 FILLER_35_2945 ();
 sg13g2_fill_2 FILLER_35_2959 ();
 sg13g2_decap_4 FILLER_35_2966 ();
 sg13g2_fill_2 FILLER_35_2970 ();
 sg13g2_fill_1 FILLER_35_2976 ();
 sg13g2_fill_2 FILLER_35_2982 ();
 sg13g2_fill_1 FILLER_35_2984 ();
 sg13g2_decap_8 FILLER_35_2993 ();
 sg13g2_decap_4 FILLER_35_3000 ();
 sg13g2_fill_2 FILLER_35_3012 ();
 sg13g2_decap_8 FILLER_35_3072 ();
 sg13g2_decap_4 FILLER_35_3079 ();
 sg13g2_fill_2 FILLER_35_3083 ();
 sg13g2_decap_8 FILLER_35_3172 ();
 sg13g2_decap_4 FILLER_35_3179 ();
 sg13g2_fill_1 FILLER_35_3183 ();
 sg13g2_decap_8 FILLER_35_3197 ();
 sg13g2_fill_1 FILLER_35_3204 ();
 sg13g2_decap_8 FILLER_35_3232 ();
 sg13g2_decap_4 FILLER_35_3244 ();
 sg13g2_fill_1 FILLER_35_3248 ();
 sg13g2_fill_2 FILLER_35_3285 ();
 sg13g2_fill_1 FILLER_35_3287 ();
 sg13g2_decap_8 FILLER_35_3310 ();
 sg13g2_decap_8 FILLER_35_3317 ();
 sg13g2_fill_1 FILLER_35_3341 ();
 sg13g2_fill_1 FILLER_35_3351 ();
 sg13g2_fill_2 FILLER_35_3358 ();
 sg13g2_fill_1 FILLER_35_3415 ();
 sg13g2_fill_2 FILLER_35_3425 ();
 sg13g2_decap_8 FILLER_35_3436 ();
 sg13g2_decap_8 FILLER_35_3443 ();
 sg13g2_decap_8 FILLER_35_3450 ();
 sg13g2_decap_8 FILLER_35_3457 ();
 sg13g2_decap_8 FILLER_35_3464 ();
 sg13g2_decap_8 FILLER_35_3471 ();
 sg13g2_decap_8 FILLER_35_3478 ();
 sg13g2_decap_8 FILLER_35_3485 ();
 sg13g2_decap_8 FILLER_35_3492 ();
 sg13g2_decap_8 FILLER_35_3499 ();
 sg13g2_decap_8 FILLER_35_3506 ();
 sg13g2_decap_8 FILLER_35_3513 ();
 sg13g2_decap_8 FILLER_35_3520 ();
 sg13g2_decap_8 FILLER_35_3527 ();
 sg13g2_decap_8 FILLER_35_3534 ();
 sg13g2_decap_8 FILLER_35_3541 ();
 sg13g2_decap_8 FILLER_35_3548 ();
 sg13g2_decap_8 FILLER_35_3555 ();
 sg13g2_decap_8 FILLER_35_3562 ();
 sg13g2_decap_8 FILLER_35_3569 ();
 sg13g2_decap_4 FILLER_35_3576 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_fill_1 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_411 ();
 sg13g2_fill_2 FILLER_36_418 ();
 sg13g2_decap_8 FILLER_36_430 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_decap_4 FILLER_36_469 ();
 sg13g2_fill_1 FILLER_36_473 ();
 sg13g2_decap_4 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_485 ();
 sg13g2_decap_8 FILLER_36_509 ();
 sg13g2_decap_8 FILLER_36_516 ();
 sg13g2_decap_8 FILLER_36_523 ();
 sg13g2_decap_4 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_534 ();
 sg13g2_fill_1 FILLER_36_540 ();
 sg13g2_fill_1 FILLER_36_558 ();
 sg13g2_decap_8 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_570 ();
 sg13g2_fill_1 FILLER_36_579 ();
 sg13g2_fill_2 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_4 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_673 ();
 sg13g2_decap_8 FILLER_36_684 ();
 sg13g2_fill_2 FILLER_36_691 ();
 sg13g2_fill_2 FILLER_36_707 ();
 sg13g2_fill_2 FILLER_36_713 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_1 FILLER_36_729 ();
 sg13g2_fill_2 FILLER_36_740 ();
 sg13g2_fill_1 FILLER_36_742 ();
 sg13g2_fill_2 FILLER_36_749 ();
 sg13g2_fill_1 FILLER_36_751 ();
 sg13g2_fill_2 FILLER_36_767 ();
 sg13g2_fill_2 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_fill_1 FILLER_36_827 ();
 sg13g2_decap_4 FILLER_36_843 ();
 sg13g2_fill_2 FILLER_36_847 ();
 sg13g2_fill_2 FILLER_36_943 ();
 sg13g2_decap_8 FILLER_36_958 ();
 sg13g2_fill_1 FILLER_36_965 ();
 sg13g2_decap_8 FILLER_36_976 ();
 sg13g2_decap_8 FILLER_36_983 ();
 sg13g2_fill_1 FILLER_36_990 ();
 sg13g2_fill_1 FILLER_36_1004 ();
 sg13g2_fill_2 FILLER_36_1011 ();
 sg13g2_fill_2 FILLER_36_1021 ();
 sg13g2_fill_1 FILLER_36_1023 ();
 sg13g2_decap_4 FILLER_36_1049 ();
 sg13g2_fill_1 FILLER_36_1053 ();
 sg13g2_decap_8 FILLER_36_1081 ();
 sg13g2_fill_2 FILLER_36_1088 ();
 sg13g2_fill_1 FILLER_36_1090 ();
 sg13g2_fill_1 FILLER_36_1104 ();
 sg13g2_decap_4 FILLER_36_1118 ();
 sg13g2_fill_1 FILLER_36_1122 ();
 sg13g2_fill_2 FILLER_36_1136 ();
 sg13g2_fill_1 FILLER_36_1151 ();
 sg13g2_fill_1 FILLER_36_1163 ();
 sg13g2_decap_4 FILLER_36_1179 ();
 sg13g2_fill_2 FILLER_36_1183 ();
 sg13g2_decap_4 FILLER_36_1198 ();
 sg13g2_decap_8 FILLER_36_1243 ();
 sg13g2_fill_2 FILLER_36_1266 ();
 sg13g2_fill_2 FILLER_36_1288 ();
 sg13g2_fill_2 FILLER_36_1305 ();
 sg13g2_decap_8 FILLER_36_1311 ();
 sg13g2_fill_1 FILLER_36_1341 ();
 sg13g2_fill_2 FILLER_36_1361 ();
 sg13g2_fill_1 FILLER_36_1363 ();
 sg13g2_fill_1 FILLER_36_1372 ();
 sg13g2_decap_8 FILLER_36_1386 ();
 sg13g2_fill_2 FILLER_36_1393 ();
 sg13g2_fill_1 FILLER_36_1403 ();
 sg13g2_decap_8 FILLER_36_1412 ();
 sg13g2_decap_4 FILLER_36_1419 ();
 sg13g2_fill_2 FILLER_36_1423 ();
 sg13g2_decap_8 FILLER_36_1480 ();
 sg13g2_decap_8 FILLER_36_1487 ();
 sg13g2_fill_1 FILLER_36_1502 ();
 sg13g2_fill_2 FILLER_36_1511 ();
 sg13g2_decap_8 FILLER_36_1516 ();
 sg13g2_fill_2 FILLER_36_1523 ();
 sg13g2_fill_1 FILLER_36_1525 ();
 sg13g2_decap_4 FILLER_36_1534 ();
 sg13g2_fill_2 FILLER_36_1538 ();
 sg13g2_fill_2 FILLER_36_1552 ();
 sg13g2_fill_1 FILLER_36_1554 ();
 sg13g2_decap_8 FILLER_36_1564 ();
 sg13g2_decap_8 FILLER_36_1571 ();
 sg13g2_decap_8 FILLER_36_1578 ();
 sg13g2_decap_4 FILLER_36_1585 ();
 sg13g2_fill_1 FILLER_36_1589 ();
 sg13g2_fill_2 FILLER_36_1618 ();
 sg13g2_fill_1 FILLER_36_1620 ();
 sg13g2_fill_1 FILLER_36_1625 ();
 sg13g2_decap_8 FILLER_36_1638 ();
 sg13g2_fill_1 FILLER_36_1663 ();
 sg13g2_fill_2 FILLER_36_1669 ();
 sg13g2_decap_8 FILLER_36_1675 ();
 sg13g2_decap_4 FILLER_36_1682 ();
 sg13g2_fill_2 FILLER_36_1686 ();
 sg13g2_fill_2 FILLER_36_1701 ();
 sg13g2_fill_1 FILLER_36_1703 ();
 sg13g2_fill_2 FILLER_36_1709 ();
 sg13g2_fill_1 FILLER_36_1711 ();
 sg13g2_fill_1 FILLER_36_1716 ();
 sg13g2_decap_4 FILLER_36_1723 ();
 sg13g2_fill_2 FILLER_36_1727 ();
 sg13g2_fill_2 FILLER_36_1734 ();
 sg13g2_decap_8 FILLER_36_1752 ();
 sg13g2_decap_4 FILLER_36_1759 ();
 sg13g2_decap_4 FILLER_36_1776 ();
 sg13g2_decap_4 FILLER_36_1788 ();
 sg13g2_fill_2 FILLER_36_1792 ();
 sg13g2_fill_1 FILLER_36_1798 ();
 sg13g2_fill_2 FILLER_36_1816 ();
 sg13g2_fill_1 FILLER_36_1818 ();
 sg13g2_fill_2 FILLER_36_1829 ();
 sg13g2_fill_1 FILLER_36_1831 ();
 sg13g2_decap_4 FILLER_36_1838 ();
 sg13g2_fill_1 FILLER_36_1842 ();
 sg13g2_decap_8 FILLER_36_1848 ();
 sg13g2_fill_2 FILLER_36_1855 ();
 sg13g2_fill_1 FILLER_36_1857 ();
 sg13g2_decap_8 FILLER_36_1883 ();
 sg13g2_fill_2 FILLER_36_1912 ();
 sg13g2_decap_4 FILLER_36_1934 ();
 sg13g2_decap_4 FILLER_36_1963 ();
 sg13g2_decap_4 FILLER_36_1982 ();
 sg13g2_fill_2 FILLER_36_1986 ();
 sg13g2_fill_1 FILLER_36_1996 ();
 sg13g2_decap_8 FILLER_36_2002 ();
 sg13g2_fill_2 FILLER_36_2009 ();
 sg13g2_fill_1 FILLER_36_2011 ();
 sg13g2_fill_2 FILLER_36_2051 ();
 sg13g2_fill_2 FILLER_36_2058 ();
 sg13g2_decap_8 FILLER_36_2066 ();
 sg13g2_decap_8 FILLER_36_2073 ();
 sg13g2_fill_2 FILLER_36_2098 ();
 sg13g2_fill_1 FILLER_36_2100 ();
 sg13g2_fill_2 FILLER_36_2109 ();
 sg13g2_fill_1 FILLER_36_2120 ();
 sg13g2_decap_4 FILLER_36_2148 ();
 sg13g2_fill_2 FILLER_36_2152 ();
 sg13g2_fill_1 FILLER_36_2167 ();
 sg13g2_fill_2 FILLER_36_2186 ();
 sg13g2_fill_1 FILLER_36_2188 ();
 sg13g2_fill_2 FILLER_36_2197 ();
 sg13g2_fill_1 FILLER_36_2199 ();
 sg13g2_decap_4 FILLER_36_2213 ();
 sg13g2_decap_4 FILLER_36_2232 ();
 sg13g2_decap_8 FILLER_36_2250 ();
 sg13g2_decap_8 FILLER_36_2257 ();
 sg13g2_decap_4 FILLER_36_2264 ();
 sg13g2_fill_1 FILLER_36_2268 ();
 sg13g2_decap_8 FILLER_36_2296 ();
 sg13g2_fill_1 FILLER_36_2303 ();
 sg13g2_decap_8 FILLER_36_2322 ();
 sg13g2_decap_4 FILLER_36_2333 ();
 sg13g2_decap_4 FILLER_36_2350 ();
 sg13g2_fill_1 FILLER_36_2354 ();
 sg13g2_fill_2 FILLER_36_2359 ();
 sg13g2_fill_1 FILLER_36_2361 ();
 sg13g2_decap_8 FILLER_36_2368 ();
 sg13g2_decap_8 FILLER_36_2375 ();
 sg13g2_fill_1 FILLER_36_2382 ();
 sg13g2_fill_2 FILLER_36_2396 ();
 sg13g2_fill_1 FILLER_36_2398 ();
 sg13g2_decap_8 FILLER_36_2406 ();
 sg13g2_fill_1 FILLER_36_2413 ();
 sg13g2_decap_8 FILLER_36_2428 ();
 sg13g2_decap_8 FILLER_36_2435 ();
 sg13g2_decap_4 FILLER_36_2442 ();
 sg13g2_decap_8 FILLER_36_2451 ();
 sg13g2_fill_2 FILLER_36_2458 ();
 sg13g2_fill_1 FILLER_36_2460 ();
 sg13g2_fill_2 FILLER_36_2485 ();
 sg13g2_fill_2 FILLER_36_2497 ();
 sg13g2_fill_1 FILLER_36_2499 ();
 sg13g2_fill_2 FILLER_36_2519 ();
 sg13g2_fill_1 FILLER_36_2521 ();
 sg13g2_fill_1 FILLER_36_2535 ();
 sg13g2_decap_4 FILLER_36_2550 ();
 sg13g2_fill_2 FILLER_36_2554 ();
 sg13g2_decap_8 FILLER_36_2574 ();
 sg13g2_decap_4 FILLER_36_2581 ();
 sg13g2_fill_1 FILLER_36_2585 ();
 sg13g2_fill_2 FILLER_36_2603 ();
 sg13g2_fill_1 FILLER_36_2605 ();
 sg13g2_fill_2 FILLER_36_2628 ();
 sg13g2_fill_1 FILLER_36_2630 ();
 sg13g2_decap_4 FILLER_36_2653 ();
 sg13g2_fill_2 FILLER_36_2657 ();
 sg13g2_decap_8 FILLER_36_2675 ();
 sg13g2_decap_4 FILLER_36_2682 ();
 sg13g2_fill_2 FILLER_36_2686 ();
 sg13g2_decap_8 FILLER_36_2715 ();
 sg13g2_fill_2 FILLER_36_2728 ();
 sg13g2_fill_1 FILLER_36_2730 ();
 sg13g2_decap_8 FILLER_36_2743 ();
 sg13g2_decap_4 FILLER_36_2750 ();
 sg13g2_fill_1 FILLER_36_2754 ();
 sg13g2_fill_1 FILLER_36_2763 ();
 sg13g2_fill_2 FILLER_36_2787 ();
 sg13g2_decap_4 FILLER_36_2807 ();
 sg13g2_fill_1 FILLER_36_2834 ();
 sg13g2_fill_1 FILLER_36_2866 ();
 sg13g2_decap_4 FILLER_36_2880 ();
 sg13g2_fill_1 FILLER_36_2884 ();
 sg13g2_decap_4 FILLER_36_2893 ();
 sg13g2_decap_8 FILLER_36_2902 ();
 sg13g2_decap_8 FILLER_36_2909 ();
 sg13g2_decap_8 FILLER_36_2942 ();
 sg13g2_fill_2 FILLER_36_2957 ();
 sg13g2_decap_8 FILLER_36_2969 ();
 sg13g2_decap_4 FILLER_36_2976 ();
 sg13g2_fill_1 FILLER_36_2980 ();
 sg13g2_decap_8 FILLER_36_2991 ();
 sg13g2_decap_4 FILLER_36_2998 ();
 sg13g2_fill_2 FILLER_36_3002 ();
 sg13g2_fill_1 FILLER_36_3025 ();
 sg13g2_fill_2 FILLER_36_3038 ();
 sg13g2_fill_2 FILLER_36_3090 ();
 sg13g2_decap_4 FILLER_36_3096 ();
 sg13g2_fill_2 FILLER_36_3100 ();
 sg13g2_fill_2 FILLER_36_3120 ();
 sg13g2_decap_8 FILLER_36_3198 ();
 sg13g2_fill_1 FILLER_36_3205 ();
 sg13g2_decap_8 FILLER_36_3224 ();
 sg13g2_decap_4 FILLER_36_3231 ();
 sg13g2_fill_1 FILLER_36_3235 ();
 sg13g2_fill_2 FILLER_36_3279 ();
 sg13g2_decap_8 FILLER_36_3312 ();
 sg13g2_fill_2 FILLER_36_3356 ();
 sg13g2_fill_1 FILLER_36_3367 ();
 sg13g2_fill_1 FILLER_36_3382 ();
 sg13g2_fill_1 FILLER_36_3401 ();
 sg13g2_fill_2 FILLER_36_3416 ();
 sg13g2_decap_8 FILLER_36_3446 ();
 sg13g2_decap_8 FILLER_36_3453 ();
 sg13g2_decap_8 FILLER_36_3460 ();
 sg13g2_decap_8 FILLER_36_3467 ();
 sg13g2_decap_8 FILLER_36_3474 ();
 sg13g2_decap_8 FILLER_36_3481 ();
 sg13g2_decap_8 FILLER_36_3488 ();
 sg13g2_decap_8 FILLER_36_3495 ();
 sg13g2_decap_8 FILLER_36_3502 ();
 sg13g2_decap_8 FILLER_36_3509 ();
 sg13g2_decap_8 FILLER_36_3516 ();
 sg13g2_decap_8 FILLER_36_3523 ();
 sg13g2_decap_8 FILLER_36_3530 ();
 sg13g2_decap_8 FILLER_36_3537 ();
 sg13g2_decap_8 FILLER_36_3544 ();
 sg13g2_decap_8 FILLER_36_3551 ();
 sg13g2_decap_8 FILLER_36_3558 ();
 sg13g2_decap_8 FILLER_36_3565 ();
 sg13g2_decap_8 FILLER_36_3572 ();
 sg13g2_fill_1 FILLER_36_3579 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_370 ();
 sg13g2_fill_2 FILLER_37_394 ();
 sg13g2_fill_1 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_409 ();
 sg13g2_fill_2 FILLER_37_437 ();
 sg13g2_fill_1 FILLER_37_457 ();
 sg13g2_fill_2 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_465 ();
 sg13g2_decap_8 FILLER_37_520 ();
 sg13g2_fill_2 FILLER_37_527 ();
 sg13g2_decap_4 FILLER_37_537 ();
 sg13g2_fill_2 FILLER_37_541 ();
 sg13g2_fill_1 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_587 ();
 sg13g2_fill_1 FILLER_37_609 ();
 sg13g2_fill_1 FILLER_37_636 ();
 sg13g2_fill_1 FILLER_37_673 ();
 sg13g2_decap_8 FILLER_37_702 ();
 sg13g2_decap_4 FILLER_37_715 ();
 sg13g2_fill_1 FILLER_37_719 ();
 sg13g2_fill_2 FILLER_37_726 ();
 sg13g2_fill_1 FILLER_37_728 ();
 sg13g2_decap_4 FILLER_37_764 ();
 sg13g2_fill_2 FILLER_37_768 ();
 sg13g2_decap_4 FILLER_37_798 ();
 sg13g2_fill_2 FILLER_37_852 ();
 sg13g2_fill_1 FILLER_37_854 ();
 sg13g2_fill_2 FILLER_37_861 ();
 sg13g2_fill_2 FILLER_37_876 ();
 sg13g2_fill_1 FILLER_37_878 ();
 sg13g2_decap_8 FILLER_37_892 ();
 sg13g2_decap_4 FILLER_37_899 ();
 sg13g2_fill_2 FILLER_37_903 ();
 sg13g2_fill_1 FILLER_37_911 ();
 sg13g2_decap_4 FILLER_37_915 ();
 sg13g2_fill_1 FILLER_37_919 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_fill_2 FILLER_37_943 ();
 sg13g2_fill_1 FILLER_37_945 ();
 sg13g2_fill_1 FILLER_37_954 ();
 sg13g2_decap_8 FILLER_37_984 ();
 sg13g2_fill_1 FILLER_37_991 ();
 sg13g2_fill_2 FILLER_37_1010 ();
 sg13g2_fill_1 FILLER_37_1012 ();
 sg13g2_fill_2 FILLER_37_1030 ();
 sg13g2_decap_8 FILLER_37_1045 ();
 sg13g2_fill_2 FILLER_37_1052 ();
 sg13g2_decap_4 FILLER_37_1079 ();
 sg13g2_fill_1 FILLER_37_1083 ();
 sg13g2_fill_2 FILLER_37_1101 ();
 sg13g2_fill_1 FILLER_37_1103 ();
 sg13g2_decap_8 FILLER_37_1116 ();
 sg13g2_fill_1 FILLER_37_1123 ();
 sg13g2_decap_8 FILLER_37_1145 ();
 sg13g2_fill_1 FILLER_37_1152 ();
 sg13g2_decap_8 FILLER_37_1173 ();
 sg13g2_decap_4 FILLER_37_1180 ();
 sg13g2_fill_1 FILLER_37_1184 ();
 sg13g2_fill_1 FILLER_37_1193 ();
 sg13g2_decap_4 FILLER_37_1202 ();
 sg13g2_fill_1 FILLER_37_1206 ();
 sg13g2_decap_8 FILLER_37_1237 ();
 sg13g2_fill_2 FILLER_37_1244 ();
 sg13g2_decap_4 FILLER_37_1264 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_fill_1 FILLER_37_1288 ();
 sg13g2_fill_2 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1315 ();
 sg13g2_fill_2 FILLER_37_1329 ();
 sg13g2_decap_4 FILLER_37_1335 ();
 sg13g2_decap_8 FILLER_37_1352 ();
 sg13g2_decap_4 FILLER_37_1367 ();
 sg13g2_decap_8 FILLER_37_1379 ();
 sg13g2_fill_2 FILLER_37_1407 ();
 sg13g2_fill_1 FILLER_37_1409 ();
 sg13g2_fill_2 FILLER_37_1421 ();
 sg13g2_fill_1 FILLER_37_1434 ();
 sg13g2_decap_8 FILLER_37_1439 ();
 sg13g2_decap_4 FILLER_37_1446 ();
 sg13g2_fill_1 FILLER_37_1450 ();
 sg13g2_decap_4 FILLER_37_1455 ();
 sg13g2_fill_1 FILLER_37_1459 ();
 sg13g2_fill_2 FILLER_37_1473 ();
 sg13g2_fill_1 FILLER_37_1475 ();
 sg13g2_decap_8 FILLER_37_1480 ();
 sg13g2_decap_4 FILLER_37_1487 ();
 sg13g2_fill_1 FILLER_37_1491 ();
 sg13g2_fill_2 FILLER_37_1514 ();
 sg13g2_fill_1 FILLER_37_1542 ();
 sg13g2_fill_1 FILLER_37_1555 ();
 sg13g2_decap_8 FILLER_37_1589 ();
 sg13g2_decap_4 FILLER_37_1596 ();
 sg13g2_decap_8 FILLER_37_1612 ();
 sg13g2_decap_4 FILLER_37_1619 ();
 sg13g2_fill_1 FILLER_37_1623 ();
 sg13g2_decap_4 FILLER_37_1632 ();
 sg13g2_fill_2 FILLER_37_1656 ();
 sg13g2_fill_1 FILLER_37_1658 ();
 sg13g2_fill_1 FILLER_37_1684 ();
 sg13g2_decap_8 FILLER_37_1693 ();
 sg13g2_fill_2 FILLER_37_1700 ();
 sg13g2_fill_2 FILLER_37_1710 ();
 sg13g2_fill_1 FILLER_37_1712 ();
 sg13g2_fill_2 FILLER_37_1736 ();
 sg13g2_fill_1 FILLER_37_1738 ();
 sg13g2_decap_8 FILLER_37_1742 ();
 sg13g2_fill_2 FILLER_37_1763 ();
 sg13g2_fill_2 FILLER_37_1804 ();
 sg13g2_fill_2 FILLER_37_1811 ();
 sg13g2_decap_8 FILLER_37_1828 ();
 sg13g2_decap_4 FILLER_37_1861 ();
 sg13g2_fill_1 FILLER_37_1870 ();
 sg13g2_fill_2 FILLER_37_1877 ();
 sg13g2_decap_8 FILLER_37_1895 ();
 sg13g2_fill_2 FILLER_37_1962 ();
 sg13g2_fill_1 FILLER_37_1964 ();
 sg13g2_decap_8 FILLER_37_1985 ();
 sg13g2_decap_4 FILLER_37_1992 ();
 sg13g2_decap_8 FILLER_37_2004 ();
 sg13g2_fill_1 FILLER_37_2031 ();
 sg13g2_fill_2 FILLER_37_2040 ();
 sg13g2_fill_1 FILLER_37_2042 ();
 sg13g2_fill_1 FILLER_37_2051 ();
 sg13g2_decap_8 FILLER_37_2069 ();
 sg13g2_decap_8 FILLER_37_2076 ();
 sg13g2_fill_1 FILLER_37_2083 ();
 sg13g2_fill_2 FILLER_37_2093 ();
 sg13g2_fill_1 FILLER_37_2095 ();
 sg13g2_decap_8 FILLER_37_2123 ();
 sg13g2_decap_4 FILLER_37_2130 ();
 sg13g2_fill_1 FILLER_37_2134 ();
 sg13g2_fill_2 FILLER_37_2143 ();
 sg13g2_fill_1 FILLER_37_2154 ();
 sg13g2_fill_1 FILLER_37_2215 ();
 sg13g2_decap_8 FILLER_37_2264 ();
 sg13g2_fill_2 FILLER_37_2271 ();
 sg13g2_fill_1 FILLER_37_2273 ();
 sg13g2_decap_8 FILLER_37_2300 ();
 sg13g2_fill_1 FILLER_37_2349 ();
 sg13g2_decap_4 FILLER_37_2387 ();
 sg13g2_fill_2 FILLER_37_2391 ();
 sg13g2_fill_1 FILLER_37_2396 ();
 sg13g2_fill_2 FILLER_37_2425 ();
 sg13g2_fill_1 FILLER_37_2427 ();
 sg13g2_fill_2 FILLER_37_2436 ();
 sg13g2_fill_1 FILLER_37_2438 ();
 sg13g2_fill_2 FILLER_37_2470 ();
 sg13g2_decap_8 FILLER_37_2484 ();
 sg13g2_fill_2 FILLER_37_2491 ();
 sg13g2_fill_2 FILLER_37_2506 ();
 sg13g2_fill_1 FILLER_37_2508 ();
 sg13g2_decap_4 FILLER_37_2526 ();
 sg13g2_decap_8 FILLER_37_2556 ();
 sg13g2_decap_4 FILLER_37_2563 ();
 sg13g2_fill_1 FILLER_37_2594 ();
 sg13g2_fill_2 FILLER_37_2611 ();
 sg13g2_decap_8 FILLER_37_2622 ();
 sg13g2_fill_1 FILLER_37_2629 ();
 sg13g2_fill_2 FILLER_37_2635 ();
 sg13g2_fill_2 FILLER_37_2642 ();
 sg13g2_fill_1 FILLER_37_2644 ();
 sg13g2_fill_2 FILLER_37_2650 ();
 sg13g2_decap_8 FILLER_37_2672 ();
 sg13g2_decap_8 FILLER_37_2679 ();
 sg13g2_decap_4 FILLER_37_2686 ();
 sg13g2_fill_1 FILLER_37_2690 ();
 sg13g2_decap_8 FILLER_37_2713 ();
 sg13g2_fill_1 FILLER_37_2720 ();
 sg13g2_decap_8 FILLER_37_2747 ();
 sg13g2_decap_8 FILLER_37_2754 ();
 sg13g2_decap_4 FILLER_37_2781 ();
 sg13g2_fill_1 FILLER_37_2785 ();
 sg13g2_decap_8 FILLER_37_2798 ();
 sg13g2_decap_4 FILLER_37_2805 ();
 sg13g2_fill_1 FILLER_37_2809 ();
 sg13g2_fill_1 FILLER_37_2829 ();
 sg13g2_fill_1 FILLER_37_2875 ();
 sg13g2_fill_2 FILLER_37_2921 ();
 sg13g2_fill_2 FILLER_37_2952 ();
 sg13g2_fill_1 FILLER_37_2954 ();
 sg13g2_fill_1 FILLER_37_2978 ();
 sg13g2_fill_1 FILLER_37_3021 ();
 sg13g2_fill_2 FILLER_37_3049 ();
 sg13g2_fill_1 FILLER_37_3051 ();
 sg13g2_fill_1 FILLER_37_3056 ();
 sg13g2_decap_8 FILLER_37_3070 ();
 sg13g2_fill_1 FILLER_37_3077 ();
 sg13g2_fill_1 FILLER_37_3105 ();
 sg13g2_fill_2 FILLER_37_3111 ();
 sg13g2_fill_1 FILLER_37_3113 ();
 sg13g2_fill_2 FILLER_37_3128 ();
 sg13g2_fill_1 FILLER_37_3153 ();
 sg13g2_decap_4 FILLER_37_3163 ();
 sg13g2_fill_1 FILLER_37_3167 ();
 sg13g2_decap_8 FILLER_37_3187 ();
 sg13g2_fill_2 FILLER_37_3194 ();
 sg13g2_decap_4 FILLER_37_3232 ();
 sg13g2_fill_2 FILLER_37_3236 ();
 sg13g2_fill_2 FILLER_37_3294 ();
 sg13g2_decap_4 FILLER_37_3312 ();
 sg13g2_decap_4 FILLER_37_3320 ();
 sg13g2_decap_8 FILLER_37_3329 ();
 sg13g2_decap_8 FILLER_37_3336 ();
 sg13g2_fill_1 FILLER_37_3343 ();
 sg13g2_fill_2 FILLER_37_3373 ();
 sg13g2_fill_1 FILLER_37_3394 ();
 sg13g2_decap_8 FILLER_37_3427 ();
 sg13g2_decap_8 FILLER_37_3434 ();
 sg13g2_decap_8 FILLER_37_3441 ();
 sg13g2_decap_8 FILLER_37_3448 ();
 sg13g2_decap_8 FILLER_37_3455 ();
 sg13g2_decap_8 FILLER_37_3462 ();
 sg13g2_decap_8 FILLER_37_3469 ();
 sg13g2_decap_8 FILLER_37_3476 ();
 sg13g2_decap_8 FILLER_37_3483 ();
 sg13g2_decap_8 FILLER_37_3490 ();
 sg13g2_decap_8 FILLER_37_3497 ();
 sg13g2_decap_8 FILLER_37_3504 ();
 sg13g2_decap_8 FILLER_37_3511 ();
 sg13g2_decap_8 FILLER_37_3518 ();
 sg13g2_decap_8 FILLER_37_3525 ();
 sg13g2_decap_8 FILLER_37_3532 ();
 sg13g2_decap_8 FILLER_37_3539 ();
 sg13g2_decap_8 FILLER_37_3546 ();
 sg13g2_decap_8 FILLER_37_3553 ();
 sg13g2_decap_8 FILLER_37_3560 ();
 sg13g2_decap_8 FILLER_37_3567 ();
 sg13g2_decap_4 FILLER_37_3574 ();
 sg13g2_fill_2 FILLER_37_3578 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_339 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_decap_4 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_2 FILLER_38_413 ();
 sg13g2_fill_1 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_4 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_431 ();
 sg13g2_decap_4 FILLER_38_436 ();
 sg13g2_fill_2 FILLER_38_440 ();
 sg13g2_fill_2 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_491 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_fill_2 FILLER_38_538 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_decap_4 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_561 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_4 FILLER_38_581 ();
 sg13g2_fill_2 FILLER_38_585 ();
 sg13g2_decap_8 FILLER_38_590 ();
 sg13g2_fill_1 FILLER_38_597 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_fill_2 FILLER_38_659 ();
 sg13g2_fill_2 FILLER_38_680 ();
 sg13g2_fill_1 FILLER_38_682 ();
 sg13g2_decap_4 FILLER_38_700 ();
 sg13g2_fill_2 FILLER_38_707 ();
 sg13g2_decap_4 FILLER_38_718 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_fill_1 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_769 ();
 sg13g2_fill_1 FILLER_38_776 ();
 sg13g2_fill_1 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_785 ();
 sg13g2_fill_2 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_4 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_fill_2 FILLER_38_835 ();
 sg13g2_decap_4 FILLER_38_841 ();
 sg13g2_fill_2 FILLER_38_845 ();
 sg13g2_fill_1 FILLER_38_905 ();
 sg13g2_decap_4 FILLER_38_934 ();
 sg13g2_fill_2 FILLER_38_938 ();
 sg13g2_fill_2 FILLER_38_953 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_4 FILLER_38_966 ();
 sg13g2_fill_1 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_fill_1 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1024 ();
 sg13g2_fill_1 FILLER_38_1031 ();
 sg13g2_decap_4 FILLER_38_1048 ();
 sg13g2_decap_8 FILLER_38_1056 ();
 sg13g2_decap_8 FILLER_38_1063 ();
 sg13g2_fill_1 FILLER_38_1076 ();
 sg13g2_decap_8 FILLER_38_1081 ();
 sg13g2_fill_2 FILLER_38_1088 ();
 sg13g2_decap_4 FILLER_38_1120 ();
 sg13g2_fill_1 FILLER_38_1124 ();
 sg13g2_decap_4 FILLER_38_1138 ();
 sg13g2_fill_1 FILLER_38_1142 ();
 sg13g2_decap_8 FILLER_38_1156 ();
 sg13g2_fill_1 FILLER_38_1163 ();
 sg13g2_decap_8 FILLER_38_1181 ();
 sg13g2_decap_8 FILLER_38_1204 ();
 sg13g2_decap_4 FILLER_38_1211 ();
 sg13g2_fill_2 FILLER_38_1215 ();
 sg13g2_fill_2 FILLER_38_1222 ();
 sg13g2_fill_1 FILLER_38_1224 ();
 sg13g2_decap_8 FILLER_38_1281 ();
 sg13g2_decap_4 FILLER_38_1288 ();
 sg13g2_fill_1 FILLER_38_1292 ();
 sg13g2_fill_2 FILLER_38_1306 ();
 sg13g2_fill_1 FILLER_38_1312 ();
 sg13g2_fill_1 FILLER_38_1330 ();
 sg13g2_fill_2 FILLER_38_1346 ();
 sg13g2_fill_2 FILLER_38_1360 ();
 sg13g2_decap_8 FILLER_38_1380 ();
 sg13g2_decap_4 FILLER_38_1387 ();
 sg13g2_fill_1 FILLER_38_1402 ();
 sg13g2_decap_4 FILLER_38_1409 ();
 sg13g2_fill_1 FILLER_38_1433 ();
 sg13g2_fill_2 FILLER_38_1455 ();
 sg13g2_fill_2 FILLER_38_1469 ();
 sg13g2_fill_2 FILLER_38_1479 ();
 sg13g2_fill_1 FILLER_38_1481 ();
 sg13g2_fill_1 FILLER_38_1508 ();
 sg13g2_fill_2 FILLER_38_1528 ();
 sg13g2_fill_1 FILLER_38_1530 ();
 sg13g2_fill_1 FILLER_38_1536 ();
 sg13g2_decap_4 FILLER_38_1545 ();
 sg13g2_decap_8 FILLER_38_1602 ();
 sg13g2_decap_8 FILLER_38_1609 ();
 sg13g2_fill_2 FILLER_38_1616 ();
 sg13g2_fill_1 FILLER_38_1618 ();
 sg13g2_fill_1 FILLER_38_1632 ();
 sg13g2_fill_2 FILLER_38_1643 ();
 sg13g2_decap_4 FILLER_38_1661 ();
 sg13g2_fill_2 FILLER_38_1680 ();
 sg13g2_fill_1 FILLER_38_1682 ();
 sg13g2_decap_4 FILLER_38_1707 ();
 sg13g2_fill_2 FILLER_38_1711 ();
 sg13g2_fill_2 FILLER_38_1717 ();
 sg13g2_fill_1 FILLER_38_1719 ();
 sg13g2_decap_8 FILLER_38_1739 ();
 sg13g2_fill_2 FILLER_38_1746 ();
 sg13g2_fill_1 FILLER_38_1748 ();
 sg13g2_decap_8 FILLER_38_1779 ();
 sg13g2_decap_8 FILLER_38_1790 ();
 sg13g2_decap_8 FILLER_38_1821 ();
 sg13g2_fill_2 FILLER_38_1828 ();
 sg13g2_decap_8 FILLER_38_1843 ();
 sg13g2_fill_2 FILLER_38_1850 ();
 sg13g2_fill_2 FILLER_38_1873 ();
 sg13g2_fill_1 FILLER_38_1875 ();
 sg13g2_fill_2 FILLER_38_1885 ();
 sg13g2_decap_8 FILLER_38_1891 ();
 sg13g2_decap_4 FILLER_38_1898 ();
 sg13g2_decap_4 FILLER_38_1932 ();
 sg13g2_fill_1 FILLER_38_1936 ();
 sg13g2_decap_8 FILLER_38_1955 ();
 sg13g2_fill_2 FILLER_38_1962 ();
 sg13g2_decap_8 FILLER_38_1967 ();
 sg13g2_fill_1 FILLER_38_1974 ();
 sg13g2_decap_8 FILLER_38_2002 ();
 sg13g2_fill_2 FILLER_38_2009 ();
 sg13g2_fill_2 FILLER_38_2032 ();
 sg13g2_fill_1 FILLER_38_2034 ();
 sg13g2_fill_1 FILLER_38_2104 ();
 sg13g2_fill_2 FILLER_38_2110 ();
 sg13g2_fill_1 FILLER_38_2112 ();
 sg13g2_decap_8 FILLER_38_2117 ();
 sg13g2_decap_4 FILLER_38_2124 ();
 sg13g2_fill_1 FILLER_38_2155 ();
 sg13g2_fill_2 FILLER_38_2200 ();
 sg13g2_fill_2 FILLER_38_2229 ();
 sg13g2_fill_1 FILLER_38_2293 ();
 sg13g2_decap_4 FILLER_38_2301 ();
 sg13g2_fill_1 FILLER_38_2305 ();
 sg13g2_fill_1 FILLER_38_2319 ();
 sg13g2_decap_8 FILLER_38_2326 ();
 sg13g2_decap_8 FILLER_38_2333 ();
 sg13g2_fill_2 FILLER_38_2363 ();
 sg13g2_fill_1 FILLER_38_2365 ();
 sg13g2_fill_2 FILLER_38_2383 ();
 sg13g2_fill_1 FILLER_38_2385 ();
 sg13g2_decap_8 FILLER_38_2410 ();
 sg13g2_fill_2 FILLER_38_2417 ();
 sg13g2_fill_1 FILLER_38_2431 ();
 sg13g2_decap_8 FILLER_38_2438 ();
 sg13g2_decap_4 FILLER_38_2445 ();
 sg13g2_fill_1 FILLER_38_2449 ();
 sg13g2_decap_4 FILLER_38_2459 ();
 sg13g2_fill_2 FILLER_38_2463 ();
 sg13g2_decap_8 FILLER_38_2486 ();
 sg13g2_decap_4 FILLER_38_2493 ();
 sg13g2_decap_8 FILLER_38_2507 ();
 sg13g2_fill_2 FILLER_38_2514 ();
 sg13g2_fill_1 FILLER_38_2516 ();
 sg13g2_decap_8 FILLER_38_2522 ();
 sg13g2_decap_4 FILLER_38_2529 ();
 sg13g2_decap_8 FILLER_38_2546 ();
 sg13g2_decap_4 FILLER_38_2553 ();
 sg13g2_fill_2 FILLER_38_2557 ();
 sg13g2_fill_1 FILLER_38_2564 ();
 sg13g2_decap_8 FILLER_38_2569 ();
 sg13g2_decap_4 FILLER_38_2576 ();
 sg13g2_fill_2 FILLER_38_2580 ();
 sg13g2_fill_2 FILLER_38_2604 ();
 sg13g2_fill_2 FILLER_38_2616 ();
 sg13g2_fill_2 FILLER_38_2635 ();
 sg13g2_fill_1 FILLER_38_2637 ();
 sg13g2_fill_2 FILLER_38_2656 ();
 sg13g2_fill_1 FILLER_38_2658 ();
 sg13g2_fill_2 FILLER_38_2718 ();
 sg13g2_decap_4 FILLER_38_2740 ();
 sg13g2_fill_2 FILLER_38_2744 ();
 sg13g2_fill_2 FILLER_38_2750 ();
 sg13g2_decap_4 FILLER_38_2757 ();
 sg13g2_fill_1 FILLER_38_2777 ();
 sg13g2_decap_8 FILLER_38_2792 ();
 sg13g2_decap_8 FILLER_38_2799 ();
 sg13g2_fill_2 FILLER_38_2819 ();
 sg13g2_fill_1 FILLER_38_2821 ();
 sg13g2_fill_1 FILLER_38_2835 ();
 sg13g2_decap_4 FILLER_38_2840 ();
 sg13g2_fill_2 FILLER_38_2844 ();
 sg13g2_fill_2 FILLER_38_2857 ();
 sg13g2_decap_8 FILLER_38_2864 ();
 sg13g2_decap_8 FILLER_38_2871 ();
 sg13g2_decap_4 FILLER_38_2878 ();
 sg13g2_fill_1 FILLER_38_2882 ();
 sg13g2_fill_2 FILLER_38_2886 ();
 sg13g2_fill_1 FILLER_38_2888 ();
 sg13g2_decap_8 FILLER_38_2894 ();
 sg13g2_decap_8 FILLER_38_2901 ();
 sg13g2_decap_8 FILLER_38_2908 ();
 sg13g2_fill_1 FILLER_38_2919 ();
 sg13g2_fill_2 FILLER_38_2946 ();
 sg13g2_decap_4 FILLER_38_2984 ();
 sg13g2_fill_1 FILLER_38_2988 ();
 sg13g2_fill_1 FILLER_38_3016 ();
 sg13g2_decap_8 FILLER_38_3044 ();
 sg13g2_decap_8 FILLER_38_3087 ();
 sg13g2_fill_2 FILLER_38_3094 ();
 sg13g2_fill_1 FILLER_38_3096 ();
 sg13g2_fill_2 FILLER_38_3115 ();
 sg13g2_fill_1 FILLER_38_3117 ();
 sg13g2_fill_2 FILLER_38_3123 ();
 sg13g2_fill_2 FILLER_38_3170 ();
 sg13g2_fill_1 FILLER_38_3172 ();
 sg13g2_decap_8 FILLER_38_3233 ();
 sg13g2_fill_2 FILLER_38_3240 ();
 sg13g2_fill_1 FILLER_38_3242 ();
 sg13g2_decap_8 FILLER_38_3256 ();
 sg13g2_decap_4 FILLER_38_3263 ();
 sg13g2_fill_1 FILLER_38_3267 ();
 sg13g2_decap_4 FILLER_38_3278 ();
 sg13g2_fill_2 FILLER_38_3282 ();
 sg13g2_decap_4 FILLER_38_3291 ();
 sg13g2_fill_2 FILLER_38_3295 ();
 sg13g2_decap_8 FILLER_38_3305 ();
 sg13g2_decap_4 FILLER_38_3312 ();
 sg13g2_fill_2 FILLER_38_3316 ();
 sg13g2_fill_2 FILLER_38_3328 ();
 sg13g2_fill_1 FILLER_38_3330 ();
 sg13g2_decap_4 FILLER_38_3344 ();
 sg13g2_fill_1 FILLER_38_3348 ();
 sg13g2_decap_8 FILLER_38_3361 ();
 sg13g2_fill_2 FILLER_38_3368 ();
 sg13g2_fill_1 FILLER_38_3370 ();
 sg13g2_decap_4 FILLER_38_3375 ();
 sg13g2_fill_1 FILLER_38_3379 ();
 sg13g2_decap_8 FILLER_38_3393 ();
 sg13g2_decap_8 FILLER_38_3413 ();
 sg13g2_decap_8 FILLER_38_3420 ();
 sg13g2_fill_2 FILLER_38_3433 ();
 sg13g2_decap_8 FILLER_38_3462 ();
 sg13g2_decap_8 FILLER_38_3469 ();
 sg13g2_decap_8 FILLER_38_3476 ();
 sg13g2_decap_8 FILLER_38_3483 ();
 sg13g2_decap_8 FILLER_38_3490 ();
 sg13g2_decap_8 FILLER_38_3497 ();
 sg13g2_decap_8 FILLER_38_3504 ();
 sg13g2_decap_8 FILLER_38_3511 ();
 sg13g2_decap_8 FILLER_38_3518 ();
 sg13g2_decap_8 FILLER_38_3525 ();
 sg13g2_decap_8 FILLER_38_3532 ();
 sg13g2_decap_8 FILLER_38_3539 ();
 sg13g2_decap_8 FILLER_38_3546 ();
 sg13g2_decap_8 FILLER_38_3553 ();
 sg13g2_decap_8 FILLER_38_3560 ();
 sg13g2_decap_8 FILLER_38_3567 ();
 sg13g2_decap_4 FILLER_38_3574 ();
 sg13g2_fill_2 FILLER_38_3578 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_124 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_154 ();
 sg13g2_decap_4 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_223 ();
 sg13g2_decap_8 FILLER_39_230 ();
 sg13g2_decap_8 FILLER_39_237 ();
 sg13g2_fill_2 FILLER_39_244 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_fill_2 FILLER_39_280 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_fill_1 FILLER_39_323 ();
 sg13g2_fill_1 FILLER_39_338 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_39_414 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_fill_1 FILLER_39_448 ();
 sg13g2_fill_1 FILLER_39_454 ();
 sg13g2_fill_2 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_472 ();
 sg13g2_fill_1 FILLER_39_479 ();
 sg13g2_decap_8 FILLER_39_484 ();
 sg13g2_fill_1 FILLER_39_491 ();
 sg13g2_fill_2 FILLER_39_497 ();
 sg13g2_fill_1 FILLER_39_521 ();
 sg13g2_fill_1 FILLER_39_534 ();
 sg13g2_fill_2 FILLER_39_552 ();
 sg13g2_fill_1 FILLER_39_554 ();
 sg13g2_fill_2 FILLER_39_564 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_613 ();
 sg13g2_fill_1 FILLER_39_620 ();
 sg13g2_decap_4 FILLER_39_723 ();
 sg13g2_fill_2 FILLER_39_727 ();
 sg13g2_fill_2 FILLER_39_733 ();
 sg13g2_fill_1 FILLER_39_735 ();
 sg13g2_fill_2 FILLER_39_765 ();
 sg13g2_fill_1 FILLER_39_767 ();
 sg13g2_decap_4 FILLER_39_787 ();
 sg13g2_fill_1 FILLER_39_791 ();
 sg13g2_fill_1 FILLER_39_820 ();
 sg13g2_fill_1 FILLER_39_830 ();
 sg13g2_fill_2 FILLER_39_888 ();
 sg13g2_decap_4 FILLER_39_899 ();
 sg13g2_fill_2 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_921 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_fill_2 FILLER_39_935 ();
 sg13g2_fill_1 FILLER_39_947 ();
 sg13g2_decap_4 FILLER_39_951 ();
 sg13g2_fill_2 FILLER_39_955 ();
 sg13g2_decap_4 FILLER_39_960 ();
 sg13g2_fill_2 FILLER_39_964 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_fill_2 FILLER_39_994 ();
 sg13g2_decap_4 FILLER_39_1016 ();
 sg13g2_fill_2 FILLER_39_1020 ();
 sg13g2_fill_2 FILLER_39_1032 ();
 sg13g2_fill_1 FILLER_39_1039 ();
 sg13g2_decap_8 FILLER_39_1060 ();
 sg13g2_decap_4 FILLER_39_1088 ();
 sg13g2_fill_1 FILLER_39_1092 ();
 sg13g2_fill_2 FILLER_39_1100 ();
 sg13g2_fill_1 FILLER_39_1102 ();
 sg13g2_decap_4 FILLER_39_1129 ();
 sg13g2_fill_1 FILLER_39_1133 ();
 sg13g2_fill_1 FILLER_39_1147 ();
 sg13g2_fill_1 FILLER_39_1152 ();
 sg13g2_fill_2 FILLER_39_1158 ();
 sg13g2_decap_8 FILLER_39_1176 ();
 sg13g2_fill_2 FILLER_39_1183 ();
 sg13g2_fill_1 FILLER_39_1185 ();
 sg13g2_fill_2 FILLER_39_1207 ();
 sg13g2_fill_1 FILLER_39_1209 ();
 sg13g2_decap_8 FILLER_39_1231 ();
 sg13g2_decap_4 FILLER_39_1243 ();
 sg13g2_fill_2 FILLER_39_1247 ();
 sg13g2_decap_8 FILLER_39_1255 ();
 sg13g2_decap_4 FILLER_39_1262 ();
 sg13g2_fill_1 FILLER_39_1266 ();
 sg13g2_decap_4 FILLER_39_1312 ();
 sg13g2_fill_1 FILLER_39_1316 ();
 sg13g2_decap_4 FILLER_39_1346 ();
 sg13g2_decap_8 FILLER_39_1358 ();
 sg13g2_fill_2 FILLER_39_1365 ();
 sg13g2_fill_1 FILLER_39_1372 ();
 sg13g2_decap_8 FILLER_39_1385 ();
 sg13g2_fill_1 FILLER_39_1392 ();
 sg13g2_decap_4 FILLER_39_1406 ();
 sg13g2_decap_8 FILLER_39_1437 ();
 sg13g2_decap_4 FILLER_39_1444 ();
 sg13g2_fill_2 FILLER_39_1448 ();
 sg13g2_fill_2 FILLER_39_1486 ();
 sg13g2_fill_1 FILLER_39_1488 ();
 sg13g2_decap_4 FILLER_39_1510 ();
 sg13g2_fill_2 FILLER_39_1534 ();
 sg13g2_decap_4 FILLER_39_1549 ();
 sg13g2_fill_1 FILLER_39_1561 ();
 sg13g2_fill_2 FILLER_39_1572 ();
 sg13g2_decap_4 FILLER_39_1591 ();
 sg13g2_fill_1 FILLER_39_1595 ();
 sg13g2_decap_8 FILLER_39_1608 ();
 sg13g2_fill_2 FILLER_39_1615 ();
 sg13g2_fill_1 FILLER_39_1617 ();
 sg13g2_decap_8 FILLER_39_1632 ();
 sg13g2_decap_8 FILLER_39_1639 ();
 sg13g2_fill_2 FILLER_39_1650 ();
 sg13g2_fill_1 FILLER_39_1652 ();
 sg13g2_fill_1 FILLER_39_1662 ();
 sg13g2_fill_1 FILLER_39_1672 ();
 sg13g2_decap_8 FILLER_39_1687 ();
 sg13g2_fill_1 FILLER_39_1694 ();
 sg13g2_fill_2 FILLER_39_1711 ();
 sg13g2_fill_1 FILLER_39_1713 ();
 sg13g2_fill_2 FILLER_39_1745 ();
 sg13g2_fill_1 FILLER_39_1747 ();
 sg13g2_decap_8 FILLER_39_1783 ();
 sg13g2_decap_8 FILLER_39_1790 ();
 sg13g2_fill_2 FILLER_39_1797 ();
 sg13g2_fill_1 FILLER_39_1799 ();
 sg13g2_fill_2 FILLER_39_1809 ();
 sg13g2_fill_1 FILLER_39_1811 ();
 sg13g2_fill_1 FILLER_39_1817 ();
 sg13g2_decap_8 FILLER_39_1823 ();
 sg13g2_decap_4 FILLER_39_1834 ();
 sg13g2_fill_1 FILLER_39_1838 ();
 sg13g2_decap_8 FILLER_39_1852 ();
 sg13g2_decap_8 FILLER_39_1890 ();
 sg13g2_decap_4 FILLER_39_1897 ();
 sg13g2_fill_2 FILLER_39_1905 ();
 sg13g2_fill_1 FILLER_39_1907 ();
 sg13g2_fill_2 FILLER_39_1913 ();
 sg13g2_decap_4 FILLER_39_1942 ();
 sg13g2_fill_2 FILLER_39_1987 ();
 sg13g2_fill_2 FILLER_39_1996 ();
 sg13g2_decap_4 FILLER_39_2007 ();
 sg13g2_fill_2 FILLER_39_2019 ();
 sg13g2_decap_8 FILLER_39_2079 ();
 sg13g2_decap_8 FILLER_39_2086 ();
 sg13g2_decap_8 FILLER_39_2093 ();
 sg13g2_fill_1 FILLER_39_2100 ();
 sg13g2_fill_2 FILLER_39_2137 ();
 sg13g2_decap_8 FILLER_39_2157 ();
 sg13g2_decap_8 FILLER_39_2164 ();
 sg13g2_fill_2 FILLER_39_2171 ();
 sg13g2_decap_8 FILLER_39_2186 ();
 sg13g2_decap_8 FILLER_39_2193 ();
 sg13g2_fill_2 FILLER_39_2200 ();
 sg13g2_decap_8 FILLER_39_2216 ();
 sg13g2_fill_2 FILLER_39_2223 ();
 sg13g2_fill_2 FILLER_39_2259 ();
 sg13g2_decap_8 FILLER_39_2283 ();
 sg13g2_fill_2 FILLER_39_2290 ();
 sg13g2_fill_1 FILLER_39_2364 ();
 sg13g2_fill_2 FILLER_39_2372 ();
 sg13g2_decap_8 FILLER_39_2400 ();
 sg13g2_decap_8 FILLER_39_2407 ();
 sg13g2_decap_4 FILLER_39_2414 ();
 sg13g2_decap_4 FILLER_39_2423 ();
 sg13g2_fill_1 FILLER_39_2445 ();
 sg13g2_decap_4 FILLER_39_2468 ();
 sg13g2_fill_2 FILLER_39_2472 ();
 sg13g2_decap_4 FILLER_39_2488 ();
 sg13g2_fill_1 FILLER_39_2492 ();
 sg13g2_decap_4 FILLER_39_2525 ();
 sg13g2_decap_4 FILLER_39_2600 ();
 sg13g2_fill_1 FILLER_39_2626 ();
 sg13g2_decap_4 FILLER_39_2632 ();
 sg13g2_fill_2 FILLER_39_2641 ();
 sg13g2_fill_1 FILLER_39_2648 ();
 sg13g2_fill_1 FILLER_39_2653 ();
 sg13g2_decap_8 FILLER_39_2675 ();
 sg13g2_fill_2 FILLER_39_2682 ();
 sg13g2_decap_8 FILLER_39_2688 ();
 sg13g2_fill_2 FILLER_39_2695 ();
 sg13g2_fill_1 FILLER_39_2722 ();
 sg13g2_decap_8 FILLER_39_2731 ();
 sg13g2_fill_2 FILLER_39_2738 ();
 sg13g2_fill_1 FILLER_39_2740 ();
 sg13g2_fill_1 FILLER_39_2765 ();
 sg13g2_decap_8 FILLER_39_2771 ();
 sg13g2_decap_4 FILLER_39_2778 ();
 sg13g2_fill_2 FILLER_39_2782 ();
 sg13g2_decap_8 FILLER_39_2801 ();
 sg13g2_decap_4 FILLER_39_2808 ();
 sg13g2_decap_8 FILLER_39_2830 ();
 sg13g2_fill_2 FILLER_39_2837 ();
 sg13g2_decap_4 FILLER_39_2844 ();
 sg13g2_fill_1 FILLER_39_2848 ();
 sg13g2_decap_4 FILLER_39_2852 ();
 sg13g2_fill_2 FILLER_39_2892 ();
 sg13g2_fill_1 FILLER_39_2907 ();
 sg13g2_fill_2 FILLER_39_2940 ();
 sg13g2_fill_2 FILLER_39_2946 ();
 sg13g2_fill_1 FILLER_39_2948 ();
 sg13g2_fill_1 FILLER_39_2971 ();
 sg13g2_decap_8 FILLER_39_3002 ();
 sg13g2_decap_4 FILLER_39_3009 ();
 sg13g2_decap_4 FILLER_39_3025 ();
 sg13g2_fill_1 FILLER_39_3029 ();
 sg13g2_fill_1 FILLER_39_3048 ();
 sg13g2_fill_1 FILLER_39_3068 ();
 sg13g2_decap_4 FILLER_39_3082 ();
 sg13g2_fill_2 FILLER_39_3086 ();
 sg13g2_decap_8 FILLER_39_3097 ();
 sg13g2_decap_4 FILLER_39_3104 ();
 sg13g2_decap_4 FILLER_39_3172 ();
 sg13g2_fill_2 FILLER_39_3176 ();
 sg13g2_decap_8 FILLER_39_3223 ();
 sg13g2_decap_4 FILLER_39_3230 ();
 sg13g2_fill_2 FILLER_39_3262 ();
 sg13g2_decap_8 FILLER_39_3304 ();
 sg13g2_fill_2 FILLER_39_3311 ();
 sg13g2_fill_2 FILLER_39_3330 ();
 sg13g2_decap_8 FILLER_39_3369 ();
 sg13g2_decap_4 FILLER_39_3376 ();
 sg13g2_decap_4 FILLER_39_3385 ();
 sg13g2_fill_2 FILLER_39_3389 ();
 sg13g2_fill_2 FILLER_39_3396 ();
 sg13g2_fill_1 FILLER_39_3398 ();
 sg13g2_fill_1 FILLER_39_3422 ();
 sg13g2_fill_2 FILLER_39_3437 ();
 sg13g2_decap_8 FILLER_39_3452 ();
 sg13g2_decap_8 FILLER_39_3459 ();
 sg13g2_decap_8 FILLER_39_3466 ();
 sg13g2_decap_8 FILLER_39_3473 ();
 sg13g2_decap_8 FILLER_39_3480 ();
 sg13g2_decap_8 FILLER_39_3487 ();
 sg13g2_decap_8 FILLER_39_3494 ();
 sg13g2_decap_8 FILLER_39_3501 ();
 sg13g2_decap_8 FILLER_39_3508 ();
 sg13g2_decap_8 FILLER_39_3515 ();
 sg13g2_decap_8 FILLER_39_3522 ();
 sg13g2_decap_8 FILLER_39_3529 ();
 sg13g2_decap_8 FILLER_39_3536 ();
 sg13g2_decap_8 FILLER_39_3543 ();
 sg13g2_decap_8 FILLER_39_3550 ();
 sg13g2_decap_8 FILLER_39_3557 ();
 sg13g2_decap_8 FILLER_39_3564 ();
 sg13g2_decap_8 FILLER_39_3571 ();
 sg13g2_fill_2 FILLER_39_3578 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_112 ();
 sg13g2_fill_1 FILLER_40_114 ();
 sg13g2_fill_2 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_145 ();
 sg13g2_decap_8 FILLER_40_178 ();
 sg13g2_fill_1 FILLER_40_185 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_decap_8 FILLER_40_270 ();
 sg13g2_decap_4 FILLER_40_277 ();
 sg13g2_decap_8 FILLER_40_291 ();
 sg13g2_fill_2 FILLER_40_298 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_fill_2 FILLER_40_349 ();
 sg13g2_fill_2 FILLER_40_371 ();
 sg13g2_fill_2 FILLER_40_395 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_fill_2 FILLER_40_417 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_decap_4 FILLER_40_485 ();
 sg13g2_fill_2 FILLER_40_512 ();
 sg13g2_fill_1 FILLER_40_514 ();
 sg13g2_fill_2 FILLER_40_539 ();
 sg13g2_fill_1 FILLER_40_541 ();
 sg13g2_fill_2 FILLER_40_567 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_fill_2 FILLER_40_583 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_decap_4 FILLER_40_590 ();
 sg13g2_fill_2 FILLER_40_594 ();
 sg13g2_decap_8 FILLER_40_614 ();
 sg13g2_fill_2 FILLER_40_634 ();
 sg13g2_fill_2 FILLER_40_640 ();
 sg13g2_fill_1 FILLER_40_642 ();
 sg13g2_fill_2 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_650 ();
 sg13g2_decap_8 FILLER_40_656 ();
 sg13g2_fill_2 FILLER_40_663 ();
 sg13g2_fill_2 FILLER_40_693 ();
 sg13g2_fill_1 FILLER_40_695 ();
 sg13g2_decap_4 FILLER_40_718 ();
 sg13g2_fill_2 FILLER_40_722 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_fill_2 FILLER_40_785 ();
 sg13g2_fill_1 FILLER_40_787 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_4 FILLER_40_810 ();
 sg13g2_fill_2 FILLER_40_814 ();
 sg13g2_fill_2 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_fill_2 FILLER_40_852 ();
 sg13g2_fill_1 FILLER_40_854 ();
 sg13g2_decap_4 FILLER_40_878 ();
 sg13g2_fill_1 FILLER_40_882 ();
 sg13g2_fill_1 FILLER_40_888 ();
 sg13g2_decap_4 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_fill_2 FILLER_40_966 ();
 sg13g2_decap_4 FILLER_40_1011 ();
 sg13g2_fill_1 FILLER_40_1015 ();
 sg13g2_decap_4 FILLER_40_1032 ();
 sg13g2_fill_1 FILLER_40_1046 ();
 sg13g2_decap_8 FILLER_40_1052 ();
 sg13g2_decap_4 FILLER_40_1059 ();
 sg13g2_fill_2 FILLER_40_1063 ();
 sg13g2_fill_1 FILLER_40_1074 ();
 sg13g2_decap_4 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1091 ();
 sg13g2_decap_4 FILLER_40_1100 ();
 sg13g2_fill_1 FILLER_40_1109 ();
 sg13g2_fill_2 FILLER_40_1121 ();
 sg13g2_decap_4 FILLER_40_1156 ();
 sg13g2_fill_2 FILLER_40_1160 ();
 sg13g2_decap_4 FILLER_40_1209 ();
 sg13g2_fill_1 FILLER_40_1213 ();
 sg13g2_fill_2 FILLER_40_1231 ();
 sg13g2_fill_1 FILLER_40_1233 ();
 sg13g2_decap_8 FILLER_40_1283 ();
 sg13g2_decap_4 FILLER_40_1290 ();
 sg13g2_decap_4 FILLER_40_1302 ();
 sg13g2_fill_2 FILLER_40_1306 ();
 sg13g2_decap_8 FILLER_40_1317 ();
 sg13g2_fill_2 FILLER_40_1324 ();
 sg13g2_fill_1 FILLER_40_1326 ();
 sg13g2_decap_8 FILLER_40_1337 ();
 sg13g2_decap_4 FILLER_40_1344 ();
 sg13g2_fill_2 FILLER_40_1348 ();
 sg13g2_fill_1 FILLER_40_1409 ();
 sg13g2_fill_1 FILLER_40_1428 ();
 sg13g2_decap_8 FILLER_40_1436 ();
 sg13g2_decap_8 FILLER_40_1443 ();
 sg13g2_fill_2 FILLER_40_1477 ();
 sg13g2_fill_1 FILLER_40_1479 ();
 sg13g2_decap_8 FILLER_40_1485 ();
 sg13g2_decap_4 FILLER_40_1492 ();
 sg13g2_fill_2 FILLER_40_1496 ();
 sg13g2_decap_4 FILLER_40_1536 ();
 sg13g2_fill_2 FILLER_40_1540 ();
 sg13g2_fill_2 FILLER_40_1547 ();
 sg13g2_fill_1 FILLER_40_1549 ();
 sg13g2_decap_4 FILLER_40_1555 ();
 sg13g2_fill_1 FILLER_40_1559 ();
 sg13g2_fill_2 FILLER_40_1565 ();
 sg13g2_fill_2 FILLER_40_1571 ();
 sg13g2_fill_1 FILLER_40_1573 ();
 sg13g2_decap_4 FILLER_40_1579 ();
 sg13g2_fill_1 FILLER_40_1587 ();
 sg13g2_fill_2 FILLER_40_1596 ();
 sg13g2_fill_1 FILLER_40_1658 ();
 sg13g2_fill_1 FILLER_40_1687 ();
 sg13g2_decap_8 FILLER_40_1693 ();
 sg13g2_decap_8 FILLER_40_1700 ();
 sg13g2_decap_4 FILLER_40_1707 ();
 sg13g2_fill_2 FILLER_40_1716 ();
 sg13g2_fill_1 FILLER_40_1812 ();
 sg13g2_fill_1 FILLER_40_1822 ();
 sg13g2_fill_2 FILLER_40_1831 ();
 sg13g2_fill_1 FILLER_40_1833 ();
 sg13g2_fill_2 FILLER_40_1879 ();
 sg13g2_fill_1 FILLER_40_1884 ();
 sg13g2_fill_1 FILLER_40_1912 ();
 sg13g2_fill_2 FILLER_40_1922 ();
 sg13g2_fill_2 FILLER_40_1929 ();
 sg13g2_fill_1 FILLER_40_1945 ();
 sg13g2_fill_2 FILLER_40_1959 ();
 sg13g2_fill_1 FILLER_40_1961 ();
 sg13g2_decap_4 FILLER_40_1965 ();
 sg13g2_fill_1 FILLER_40_1969 ();
 sg13g2_fill_1 FILLER_40_2046 ();
 sg13g2_fill_1 FILLER_40_2065 ();
 sg13g2_decap_8 FILLER_40_2094 ();
 sg13g2_decap_8 FILLER_40_2123 ();
 sg13g2_decap_4 FILLER_40_2130 ();
 sg13g2_fill_1 FILLER_40_2174 ();
 sg13g2_fill_2 FILLER_40_2179 ();
 sg13g2_decap_8 FILLER_40_2219 ();
 sg13g2_fill_2 FILLER_40_2226 ();
 sg13g2_fill_1 FILLER_40_2238 ();
 sg13g2_decap_8 FILLER_40_2297 ();
 sg13g2_decap_8 FILLER_40_2308 ();
 sg13g2_decap_4 FILLER_40_2315 ();
 sg13g2_fill_2 FILLER_40_2319 ();
 sg13g2_decap_4 FILLER_40_2328 ();
 sg13g2_fill_2 FILLER_40_2332 ();
 sg13g2_decap_4 FILLER_40_2339 ();
 sg13g2_decap_8 FILLER_40_2359 ();
 sg13g2_decap_8 FILLER_40_2366 ();
 sg13g2_fill_1 FILLER_40_2378 ();
 sg13g2_fill_1 FILLER_40_2385 ();
 sg13g2_decap_8 FILLER_40_2398 ();
 sg13g2_decap_4 FILLER_40_2405 ();
 sg13g2_fill_2 FILLER_40_2409 ();
 sg13g2_fill_2 FILLER_40_2429 ();
 sg13g2_fill_1 FILLER_40_2431 ();
 sg13g2_fill_1 FILLER_40_2448 ();
 sg13g2_fill_1 FILLER_40_2454 ();
 sg13g2_fill_1 FILLER_40_2460 ();
 sg13g2_fill_2 FILLER_40_2465 ();
 sg13g2_decap_8 FILLER_40_2484 ();
 sg13g2_fill_2 FILLER_40_2491 ();
 sg13g2_fill_2 FILLER_40_2499 ();
 sg13g2_decap_8 FILLER_40_2546 ();
 sg13g2_decap_4 FILLER_40_2553 ();
 sg13g2_decap_8 FILLER_40_2588 ();
 sg13g2_fill_1 FILLER_40_2595 ();
 sg13g2_fill_2 FILLER_40_2607 ();
 sg13g2_fill_2 FILLER_40_2619 ();
 sg13g2_decap_4 FILLER_40_2626 ();
 sg13g2_decap_4 FILLER_40_2636 ();
 sg13g2_fill_1 FILLER_40_2649 ();
 sg13g2_decap_4 FILLER_40_2658 ();
 sg13g2_fill_2 FILLER_40_2670 ();
 sg13g2_fill_1 FILLER_40_2672 ();
 sg13g2_decap_4 FILLER_40_2680 ();
 sg13g2_fill_2 FILLER_40_2684 ();
 sg13g2_fill_2 FILLER_40_2699 ();
 sg13g2_fill_1 FILLER_40_2701 ();
 sg13g2_fill_2 FILLER_40_2751 ();
 sg13g2_fill_1 FILLER_40_2753 ();
 sg13g2_fill_1 FILLER_40_2765 ();
 sg13g2_decap_8 FILLER_40_2778 ();
 sg13g2_decap_4 FILLER_40_2785 ();
 sg13g2_decap_8 FILLER_40_2802 ();
 sg13g2_decap_8 FILLER_40_2858 ();
 sg13g2_fill_2 FILLER_40_2865 ();
 sg13g2_decap_4 FILLER_40_2875 ();
 sg13g2_decap_8 FILLER_40_2915 ();
 sg13g2_decap_4 FILLER_40_2922 ();
 sg13g2_fill_1 FILLER_40_2926 ();
 sg13g2_decap_8 FILLER_40_2932 ();
 sg13g2_decap_8 FILLER_40_2939 ();
 sg13g2_fill_2 FILLER_40_2946 ();
 sg13g2_decap_8 FILLER_40_2985 ();
 sg13g2_fill_2 FILLER_40_2992 ();
 sg13g2_fill_1 FILLER_40_2998 ();
 sg13g2_decap_8 FILLER_40_3008 ();
 sg13g2_fill_1 FILLER_40_3019 ();
 sg13g2_fill_2 FILLER_40_3091 ();
 sg13g2_fill_1 FILLER_40_3093 ();
 sg13g2_fill_1 FILLER_40_3103 ();
 sg13g2_fill_2 FILLER_40_3108 ();
 sg13g2_fill_2 FILLER_40_3119 ();
 sg13g2_fill_1 FILLER_40_3121 ();
 sg13g2_decap_4 FILLER_40_3180 ();
 sg13g2_fill_2 FILLER_40_3230 ();
 sg13g2_fill_1 FILLER_40_3232 ();
 sg13g2_fill_2 FILLER_40_3270 ();
 sg13g2_fill_2 FILLER_40_3276 ();
 sg13g2_fill_2 FILLER_40_3286 ();
 sg13g2_fill_1 FILLER_40_3288 ();
 sg13g2_fill_2 FILLER_40_3293 ();
 sg13g2_fill_1 FILLER_40_3295 ();
 sg13g2_decap_8 FILLER_40_3304 ();
 sg13g2_decap_8 FILLER_40_3311 ();
 sg13g2_decap_8 FILLER_40_3327 ();
 sg13g2_decap_8 FILLER_40_3334 ();
 sg13g2_fill_1 FILLER_40_3341 ();
 sg13g2_decap_4 FILLER_40_3347 ();
 sg13g2_fill_2 FILLER_40_3358 ();
 sg13g2_decap_8 FILLER_40_3365 ();
 sg13g2_fill_1 FILLER_40_3372 ();
 sg13g2_fill_2 FILLER_40_3413 ();
 sg13g2_decap_8 FILLER_40_3419 ();
 sg13g2_decap_4 FILLER_40_3426 ();
 sg13g2_decap_4 FILLER_40_3438 ();
 sg13g2_fill_1 FILLER_40_3442 ();
 sg13g2_decap_8 FILLER_40_3471 ();
 sg13g2_decap_8 FILLER_40_3478 ();
 sg13g2_decap_8 FILLER_40_3485 ();
 sg13g2_decap_8 FILLER_40_3492 ();
 sg13g2_decap_8 FILLER_40_3499 ();
 sg13g2_decap_8 FILLER_40_3506 ();
 sg13g2_decap_8 FILLER_40_3513 ();
 sg13g2_decap_8 FILLER_40_3520 ();
 sg13g2_decap_8 FILLER_40_3527 ();
 sg13g2_decap_8 FILLER_40_3534 ();
 sg13g2_decap_8 FILLER_40_3541 ();
 sg13g2_decap_8 FILLER_40_3548 ();
 sg13g2_decap_8 FILLER_40_3555 ();
 sg13g2_decap_8 FILLER_40_3562 ();
 sg13g2_decap_8 FILLER_40_3569 ();
 sg13g2_decap_4 FILLER_40_3576 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_fill_2 FILLER_41_120 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_decap_8 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_fill_2 FILLER_41_166 ();
 sg13g2_decap_4 FILLER_41_182 ();
 sg13g2_fill_1 FILLER_41_186 ();
 sg13g2_fill_1 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_decap_4 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_decap_4 FILLER_41_443 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_4 FILLER_41_471 ();
 sg13g2_decap_4 FILLER_41_483 ();
 sg13g2_fill_1 FILLER_41_487 ();
 sg13g2_decap_8 FILLER_41_512 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_fill_1 FILLER_41_523 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_decap_8 FILLER_41_575 ();
 sg13g2_decap_4 FILLER_41_582 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_fill_2 FILLER_41_601 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_fill_2 FILLER_41_722 ();
 sg13g2_fill_1 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_4 FILLER_41_749 ();
 sg13g2_fill_1 FILLER_41_753 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_4 FILLER_41_766 ();
 sg13g2_fill_1 FILLER_41_770 ();
 sg13g2_fill_1 FILLER_41_796 ();
 sg13g2_fill_2 FILLER_41_801 ();
 sg13g2_fill_2 FILLER_41_817 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_846 ();
 sg13g2_fill_1 FILLER_41_848 ();
 sg13g2_decap_8 FILLER_41_863 ();
 sg13g2_decap_4 FILLER_41_870 ();
 sg13g2_fill_1 FILLER_41_874 ();
 sg13g2_fill_2 FILLER_41_900 ();
 sg13g2_fill_1 FILLER_41_902 ();
 sg13g2_decap_8 FILLER_41_911 ();
 sg13g2_decap_8 FILLER_41_918 ();
 sg13g2_decap_8 FILLER_41_925 ();
 sg13g2_decap_4 FILLER_41_932 ();
 sg13g2_fill_1 FILLER_41_936 ();
 sg13g2_decap_4 FILLER_41_953 ();
 sg13g2_fill_2 FILLER_41_957 ();
 sg13g2_decap_8 FILLER_41_963 ();
 sg13g2_decap_4 FILLER_41_970 ();
 sg13g2_decap_8 FILLER_41_983 ();
 sg13g2_fill_2 FILLER_41_990 ();
 sg13g2_decap_4 FILLER_41_1019 ();
 sg13g2_decap_4 FILLER_41_1027 ();
 sg13g2_decap_8 FILLER_41_1063 ();
 sg13g2_fill_1 FILLER_41_1075 ();
 sg13g2_decap_8 FILLER_41_1085 ();
 sg13g2_fill_2 FILLER_41_1092 ();
 sg13g2_fill_1 FILLER_41_1094 ();
 sg13g2_fill_1 FILLER_41_1123 ();
 sg13g2_decap_8 FILLER_41_1146 ();
 sg13g2_decap_4 FILLER_41_1153 ();
 sg13g2_fill_2 FILLER_41_1169 ();
 sg13g2_decap_8 FILLER_41_1181 ();
 sg13g2_fill_2 FILLER_41_1188 ();
 sg13g2_fill_1 FILLER_41_1190 ();
 sg13g2_fill_2 FILLER_41_1195 ();
 sg13g2_fill_2 FILLER_41_1237 ();
 sg13g2_fill_1 FILLER_41_1239 ();
 sg13g2_fill_2 FILLER_41_1245 ();
 sg13g2_fill_1 FILLER_41_1247 ();
 sg13g2_fill_1 FILLER_41_1288 ();
 sg13g2_decap_4 FILLER_41_1348 ();
 sg13g2_fill_2 FILLER_41_1352 ();
 sg13g2_fill_2 FILLER_41_1359 ();
 sg13g2_fill_2 FILLER_41_1374 ();
 sg13g2_decap_8 FILLER_41_1385 ();
 sg13g2_fill_2 FILLER_41_1392 ();
 sg13g2_fill_1 FILLER_41_1394 ();
 sg13g2_decap_8 FILLER_41_1454 ();
 sg13g2_decap_4 FILLER_41_1461 ();
 sg13g2_fill_1 FILLER_41_1465 ();
 sg13g2_fill_2 FILLER_41_1506 ();
 sg13g2_decap_4 FILLER_41_1521 ();
 sg13g2_fill_1 FILLER_41_1570 ();
 sg13g2_fill_2 FILLER_41_1599 ();
 sg13g2_fill_1 FILLER_41_1611 ();
 sg13g2_decap_8 FILLER_41_1638 ();
 sg13g2_decap_4 FILLER_41_1658 ();
 sg13g2_fill_2 FILLER_41_1662 ();
 sg13g2_decap_4 FILLER_41_1673 ();
 sg13g2_fill_2 FILLER_41_1677 ();
 sg13g2_decap_4 FILLER_41_1723 ();
 sg13g2_fill_1 FILLER_41_1727 ();
 sg13g2_decap_8 FILLER_41_1737 ();
 sg13g2_decap_8 FILLER_41_1744 ();
 sg13g2_decap_8 FILLER_41_1751 ();
 sg13g2_fill_1 FILLER_41_1758 ();
 sg13g2_fill_2 FILLER_41_1768 ();
 sg13g2_fill_1 FILLER_41_1770 ();
 sg13g2_decap_8 FILLER_41_1788 ();
 sg13g2_fill_1 FILLER_41_1795 ();
 sg13g2_fill_1 FILLER_41_1823 ();
 sg13g2_fill_2 FILLER_41_1860 ();
 sg13g2_fill_1 FILLER_41_1862 ();
 sg13g2_decap_4 FILLER_41_1930 ();
 sg13g2_fill_2 FILLER_41_1987 ();
 sg13g2_decap_4 FILLER_41_2007 ();
 sg13g2_decap_8 FILLER_41_2020 ();
 sg13g2_decap_4 FILLER_41_2027 ();
 sg13g2_fill_2 FILLER_41_2031 ();
 sg13g2_decap_4 FILLER_41_2097 ();
 sg13g2_fill_1 FILLER_41_2101 ();
 sg13g2_decap_4 FILLER_41_2138 ();
 sg13g2_fill_2 FILLER_41_2151 ();
 sg13g2_decap_4 FILLER_41_2162 ();
 sg13g2_fill_2 FILLER_41_2206 ();
 sg13g2_decap_4 FILLER_41_2235 ();
 sg13g2_fill_1 FILLER_41_2239 ();
 sg13g2_decap_8 FILLER_41_2281 ();
 sg13g2_decap_8 FILLER_41_2288 ();
 sg13g2_decap_4 FILLER_41_2295 ();
 sg13g2_fill_1 FILLER_41_2344 ();
 sg13g2_fill_2 FILLER_41_2353 ();
 sg13g2_fill_2 FILLER_41_2376 ();
 sg13g2_decap_4 FILLER_41_2396 ();
 sg13g2_decap_4 FILLER_41_2406 ();
 sg13g2_fill_2 FILLER_41_2410 ();
 sg13g2_fill_2 FILLER_41_2425 ();
 sg13g2_decap_4 FILLER_41_2440 ();
 sg13g2_fill_1 FILLER_41_2444 ();
 sg13g2_fill_2 FILLER_41_2449 ();
 sg13g2_decap_8 FILLER_41_2456 ();
 sg13g2_decap_8 FILLER_41_2463 ();
 sg13g2_fill_1 FILLER_41_2498 ();
 sg13g2_decap_4 FILLER_41_2555 ();
 sg13g2_fill_1 FILLER_41_2564 ();
 sg13g2_decap_8 FILLER_41_2593 ();
 sg13g2_fill_1 FILLER_41_2605 ();
 sg13g2_decap_4 FILLER_41_2611 ();
 sg13g2_fill_1 FILLER_41_2615 ();
 sg13g2_decap_4 FILLER_41_2632 ();
 sg13g2_fill_2 FILLER_41_2636 ();
 sg13g2_fill_2 FILLER_41_2661 ();
 sg13g2_fill_2 FILLER_41_2669 ();
 sg13g2_fill_1 FILLER_41_2671 ();
 sg13g2_fill_1 FILLER_41_2700 ();
 sg13g2_decap_8 FILLER_41_2744 ();
 sg13g2_fill_2 FILLER_41_2751 ();
 sg13g2_fill_1 FILLER_41_2753 ();
 sg13g2_fill_2 FILLER_41_2817 ();
 sg13g2_decap_4 FILLER_41_2832 ();
 sg13g2_fill_1 FILLER_41_2836 ();
 sg13g2_fill_2 FILLER_41_2841 ();
 sg13g2_fill_1 FILLER_41_2843 ();
 sg13g2_fill_2 FILLER_41_2903 ();
 sg13g2_fill_1 FILLER_41_2905 ();
 sg13g2_decap_8 FILLER_41_2909 ();
 sg13g2_decap_8 FILLER_41_2916 ();
 sg13g2_fill_2 FILLER_41_3017 ();
 sg13g2_fill_1 FILLER_41_3019 ();
 sg13g2_fill_1 FILLER_41_3025 ();
 sg13g2_fill_2 FILLER_41_3030 ();
 sg13g2_fill_1 FILLER_41_3032 ();
 sg13g2_decap_8 FILLER_41_3046 ();
 sg13g2_decap_8 FILLER_41_3053 ();
 sg13g2_fill_1 FILLER_41_3060 ();
 sg13g2_fill_1 FILLER_41_3103 ();
 sg13g2_fill_2 FILLER_41_3136 ();
 sg13g2_fill_1 FILLER_41_3138 ();
 sg13g2_decap_4 FILLER_41_3161 ();
 sg13g2_fill_2 FILLER_41_3202 ();
 sg13g2_decap_4 FILLER_41_3231 ();
 sg13g2_fill_2 FILLER_41_3235 ();
 sg13g2_fill_2 FILLER_41_3242 ();
 sg13g2_fill_1 FILLER_41_3244 ();
 sg13g2_decap_4 FILLER_41_3267 ();
 sg13g2_fill_1 FILLER_41_3271 ();
 sg13g2_fill_1 FILLER_41_3285 ();
 sg13g2_fill_1 FILLER_41_3291 ();
 sg13g2_decap_4 FILLER_41_3298 ();
 sg13g2_fill_1 FILLER_41_3307 ();
 sg13g2_fill_2 FILLER_41_3325 ();
 sg13g2_fill_1 FILLER_41_3327 ();
 sg13g2_decap_4 FILLER_41_3336 ();
 sg13g2_decap_4 FILLER_41_3353 ();
 sg13g2_decap_4 FILLER_41_3361 ();
 sg13g2_fill_1 FILLER_41_3365 ();
 sg13g2_fill_1 FILLER_41_3371 ();
 sg13g2_fill_1 FILLER_41_3380 ();
 sg13g2_decap_8 FILLER_41_3390 ();
 sg13g2_decap_4 FILLER_41_3397 ();
 sg13g2_fill_2 FILLER_41_3401 ();
 sg13g2_fill_2 FILLER_41_3415 ();
 sg13g2_fill_1 FILLER_41_3417 ();
 sg13g2_fill_1 FILLER_41_3428 ();
 sg13g2_fill_1 FILLER_41_3455 ();
 sg13g2_decap_8 FILLER_41_3465 ();
 sg13g2_decap_8 FILLER_41_3472 ();
 sg13g2_decap_8 FILLER_41_3479 ();
 sg13g2_decap_8 FILLER_41_3486 ();
 sg13g2_decap_8 FILLER_41_3493 ();
 sg13g2_decap_8 FILLER_41_3500 ();
 sg13g2_decap_8 FILLER_41_3507 ();
 sg13g2_decap_8 FILLER_41_3514 ();
 sg13g2_decap_8 FILLER_41_3521 ();
 sg13g2_decap_8 FILLER_41_3528 ();
 sg13g2_decap_8 FILLER_41_3535 ();
 sg13g2_decap_8 FILLER_41_3542 ();
 sg13g2_decap_8 FILLER_41_3549 ();
 sg13g2_decap_8 FILLER_41_3556 ();
 sg13g2_decap_8 FILLER_41_3563 ();
 sg13g2_decap_8 FILLER_41_3570 ();
 sg13g2_fill_2 FILLER_41_3577 ();
 sg13g2_fill_1 FILLER_41_3579 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_4 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_95 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_decap_4 FILLER_42_186 ();
 sg13g2_decap_4 FILLER_42_193 ();
 sg13g2_decap_4 FILLER_42_209 ();
 sg13g2_fill_2 FILLER_42_213 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_296 ();
 sg13g2_decap_4 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_fill_1 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_4 FILLER_42_469 ();
 sg13g2_fill_1 FILLER_42_473 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_fill_2 FILLER_42_490 ();
 sg13g2_fill_1 FILLER_42_519 ();
 sg13g2_fill_2 FILLER_42_527 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_decap_4 FILLER_42_549 ();
 sg13g2_fill_1 FILLER_42_553 ();
 sg13g2_fill_1 FILLER_42_559 ();
 sg13g2_fill_2 FILLER_42_565 ();
 sg13g2_fill_1 FILLER_42_567 ();
 sg13g2_decap_4 FILLER_42_572 ();
 sg13g2_fill_1 FILLER_42_576 ();
 sg13g2_fill_2 FILLER_42_585 ();
 sg13g2_fill_2 FILLER_42_610 ();
 sg13g2_fill_1 FILLER_42_612 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_fill_2 FILLER_42_637 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_decap_8 FILLER_42_653 ();
 sg13g2_decap_8 FILLER_42_660 ();
 sg13g2_fill_2 FILLER_42_703 ();
 sg13g2_fill_2 FILLER_42_732 ();
 sg13g2_fill_1 FILLER_42_734 ();
 sg13g2_decap_8 FILLER_42_771 ();
 sg13g2_fill_2 FILLER_42_778 ();
 sg13g2_fill_1 FILLER_42_798 ();
 sg13g2_decap_4 FILLER_42_808 ();
 sg13g2_fill_1 FILLER_42_812 ();
 sg13g2_fill_1 FILLER_42_817 ();
 sg13g2_fill_1 FILLER_42_822 ();
 sg13g2_fill_2 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_837 ();
 sg13g2_fill_1 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_873 ();
 sg13g2_fill_2 FILLER_42_880 ();
 sg13g2_decap_8 FILLER_42_895 ();
 sg13g2_decap_4 FILLER_42_902 ();
 sg13g2_fill_2 FILLER_42_906 ();
 sg13g2_fill_1 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_932 ();
 sg13g2_fill_2 FILLER_42_939 ();
 sg13g2_fill_1 FILLER_42_941 ();
 sg13g2_decap_4 FILLER_42_945 ();
 sg13g2_decap_4 FILLER_42_985 ();
 sg13g2_fill_2 FILLER_42_989 ();
 sg13g2_fill_1 FILLER_42_1000 ();
 sg13g2_fill_1 FILLER_42_1004 ();
 sg13g2_fill_2 FILLER_42_1026 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_4 FILLER_42_1038 ();
 sg13g2_decap_4 FILLER_42_1054 ();
 sg13g2_fill_1 FILLER_42_1058 ();
 sg13g2_decap_8 FILLER_42_1087 ();
 sg13g2_fill_1 FILLER_42_1094 ();
 sg13g2_decap_8 FILLER_42_1103 ();
 sg13g2_decap_4 FILLER_42_1138 ();
 sg13g2_fill_1 FILLER_42_1142 ();
 sg13g2_fill_2 FILLER_42_1170 ();
 sg13g2_fill_1 FILLER_42_1172 ();
 sg13g2_decap_8 FILLER_42_1200 ();
 sg13g2_decap_4 FILLER_42_1207 ();
 sg13g2_fill_1 FILLER_42_1211 ();
 sg13g2_fill_2 FILLER_42_1230 ();
 sg13g2_decap_4 FILLER_42_1289 ();
 sg13g2_fill_1 FILLER_42_1293 ();
 sg13g2_fill_2 FILLER_42_1310 ();
 sg13g2_fill_1 FILLER_42_1321 ();
 sg13g2_fill_2 FILLER_42_1340 ();
 sg13g2_fill_2 FILLER_42_1356 ();
 sg13g2_fill_1 FILLER_42_1358 ();
 sg13g2_decap_4 FILLER_42_1380 ();
 sg13g2_fill_2 FILLER_42_1384 ();
 sg13g2_fill_2 FILLER_42_1404 ();
 sg13g2_fill_1 FILLER_42_1406 ();
 sg13g2_decap_8 FILLER_42_1420 ();
 sg13g2_decap_8 FILLER_42_1427 ();
 sg13g2_decap_8 FILLER_42_1434 ();
 sg13g2_fill_2 FILLER_42_1441 ();
 sg13g2_fill_2 FILLER_42_1457 ();
 sg13g2_decap_8 FILLER_42_1481 ();
 sg13g2_decap_8 FILLER_42_1488 ();
 sg13g2_decap_8 FILLER_42_1495 ();
 sg13g2_fill_1 FILLER_42_1524 ();
 sg13g2_fill_1 FILLER_42_1556 ();
 sg13g2_fill_2 FILLER_42_1579 ();
 sg13g2_fill_1 FILLER_42_1581 ();
 sg13g2_fill_1 FILLER_42_1627 ();
 sg13g2_fill_2 FILLER_42_1700 ();
 sg13g2_fill_2 FILLER_42_1711 ();
 sg13g2_fill_1 FILLER_42_1799 ();
 sg13g2_fill_2 FILLER_42_1827 ();
 sg13g2_decap_4 FILLER_42_1869 ();
 sg13g2_fill_2 FILLER_42_1873 ();
 sg13g2_fill_2 FILLER_42_1910 ();
 sg13g2_fill_1 FILLER_42_1912 ();
 sg13g2_decap_4 FILLER_42_1949 ();
 sg13g2_fill_1 FILLER_42_1953 ();
 sg13g2_fill_2 FILLER_42_1999 ();
 sg13g2_fill_1 FILLER_42_2037 ();
 sg13g2_decap_8 FILLER_42_2043 ();
 sg13g2_fill_2 FILLER_42_2050 ();
 sg13g2_fill_2 FILLER_42_2061 ();
 sg13g2_fill_1 FILLER_42_2077 ();
 sg13g2_fill_1 FILLER_42_2096 ();
 sg13g2_fill_1 FILLER_42_2102 ();
 sg13g2_decap_4 FILLER_42_2121 ();
 sg13g2_fill_2 FILLER_42_2125 ();
 sg13g2_fill_1 FILLER_42_2177 ();
 sg13g2_decap_4 FILLER_42_2192 ();
 sg13g2_fill_1 FILLER_42_2200 ();
 sg13g2_decap_4 FILLER_42_2219 ();
 sg13g2_fill_2 FILLER_42_2223 ();
 sg13g2_decap_4 FILLER_42_2239 ();
 sg13g2_fill_2 FILLER_42_2247 ();
 sg13g2_fill_1 FILLER_42_2249 ();
 sg13g2_fill_1 FILLER_42_2263 ();
 sg13g2_decap_4 FILLER_42_2291 ();
 sg13g2_fill_1 FILLER_42_2295 ();
 sg13g2_fill_2 FILLER_42_2309 ();
 sg13g2_fill_1 FILLER_42_2311 ();
 sg13g2_fill_1 FILLER_42_2343 ();
 sg13g2_fill_2 FILLER_42_2349 ();
 sg13g2_fill_1 FILLER_42_2351 ();
 sg13g2_fill_2 FILLER_42_2357 ();
 sg13g2_fill_2 FILLER_42_2384 ();
 sg13g2_decap_4 FILLER_42_2406 ();
 sg13g2_fill_2 FILLER_42_2423 ();
 sg13g2_fill_1 FILLER_42_2428 ();
 sg13g2_fill_2 FILLER_42_2434 ();
 sg13g2_fill_1 FILLER_42_2444 ();
 sg13g2_decap_4 FILLER_42_2466 ();
 sg13g2_decap_4 FILLER_42_2492 ();
 sg13g2_fill_1 FILLER_42_2496 ();
 sg13g2_fill_2 FILLER_42_2500 ();
 sg13g2_fill_2 FILLER_42_2509 ();
 sg13g2_decap_4 FILLER_42_2537 ();
 sg13g2_fill_1 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2568 ();
 sg13g2_decap_8 FILLER_42_2575 ();
 sg13g2_decap_8 FILLER_42_2582 ();
 sg13g2_fill_2 FILLER_42_2589 ();
 sg13g2_decap_8 FILLER_42_2604 ();
 sg13g2_decap_4 FILLER_42_2611 ();
 sg13g2_fill_2 FILLER_42_2620 ();
 sg13g2_fill_1 FILLER_42_2622 ();
 sg13g2_decap_8 FILLER_42_2628 ();
 sg13g2_decap_8 FILLER_42_2635 ();
 sg13g2_fill_2 FILLER_42_2642 ();
 sg13g2_fill_2 FILLER_42_2665 ();
 sg13g2_fill_1 FILLER_42_2676 ();
 sg13g2_decap_8 FILLER_42_2681 ();
 sg13g2_decap_4 FILLER_42_2688 ();
 sg13g2_fill_2 FILLER_42_2695 ();
 sg13g2_decap_4 FILLER_42_2764 ();
 sg13g2_fill_2 FILLER_42_2768 ();
 sg13g2_fill_1 FILLER_42_2791 ();
 sg13g2_fill_2 FILLER_42_2864 ();
 sg13g2_decap_4 FILLER_42_2879 ();
 sg13g2_fill_1 FILLER_42_2883 ();
 sg13g2_fill_2 FILLER_42_2893 ();
 sg13g2_fill_1 FILLER_42_2895 ();
 sg13g2_decap_4 FILLER_42_2923 ();
 sg13g2_fill_2 FILLER_42_2934 ();
 sg13g2_decap_8 FILLER_42_2985 ();
 sg13g2_decap_8 FILLER_42_2992 ();
 sg13g2_decap_8 FILLER_42_2999 ();
 sg13g2_decap_8 FILLER_42_3006 ();
 sg13g2_fill_1 FILLER_42_3013 ();
 sg13g2_fill_1 FILLER_42_3055 ();
 sg13g2_fill_2 FILLER_42_3097 ();
 sg13g2_fill_2 FILLER_42_3118 ();
 sg13g2_fill_1 FILLER_42_3170 ();
 sg13g2_decap_8 FILLER_42_3184 ();
 sg13g2_decap_8 FILLER_42_3191 ();
 sg13g2_fill_2 FILLER_42_3208 ();
 sg13g2_fill_1 FILLER_42_3210 ();
 sg13g2_decap_4 FILLER_42_3238 ();
 sg13g2_fill_2 FILLER_42_3247 ();
 sg13g2_decap_8 FILLER_42_3260 ();
 sg13g2_decap_4 FILLER_42_3281 ();
 sg13g2_fill_2 FILLER_42_3289 ();
 sg13g2_fill_1 FILLER_42_3291 ();
 sg13g2_fill_2 FILLER_42_3312 ();
 sg13g2_fill_1 FILLER_42_3314 ();
 sg13g2_decap_8 FILLER_42_3327 ();
 sg13g2_decap_4 FILLER_42_3334 ();
 sg13g2_decap_8 FILLER_42_3352 ();
 sg13g2_decap_4 FILLER_42_3359 ();
 sg13g2_fill_2 FILLER_42_3371 ();
 sg13g2_decap_8 FILLER_42_3394 ();
 sg13g2_fill_1 FILLER_42_3401 ();
 sg13g2_decap_8 FILLER_42_3417 ();
 sg13g2_fill_2 FILLER_42_3424 ();
 sg13g2_decap_8 FILLER_42_3464 ();
 sg13g2_decap_8 FILLER_42_3471 ();
 sg13g2_decap_8 FILLER_42_3478 ();
 sg13g2_decap_8 FILLER_42_3485 ();
 sg13g2_decap_8 FILLER_42_3492 ();
 sg13g2_decap_8 FILLER_42_3499 ();
 sg13g2_decap_8 FILLER_42_3506 ();
 sg13g2_decap_8 FILLER_42_3513 ();
 sg13g2_decap_8 FILLER_42_3520 ();
 sg13g2_decap_8 FILLER_42_3527 ();
 sg13g2_decap_8 FILLER_42_3534 ();
 sg13g2_decap_8 FILLER_42_3541 ();
 sg13g2_decap_8 FILLER_42_3548 ();
 sg13g2_decap_8 FILLER_42_3555 ();
 sg13g2_decap_8 FILLER_42_3562 ();
 sg13g2_decap_8 FILLER_42_3569 ();
 sg13g2_decap_4 FILLER_42_3576 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_136 ();
 sg13g2_fill_2 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_211 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_decap_4 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_4 FILLER_43_364 ();
 sg13g2_fill_2 FILLER_43_368 ();
 sg13g2_decap_4 FILLER_43_387 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_409 ();
 sg13g2_decap_8 FILLER_43_424 ();
 sg13g2_decap_8 FILLER_43_431 ();
 sg13g2_fill_1 FILLER_43_438 ();
 sg13g2_fill_1 FILLER_43_466 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_566 ();
 sg13g2_fill_1 FILLER_43_591 ();
 sg13g2_fill_2 FILLER_43_668 ();
 sg13g2_fill_2 FILLER_43_687 ();
 sg13g2_fill_1 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_733 ();
 sg13g2_fill_2 FILLER_43_754 ();
 sg13g2_fill_1 FILLER_43_756 ();
 sg13g2_decap_4 FILLER_43_766 ();
 sg13g2_decap_4 FILLER_43_816 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_4 FILLER_43_839 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_864 ();
 sg13g2_decap_8 FILLER_43_871 ();
 sg13g2_fill_2 FILLER_43_878 ();
 sg13g2_fill_1 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_888 ();
 sg13g2_fill_1 FILLER_43_895 ();
 sg13g2_decap_4 FILLER_43_964 ();
 sg13g2_fill_1 FILLER_43_968 ();
 sg13g2_fill_2 FILLER_43_1009 ();
 sg13g2_decap_8 FILLER_43_1047 ();
 sg13g2_decap_8 FILLER_43_1054 ();
 sg13g2_fill_2 FILLER_43_1061 ();
 sg13g2_fill_1 FILLER_43_1063 ();
 sg13g2_decap_8 FILLER_43_1080 ();
 sg13g2_fill_1 FILLER_43_1105 ();
 sg13g2_decap_8 FILLER_43_1110 ();
 sg13g2_fill_2 FILLER_43_1126 ();
 sg13g2_fill_1 FILLER_43_1128 ();
 sg13g2_fill_1 FILLER_43_1146 ();
 sg13g2_fill_1 FILLER_43_1173 ();
 sg13g2_fill_2 FILLER_43_1187 ();
 sg13g2_fill_1 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1230 ();
 sg13g2_decap_4 FILLER_43_1424 ();
 sg13g2_fill_1 FILLER_43_1428 ();
 sg13g2_decap_8 FILLER_43_1436 ();
 sg13g2_decap_4 FILLER_43_1443 ();
 sg13g2_fill_1 FILLER_43_1474 ();
 sg13g2_fill_1 FILLER_43_1538 ();
 sg13g2_fill_2 FILLER_43_1569 ();
 sg13g2_fill_2 FILLER_43_1615 ();
 sg13g2_fill_1 FILLER_43_1617 ();
 sg13g2_decap_8 FILLER_43_1663 ();
 sg13g2_decap_4 FILLER_43_1670 ();
 sg13g2_fill_1 FILLER_43_1674 ();
 sg13g2_fill_2 FILLER_43_1688 ();
 sg13g2_decap_8 FILLER_43_1726 ();
 sg13g2_decap_8 FILLER_43_1733 ();
 sg13g2_decap_8 FILLER_43_1744 ();
 sg13g2_decap_8 FILLER_43_1751 ();
 sg13g2_decap_8 FILLER_43_1758 ();
 sg13g2_fill_1 FILLER_43_1765 ();
 sg13g2_decap_8 FILLER_43_1779 ();
 sg13g2_fill_1 FILLER_43_1786 ();
 sg13g2_fill_1 FILLER_43_1830 ();
 sg13g2_fill_2 FILLER_43_1854 ();
 sg13g2_fill_1 FILLER_43_1856 ();
 sg13g2_fill_2 FILLER_43_1914 ();
 sg13g2_fill_2 FILLER_43_1948 ();
 sg13g2_fill_2 FILLER_43_2007 ();
 sg13g2_fill_1 FILLER_43_2009 ();
 sg13g2_fill_1 FILLER_43_2046 ();
 sg13g2_decap_8 FILLER_43_2056 ();
 sg13g2_fill_2 FILLER_43_2063 ();
 sg13g2_decap_4 FILLER_43_2096 ();
 sg13g2_decap_4 FILLER_43_2113 ();
 sg13g2_fill_1 FILLER_43_2117 ();
 sg13g2_fill_2 FILLER_43_2150 ();
 sg13g2_fill_1 FILLER_43_2152 ();
 sg13g2_fill_2 FILLER_43_2184 ();
 sg13g2_fill_1 FILLER_43_2227 ();
 sg13g2_decap_4 FILLER_43_2255 ();
 sg13g2_decap_8 FILLER_43_2268 ();
 sg13g2_decap_4 FILLER_43_2275 ();
 sg13g2_fill_2 FILLER_43_2279 ();
 sg13g2_fill_2 FILLER_43_2298 ();
 sg13g2_fill_2 FILLER_43_2313 ();
 sg13g2_fill_1 FILLER_43_2315 ();
 sg13g2_decap_8 FILLER_43_2335 ();
 sg13g2_fill_2 FILLER_43_2342 ();
 sg13g2_fill_1 FILLER_43_2344 ();
 sg13g2_decap_8 FILLER_43_2349 ();
 sg13g2_decap_4 FILLER_43_2356 ();
 sg13g2_fill_1 FILLER_43_2360 ();
 sg13g2_fill_2 FILLER_43_2377 ();
 sg13g2_decap_4 FILLER_43_2384 ();
 sg13g2_fill_2 FILLER_43_2388 ();
 sg13g2_decap_8 FILLER_43_2408 ();
 sg13g2_fill_2 FILLER_43_2415 ();
 sg13g2_fill_1 FILLER_43_2417 ();
 sg13g2_fill_1 FILLER_43_2427 ();
 sg13g2_fill_2 FILLER_43_2453 ();
 sg13g2_fill_1 FILLER_43_2455 ();
 sg13g2_decap_8 FILLER_43_2464 ();
 sg13g2_fill_2 FILLER_43_2471 ();
 sg13g2_fill_2 FILLER_43_2559 ();
 sg13g2_fill_1 FILLER_43_2561 ();
 sg13g2_fill_2 FILLER_43_2617 ();
 sg13g2_decap_8 FILLER_43_2679 ();
 sg13g2_decap_8 FILLER_43_2733 ();
 sg13g2_decap_8 FILLER_43_2757 ();
 sg13g2_decap_8 FILLER_43_2764 ();
 sg13g2_decap_4 FILLER_43_2771 ();
 sg13g2_fill_1 FILLER_43_2802 ();
 sg13g2_fill_1 FILLER_43_2829 ();
 sg13g2_fill_2 FILLER_43_2853 ();
 sg13g2_fill_1 FILLER_43_2873 ();
 sg13g2_fill_1 FILLER_43_2878 ();
 sg13g2_decap_4 FILLER_43_2897 ();
 sg13g2_decap_4 FILLER_43_2909 ();
 sg13g2_fill_2 FILLER_43_2935 ();
 sg13g2_fill_2 FILLER_43_2950 ();
 sg13g2_fill_1 FILLER_43_2952 ();
 sg13g2_decap_4 FILLER_43_2985 ();
 sg13g2_fill_2 FILLER_43_2993 ();
 sg13g2_decap_8 FILLER_43_3023 ();
 sg13g2_fill_2 FILLER_43_3030 ();
 sg13g2_fill_1 FILLER_43_3032 ();
 sg13g2_fill_1 FILLER_43_3043 ();
 sg13g2_fill_2 FILLER_43_3070 ();
 sg13g2_fill_2 FILLER_43_3114 ();
 sg13g2_fill_1 FILLER_43_3116 ();
 sg13g2_fill_1 FILLER_43_3130 ();
 sg13g2_fill_2 FILLER_43_3158 ();
 sg13g2_decap_4 FILLER_43_3207 ();
 sg13g2_fill_2 FILLER_43_3211 ();
 sg13g2_decap_8 FILLER_43_3231 ();
 sg13g2_fill_1 FILLER_43_3238 ();
 sg13g2_fill_1 FILLER_43_3282 ();
 sg13g2_fill_2 FILLER_43_3327 ();
 sg13g2_decap_4 FILLER_43_3334 ();
 sg13g2_fill_2 FILLER_43_3338 ();
 sg13g2_decap_8 FILLER_43_3352 ();
 sg13g2_fill_1 FILLER_43_3359 ();
 sg13g2_decap_4 FILLER_43_3376 ();
 sg13g2_decap_4 FILLER_43_3390 ();
 sg13g2_fill_2 FILLER_43_3394 ();
 sg13g2_decap_8 FILLER_43_3425 ();
 sg13g2_decap_8 FILLER_43_3432 ();
 sg13g2_fill_2 FILLER_43_3439 ();
 sg13g2_decap_8 FILLER_43_3445 ();
 sg13g2_decap_8 FILLER_43_3452 ();
 sg13g2_decap_8 FILLER_43_3459 ();
 sg13g2_decap_8 FILLER_43_3466 ();
 sg13g2_decap_8 FILLER_43_3473 ();
 sg13g2_decap_8 FILLER_43_3480 ();
 sg13g2_decap_8 FILLER_43_3487 ();
 sg13g2_decap_8 FILLER_43_3494 ();
 sg13g2_decap_8 FILLER_43_3501 ();
 sg13g2_decap_8 FILLER_43_3508 ();
 sg13g2_decap_8 FILLER_43_3515 ();
 sg13g2_decap_8 FILLER_43_3522 ();
 sg13g2_decap_8 FILLER_43_3529 ();
 sg13g2_decap_8 FILLER_43_3536 ();
 sg13g2_decap_8 FILLER_43_3543 ();
 sg13g2_decap_8 FILLER_43_3550 ();
 sg13g2_decap_8 FILLER_43_3557 ();
 sg13g2_decap_8 FILLER_43_3564 ();
 sg13g2_decap_8 FILLER_43_3571 ();
 sg13g2_fill_2 FILLER_43_3578 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_4 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_93 ();
 sg13g2_decap_8 FILLER_44_100 ();
 sg13g2_decap_8 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_116 ();
 sg13g2_decap_4 FILLER_44_155 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_decap_4 FILLER_44_228 ();
 sg13g2_fill_2 FILLER_44_232 ();
 sg13g2_fill_1 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_254 ();
 sg13g2_decap_4 FILLER_44_261 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_decap_4 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_285 ();
 sg13g2_decap_4 FILLER_44_309 ();
 sg13g2_fill_2 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_fill_2 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_428 ();
 sg13g2_decap_4 FILLER_44_435 ();
 sg13g2_decap_8 FILLER_44_444 ();
 sg13g2_decap_4 FILLER_44_495 ();
 sg13g2_fill_2 FILLER_44_504 ();
 sg13g2_fill_1 FILLER_44_506 ();
 sg13g2_fill_2 FILLER_44_520 ();
 sg13g2_fill_1 FILLER_44_555 ();
 sg13g2_fill_2 FILLER_44_565 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_2 FILLER_44_622 ();
 sg13g2_fill_1 FILLER_44_624 ();
 sg13g2_fill_1 FILLER_44_639 ();
 sg13g2_fill_1 FILLER_44_654 ();
 sg13g2_fill_2 FILLER_44_725 ();
 sg13g2_fill_1 FILLER_44_727 ();
 sg13g2_fill_2 FILLER_44_774 ();
 sg13g2_fill_1 FILLER_44_776 ();
 sg13g2_decap_4 FILLER_44_787 ();
 sg13g2_fill_2 FILLER_44_791 ();
 sg13g2_fill_2 FILLER_44_797 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_950 ();
 sg13g2_decap_8 FILLER_44_957 ();
 sg13g2_fill_2 FILLER_44_964 ();
 sg13g2_fill_2 FILLER_44_970 ();
 sg13g2_fill_2 FILLER_44_1010 ();
 sg13g2_decap_4 FILLER_44_1058 ();
 sg13g2_decap_4 FILLER_44_1093 ();
 sg13g2_fill_1 FILLER_44_1097 ();
 sg13g2_fill_2 FILLER_44_1126 ();
 sg13g2_fill_2 FILLER_44_1173 ();
 sg13g2_fill_2 FILLER_44_1180 ();
 sg13g2_fill_1 FILLER_44_1182 ();
 sg13g2_fill_1 FILLER_44_1228 ();
 sg13g2_decap_8 FILLER_44_1256 ();
 sg13g2_fill_1 FILLER_44_1263 ();
 sg13g2_fill_2 FILLER_44_1290 ();
 sg13g2_fill_1 FILLER_44_1292 ();
 sg13g2_fill_2 FILLER_44_1298 ();
 sg13g2_fill_1 FILLER_44_1300 ();
 sg13g2_decap_8 FILLER_44_1314 ();
 sg13g2_decap_8 FILLER_44_1321 ();
 sg13g2_fill_2 FILLER_44_1328 ();
 sg13g2_fill_1 FILLER_44_1330 ();
 sg13g2_fill_2 FILLER_44_1335 ();
 sg13g2_fill_1 FILLER_44_1337 ();
 sg13g2_fill_2 FILLER_44_1426 ();
 sg13g2_fill_1 FILLER_44_1428 ();
 sg13g2_decap_4 FILLER_44_1456 ();
 sg13g2_fill_2 FILLER_44_1478 ();
 sg13g2_fill_1 FILLER_44_1480 ();
 sg13g2_decap_8 FILLER_44_1503 ();
 sg13g2_fill_2 FILLER_44_1560 ();
 sg13g2_decap_8 FILLER_44_1571 ();
 sg13g2_decap_8 FILLER_44_1578 ();
 sg13g2_decap_4 FILLER_44_1585 ();
 sg13g2_fill_2 FILLER_44_1589 ();
 sg13g2_decap_8 FILLER_44_1711 ();
 sg13g2_decap_8 FILLER_44_1718 ();
 sg13g2_decap_8 FILLER_44_1725 ();
 sg13g2_fill_1 FILLER_44_1732 ();
 sg13g2_fill_2 FILLER_44_1761 ();
 sg13g2_fill_1 FILLER_44_1763 ();
 sg13g2_decap_8 FILLER_44_1769 ();
 sg13g2_fill_2 FILLER_44_1776 ();
 sg13g2_fill_1 FILLER_44_1778 ();
 sg13g2_fill_2 FILLER_44_1834 ();
 sg13g2_fill_2 FILLER_44_1903 ();
 sg13g2_decap_4 FILLER_44_1936 ();
 sg13g2_decap_8 FILLER_44_1949 ();
 sg13g2_decap_8 FILLER_44_1956 ();
 sg13g2_decap_4 FILLER_44_1963 ();
 sg13g2_fill_1 FILLER_44_1967 ();
 sg13g2_fill_2 FILLER_44_2000 ();
 sg13g2_decap_4 FILLER_44_2038 ();
 sg13g2_fill_2 FILLER_44_2078 ();
 sg13g2_fill_1 FILLER_44_2080 ();
 sg13g2_decap_4 FILLER_44_2094 ();
 sg13g2_fill_1 FILLER_44_2098 ();
 sg13g2_fill_2 FILLER_44_2142 ();
 sg13g2_fill_1 FILLER_44_2144 ();
 sg13g2_decap_8 FILLER_44_2154 ();
 sg13g2_decap_4 FILLER_44_2161 ();
 sg13g2_fill_1 FILLER_44_2165 ();
 sg13g2_fill_2 FILLER_44_2179 ();
 sg13g2_fill_2 FILLER_44_2190 ();
 sg13g2_fill_1 FILLER_44_2192 ();
 sg13g2_fill_2 FILLER_44_2206 ();
 sg13g2_fill_1 FILLER_44_2208 ();
 sg13g2_fill_1 FILLER_44_2218 ();
 sg13g2_fill_2 FILLER_44_2241 ();
 sg13g2_fill_1 FILLER_44_2243 ();
 sg13g2_fill_1 FILLER_44_2276 ();
 sg13g2_fill_1 FILLER_44_2294 ();
 sg13g2_decap_4 FILLER_44_2347 ();
 sg13g2_decap_4 FILLER_44_2359 ();
 sg13g2_fill_1 FILLER_44_2363 ();
 sg13g2_fill_1 FILLER_44_2380 ();
 sg13g2_fill_2 FILLER_44_2386 ();
 sg13g2_fill_1 FILLER_44_2388 ();
 sg13g2_decap_8 FILLER_44_2396 ();
 sg13g2_decap_8 FILLER_44_2403 ();
 sg13g2_decap_8 FILLER_44_2410 ();
 sg13g2_fill_1 FILLER_44_2425 ();
 sg13g2_fill_2 FILLER_44_2456 ();
 sg13g2_decap_8 FILLER_44_2469 ();
 sg13g2_decap_8 FILLER_44_2503 ();
 sg13g2_decap_8 FILLER_44_2510 ();
 sg13g2_fill_2 FILLER_44_2517 ();
 sg13g2_fill_1 FILLER_44_2519 ();
 sg13g2_fill_2 FILLER_44_2524 ();
 sg13g2_fill_2 FILLER_44_2544 ();
 sg13g2_fill_1 FILLER_44_2546 ();
 sg13g2_fill_2 FILLER_44_2563 ();
 sg13g2_fill_2 FILLER_44_2574 ();
 sg13g2_fill_1 FILLER_44_2589 ();
 sg13g2_fill_2 FILLER_44_2607 ();
 sg13g2_decap_8 FILLER_44_2641 ();
 sg13g2_decap_8 FILLER_44_2648 ();
 sg13g2_decap_8 FILLER_44_2655 ();
 sg13g2_decap_4 FILLER_44_2662 ();
 sg13g2_fill_2 FILLER_44_2714 ();
 sg13g2_fill_2 FILLER_44_2788 ();
 sg13g2_decap_4 FILLER_44_2816 ();
 sg13g2_fill_2 FILLER_44_2820 ();
 sg13g2_decap_4 FILLER_44_2831 ();
 sg13g2_decap_4 FILLER_44_2884 ();
 sg13g2_fill_1 FILLER_44_2888 ();
 sg13g2_fill_2 FILLER_44_2916 ();
 sg13g2_fill_1 FILLER_44_2945 ();
 sg13g2_fill_2 FILLER_44_2973 ();
 sg13g2_fill_2 FILLER_44_3002 ();
 sg13g2_fill_2 FILLER_44_3026 ();
 sg13g2_fill_1 FILLER_44_3028 ();
 sg13g2_decap_8 FILLER_44_3033 ();
 sg13g2_decap_4 FILLER_44_3040 ();
 sg13g2_fill_2 FILLER_44_3044 ();
 sg13g2_fill_2 FILLER_44_3059 ();
 sg13g2_fill_1 FILLER_44_3061 ();
 sg13g2_fill_1 FILLER_44_3136 ();
 sg13g2_decap_8 FILLER_44_3155 ();
 sg13g2_decap_8 FILLER_44_3162 ();
 sg13g2_fill_2 FILLER_44_3169 ();
 sg13g2_decap_8 FILLER_44_3193 ();
 sg13g2_decap_4 FILLER_44_3200 ();
 sg13g2_fill_1 FILLER_44_3204 ();
 sg13g2_decap_8 FILLER_44_3232 ();
 sg13g2_decap_4 FILLER_44_3239 ();
 sg13g2_fill_1 FILLER_44_3243 ();
 sg13g2_decap_8 FILLER_44_3248 ();
 sg13g2_decap_8 FILLER_44_3255 ();
 sg13g2_fill_1 FILLER_44_3296 ();
 sg13g2_decap_8 FILLER_44_3315 ();
 sg13g2_fill_2 FILLER_44_3322 ();
 sg13g2_fill_1 FILLER_44_3324 ();
 sg13g2_decap_4 FILLER_44_3333 ();
 sg13g2_fill_2 FILLER_44_3337 ();
 sg13g2_fill_2 FILLER_44_3352 ();
 sg13g2_fill_1 FILLER_44_3354 ();
 sg13g2_decap_4 FILLER_44_3372 ();
 sg13g2_fill_2 FILLER_44_3393 ();
 sg13g2_decap_4 FILLER_44_3410 ();
 sg13g2_fill_2 FILLER_44_3427 ();
 sg13g2_fill_1 FILLER_44_3429 ();
 sg13g2_decap_8 FILLER_44_3457 ();
 sg13g2_decap_8 FILLER_44_3464 ();
 sg13g2_decap_8 FILLER_44_3471 ();
 sg13g2_decap_8 FILLER_44_3478 ();
 sg13g2_decap_8 FILLER_44_3485 ();
 sg13g2_decap_8 FILLER_44_3492 ();
 sg13g2_decap_8 FILLER_44_3499 ();
 sg13g2_decap_8 FILLER_44_3506 ();
 sg13g2_decap_8 FILLER_44_3513 ();
 sg13g2_decap_8 FILLER_44_3520 ();
 sg13g2_decap_8 FILLER_44_3527 ();
 sg13g2_decap_8 FILLER_44_3534 ();
 sg13g2_decap_8 FILLER_44_3541 ();
 sg13g2_decap_8 FILLER_44_3548 ();
 sg13g2_decap_8 FILLER_44_3555 ();
 sg13g2_decap_8 FILLER_44_3562 ();
 sg13g2_decap_8 FILLER_44_3569 ();
 sg13g2_decap_4 FILLER_44_3576 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_112 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_181 ();
 sg13g2_decap_8 FILLER_45_188 ();
 sg13g2_fill_2 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_2 FILLER_45_202 ();
 sg13g2_fill_1 FILLER_45_204 ();
 sg13g2_decap_4 FILLER_45_210 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_230 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_decap_4 FILLER_45_366 ();
 sg13g2_decap_4 FILLER_45_375 ();
 sg13g2_fill_2 FILLER_45_410 ();
 sg13g2_fill_1 FILLER_45_416 ();
 sg13g2_decap_4 FILLER_45_462 ();
 sg13g2_fill_1 FILLER_45_488 ();
 sg13g2_decap_8 FILLER_45_543 ();
 sg13g2_decap_8 FILLER_45_646 ();
 sg13g2_decap_8 FILLER_45_653 ();
 sg13g2_decap_4 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_674 ();
 sg13g2_fill_2 FILLER_45_697 ();
 sg13g2_fill_2 FILLER_45_736 ();
 sg13g2_decap_4 FILLER_45_769 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_864 ();
 sg13g2_fill_1 FILLER_45_871 ();
 sg13g2_fill_2 FILLER_45_881 ();
 sg13g2_fill_1 FILLER_45_883 ();
 sg13g2_fill_2 FILLER_45_924 ();
 sg13g2_fill_1 FILLER_45_926 ();
 sg13g2_fill_2 FILLER_45_968 ();
 sg13g2_fill_1 FILLER_45_970 ();
 sg13g2_fill_2 FILLER_45_999 ();
 sg13g2_fill_1 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1052 ();
 sg13g2_decap_4 FILLER_45_1059 ();
 sg13g2_fill_2 FILLER_45_1063 ();
 sg13g2_fill_2 FILLER_45_1088 ();
 sg13g2_fill_1 FILLER_45_1090 ();
 sg13g2_fill_1 FILLER_45_1146 ();
 sg13g2_fill_2 FILLER_45_1161 ();
 sg13g2_fill_1 FILLER_45_1163 ();
 sg13g2_decap_8 FILLER_45_1200 ();
 sg13g2_fill_2 FILLER_45_1207 ();
 sg13g2_fill_2 FILLER_45_1214 ();
 sg13g2_decap_4 FILLER_45_1234 ();
 sg13g2_fill_1 FILLER_45_1257 ();
 sg13g2_fill_2 FILLER_45_1272 ();
 sg13g2_fill_1 FILLER_45_1274 ();
 sg13g2_decap_4 FILLER_45_1294 ();
 sg13g2_fill_1 FILLER_45_1298 ();
 sg13g2_fill_1 FILLER_45_1331 ();
 sg13g2_fill_2 FILLER_45_1336 ();
 sg13g2_fill_1 FILLER_45_1338 ();
 sg13g2_decap_4 FILLER_45_1371 ();
 sg13g2_fill_2 FILLER_45_1375 ();
 sg13g2_fill_1 FILLER_45_1382 ();
 sg13g2_fill_2 FILLER_45_1442 ();
 sg13g2_fill_1 FILLER_45_1444 ();
 sg13g2_fill_1 FILLER_45_1459 ();
 sg13g2_fill_1 FILLER_45_1487 ();
 sg13g2_fill_1 FILLER_45_1539 ();
 sg13g2_fill_2 FILLER_45_1578 ();
 sg13g2_decap_8 FILLER_45_1608 ();
 sg13g2_decap_8 FILLER_45_1615 ();
 sg13g2_fill_2 FILLER_45_1622 ();
 sg13g2_fill_1 FILLER_45_1624 ();
 sg13g2_decap_4 FILLER_45_1630 ();
 sg13g2_fill_1 FILLER_45_1634 ();
 sg13g2_decap_8 FILLER_45_1639 ();
 sg13g2_fill_1 FILLER_45_1646 ();
 sg13g2_decap_4 FILLER_45_1656 ();
 sg13g2_decap_8 FILLER_45_1673 ();
 sg13g2_decap_4 FILLER_45_1707 ();
 sg13g2_fill_1 FILLER_45_1711 ();
 sg13g2_fill_2 FILLER_45_1739 ();
 sg13g2_fill_2 FILLER_45_1782 ();
 sg13g2_decap_8 FILLER_45_1797 ();
 sg13g2_fill_1 FILLER_45_1804 ();
 sg13g2_decap_8 FILLER_45_1814 ();
 sg13g2_fill_2 FILLER_45_1854 ();
 sg13g2_fill_1 FILLER_45_1878 ();
 sg13g2_fill_2 FILLER_45_1884 ();
 sg13g2_fill_1 FILLER_45_1895 ();
 sg13g2_decap_4 FILLER_45_1910 ();
 sg13g2_fill_2 FILLER_45_1929 ();
 sg13g2_fill_1 FILLER_45_1931 ();
 sg13g2_decap_8 FILLER_45_1941 ();
 sg13g2_decap_8 FILLER_45_1948 ();
 sg13g2_fill_2 FILLER_45_1955 ();
 sg13g2_decap_4 FILLER_45_1961 ();
 sg13g2_fill_1 FILLER_45_1965 ();
 sg13g2_decap_8 FILLER_45_1971 ();
 sg13g2_decap_4 FILLER_45_1982 ();
 sg13g2_fill_1 FILLER_45_1986 ();
 sg13g2_fill_2 FILLER_45_2000 ();
 sg13g2_decap_8 FILLER_45_2010 ();
 sg13g2_fill_2 FILLER_45_2017 ();
 sg13g2_decap_4 FILLER_45_2028 ();
 sg13g2_decap_8 FILLER_45_2037 ();
 sg13g2_fill_1 FILLER_45_2044 ();
 sg13g2_fill_1 FILLER_45_2050 ();
 sg13g2_fill_1 FILLER_45_2061 ();
 sg13g2_fill_2 FILLER_45_2076 ();
 sg13g2_fill_1 FILLER_45_2078 ();
 sg13g2_fill_1 FILLER_45_2133 ();
 sg13g2_fill_1 FILLER_45_2188 ();
 sg13g2_fill_2 FILLER_45_2217 ();
 sg13g2_fill_1 FILLER_45_2259 ();
 sg13g2_decap_8 FILLER_45_2314 ();
 sg13g2_fill_2 FILLER_45_2334 ();
 sg13g2_fill_1 FILLER_45_2336 ();
 sg13g2_decap_8 FILLER_45_2365 ();
 sg13g2_decap_8 FILLER_45_2372 ();
 sg13g2_decap_4 FILLER_45_2379 ();
 sg13g2_fill_1 FILLER_45_2383 ();
 sg13g2_decap_4 FILLER_45_2412 ();
 sg13g2_fill_2 FILLER_45_2422 ();
 sg13g2_decap_8 FILLER_45_2441 ();
 sg13g2_fill_1 FILLER_45_2448 ();
 sg13g2_fill_2 FILLER_45_2454 ();
 sg13g2_fill_1 FILLER_45_2456 ();
 sg13g2_fill_2 FILLER_45_2494 ();
 sg13g2_fill_1 FILLER_45_2496 ();
 sg13g2_decap_4 FILLER_45_2506 ();
 sg13g2_fill_2 FILLER_45_2515 ();
 sg13g2_fill_1 FILLER_45_2557 ();
 sg13g2_decap_4 FILLER_45_2599 ();
 sg13g2_fill_2 FILLER_45_2603 ();
 sg13g2_fill_2 FILLER_45_2679 ();
 sg13g2_decap_4 FILLER_45_2685 ();
 sg13g2_fill_2 FILLER_45_2689 ();
 sg13g2_decap_8 FILLER_45_2731 ();
 sg13g2_fill_2 FILLER_45_2751 ();
 sg13g2_fill_2 FILLER_45_2756 ();
 sg13g2_fill_1 FILLER_45_2758 ();
 sg13g2_decap_4 FILLER_45_2764 ();
 sg13g2_fill_2 FILLER_45_2768 ();
 sg13g2_fill_1 FILLER_45_2802 ();
 sg13g2_fill_2 FILLER_45_2862 ();
 sg13g2_fill_2 FILLER_45_2967 ();
 sg13g2_decap_4 FILLER_45_3002 ();
 sg13g2_fill_1 FILLER_45_3006 ();
 sg13g2_fill_1 FILLER_45_3037 ();
 sg13g2_decap_8 FILLER_45_3048 ();
 sg13g2_decap_8 FILLER_45_3159 ();
 sg13g2_fill_2 FILLER_45_3166 ();
 sg13g2_fill_1 FILLER_45_3168 ();
 sg13g2_fill_2 FILLER_45_3228 ();
 sg13g2_fill_1 FILLER_45_3230 ();
 sg13g2_fill_2 FILLER_45_3241 ();
 sg13g2_decap_4 FILLER_45_3252 ();
 sg13g2_decap_4 FILLER_45_3261 ();
 sg13g2_fill_2 FILLER_45_3265 ();
 sg13g2_decap_8 FILLER_45_3280 ();
 sg13g2_fill_1 FILLER_45_3287 ();
 sg13g2_decap_4 FILLER_45_3293 ();
 sg13g2_fill_2 FILLER_45_3297 ();
 sg13g2_decap_8 FILLER_45_3334 ();
 sg13g2_fill_1 FILLER_45_3341 ();
 sg13g2_decap_8 FILLER_45_3369 ();
 sg13g2_decap_8 FILLER_45_3376 ();
 sg13g2_fill_2 FILLER_45_3394 ();
 sg13g2_fill_1 FILLER_45_3413 ();
 sg13g2_decap_8 FILLER_45_3446 ();
 sg13g2_decap_8 FILLER_45_3453 ();
 sg13g2_decap_8 FILLER_45_3460 ();
 sg13g2_decap_8 FILLER_45_3467 ();
 sg13g2_decap_8 FILLER_45_3474 ();
 sg13g2_decap_8 FILLER_45_3481 ();
 sg13g2_decap_8 FILLER_45_3488 ();
 sg13g2_decap_8 FILLER_45_3495 ();
 sg13g2_decap_8 FILLER_45_3502 ();
 sg13g2_decap_8 FILLER_45_3509 ();
 sg13g2_decap_8 FILLER_45_3516 ();
 sg13g2_decap_8 FILLER_45_3523 ();
 sg13g2_decap_8 FILLER_45_3530 ();
 sg13g2_decap_8 FILLER_45_3537 ();
 sg13g2_decap_8 FILLER_45_3544 ();
 sg13g2_decap_8 FILLER_45_3551 ();
 sg13g2_decap_8 FILLER_45_3558 ();
 sg13g2_decap_8 FILLER_45_3565 ();
 sg13g2_decap_8 FILLER_45_3572 ();
 sg13g2_fill_1 FILLER_45_3579 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_fill_1 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_121 ();
 sg13g2_decap_8 FILLER_46_163 ();
 sg13g2_decap_4 FILLER_46_170 ();
 sg13g2_fill_1 FILLER_46_183 ();
 sg13g2_fill_2 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_195 ();
 sg13g2_fill_2 FILLER_46_209 ();
 sg13g2_fill_1 FILLER_46_211 ();
 sg13g2_fill_1 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_272 ();
 sg13g2_decap_8 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_286 ();
 sg13g2_fill_1 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_fill_2 FILLER_46_360 ();
 sg13g2_fill_2 FILLER_46_425 ();
 sg13g2_decap_8 FILLER_46_467 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_502 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_decap_4 FILLER_46_523 ();
 sg13g2_decap_4 FILLER_46_531 ();
 sg13g2_fill_2 FILLER_46_535 ();
 sg13g2_fill_1 FILLER_46_541 ();
 sg13g2_fill_2 FILLER_46_551 ();
 sg13g2_fill_1 FILLER_46_575 ();
 sg13g2_fill_2 FILLER_46_589 ();
 sg13g2_decap_8 FILLER_46_633 ();
 sg13g2_fill_2 FILLER_46_640 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_fill_2 FILLER_46_735 ();
 sg13g2_fill_1 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_fill_1 FILLER_46_895 ();
 sg13g2_fill_2 FILLER_46_914 ();
 sg13g2_fill_1 FILLER_46_916 ();
 sg13g2_fill_2 FILLER_46_962 ();
 sg13g2_fill_1 FILLER_46_981 ();
 sg13g2_fill_1 FILLER_46_991 ();
 sg13g2_decap_4 FILLER_46_1012 ();
 sg13g2_fill_2 FILLER_46_1048 ();
 sg13g2_fill_1 FILLER_46_1087 ();
 sg13g2_fill_1 FILLER_46_1124 ();
 sg13g2_fill_1 FILLER_46_1139 ();
 sg13g2_fill_1 FILLER_46_1181 ();
 sg13g2_fill_2 FILLER_46_1187 ();
 sg13g2_fill_1 FILLER_46_1189 ();
 sg13g2_decap_4 FILLER_46_1212 ();
 sg13g2_fill_2 FILLER_46_1216 ();
 sg13g2_fill_1 FILLER_46_1264 ();
 sg13g2_decap_4 FILLER_46_1278 ();
 sg13g2_fill_2 FILLER_46_1333 ();
 sg13g2_fill_1 FILLER_46_1335 ();
 sg13g2_decap_4 FILLER_46_1350 ();
 sg13g2_fill_2 FILLER_46_1354 ();
 sg13g2_fill_2 FILLER_46_1388 ();
 sg13g2_fill_1 FILLER_46_1390 ();
 sg13g2_fill_1 FILLER_46_1432 ();
 sg13g2_fill_2 FILLER_46_1447 ();
 sg13g2_decap_8 FILLER_46_1481 ();
 sg13g2_fill_2 FILLER_46_1524 ();
 sg13g2_fill_2 FILLER_46_1535 ();
 sg13g2_fill_1 FILLER_46_1537 ();
 sg13g2_fill_2 FILLER_46_1547 ();
 sg13g2_decap_4 FILLER_46_1640 ();
 sg13g2_fill_1 FILLER_46_1644 ();
 sg13g2_fill_2 FILLER_46_1682 ();
 sg13g2_decap_8 FILLER_46_1688 ();
 sg13g2_fill_2 FILLER_46_1695 ();
 sg13g2_fill_1 FILLER_46_1697 ();
 sg13g2_fill_2 FILLER_46_1734 ();
 sg13g2_fill_1 FILLER_46_1736 ();
 sg13g2_fill_1 FILLER_46_1756 ();
 sg13g2_fill_1 FILLER_46_1770 ();
 sg13g2_decap_4 FILLER_46_1776 ();
 sg13g2_fill_2 FILLER_46_1780 ();
 sg13g2_fill_2 FILLER_46_1787 ();
 sg13g2_fill_2 FILLER_46_1802 ();
 sg13g2_fill_1 FILLER_46_1804 ();
 sg13g2_decap_8 FILLER_46_1833 ();
 sg13g2_fill_2 FILLER_46_1840 ();
 sg13g2_fill_1 FILLER_46_1869 ();
 sg13g2_fill_2 FILLER_46_1902 ();
 sg13g2_fill_1 FILLER_46_1904 ();
 sg13g2_fill_2 FILLER_46_1933 ();
 sg13g2_decap_8 FILLER_46_1981 ();
 sg13g2_fill_1 FILLER_46_1988 ();
 sg13g2_fill_1 FILLER_46_2003 ();
 sg13g2_fill_1 FILLER_46_2031 ();
 sg13g2_fill_2 FILLER_46_2058 ();
 sg13g2_fill_1 FILLER_46_2060 ();
 sg13g2_decap_4 FILLER_46_2089 ();
 sg13g2_fill_2 FILLER_46_2102 ();
 sg13g2_fill_1 FILLER_46_2113 ();
 sg13g2_fill_2 FILLER_46_2146 ();
 sg13g2_fill_1 FILLER_46_2148 ();
 sg13g2_fill_2 FILLER_46_2200 ();
 sg13g2_fill_1 FILLER_46_2202 ();
 sg13g2_decap_8 FILLER_46_2212 ();
 sg13g2_decap_4 FILLER_46_2219 ();
 sg13g2_fill_2 FILLER_46_2241 ();
 sg13g2_fill_2 FILLER_46_2271 ();
 sg13g2_fill_1 FILLER_46_2352 ();
 sg13g2_fill_2 FILLER_46_2413 ();
 sg13g2_fill_2 FILLER_46_2446 ();
 sg13g2_fill_1 FILLER_46_2448 ();
 sg13g2_fill_1 FILLER_46_2458 ();
 sg13g2_decap_8 FILLER_46_2472 ();
 sg13g2_decap_4 FILLER_46_2479 ();
 sg13g2_fill_2 FILLER_46_2483 ();
 sg13g2_fill_2 FILLER_46_2504 ();
 sg13g2_fill_1 FILLER_46_2506 ();
 sg13g2_fill_2 FILLER_46_2621 ();
 sg13g2_fill_1 FILLER_46_2623 ();
 sg13g2_decap_8 FILLER_46_2641 ();
 sg13g2_decap_8 FILLER_46_2665 ();
 sg13g2_fill_1 FILLER_46_2708 ();
 sg13g2_fill_1 FILLER_46_2791 ();
 sg13g2_decap_4 FILLER_46_2801 ();
 sg13g2_fill_1 FILLER_46_2805 ();
 sg13g2_fill_2 FILLER_46_2846 ();
 sg13g2_fill_1 FILLER_46_2897 ();
 sg13g2_fill_1 FILLER_46_2921 ();
 sg13g2_fill_2 FILLER_46_2932 ();
 sg13g2_fill_1 FILLER_46_2934 ();
 sg13g2_fill_2 FILLER_46_2945 ();
 sg13g2_fill_2 FILLER_46_3001 ();
 sg13g2_fill_1 FILLER_46_3003 ();
 sg13g2_fill_1 FILLER_46_3027 ();
 sg13g2_fill_1 FILLER_46_3073 ();
 sg13g2_fill_2 FILLER_46_3106 ();
 sg13g2_fill_1 FILLER_46_3108 ();
 sg13g2_fill_1 FILLER_46_3151 ();
 sg13g2_fill_2 FILLER_46_3202 ();
 sg13g2_fill_1 FILLER_46_3204 ();
 sg13g2_fill_1 FILLER_46_3215 ();
 sg13g2_fill_1 FILLER_46_3243 ();
 sg13g2_fill_2 FILLER_46_3285 ();
 sg13g2_fill_2 FILLER_46_3309 ();
 sg13g2_fill_2 FILLER_46_3315 ();
 sg13g2_decap_8 FILLER_46_3326 ();
 sg13g2_fill_2 FILLER_46_3333 ();
 sg13g2_decap_8 FILLER_46_3363 ();
 sg13g2_decap_4 FILLER_46_3375 ();
 sg13g2_fill_2 FILLER_46_3383 ();
 sg13g2_fill_1 FILLER_46_3385 ();
 sg13g2_fill_2 FILLER_46_3399 ();
 sg13g2_fill_2 FILLER_46_3413 ();
 sg13g2_fill_1 FILLER_46_3415 ();
 sg13g2_decap_8 FILLER_46_3429 ();
 sg13g2_decap_8 FILLER_46_3436 ();
 sg13g2_decap_8 FILLER_46_3443 ();
 sg13g2_decap_8 FILLER_46_3450 ();
 sg13g2_decap_8 FILLER_46_3457 ();
 sg13g2_decap_8 FILLER_46_3464 ();
 sg13g2_decap_8 FILLER_46_3471 ();
 sg13g2_decap_8 FILLER_46_3478 ();
 sg13g2_decap_8 FILLER_46_3485 ();
 sg13g2_decap_8 FILLER_46_3492 ();
 sg13g2_decap_8 FILLER_46_3499 ();
 sg13g2_decap_8 FILLER_46_3506 ();
 sg13g2_decap_8 FILLER_46_3513 ();
 sg13g2_decap_8 FILLER_46_3520 ();
 sg13g2_decap_8 FILLER_46_3527 ();
 sg13g2_decap_8 FILLER_46_3534 ();
 sg13g2_decap_8 FILLER_46_3541 ();
 sg13g2_decap_8 FILLER_46_3548 ();
 sg13g2_decap_8 FILLER_46_3555 ();
 sg13g2_decap_8 FILLER_46_3562 ();
 sg13g2_decap_8 FILLER_46_3569 ();
 sg13g2_decap_4 FILLER_46_3576 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_decap_8 FILLER_47_94 ();
 sg13g2_decap_8 FILLER_47_101 ();
 sg13g2_decap_4 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_144 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_decap_8 FILLER_47_171 ();
 sg13g2_decap_8 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_210 ();
 sg13g2_fill_2 FILLER_47_216 ();
 sg13g2_fill_1 FILLER_47_218 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_fill_1 FILLER_47_267 ();
 sg13g2_decap_4 FILLER_47_295 ();
 sg13g2_fill_1 FILLER_47_299 ();
 sg13g2_fill_2 FILLER_47_320 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_fill_1 FILLER_47_433 ();
 sg13g2_fill_2 FILLER_47_496 ();
 sg13g2_fill_1 FILLER_47_498 ();
 sg13g2_decap_8 FILLER_47_562 ();
 sg13g2_decap_8 FILLER_47_569 ();
 sg13g2_decap_8 FILLER_47_576 ();
 sg13g2_decap_8 FILLER_47_583 ();
 sg13g2_decap_4 FILLER_47_622 ();
 sg13g2_fill_1 FILLER_47_626 ();
 sg13g2_decap_4 FILLER_47_666 ();
 sg13g2_decap_4 FILLER_47_711 ();
 sg13g2_fill_1 FILLER_47_715 ();
 sg13g2_fill_1 FILLER_47_726 ();
 sg13g2_decap_4 FILLER_47_759 ();
 sg13g2_fill_2 FILLER_47_763 ();
 sg13g2_fill_1 FILLER_47_801 ();
 sg13g2_fill_2 FILLER_47_835 ();
 sg13g2_fill_1 FILLER_47_837 ();
 sg13g2_fill_2 FILLER_47_865 ();
 sg13g2_fill_2 FILLER_47_886 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_fill_2 FILLER_47_927 ();
 sg13g2_fill_1 FILLER_47_951 ();
 sg13g2_fill_2 FILLER_47_976 ();
 sg13g2_fill_1 FILLER_47_978 ();
 sg13g2_fill_1 FILLER_47_988 ();
 sg13g2_fill_1 FILLER_47_1007 ();
 sg13g2_decap_4 FILLER_47_1034 ();
 sg13g2_fill_2 FILLER_47_1038 ();
 sg13g2_fill_2 FILLER_47_1077 ();
 sg13g2_decap_8 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1096 ();
 sg13g2_fill_1 FILLER_47_1140 ();
 sg13g2_fill_2 FILLER_47_1155 ();
 sg13g2_fill_2 FILLER_47_1174 ();
 sg13g2_fill_1 FILLER_47_1239 ();
 sg13g2_decap_4 FILLER_47_1244 ();
 sg13g2_fill_1 FILLER_47_1248 ();
 sg13g2_decap_8 FILLER_47_1289 ();
 sg13g2_fill_2 FILLER_47_1296 ();
 sg13g2_fill_2 FILLER_47_1351 ();
 sg13g2_fill_1 FILLER_47_1367 ();
 sg13g2_fill_2 FILLER_47_1387 ();
 sg13g2_fill_1 FILLER_47_1389 ();
 sg13g2_fill_1 FILLER_47_1417 ();
 sg13g2_fill_1 FILLER_47_1447 ();
 sg13g2_fill_2 FILLER_47_1461 ();
 sg13g2_decap_8 FILLER_47_1489 ();
 sg13g2_decap_4 FILLER_47_1501 ();
 sg13g2_fill_1 FILLER_47_1515 ();
 sg13g2_fill_2 FILLER_47_1548 ();
 sg13g2_fill_1 FILLER_47_1550 ();
 sg13g2_fill_1 FILLER_47_1561 ();
 sg13g2_fill_2 FILLER_47_1576 ();
 sg13g2_fill_1 FILLER_47_1578 ();
 sg13g2_fill_1 FILLER_47_1608 ();
 sg13g2_fill_2 FILLER_47_1618 ();
 sg13g2_fill_2 FILLER_47_1662 ();
 sg13g2_fill_1 FILLER_47_1664 ();
 sg13g2_fill_1 FILLER_47_1674 ();
 sg13g2_fill_1 FILLER_47_1707 ();
 sg13g2_fill_2 FILLER_47_1771 ();
 sg13g2_fill_1 FILLER_47_1773 ();
 sg13g2_fill_1 FILLER_47_1807 ();
 sg13g2_decap_8 FILLER_47_1817 ();
 sg13g2_decap_4 FILLER_47_1829 ();
 sg13g2_fill_2 FILLER_47_1856 ();
 sg13g2_fill_2 FILLER_47_1885 ();
 sg13g2_fill_2 FILLER_47_1901 ();
 sg13g2_fill_1 FILLER_47_1903 ();
 sg13g2_fill_1 FILLER_47_1917 ();
 sg13g2_fill_2 FILLER_47_1973 ();
 sg13g2_fill_1 FILLER_47_1975 ();
 sg13g2_fill_1 FILLER_47_2008 ();
 sg13g2_decap_4 FILLER_47_2013 ();
 sg13g2_fill_1 FILLER_47_2017 ();
 sg13g2_fill_1 FILLER_47_2027 ();
 sg13g2_fill_2 FILLER_47_2032 ();
 sg13g2_decap_8 FILLER_47_2039 ();
 sg13g2_decap_4 FILLER_47_2046 ();
 sg13g2_fill_1 FILLER_47_2050 ();
 sg13g2_fill_1 FILLER_47_2068 ();
 sg13g2_fill_2 FILLER_47_2096 ();
 sg13g2_fill_1 FILLER_47_2098 ();
 sg13g2_decap_4 FILLER_47_2123 ();
 sg13g2_fill_2 FILLER_47_2132 ();
 sg13g2_fill_2 FILLER_47_2144 ();
 sg13g2_fill_2 FILLER_47_2168 ();
 sg13g2_fill_2 FILLER_47_2188 ();
 sg13g2_fill_1 FILLER_47_2199 ();
 sg13g2_fill_1 FILLER_47_2246 ();
 sg13g2_fill_2 FILLER_47_2256 ();
 sg13g2_fill_1 FILLER_47_2258 ();
 sg13g2_decap_4 FILLER_47_2268 ();
 sg13g2_decap_8 FILLER_47_2317 ();
 sg13g2_decap_8 FILLER_47_2324 ();
 sg13g2_fill_1 FILLER_47_2353 ();
 sg13g2_fill_1 FILLER_47_2382 ();
 sg13g2_fill_2 FILLER_47_2388 ();
 sg13g2_decap_4 FILLER_47_2418 ();
 sg13g2_fill_1 FILLER_47_2422 ();
 sg13g2_decap_8 FILLER_47_2427 ();
 sg13g2_fill_1 FILLER_47_2587 ();
 sg13g2_decap_4 FILLER_47_2593 ();
 sg13g2_fill_1 FILLER_47_2597 ();
 sg13g2_decap_8 FILLER_47_2605 ();
 sg13g2_decap_4 FILLER_47_2612 ();
 sg13g2_fill_1 FILLER_47_2616 ();
 sg13g2_fill_2 FILLER_47_2630 ();
 sg13g2_fill_1 FILLER_47_2637 ();
 sg13g2_decap_8 FILLER_47_2680 ();
 sg13g2_decap_4 FILLER_47_2687 ();
 sg13g2_fill_2 FILLER_47_2700 ();
 sg13g2_fill_1 FILLER_47_2702 ();
 sg13g2_fill_1 FILLER_47_2716 ();
 sg13g2_decap_4 FILLER_47_2735 ();
 sg13g2_fill_2 FILLER_47_2739 ();
 sg13g2_fill_2 FILLER_47_2750 ();
 sg13g2_fill_1 FILLER_47_2752 ();
 sg13g2_fill_2 FILLER_47_2766 ();
 sg13g2_fill_1 FILLER_47_2768 ();
 sg13g2_fill_2 FILLER_47_2796 ();
 sg13g2_fill_1 FILLER_47_2798 ();
 sg13g2_fill_2 FILLER_47_2880 ();
 sg13g2_fill_1 FILLER_47_2882 ();
 sg13g2_fill_2 FILLER_47_2934 ();
 sg13g2_fill_1 FILLER_47_2936 ();
 sg13g2_decap_8 FILLER_47_2942 ();
 sg13g2_fill_2 FILLER_47_2962 ();
 sg13g2_fill_1 FILLER_47_2964 ();
 sg13g2_decap_8 FILLER_47_2992 ();
 sg13g2_fill_2 FILLER_47_3004 ();
 sg13g2_fill_1 FILLER_47_3006 ();
 sg13g2_fill_2 FILLER_47_3094 ();
 sg13g2_fill_2 FILLER_47_3113 ();
 sg13g2_fill_2 FILLER_47_3127 ();
 sg13g2_fill_1 FILLER_47_3129 ();
 sg13g2_fill_2 FILLER_47_3165 ();
 sg13g2_fill_2 FILLER_47_3180 ();
 sg13g2_decap_8 FILLER_47_3273 ();
 sg13g2_fill_2 FILLER_47_3280 ();
 sg13g2_fill_1 FILLER_47_3323 ();
 sg13g2_fill_2 FILLER_47_3330 ();
 sg13g2_fill_1 FILLER_47_3332 ();
 sg13g2_fill_1 FILLER_47_3351 ();
 sg13g2_fill_1 FILLER_47_3361 ();
 sg13g2_decap_8 FILLER_47_3456 ();
 sg13g2_decap_8 FILLER_47_3463 ();
 sg13g2_decap_8 FILLER_47_3470 ();
 sg13g2_decap_8 FILLER_47_3477 ();
 sg13g2_decap_8 FILLER_47_3484 ();
 sg13g2_decap_8 FILLER_47_3491 ();
 sg13g2_decap_8 FILLER_47_3498 ();
 sg13g2_decap_8 FILLER_47_3505 ();
 sg13g2_decap_8 FILLER_47_3512 ();
 sg13g2_decap_8 FILLER_47_3519 ();
 sg13g2_decap_8 FILLER_47_3526 ();
 sg13g2_decap_8 FILLER_47_3533 ();
 sg13g2_decap_8 FILLER_47_3540 ();
 sg13g2_decap_8 FILLER_47_3547 ();
 sg13g2_decap_8 FILLER_47_3554 ();
 sg13g2_decap_8 FILLER_47_3561 ();
 sg13g2_decap_8 FILLER_47_3568 ();
 sg13g2_decap_4 FILLER_47_3575 ();
 sg13g2_fill_1 FILLER_47_3579 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_77 ();
 sg13g2_fill_1 FILLER_48_79 ();
 sg13g2_decap_4 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_121 ();
 sg13g2_fill_2 FILLER_48_165 ();
 sg13g2_decap_4 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_175 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_1 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_decap_8 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_241 ();
 sg13g2_fill_2 FILLER_48_259 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_decap_4 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_301 ();
 sg13g2_decap_4 FILLER_48_330 ();
 sg13g2_fill_2 FILLER_48_334 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_4 FILLER_48_397 ();
 sg13g2_fill_2 FILLER_48_401 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_2 FILLER_48_464 ();
 sg13g2_decap_8 FILLER_48_512 ();
 sg13g2_fill_2 FILLER_48_528 ();
 sg13g2_fill_2 FILLER_48_544 ();
 sg13g2_fill_1 FILLER_48_546 ();
 sg13g2_fill_2 FILLER_48_605 ();
 sg13g2_decap_8 FILLER_48_674 ();
 sg13g2_decap_4 FILLER_48_721 ();
 sg13g2_fill_2 FILLER_48_776 ();
 sg13g2_fill_1 FILLER_48_791 ();
 sg13g2_fill_2 FILLER_48_809 ();
 sg13g2_fill_1 FILLER_48_852 ();
 sg13g2_decap_8 FILLER_48_880 ();
 sg13g2_decap_8 FILLER_48_887 ();
 sg13g2_fill_2 FILLER_48_934 ();
 sg13g2_fill_1 FILLER_48_936 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_fill_1 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_48_1069 ();
 sg13g2_decap_4 FILLER_48_1076 ();
 sg13g2_decap_8 FILLER_48_1107 ();
 sg13g2_fill_2 FILLER_48_1114 ();
 sg13g2_fill_2 FILLER_48_1142 ();
 sg13g2_decap_4 FILLER_48_1193 ();
 sg13g2_fill_2 FILLER_48_1197 ();
 sg13g2_decap_8 FILLER_48_1212 ();
 sg13g2_fill_1 FILLER_48_1229 ();
 sg13g2_fill_1 FILLER_48_1285 ();
 sg13g2_decap_8 FILLER_48_1296 ();
 sg13g2_decap_8 FILLER_48_1303 ();
 sg13g2_decap_8 FILLER_48_1310 ();
 sg13g2_decap_4 FILLER_48_1317 ();
 sg13g2_fill_2 FILLER_48_1376 ();
 sg13g2_fill_1 FILLER_48_1378 ();
 sg13g2_fill_1 FILLER_48_1388 ();
 sg13g2_fill_2 FILLER_48_1416 ();
 sg13g2_fill_1 FILLER_48_1418 ();
 sg13g2_fill_2 FILLER_48_1432 ();
 sg13g2_decap_4 FILLER_48_1470 ();
 sg13g2_fill_2 FILLER_48_1474 ();
 sg13g2_decap_8 FILLER_48_1503 ();
 sg13g2_fill_1 FILLER_48_1510 ();
 sg13g2_decap_4 FILLER_48_1538 ();
 sg13g2_decap_4 FILLER_48_1596 ();
 sg13g2_fill_2 FILLER_48_1600 ();
 sg13g2_fill_1 FILLER_48_1629 ();
 sg13g2_decap_8 FILLER_48_1671 ();
 sg13g2_fill_2 FILLER_48_1678 ();
 sg13g2_fill_2 FILLER_48_1690 ();
 sg13g2_fill_1 FILLER_48_1719 ();
 sg13g2_fill_2 FILLER_48_1725 ();
 sg13g2_fill_1 FILLER_48_1727 ();
 sg13g2_fill_2 FILLER_48_1737 ();
 sg13g2_fill_1 FILLER_48_1739 ();
 sg13g2_fill_1 FILLER_48_1753 ();
 sg13g2_decap_8 FILLER_48_1763 ();
 sg13g2_decap_4 FILLER_48_1770 ();
 sg13g2_fill_1 FILLER_48_1774 ();
 sg13g2_fill_2 FILLER_48_1788 ();
 sg13g2_fill_2 FILLER_48_1875 ();
 sg13g2_fill_2 FILLER_48_1882 ();
 sg13g2_fill_1 FILLER_48_1884 ();
 sg13g2_fill_1 FILLER_48_1895 ();
 sg13g2_fill_1 FILLER_48_1914 ();
 sg13g2_fill_1 FILLER_48_1924 ();
 sg13g2_fill_2 FILLER_48_1930 ();
 sg13g2_fill_1 FILLER_48_1932 ();
 sg13g2_decap_4 FILLER_48_1946 ();
 sg13g2_fill_2 FILLER_48_1950 ();
 sg13g2_fill_2 FILLER_48_1972 ();
 sg13g2_fill_1 FILLER_48_2001 ();
 sg13g2_fill_2 FILLER_48_2029 ();
 sg13g2_fill_2 FILLER_48_2036 ();
 sg13g2_fill_1 FILLER_48_2038 ();
 sg13g2_decap_8 FILLER_48_2043 ();
 sg13g2_fill_1 FILLER_48_2050 ();
 sg13g2_fill_2 FILLER_48_2060 ();
 sg13g2_fill_2 FILLER_48_2099 ();
 sg13g2_decap_4 FILLER_48_2118 ();
 sg13g2_fill_2 FILLER_48_2131 ();
 sg13g2_fill_2 FILLER_48_2137 ();
 sg13g2_decap_8 FILLER_48_2171 ();
 sg13g2_fill_1 FILLER_48_2178 ();
 sg13g2_fill_1 FILLER_48_2215 ();
 sg13g2_fill_2 FILLER_48_2261 ();
 sg13g2_fill_1 FILLER_48_2263 ();
 sg13g2_decap_4 FILLER_48_2297 ();
 sg13g2_fill_2 FILLER_48_2301 ();
 sg13g2_fill_1 FILLER_48_2312 ();
 sg13g2_fill_2 FILLER_48_2331 ();
 sg13g2_fill_1 FILLER_48_2333 ();
 sg13g2_fill_1 FILLER_48_2352 ();
 sg13g2_fill_2 FILLER_48_2380 ();
 sg13g2_fill_1 FILLER_48_2382 ();
 sg13g2_fill_1 FILLER_48_2388 ();
 sg13g2_fill_1 FILLER_48_2407 ();
 sg13g2_decap_4 FILLER_48_2458 ();
 sg13g2_fill_1 FILLER_48_2462 ();
 sg13g2_fill_2 FILLER_48_2472 ();
 sg13g2_decap_8 FILLER_48_2478 ();
 sg13g2_decap_8 FILLER_48_2485 ();
 sg13g2_fill_2 FILLER_48_2496 ();
 sg13g2_decap_4 FILLER_48_2511 ();
 sg13g2_decap_4 FILLER_48_2524 ();
 sg13g2_fill_1 FILLER_48_2528 ();
 sg13g2_decap_4 FILLER_48_2540 ();
 sg13g2_fill_2 FILLER_48_2544 ();
 sg13g2_fill_1 FILLER_48_2558 ();
 sg13g2_decap_8 FILLER_48_2590 ();
 sg13g2_fill_2 FILLER_48_2597 ();
 sg13g2_fill_1 FILLER_48_2599 ();
 sg13g2_fill_2 FILLER_48_2628 ();
 sg13g2_fill_2 FILLER_48_2652 ();
 sg13g2_fill_1 FILLER_48_2687 ();
 sg13g2_fill_1 FILLER_48_2710 ();
 sg13g2_fill_1 FILLER_48_2719 ();
 sg13g2_fill_2 FILLER_48_2738 ();
 sg13g2_fill_1 FILLER_48_2740 ();
 sg13g2_decap_8 FILLER_48_2763 ();
 sg13g2_decap_4 FILLER_48_2775 ();
 sg13g2_decap_8 FILLER_48_2803 ();
 sg13g2_fill_1 FILLER_48_2819 ();
 sg13g2_decap_8 FILLER_48_2829 ();
 sg13g2_decap_8 FILLER_48_2836 ();
 sg13g2_fill_2 FILLER_48_2843 ();
 sg13g2_fill_1 FILLER_48_2845 ();
 sg13g2_fill_2 FILLER_48_2901 ();
 sg13g2_fill_1 FILLER_48_2917 ();
 sg13g2_decap_4 FILLER_48_2935 ();
 sg13g2_fill_2 FILLER_48_2939 ();
 sg13g2_fill_1 FILLER_48_2959 ();
 sg13g2_fill_1 FILLER_48_2983 ();
 sg13g2_decap_8 FILLER_48_2988 ();
 sg13g2_fill_2 FILLER_48_3000 ();
 sg13g2_decap_4 FILLER_48_3067 ();
 sg13g2_fill_2 FILLER_48_3071 ();
 sg13g2_fill_2 FILLER_48_3082 ();
 sg13g2_fill_2 FILLER_48_3097 ();
 sg13g2_fill_1 FILLER_48_3099 ();
 sg13g2_fill_1 FILLER_48_3104 ();
 sg13g2_fill_1 FILLER_48_3152 ();
 sg13g2_decap_8 FILLER_48_3181 ();
 sg13g2_decap_4 FILLER_48_3188 ();
 sg13g2_fill_1 FILLER_48_3192 ();
 sg13g2_decap_8 FILLER_48_3248 ();
 sg13g2_fill_2 FILLER_48_3255 ();
 sg13g2_fill_1 FILLER_48_3298 ();
 sg13g2_fill_2 FILLER_48_3307 ();
 sg13g2_fill_1 FILLER_48_3309 ();
 sg13g2_fill_2 FILLER_48_3327 ();
 sg13g2_fill_1 FILLER_48_3329 ();
 sg13g2_fill_1 FILLER_48_3343 ();
 sg13g2_fill_1 FILLER_48_3348 ();
 sg13g2_decap_4 FILLER_48_3357 ();
 sg13g2_fill_2 FILLER_48_3378 ();
 sg13g2_decap_8 FILLER_48_3415 ();
 sg13g2_decap_4 FILLER_48_3422 ();
 sg13g2_decap_8 FILLER_48_3439 ();
 sg13g2_decap_8 FILLER_48_3446 ();
 sg13g2_decap_8 FILLER_48_3453 ();
 sg13g2_decap_8 FILLER_48_3460 ();
 sg13g2_decap_8 FILLER_48_3467 ();
 sg13g2_decap_8 FILLER_48_3474 ();
 sg13g2_decap_8 FILLER_48_3481 ();
 sg13g2_decap_8 FILLER_48_3488 ();
 sg13g2_decap_8 FILLER_48_3495 ();
 sg13g2_decap_8 FILLER_48_3502 ();
 sg13g2_decap_8 FILLER_48_3509 ();
 sg13g2_decap_8 FILLER_48_3516 ();
 sg13g2_decap_8 FILLER_48_3523 ();
 sg13g2_decap_8 FILLER_48_3530 ();
 sg13g2_decap_8 FILLER_48_3537 ();
 sg13g2_decap_8 FILLER_48_3544 ();
 sg13g2_decap_8 FILLER_48_3551 ();
 sg13g2_decap_8 FILLER_48_3558 ();
 sg13g2_decap_8 FILLER_48_3565 ();
 sg13g2_decap_8 FILLER_48_3572 ();
 sg13g2_fill_1 FILLER_48_3579 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_90 ();
 sg13g2_decap_8 FILLER_49_97 ();
 sg13g2_decap_8 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_153 ();
 sg13g2_fill_2 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_decap_8 FILLER_49_243 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_4 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_fill_2 FILLER_49_291 ();
 sg13g2_decap_4 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_333 ();
 sg13g2_fill_2 FILLER_49_405 ();
 sg13g2_fill_2 FILLER_49_456 ();
 sg13g2_fill_2 FILLER_49_463 ();
 sg13g2_fill_1 FILLER_49_465 ();
 sg13g2_fill_2 FILLER_49_497 ();
 sg13g2_fill_1 FILLER_49_499 ();
 sg13g2_decap_8 FILLER_49_509 ();
 sg13g2_decap_8 FILLER_49_516 ();
 sg13g2_decap_4 FILLER_49_523 ();
 sg13g2_fill_2 FILLER_49_527 ();
 sg13g2_decap_4 FILLER_49_560 ();
 sg13g2_fill_2 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_575 ();
 sg13g2_fill_2 FILLER_49_580 ();
 sg13g2_fill_2 FILLER_49_594 ();
 sg13g2_decap_8 FILLER_49_617 ();
 sg13g2_decap_8 FILLER_49_624 ();
 sg13g2_decap_4 FILLER_49_668 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_730 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_4 FILLER_49_753 ();
 sg13g2_fill_1 FILLER_49_757 ();
 sg13g2_fill_2 FILLER_49_858 ();
 sg13g2_fill_2 FILLER_49_870 ();
 sg13g2_fill_1 FILLER_49_951 ();
 sg13g2_fill_2 FILLER_49_996 ();
 sg13g2_decap_8 FILLER_49_1002 ();
 sg13g2_decap_8 FILLER_49_1009 ();
 sg13g2_decap_8 FILLER_49_1016 ();
 sg13g2_fill_2 FILLER_49_1023 ();
 sg13g2_decap_8 FILLER_49_1038 ();
 sg13g2_fill_2 FILLER_49_1045 ();
 sg13g2_fill_1 FILLER_49_1061 ();
 sg13g2_decap_4 FILLER_49_1075 ();
 sg13g2_fill_1 FILLER_49_1079 ();
 sg13g2_fill_1 FILLER_49_1089 ();
 sg13g2_decap_8 FILLER_49_1109 ();
 sg13g2_decap_4 FILLER_49_1116 ();
 sg13g2_fill_1 FILLER_49_1157 ();
 sg13g2_decap_4 FILLER_49_1208 ();
 sg13g2_fill_2 FILLER_49_1212 ();
 sg13g2_decap_8 FILLER_49_1244 ();
 sg13g2_fill_1 FILLER_49_1251 ();
 sg13g2_decap_8 FILLER_49_1346 ();
 sg13g2_fill_2 FILLER_49_1353 ();
 sg13g2_fill_2 FILLER_49_1369 ();
 sg13g2_decap_8 FILLER_49_1398 ();
 sg13g2_fill_2 FILLER_49_1418 ();
 sg13g2_fill_2 FILLER_49_1447 ();
 sg13g2_decap_8 FILLER_49_1459 ();
 sg13g2_decap_4 FILLER_49_1466 ();
 sg13g2_fill_1 FILLER_49_1470 ();
 sg13g2_fill_2 FILLER_49_1494 ();
 sg13g2_decap_4 FILLER_49_1522 ();
 sg13g2_fill_2 FILLER_49_1526 ();
 sg13g2_decap_4 FILLER_49_1541 ();
 sg13g2_fill_2 FILLER_49_1545 ();
 sg13g2_fill_1 FILLER_49_1556 ();
 sg13g2_fill_2 FILLER_49_1575 ();
 sg13g2_fill_1 FILLER_49_1586 ();
 sg13g2_decap_8 FILLER_49_1601 ();
 sg13g2_decap_8 FILLER_49_1608 ();
 sg13g2_fill_1 FILLER_49_1615 ();
 sg13g2_fill_1 FILLER_49_1625 ();
 sg13g2_fill_1 FILLER_49_1639 ();
 sg13g2_decap_4 FILLER_49_1681 ();
 sg13g2_fill_2 FILLER_49_1690 ();
 sg13g2_fill_1 FILLER_49_1692 ();
 sg13g2_fill_2 FILLER_49_1741 ();
 sg13g2_fill_1 FILLER_49_1743 ();
 sg13g2_decap_8 FILLER_49_1772 ();
 sg13g2_fill_1 FILLER_49_1779 ();
 sg13g2_fill_2 FILLER_49_1824 ();
 sg13g2_fill_2 FILLER_49_1831 ();
 sg13g2_fill_1 FILLER_49_1833 ();
 sg13g2_fill_2 FILLER_49_1848 ();
 sg13g2_fill_2 FILLER_49_1859 ();
 sg13g2_fill_1 FILLER_49_1861 ();
 sg13g2_fill_2 FILLER_49_1867 ();
 sg13g2_fill_1 FILLER_49_1869 ();
 sg13g2_fill_2 FILLER_49_1883 ();
 sg13g2_fill_1 FILLER_49_1913 ();
 sg13g2_fill_2 FILLER_49_1960 ();
 sg13g2_fill_1 FILLER_49_1962 ();
 sg13g2_fill_2 FILLER_49_2064 ();
 sg13g2_fill_1 FILLER_49_2066 ();
 sg13g2_fill_1 FILLER_49_2081 ();
 sg13g2_decap_8 FILLER_49_2138 ();
 sg13g2_fill_1 FILLER_49_2145 ();
 sg13g2_fill_2 FILLER_49_2206 ();
 sg13g2_fill_1 FILLER_49_2208 ();
 sg13g2_fill_2 FILLER_49_2228 ();
 sg13g2_fill_1 FILLER_49_2230 ();
 sg13g2_decap_4 FILLER_49_2248 ();
 sg13g2_decap_8 FILLER_49_2269 ();
 sg13g2_decap_4 FILLER_49_2276 ();
 sg13g2_fill_2 FILLER_49_2280 ();
 sg13g2_fill_1 FILLER_49_2287 ();
 sg13g2_decap_4 FILLER_49_2292 ();
 sg13g2_decap_4 FILLER_49_2301 ();
 sg13g2_fill_1 FILLER_49_2305 ();
 sg13g2_fill_1 FILLER_49_2366 ();
 sg13g2_fill_1 FILLER_49_2381 ();
 sg13g2_fill_2 FILLER_49_2404 ();
 sg13g2_fill_1 FILLER_49_2406 ();
 sg13g2_fill_2 FILLER_49_2435 ();
 sg13g2_fill_1 FILLER_49_2437 ();
 sg13g2_fill_2 FILLER_49_2508 ();
 sg13g2_fill_1 FILLER_49_2510 ();
 sg13g2_decap_8 FILLER_49_2524 ();
 sg13g2_fill_2 FILLER_49_2531 ();
 sg13g2_fill_1 FILLER_49_2533 ();
 sg13g2_fill_2 FILLER_49_2554 ();
 sg13g2_fill_2 FILLER_49_2573 ();
 sg13g2_fill_1 FILLER_49_2575 ();
 sg13g2_fill_1 FILLER_49_2581 ();
 sg13g2_fill_1 FILLER_49_2633 ();
 sg13g2_fill_2 FILLER_49_2693 ();
 sg13g2_decap_4 FILLER_49_2737 ();
 sg13g2_fill_1 FILLER_49_2741 ();
 sg13g2_fill_1 FILLER_49_2778 ();
 sg13g2_decap_4 FILLER_49_2793 ();
 sg13g2_fill_2 FILLER_49_2797 ();
 sg13g2_fill_2 FILLER_49_2808 ();
 sg13g2_fill_2 FILLER_49_2847 ();
 sg13g2_fill_2 FILLER_49_2854 ();
 sg13g2_fill_1 FILLER_49_2856 ();
 sg13g2_fill_1 FILLER_49_2862 ();
 sg13g2_fill_2 FILLER_49_2867 ();
 sg13g2_fill_2 FILLER_49_2941 ();
 sg13g2_fill_1 FILLER_49_2943 ();
 sg13g2_fill_2 FILLER_49_2954 ();
 sg13g2_fill_1 FILLER_49_2965 ();
 sg13g2_fill_2 FILLER_49_3004 ();
 sg13g2_fill_1 FILLER_49_3006 ();
 sg13g2_fill_2 FILLER_49_3034 ();
 sg13g2_decap_4 FILLER_49_3073 ();
 sg13g2_fill_2 FILLER_49_3077 ();
 sg13g2_fill_2 FILLER_49_3092 ();
 sg13g2_fill_1 FILLER_49_3094 ();
 sg13g2_fill_2 FILLER_49_3100 ();
 sg13g2_fill_1 FILLER_49_3115 ();
 sg13g2_fill_1 FILLER_49_3125 ();
 sg13g2_fill_2 FILLER_49_3177 ();
 sg13g2_fill_1 FILLER_49_3179 ();
 sg13g2_decap_4 FILLER_49_3217 ();
 sg13g2_fill_1 FILLER_49_3221 ();
 sg13g2_fill_2 FILLER_49_3258 ();
 sg13g2_fill_1 FILLER_49_3260 ();
 sg13g2_decap_8 FILLER_49_3274 ();
 sg13g2_fill_2 FILLER_49_3281 ();
 sg13g2_fill_1 FILLER_49_3283 ();
 sg13g2_decap_4 FILLER_49_3297 ();
 sg13g2_fill_2 FILLER_49_3323 ();
 sg13g2_fill_1 FILLER_49_3333 ();
 sg13g2_fill_1 FILLER_49_3342 ();
 sg13g2_fill_2 FILLER_49_3346 ();
 sg13g2_fill_1 FILLER_49_3348 ();
 sg13g2_fill_2 FILLER_49_3365 ();
 sg13g2_fill_1 FILLER_49_3387 ();
 sg13g2_decap_4 FILLER_49_3423 ();
 sg13g2_fill_1 FILLER_49_3427 ();
 sg13g2_decap_8 FILLER_49_3455 ();
 sg13g2_decap_8 FILLER_49_3462 ();
 sg13g2_decap_8 FILLER_49_3469 ();
 sg13g2_decap_8 FILLER_49_3476 ();
 sg13g2_decap_8 FILLER_49_3483 ();
 sg13g2_decap_8 FILLER_49_3490 ();
 sg13g2_decap_8 FILLER_49_3497 ();
 sg13g2_decap_8 FILLER_49_3504 ();
 sg13g2_decap_8 FILLER_49_3511 ();
 sg13g2_decap_8 FILLER_49_3518 ();
 sg13g2_decap_8 FILLER_49_3525 ();
 sg13g2_decap_8 FILLER_49_3532 ();
 sg13g2_decap_8 FILLER_49_3539 ();
 sg13g2_decap_8 FILLER_49_3546 ();
 sg13g2_decap_8 FILLER_49_3553 ();
 sg13g2_decap_8 FILLER_49_3560 ();
 sg13g2_decap_8 FILLER_49_3567 ();
 sg13g2_decap_4 FILLER_49_3574 ();
 sg13g2_fill_2 FILLER_49_3578 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_4 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_decap_4 FILLER_50_145 ();
 sg13g2_decap_8 FILLER_50_165 ();
 sg13g2_decap_8 FILLER_50_172 ();
 sg13g2_decap_8 FILLER_50_179 ();
 sg13g2_decap_4 FILLER_50_186 ();
 sg13g2_fill_1 FILLER_50_206 ();
 sg13g2_fill_2 FILLER_50_211 ();
 sg13g2_decap_4 FILLER_50_217 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_244 ();
 sg13g2_fill_2 FILLER_50_251 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_decap_4 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_276 ();
 sg13g2_fill_2 FILLER_50_301 ();
 sg13g2_fill_2 FILLER_50_347 ();
 sg13g2_fill_1 FILLER_50_358 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_fill_1 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_424 ();
 sg13g2_fill_1 FILLER_50_446 ();
 sg13g2_fill_1 FILLER_50_451 ();
 sg13g2_fill_2 FILLER_50_503 ();
 sg13g2_decap_4 FILLER_50_533 ();
 sg13g2_decap_8 FILLER_50_550 ();
 sg13g2_fill_2 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_559 ();
 sg13g2_decap_8 FILLER_50_564 ();
 sg13g2_fill_1 FILLER_50_599 ();
 sg13g2_fill_2 FILLER_50_614 ();
 sg13g2_fill_1 FILLER_50_616 ();
 sg13g2_fill_2 FILLER_50_634 ();
 sg13g2_fill_2 FILLER_50_640 ();
 sg13g2_fill_1 FILLER_50_652 ();
 sg13g2_fill_2 FILLER_50_667 ();
 sg13g2_fill_1 FILLER_50_691 ();
 sg13g2_decap_8 FILLER_50_713 ();
 sg13g2_decap_4 FILLER_50_725 ();
 sg13g2_decap_8 FILLER_50_757 ();
 sg13g2_decap_8 FILLER_50_764 ();
 sg13g2_fill_1 FILLER_50_771 ();
 sg13g2_decap_8 FILLER_50_788 ();
 sg13g2_decap_8 FILLER_50_795 ();
 sg13g2_fill_1 FILLER_50_802 ();
 sg13g2_decap_8 FILLER_50_831 ();
 sg13g2_fill_1 FILLER_50_838 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_4 FILLER_50_889 ();
 sg13g2_fill_1 FILLER_50_893 ();
 sg13g2_fill_2 FILLER_50_916 ();
 sg13g2_fill_1 FILLER_50_918 ();
 sg13g2_decap_8 FILLER_50_941 ();
 sg13g2_fill_2 FILLER_50_975 ();
 sg13g2_fill_1 FILLER_50_977 ();
 sg13g2_decap_8 FILLER_50_982 ();
 sg13g2_decap_4 FILLER_50_989 ();
 sg13g2_fill_2 FILLER_50_1021 ();
 sg13g2_fill_2 FILLER_50_1032 ();
 sg13g2_decap_8 FILLER_50_1042 ();
 sg13g2_fill_1 FILLER_50_1099 ();
 sg13g2_decap_8 FILLER_50_1128 ();
 sg13g2_decap_8 FILLER_50_1158 ();
 sg13g2_decap_8 FILLER_50_1165 ();
 sg13g2_decap_8 FILLER_50_1172 ();
 sg13g2_decap_4 FILLER_50_1220 ();
 sg13g2_fill_2 FILLER_50_1247 ();
 sg13g2_fill_2 FILLER_50_1290 ();
 sg13g2_fill_1 FILLER_50_1301 ();
 sg13g2_decap_8 FILLER_50_1331 ();
 sg13g2_fill_2 FILLER_50_1338 ();
 sg13g2_fill_1 FILLER_50_1367 ();
 sg13g2_fill_2 FILLER_50_1395 ();
 sg13g2_decap_4 FILLER_50_1446 ();
 sg13g2_decap_4 FILLER_50_1505 ();
 sg13g2_fill_1 FILLER_50_1509 ();
 sg13g2_fill_2 FILLER_50_1548 ();
 sg13g2_fill_2 FILLER_50_1563 ();
 sg13g2_fill_1 FILLER_50_1593 ();
 sg13g2_decap_4 FILLER_50_1673 ();
 sg13g2_fill_2 FILLER_50_1677 ();
 sg13g2_fill_1 FILLER_50_1684 ();
 sg13g2_fill_2 FILLER_50_1690 ();
 sg13g2_fill_1 FILLER_50_1716 ();
 sg13g2_fill_2 FILLER_50_1735 ();
 sg13g2_fill_1 FILLER_50_1737 ();
 sg13g2_fill_2 FILLER_50_1785 ();
 sg13g2_fill_1 FILLER_50_1797 ();
 sg13g2_fill_1 FILLER_50_1831 ();
 sg13g2_fill_2 FILLER_50_1873 ();
 sg13g2_fill_2 FILLER_50_1884 ();
 sg13g2_fill_2 FILLER_50_1895 ();
 sg13g2_fill_2 FILLER_50_1933 ();
 sg13g2_fill_1 FILLER_50_1935 ();
 sg13g2_fill_1 FILLER_50_1959 ();
 sg13g2_fill_2 FILLER_50_1969 ();
 sg13g2_fill_1 FILLER_50_1971 ();
 sg13g2_fill_1 FILLER_50_2004 ();
 sg13g2_fill_2 FILLER_50_2014 ();
 sg13g2_decap_4 FILLER_50_2026 ();
 sg13g2_fill_2 FILLER_50_2049 ();
 sg13g2_fill_1 FILLER_50_2051 ();
 sg13g2_fill_2 FILLER_50_2103 ();
 sg13g2_fill_1 FILLER_50_2105 ();
 sg13g2_fill_1 FILLER_50_2129 ();
 sg13g2_fill_1 FILLER_50_2145 ();
 sg13g2_decap_8 FILLER_50_2164 ();
 sg13g2_fill_2 FILLER_50_2184 ();
 sg13g2_fill_1 FILLER_50_2186 ();
 sg13g2_fill_1 FILLER_50_2223 ();
 sg13g2_fill_2 FILLER_50_2233 ();
 sg13g2_fill_1 FILLER_50_2235 ();
 sg13g2_decap_4 FILLER_50_2245 ();
 sg13g2_fill_2 FILLER_50_2254 ();
 sg13g2_fill_2 FILLER_50_2266 ();
 sg13g2_fill_2 FILLER_50_2281 ();
 sg13g2_fill_1 FILLER_50_2283 ();
 sg13g2_fill_2 FILLER_50_2308 ();
 sg13g2_fill_2 FILLER_50_2345 ();
 sg13g2_fill_1 FILLER_50_2365 ();
 sg13g2_fill_1 FILLER_50_2396 ();
 sg13g2_decap_4 FILLER_50_2425 ();
 sg13g2_fill_2 FILLER_50_2429 ();
 sg13g2_fill_2 FILLER_50_2440 ();
 sg13g2_fill_1 FILLER_50_2442 ();
 sg13g2_fill_2 FILLER_50_2479 ();
 sg13g2_fill_1 FILLER_50_2481 ();
 sg13g2_fill_2 FILLER_50_2492 ();
 sg13g2_fill_1 FILLER_50_2494 ();
 sg13g2_fill_2 FILLER_50_2523 ();
 sg13g2_fill_2 FILLER_50_2535 ();
 sg13g2_fill_1 FILLER_50_2537 ();
 sg13g2_fill_1 FILLER_50_2548 ();
 sg13g2_fill_2 FILLER_50_2571 ();
 sg13g2_fill_1 FILLER_50_2573 ();
 sg13g2_fill_2 FILLER_50_2579 ();
 sg13g2_fill_1 FILLER_50_2595 ();
 sg13g2_fill_2 FILLER_50_2651 ();
 sg13g2_fill_2 FILLER_50_2662 ();
 sg13g2_fill_1 FILLER_50_2664 ();
 sg13g2_fill_1 FILLER_50_2679 ();
 sg13g2_fill_2 FILLER_50_2711 ();
 sg13g2_fill_2 FILLER_50_2783 ();
 sg13g2_fill_1 FILLER_50_2785 ();
 sg13g2_fill_1 FILLER_50_2852 ();
 sg13g2_fill_1 FILLER_50_2887 ();
 sg13g2_fill_2 FILLER_50_2923 ();
 sg13g2_fill_1 FILLER_50_2925 ();
 sg13g2_fill_2 FILLER_50_2960 ();
 sg13g2_fill_1 FILLER_50_2962 ();
 sg13g2_fill_2 FILLER_50_2980 ();
 sg13g2_fill_1 FILLER_50_2982 ();
 sg13g2_fill_2 FILLER_50_2996 ();
 sg13g2_fill_2 FILLER_50_3007 ();
 sg13g2_fill_1 FILLER_50_3047 ();
 sg13g2_fill_2 FILLER_50_3139 ();
 sg13g2_fill_1 FILLER_50_3141 ();
 sg13g2_fill_2 FILLER_50_3191 ();
 sg13g2_fill_1 FILLER_50_3211 ();
 sg13g2_fill_2 FILLER_50_3262 ();
 sg13g2_fill_1 FILLER_50_3274 ();
 sg13g2_decap_8 FILLER_50_3293 ();
 sg13g2_decap_4 FILLER_50_3308 ();
 sg13g2_fill_1 FILLER_50_3312 ();
 sg13g2_fill_1 FILLER_50_3318 ();
 sg13g2_decap_4 FILLER_50_3327 ();
 sg13g2_fill_1 FILLER_50_3342 ();
 sg13g2_fill_2 FILLER_50_3347 ();
 sg13g2_fill_1 FILLER_50_3349 ();
 sg13g2_decap_4 FILLER_50_3364 ();
 sg13g2_decap_8 FILLER_50_3385 ();
 sg13g2_decap_4 FILLER_50_3392 ();
 sg13g2_fill_1 FILLER_50_3396 ();
 sg13g2_decap_4 FILLER_50_3404 ();
 sg13g2_fill_1 FILLER_50_3433 ();
 sg13g2_decap_8 FILLER_50_3447 ();
 sg13g2_decap_8 FILLER_50_3454 ();
 sg13g2_decap_8 FILLER_50_3461 ();
 sg13g2_decap_8 FILLER_50_3468 ();
 sg13g2_decap_8 FILLER_50_3475 ();
 sg13g2_decap_8 FILLER_50_3482 ();
 sg13g2_decap_8 FILLER_50_3489 ();
 sg13g2_decap_8 FILLER_50_3496 ();
 sg13g2_decap_8 FILLER_50_3503 ();
 sg13g2_decap_8 FILLER_50_3510 ();
 sg13g2_decap_8 FILLER_50_3517 ();
 sg13g2_decap_8 FILLER_50_3524 ();
 sg13g2_decap_8 FILLER_50_3531 ();
 sg13g2_decap_8 FILLER_50_3538 ();
 sg13g2_decap_8 FILLER_50_3545 ();
 sg13g2_decap_8 FILLER_50_3552 ();
 sg13g2_decap_8 FILLER_50_3559 ();
 sg13g2_decap_8 FILLER_50_3566 ();
 sg13g2_decap_8 FILLER_50_3573 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_decap_4 FILLER_51_108 ();
 sg13g2_fill_2 FILLER_51_112 ();
 sg13g2_fill_2 FILLER_51_146 ();
 sg13g2_fill_1 FILLER_51_152 ();
 sg13g2_decap_4 FILLER_51_171 ();
 sg13g2_decap_8 FILLER_51_181 ();
 sg13g2_decap_8 FILLER_51_188 ();
 sg13g2_fill_2 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_197 ();
 sg13g2_fill_2 FILLER_51_222 ();
 sg13g2_fill_2 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_254 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_decap_4 FILLER_51_306 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_decap_4 FILLER_51_374 ();
 sg13g2_fill_2 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_fill_2 FILLER_51_418 ();
 sg13g2_fill_2 FILLER_51_447 ();
 sg13g2_fill_2 FILLER_51_454 ();
 sg13g2_fill_2 FILLER_51_482 ();
 sg13g2_decap_8 FILLER_51_519 ();
 sg13g2_decap_4 FILLER_51_526 ();
 sg13g2_fill_1 FILLER_51_530 ();
 sg13g2_decap_8 FILLER_51_544 ();
 sg13g2_decap_4 FILLER_51_551 ();
 sg13g2_fill_1 FILLER_51_583 ();
 sg13g2_decap_8 FILLER_51_607 ();
 sg13g2_fill_2 FILLER_51_614 ();
 sg13g2_fill_2 FILLER_51_625 ();
 sg13g2_fill_1 FILLER_51_627 ();
 sg13g2_fill_2 FILLER_51_689 ();
 sg13g2_fill_1 FILLER_51_758 ();
 sg13g2_fill_1 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_777 ();
 sg13g2_decap_4 FILLER_51_784 ();
 sg13g2_decap_8 FILLER_51_792 ();
 sg13g2_fill_1 FILLER_51_799 ();
 sg13g2_decap_4 FILLER_51_817 ();
 sg13g2_decap_8 FILLER_51_834 ();
 sg13g2_decap_4 FILLER_51_841 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_fill_1 FILLER_51_871 ();
 sg13g2_decap_8 FILLER_51_886 ();
 sg13g2_fill_2 FILLER_51_1001 ();
 sg13g2_fill_2 FILLER_51_1026 ();
 sg13g2_fill_1 FILLER_51_1028 ();
 sg13g2_decap_8 FILLER_51_1073 ();
 sg13g2_decap_8 FILLER_51_1080 ();
 sg13g2_decap_8 FILLER_51_1087 ();
 sg13g2_fill_1 FILLER_51_1094 ();
 sg13g2_fill_1 FILLER_51_1122 ();
 sg13g2_decap_4 FILLER_51_1127 ();
 sg13g2_fill_2 FILLER_51_1131 ();
 sg13g2_decap_4 FILLER_51_1174 ();
 sg13g2_fill_2 FILLER_51_1178 ();
 sg13g2_fill_1 FILLER_51_1184 ();
 sg13g2_decap_4 FILLER_51_1261 ();
 sg13g2_decap_4 FILLER_51_1309 ();
 sg13g2_fill_1 FILLER_51_1313 ();
 sg13g2_decap_8 FILLER_51_1341 ();
 sg13g2_decap_8 FILLER_51_1348 ();
 sg13g2_fill_2 FILLER_51_1355 ();
 sg13g2_fill_1 FILLER_51_1357 ();
 sg13g2_fill_2 FILLER_51_1372 ();
 sg13g2_decap_8 FILLER_51_1397 ();
 sg13g2_decap_4 FILLER_51_1404 ();
 sg13g2_fill_2 FILLER_51_1418 ();
 sg13g2_decap_4 FILLER_51_1434 ();
 sg13g2_decap_4 FILLER_51_1456 ();
 sg13g2_fill_2 FILLER_51_1474 ();
 sg13g2_fill_1 FILLER_51_1476 ();
 sg13g2_decap_4 FILLER_51_1482 ();
 sg13g2_decap_4 FILLER_51_1490 ();
 sg13g2_fill_2 FILLER_51_1494 ();
 sg13g2_fill_1 FILLER_51_1505 ();
 sg13g2_fill_1 FILLER_51_1519 ();
 sg13g2_fill_2 FILLER_51_1524 ();
 sg13g2_fill_1 FILLER_51_1526 ();
 sg13g2_decap_8 FILLER_51_1536 ();
 sg13g2_decap_8 FILLER_51_1543 ();
 sg13g2_decap_8 FILLER_51_1550 ();
 sg13g2_fill_2 FILLER_51_1584 ();
 sg13g2_fill_1 FILLER_51_1595 ();
 sg13g2_fill_1 FILLER_51_1605 ();
 sg13g2_fill_2 FILLER_51_1640 ();
 sg13g2_fill_2 FILLER_51_1688 ();
 sg13g2_fill_2 FILLER_51_1705 ();
 sg13g2_fill_2 FILLER_51_1772 ();
 sg13g2_fill_2 FILLER_51_1828 ();
 sg13g2_fill_1 FILLER_51_1830 ();
 sg13g2_decap_4 FILLER_51_1840 ();
 sg13g2_fill_1 FILLER_51_1872 ();
 sg13g2_fill_1 FILLER_51_1927 ();
 sg13g2_fill_2 FILLER_51_1988 ();
 sg13g2_fill_1 FILLER_51_1990 ();
 sg13g2_fill_2 FILLER_51_2018 ();
 sg13g2_fill_1 FILLER_51_2020 ();
 sg13g2_fill_2 FILLER_51_2077 ();
 sg13g2_fill_2 FILLER_51_2124 ();
 sg13g2_decap_4 FILLER_51_2140 ();
 sg13g2_fill_1 FILLER_51_2144 ();
 sg13g2_fill_2 FILLER_51_2158 ();
 sg13g2_fill_1 FILLER_51_2160 ();
 sg13g2_fill_1 FILLER_51_2198 ();
 sg13g2_decap_8 FILLER_51_2208 ();
 sg13g2_decap_8 FILLER_51_2215 ();
 sg13g2_fill_2 FILLER_51_2240 ();
 sg13g2_fill_1 FILLER_51_2242 ();
 sg13g2_decap_4 FILLER_51_2285 ();
 sg13g2_fill_1 FILLER_51_2289 ();
 sg13g2_decap_4 FILLER_51_2294 ();
 sg13g2_fill_2 FILLER_51_2298 ();
 sg13g2_fill_2 FILLER_51_2316 ();
 sg13g2_fill_1 FILLER_51_2318 ();
 sg13g2_fill_2 FILLER_51_2346 ();
 sg13g2_fill_1 FILLER_51_2348 ();
 sg13g2_fill_1 FILLER_51_2377 ();
 sg13g2_decap_4 FILLER_51_2434 ();
 sg13g2_fill_2 FILLER_51_2438 ();
 sg13g2_decap_8 FILLER_51_2502 ();
 sg13g2_decap_4 FILLER_51_2509 ();
 sg13g2_fill_2 FILLER_51_2513 ();
 sg13g2_fill_2 FILLER_51_2578 ();
 sg13g2_fill_1 FILLER_51_2580 ();
 sg13g2_fill_2 FILLER_51_2608 ();
 sg13g2_fill_1 FILLER_51_2610 ();
 sg13g2_fill_2 FILLER_51_2620 ();
 sg13g2_fill_2 FILLER_51_2700 ();
 sg13g2_fill_2 FILLER_51_2748 ();
 sg13g2_decap_8 FILLER_51_2837 ();
 sg13g2_decap_4 FILLER_51_2844 ();
 sg13g2_fill_2 FILLER_51_2889 ();
 sg13g2_fill_1 FILLER_51_2891 ();
 sg13g2_fill_2 FILLER_51_2906 ();
 sg13g2_fill_1 FILLER_51_2908 ();
 sg13g2_fill_1 FILLER_51_2919 ();
 sg13g2_fill_1 FILLER_51_2930 ();
 sg13g2_fill_2 FILLER_51_2945 ();
 sg13g2_fill_1 FILLER_51_2947 ();
 sg13g2_decap_4 FILLER_51_3051 ();
 sg13g2_fill_1 FILLER_51_3091 ();
 sg13g2_fill_2 FILLER_51_3115 ();
 sg13g2_fill_1 FILLER_51_3117 ();
 sg13g2_fill_2 FILLER_51_3127 ();
 sg13g2_fill_1 FILLER_51_3129 ();
 sg13g2_fill_1 FILLER_51_3180 ();
 sg13g2_fill_2 FILLER_51_3200 ();
 sg13g2_fill_1 FILLER_51_3202 ();
 sg13g2_fill_2 FILLER_51_3293 ();
 sg13g2_fill_1 FILLER_51_3295 ();
 sg13g2_decap_8 FILLER_51_3320 ();
 sg13g2_fill_2 FILLER_51_3327 ();
 sg13g2_fill_1 FILLER_51_3329 ();
 sg13g2_decap_4 FILLER_51_3347 ();
 sg13g2_decap_8 FILLER_51_3356 ();
 sg13g2_decap_8 FILLER_51_3363 ();
 sg13g2_decap_8 FILLER_51_3370 ();
 sg13g2_fill_1 FILLER_51_3377 ();
 sg13g2_fill_2 FILLER_51_3387 ();
 sg13g2_decap_4 FILLER_51_3393 ();
 sg13g2_fill_1 FILLER_51_3409 ();
 sg13g2_decap_4 FILLER_51_3415 ();
 sg13g2_decap_8 FILLER_51_3447 ();
 sg13g2_decap_8 FILLER_51_3454 ();
 sg13g2_decap_8 FILLER_51_3461 ();
 sg13g2_decap_8 FILLER_51_3468 ();
 sg13g2_decap_8 FILLER_51_3475 ();
 sg13g2_decap_8 FILLER_51_3482 ();
 sg13g2_decap_8 FILLER_51_3489 ();
 sg13g2_decap_8 FILLER_51_3496 ();
 sg13g2_decap_8 FILLER_51_3503 ();
 sg13g2_decap_8 FILLER_51_3510 ();
 sg13g2_decap_8 FILLER_51_3517 ();
 sg13g2_decap_8 FILLER_51_3524 ();
 sg13g2_decap_8 FILLER_51_3531 ();
 sg13g2_decap_8 FILLER_51_3538 ();
 sg13g2_decap_8 FILLER_51_3545 ();
 sg13g2_decap_8 FILLER_51_3552 ();
 sg13g2_decap_8 FILLER_51_3559 ();
 sg13g2_decap_8 FILLER_51_3566 ();
 sg13g2_decap_8 FILLER_51_3573 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_89 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_101 ();
 sg13g2_decap_4 FILLER_52_135 ();
 sg13g2_fill_1 FILLER_52_139 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_decap_8 FILLER_52_185 ();
 sg13g2_decap_4 FILLER_52_192 ();
 sg13g2_fill_2 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_205 ();
 sg13g2_decap_8 FILLER_52_216 ();
 sg13g2_fill_2 FILLER_52_223 ();
 sg13g2_fill_2 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_297 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_fill_2 FILLER_52_334 ();
 sg13g2_decap_4 FILLER_52_340 ();
 sg13g2_fill_2 FILLER_52_344 ();
 sg13g2_decap_4 FILLER_52_350 ();
 sg13g2_fill_2 FILLER_52_430 ();
 sg13g2_fill_1 FILLER_52_432 ();
 sg13g2_fill_2 FILLER_52_438 ();
 sg13g2_fill_1 FILLER_52_461 ();
 sg13g2_fill_1 FILLER_52_510 ();
 sg13g2_decap_4 FILLER_52_528 ();
 sg13g2_fill_2 FILLER_52_532 ();
 sg13g2_fill_2 FILLER_52_581 ();
 sg13g2_fill_2 FILLER_52_592 ();
 sg13g2_fill_1 FILLER_52_599 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_fill_1 FILLER_52_610 ();
 sg13g2_fill_2 FILLER_52_635 ();
 sg13g2_fill_1 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_669 ();
 sg13g2_fill_2 FILLER_52_695 ();
 sg13g2_fill_2 FILLER_52_704 ();
 sg13g2_fill_1 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_711 ();
 sg13g2_decap_4 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_725 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_fill_2 FILLER_52_742 ();
 sg13g2_fill_1 FILLER_52_744 ();
 sg13g2_fill_2 FILLER_52_749 ();
 sg13g2_fill_1 FILLER_52_751 ();
 sg13g2_decap_4 FILLER_52_836 ();
 sg13g2_fill_2 FILLER_52_873 ();
 sg13g2_fill_1 FILLER_52_875 ();
 sg13g2_decap_8 FILLER_52_917 ();
 sg13g2_decap_4 FILLER_52_924 ();
 sg13g2_fill_1 FILLER_52_941 ();
 sg13g2_decap_4 FILLER_52_946 ();
 sg13g2_fill_1 FILLER_52_950 ();
 sg13g2_fill_1 FILLER_52_978 ();
 sg13g2_decap_4 FILLER_52_982 ();
 sg13g2_fill_1 FILLER_52_1027 ();
 sg13g2_fill_2 FILLER_52_1050 ();
 sg13g2_fill_2 FILLER_52_1061 ();
 sg13g2_decap_8 FILLER_52_1071 ();
 sg13g2_fill_2 FILLER_52_1078 ();
 sg13g2_fill_1 FILLER_52_1080 ();
 sg13g2_decap_4 FILLER_52_1101 ();
 sg13g2_decap_4 FILLER_52_1159 ();
 sg13g2_fill_2 FILLER_52_1163 ();
 sg13g2_fill_1 FILLER_52_1174 ();
 sg13g2_fill_2 FILLER_52_1226 ();
 sg13g2_fill_2 FILLER_52_1248 ();
 sg13g2_fill_2 FILLER_52_1264 ();
 sg13g2_decap_8 FILLER_52_1271 ();
 sg13g2_fill_2 FILLER_52_1278 ();
 sg13g2_decap_8 FILLER_52_1334 ();
 sg13g2_decap_8 FILLER_52_1341 ();
 sg13g2_decap_4 FILLER_52_1348 ();
 sg13g2_fill_1 FILLER_52_1352 ();
 sg13g2_decap_4 FILLER_52_1366 ();
 sg13g2_fill_2 FILLER_52_1404 ();
 sg13g2_decap_4 FILLER_52_1419 ();
 sg13g2_fill_1 FILLER_52_1423 ();
 sg13g2_decap_8 FILLER_52_1465 ();
 sg13g2_fill_2 FILLER_52_1477 ();
 sg13g2_fill_1 FILLER_52_1479 ();
 sg13g2_fill_2 FILLER_52_1563 ();
 sg13g2_fill_2 FILLER_52_1606 ();
 sg13g2_decap_4 FILLER_52_1671 ();
 sg13g2_fill_1 FILLER_52_1675 ();
 sg13g2_fill_1 FILLER_52_1739 ();
 sg13g2_fill_2 FILLER_52_1749 ();
 sg13g2_fill_2 FILLER_52_1779 ();
 sg13g2_fill_1 FILLER_52_1781 ();
 sg13g2_fill_1 FILLER_52_1809 ();
 sg13g2_decap_4 FILLER_52_1842 ();
 sg13g2_fill_2 FILLER_52_1863 ();
 sg13g2_fill_2 FILLER_52_1879 ();
 sg13g2_fill_2 FILLER_52_1898 ();
 sg13g2_fill_1 FILLER_52_2035 ();
 sg13g2_fill_2 FILLER_52_2129 ();
 sg13g2_fill_1 FILLER_52_2131 ();
 sg13g2_decap_8 FILLER_52_2160 ();
 sg13g2_decap_8 FILLER_52_2167 ();
 sg13g2_decap_4 FILLER_52_2174 ();
 sg13g2_fill_2 FILLER_52_2178 ();
 sg13g2_fill_2 FILLER_52_2236 ();
 sg13g2_fill_1 FILLER_52_2238 ();
 sg13g2_decap_4 FILLER_52_2261 ();
 sg13g2_fill_2 FILLER_52_2265 ();
 sg13g2_fill_2 FILLER_52_2276 ();
 sg13g2_fill_1 FILLER_52_2278 ();
 sg13g2_fill_2 FILLER_52_2342 ();
 sg13g2_fill_1 FILLER_52_2357 ();
 sg13g2_fill_2 FILLER_52_2386 ();
 sg13g2_decap_8 FILLER_52_2397 ();
 sg13g2_fill_2 FILLER_52_2442 ();
 sg13g2_decap_8 FILLER_52_2503 ();
 sg13g2_fill_1 FILLER_52_2523 ();
 sg13g2_fill_2 FILLER_52_2562 ();
 sg13g2_fill_1 FILLER_52_2564 ();
 sg13g2_fill_1 FILLER_52_2592 ();
 sg13g2_fill_1 FILLER_52_2631 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_fill_1 FILLER_52_2670 ();
 sg13g2_fill_2 FILLER_52_2743 ();
 sg13g2_fill_2 FILLER_52_2781 ();
 sg13g2_fill_1 FILLER_52_2811 ();
 sg13g2_fill_2 FILLER_52_2849 ();
 sg13g2_fill_2 FILLER_52_2861 ();
 sg13g2_fill_1 FILLER_52_2863 ();
 sg13g2_fill_2 FILLER_52_2910 ();
 sg13g2_fill_2 FILLER_52_2957 ();
 sg13g2_fill_2 FILLER_52_2985 ();
 sg13g2_fill_2 FILLER_52_3015 ();
 sg13g2_fill_2 FILLER_52_3044 ();
 sg13g2_decap_8 FILLER_52_3069 ();
 sg13g2_fill_2 FILLER_52_3140 ();
 sg13g2_fill_2 FILLER_52_3181 ();
 sg13g2_decap_8 FILLER_52_3211 ();
 sg13g2_decap_4 FILLER_52_3218 ();
 sg13g2_fill_1 FILLER_52_3222 ();
 sg13g2_decap_8 FILLER_52_3232 ();
 sg13g2_decap_8 FILLER_52_3239 ();
 sg13g2_fill_2 FILLER_52_3246 ();
 sg13g2_fill_2 FILLER_52_3257 ();
 sg13g2_decap_8 FILLER_52_3279 ();
 sg13g2_decap_4 FILLER_52_3286 ();
 sg13g2_decap_8 FILLER_52_3308 ();
 sg13g2_decap_8 FILLER_52_3315 ();
 sg13g2_decap_8 FILLER_52_3322 ();
 sg13g2_fill_2 FILLER_52_3329 ();
 sg13g2_fill_1 FILLER_52_3331 ();
 sg13g2_fill_2 FILLER_52_3355 ();
 sg13g2_fill_1 FILLER_52_3357 ();
 sg13g2_fill_2 FILLER_52_3376 ();
 sg13g2_fill_1 FILLER_52_3378 ();
 sg13g2_fill_2 FILLER_52_3392 ();
 sg13g2_fill_1 FILLER_52_3394 ();
 sg13g2_fill_1 FILLER_52_3423 ();
 sg13g2_decap_8 FILLER_52_3428 ();
 sg13g2_decap_8 FILLER_52_3435 ();
 sg13g2_decap_8 FILLER_52_3442 ();
 sg13g2_decap_8 FILLER_52_3449 ();
 sg13g2_decap_8 FILLER_52_3456 ();
 sg13g2_decap_8 FILLER_52_3463 ();
 sg13g2_decap_8 FILLER_52_3470 ();
 sg13g2_decap_8 FILLER_52_3477 ();
 sg13g2_decap_8 FILLER_52_3484 ();
 sg13g2_decap_8 FILLER_52_3491 ();
 sg13g2_decap_8 FILLER_52_3498 ();
 sg13g2_decap_8 FILLER_52_3505 ();
 sg13g2_decap_8 FILLER_52_3512 ();
 sg13g2_decap_8 FILLER_52_3519 ();
 sg13g2_decap_8 FILLER_52_3526 ();
 sg13g2_decap_8 FILLER_52_3533 ();
 sg13g2_decap_8 FILLER_52_3540 ();
 sg13g2_decap_8 FILLER_52_3547 ();
 sg13g2_decap_8 FILLER_52_3554 ();
 sg13g2_decap_8 FILLER_52_3561 ();
 sg13g2_decap_8 FILLER_52_3568 ();
 sg13g2_decap_4 FILLER_52_3575 ();
 sg13g2_fill_1 FILLER_52_3579 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_fill_2 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_121 ();
 sg13g2_decap_4 FILLER_53_135 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_decap_4 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_214 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_1 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_292 ();
 sg13g2_fill_1 FILLER_53_296 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_decap_4 FILLER_53_386 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_461 ();
 sg13g2_fill_2 FILLER_53_467 ();
 sg13g2_fill_1 FILLER_53_469 ();
 sg13g2_decap_8 FILLER_53_528 ();
 sg13g2_fill_2 FILLER_53_535 ();
 sg13g2_fill_2 FILLER_53_542 ();
 sg13g2_fill_1 FILLER_53_544 ();
 sg13g2_fill_2 FILLER_53_562 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_decap_4 FILLER_53_633 ();
 sg13g2_decap_4 FILLER_53_641 ();
 sg13g2_fill_1 FILLER_53_661 ();
 sg13g2_fill_2 FILLER_53_671 ();
 sg13g2_fill_1 FILLER_53_673 ();
 sg13g2_decap_8 FILLER_53_683 ();
 sg13g2_decap_8 FILLER_53_690 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_decap_4 FILLER_53_839 ();
 sg13g2_fill_1 FILLER_53_886 ();
 sg13g2_decap_8 FILLER_53_896 ();
 sg13g2_decap_8 FILLER_53_903 ();
 sg13g2_fill_2 FILLER_53_941 ();
 sg13g2_fill_1 FILLER_53_943 ();
 sg13g2_decap_4 FILLER_53_963 ();
 sg13g2_fill_2 FILLER_53_967 ();
 sg13g2_fill_1 FILLER_53_993 ();
 sg13g2_decap_8 FILLER_53_998 ();
 sg13g2_fill_2 FILLER_53_1009 ();
 sg13g2_fill_1 FILLER_53_1011 ();
 sg13g2_fill_2 FILLER_53_1017 ();
 sg13g2_fill_1 FILLER_53_1019 ();
 sg13g2_fill_1 FILLER_53_1025 ();
 sg13g2_decap_4 FILLER_53_1035 ();
 sg13g2_fill_1 FILLER_53_1039 ();
 sg13g2_fill_2 FILLER_53_1061 ();
 sg13g2_decap_4 FILLER_53_1076 ();
 sg13g2_fill_1 FILLER_53_1080 ();
 sg13g2_fill_1 FILLER_53_1089 ();
 sg13g2_fill_2 FILLER_53_1099 ();
 sg13g2_fill_1 FILLER_53_1101 ();
 sg13g2_decap_4 FILLER_53_1107 ();
 sg13g2_fill_1 FILLER_53_1111 ();
 sg13g2_decap_4 FILLER_53_1125 ();
 sg13g2_fill_2 FILLER_53_1148 ();
 sg13g2_fill_1 FILLER_53_1150 ();
 sg13g2_decap_4 FILLER_53_1155 ();
 sg13g2_fill_2 FILLER_53_1159 ();
 sg13g2_fill_1 FILLER_53_1189 ();
 sg13g2_decap_8 FILLER_53_1226 ();
 sg13g2_decap_4 FILLER_53_1249 ();
 sg13g2_fill_1 FILLER_53_1253 ();
 sg13g2_fill_2 FILLER_53_1266 ();
 sg13g2_fill_2 FILLER_53_1282 ();
 sg13g2_fill_1 FILLER_53_1284 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_fill_1 FILLER_53_1306 ();
 sg13g2_fill_1 FILLER_53_1329 ();
 sg13g2_decap_4 FILLER_53_1357 ();
 sg13g2_fill_2 FILLER_53_1374 ();
 sg13g2_fill_2 FILLER_53_1399 ();
 sg13g2_fill_1 FILLER_53_1401 ();
 sg13g2_fill_2 FILLER_53_1430 ();
 sg13g2_decap_8 FILLER_53_1458 ();
 sg13g2_decap_8 FILLER_53_1480 ();
 sg13g2_decap_8 FILLER_53_1487 ();
 sg13g2_decap_4 FILLER_53_1494 ();
 sg13g2_fill_2 FILLER_53_1528 ();
 sg13g2_fill_2 FILLER_53_1536 ();
 sg13g2_decap_4 FILLER_53_1551 ();
 sg13g2_fill_1 FILLER_53_1626 ();
 sg13g2_fill_1 FILLER_53_1642 ();
 sg13g2_decap_4 FILLER_53_1687 ();
 sg13g2_fill_2 FILLER_53_1691 ();
 sg13g2_decap_8 FILLER_53_1721 ();
 sg13g2_decap_8 FILLER_53_1728 ();
 sg13g2_decap_4 FILLER_53_1776 ();
 sg13g2_decap_4 FILLER_53_1793 ();
 sg13g2_decap_8 FILLER_53_1825 ();
 sg13g2_decap_4 FILLER_53_1832 ();
 sg13g2_decap_8 FILLER_53_1937 ();
 sg13g2_fill_1 FILLER_53_1944 ();
 sg13g2_fill_2 FILLER_53_1972 ();
 sg13g2_fill_1 FILLER_53_1974 ();
 sg13g2_decap_4 FILLER_53_2038 ();
 sg13g2_fill_1 FILLER_53_2042 ();
 sg13g2_fill_2 FILLER_53_2069 ();
 sg13g2_fill_1 FILLER_53_2071 ();
 sg13g2_fill_2 FILLER_53_2090 ();
 sg13g2_fill_1 FILLER_53_2092 ();
 sg13g2_fill_1 FILLER_53_2120 ();
 sg13g2_decap_8 FILLER_53_2152 ();
 sg13g2_fill_1 FILLER_53_2159 ();
 sg13g2_decap_4 FILLER_53_2187 ();
 sg13g2_fill_1 FILLER_53_2191 ();
 sg13g2_decap_8 FILLER_53_2196 ();
 sg13g2_fill_2 FILLER_53_2272 ();
 sg13g2_decap_4 FILLER_53_2284 ();
 sg13g2_fill_2 FILLER_53_2288 ();
 sg13g2_fill_2 FILLER_53_2309 ();
 sg13g2_fill_1 FILLER_53_2311 ();
 sg13g2_fill_2 FILLER_53_2322 ();
 sg13g2_fill_2 FILLER_53_2337 ();
 sg13g2_fill_1 FILLER_53_2339 ();
 sg13g2_decap_4 FILLER_53_2370 ();
 sg13g2_fill_2 FILLER_53_2387 ();
 sg13g2_fill_2 FILLER_53_2393 ();
 sg13g2_fill_2 FILLER_53_2421 ();
 sg13g2_fill_1 FILLER_53_2423 ();
 sg13g2_fill_1 FILLER_53_2451 ();
 sg13g2_fill_2 FILLER_53_2461 ();
 sg13g2_fill_1 FILLER_53_2463 ();
 sg13g2_decap_4 FILLER_53_2520 ();
 sg13g2_fill_1 FILLER_53_2524 ();
 sg13g2_decap_8 FILLER_53_2552 ();
 sg13g2_decap_8 FILLER_53_2591 ();
 sg13g2_fill_1 FILLER_53_2598 ();
 sg13g2_decap_8 FILLER_53_2603 ();
 sg13g2_decap_8 FILLER_53_2610 ();
 sg13g2_decap_4 FILLER_53_2617 ();
 sg13g2_fill_1 FILLER_53_2652 ();
 sg13g2_fill_2 FILLER_53_2743 ();
 sg13g2_decap_8 FILLER_53_2758 ();
 sg13g2_decap_4 FILLER_53_2765 ();
 sg13g2_fill_1 FILLER_53_2769 ();
 sg13g2_fill_2 FILLER_53_2788 ();
 sg13g2_fill_1 FILLER_53_2790 ();
 sg13g2_decap_4 FILLER_53_2832 ();
 sg13g2_fill_1 FILLER_53_2836 ();
 sg13g2_fill_2 FILLER_53_2863 ();
 sg13g2_fill_2 FILLER_53_2874 ();
 sg13g2_fill_1 FILLER_53_2876 ();
 sg13g2_fill_1 FILLER_53_2891 ();
 sg13g2_fill_2 FILLER_53_2996 ();
 sg13g2_fill_1 FILLER_53_2998 ();
 sg13g2_fill_1 FILLER_53_3008 ();
 sg13g2_fill_2 FILLER_53_3041 ();
 sg13g2_decap_8 FILLER_53_3048 ();
 sg13g2_fill_2 FILLER_53_3055 ();
 sg13g2_fill_2 FILLER_53_3084 ();
 sg13g2_fill_1 FILLER_53_3086 ();
 sg13g2_decap_4 FILLER_53_3118 ();
 sg13g2_fill_2 FILLER_53_3122 ();
 sg13g2_fill_2 FILLER_53_3133 ();
 sg13g2_decap_4 FILLER_53_3200 ();
 sg13g2_fill_2 FILLER_53_3204 ();
 sg13g2_decap_4 FILLER_53_3219 ();
 sg13g2_fill_2 FILLER_53_3223 ();
 sg13g2_decap_8 FILLER_53_3239 ();
 sg13g2_fill_1 FILLER_53_3246 ();
 sg13g2_decap_4 FILLER_53_3255 ();
 sg13g2_fill_1 FILLER_53_3259 ();
 sg13g2_decap_8 FILLER_53_3273 ();
 sg13g2_fill_2 FILLER_53_3280 ();
 sg13g2_fill_1 FILLER_53_3282 ();
 sg13g2_fill_1 FILLER_53_3288 ();
 sg13g2_fill_1 FILLER_53_3317 ();
 sg13g2_fill_1 FILLER_53_3327 ();
 sg13g2_fill_2 FILLER_53_3345 ();
 sg13g2_fill_1 FILLER_53_3347 ();
 sg13g2_fill_2 FILLER_53_3361 ();
 sg13g2_fill_1 FILLER_53_3363 ();
 sg13g2_fill_2 FILLER_53_3379 ();
 sg13g2_fill_1 FILLER_53_3381 ();
 sg13g2_decap_8 FILLER_53_3391 ();
 sg13g2_fill_2 FILLER_53_3398 ();
 sg13g2_decap_8 FILLER_53_3412 ();
 sg13g2_fill_2 FILLER_53_3419 ();
 sg13g2_fill_1 FILLER_53_3421 ();
 sg13g2_decap_8 FILLER_53_3426 ();
 sg13g2_decap_8 FILLER_53_3433 ();
 sg13g2_decap_8 FILLER_53_3440 ();
 sg13g2_decap_8 FILLER_53_3447 ();
 sg13g2_decap_8 FILLER_53_3454 ();
 sg13g2_decap_8 FILLER_53_3461 ();
 sg13g2_decap_8 FILLER_53_3468 ();
 sg13g2_decap_8 FILLER_53_3475 ();
 sg13g2_decap_8 FILLER_53_3482 ();
 sg13g2_decap_8 FILLER_53_3489 ();
 sg13g2_decap_8 FILLER_53_3496 ();
 sg13g2_decap_8 FILLER_53_3503 ();
 sg13g2_decap_8 FILLER_53_3510 ();
 sg13g2_decap_8 FILLER_53_3517 ();
 sg13g2_decap_8 FILLER_53_3524 ();
 sg13g2_decap_8 FILLER_53_3531 ();
 sg13g2_decap_8 FILLER_53_3538 ();
 sg13g2_decap_8 FILLER_53_3545 ();
 sg13g2_decap_8 FILLER_53_3552 ();
 sg13g2_decap_8 FILLER_53_3559 ();
 sg13g2_decap_8 FILLER_53_3566 ();
 sg13g2_decap_8 FILLER_53_3573 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_78 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_fill_2 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_94 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_181 ();
 sg13g2_fill_2 FILLER_54_245 ();
 sg13g2_fill_1 FILLER_54_247 ();
 sg13g2_fill_2 FILLER_54_253 ();
 sg13g2_decap_4 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_264 ();
 sg13g2_decap_4 FILLER_54_297 ();
 sg13g2_fill_2 FILLER_54_301 ();
 sg13g2_decap_4 FILLER_54_356 ();
 sg13g2_fill_1 FILLER_54_405 ();
 sg13g2_fill_1 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_488 ();
 sg13g2_fill_2 FILLER_54_511 ();
 sg13g2_fill_1 FILLER_54_513 ();
 sg13g2_fill_2 FILLER_54_534 ();
 sg13g2_fill_1 FILLER_54_536 ();
 sg13g2_fill_2 FILLER_54_542 ();
 sg13g2_fill_1 FILLER_54_544 ();
 sg13g2_fill_2 FILLER_54_555 ();
 sg13g2_decap_8 FILLER_54_562 ();
 sg13g2_decap_8 FILLER_54_573 ();
 sg13g2_fill_2 FILLER_54_611 ();
 sg13g2_fill_1 FILLER_54_613 ();
 sg13g2_fill_2 FILLER_54_619 ();
 sg13g2_decap_8 FILLER_54_635 ();
 sg13g2_decap_8 FILLER_54_642 ();
 sg13g2_fill_2 FILLER_54_649 ();
 sg13g2_fill_1 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_660 ();
 sg13g2_fill_2 FILLER_54_680 ();
 sg13g2_decap_8 FILLER_54_695 ();
 sg13g2_fill_1 FILLER_54_706 ();
 sg13g2_decap_4 FILLER_54_716 ();
 sg13g2_fill_2 FILLER_54_720 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_fill_2 FILLER_54_743 ();
 sg13g2_fill_1 FILLER_54_745 ();
 sg13g2_fill_2 FILLER_54_752 ();
 sg13g2_decap_8 FILLER_54_776 ();
 sg13g2_fill_2 FILLER_54_783 ();
 sg13g2_fill_2 FILLER_54_791 ();
 sg13g2_fill_1 FILLER_54_809 ();
 sg13g2_fill_1 FILLER_54_818 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_fill_1 FILLER_54_864 ();
 sg13g2_decap_8 FILLER_54_882 ();
 sg13g2_decap_4 FILLER_54_889 ();
 sg13g2_decap_4 FILLER_54_924 ();
 sg13g2_decap_4 FILLER_54_965 ();
 sg13g2_fill_2 FILLER_54_969 ();
 sg13g2_decap_8 FILLER_54_976 ();
 sg13g2_fill_1 FILLER_54_983 ();
 sg13g2_fill_2 FILLER_54_997 ();
 sg13g2_decap_4 FILLER_54_1027 ();
 sg13g2_fill_2 FILLER_54_1031 ();
 sg13g2_decap_4 FILLER_54_1038 ();
 sg13g2_fill_2 FILLER_54_1055 ();
 sg13g2_fill_1 FILLER_54_1057 ();
 sg13g2_decap_8 FILLER_54_1072 ();
 sg13g2_decap_8 FILLER_54_1079 ();
 sg13g2_decap_8 FILLER_54_1160 ();
 sg13g2_fill_2 FILLER_54_1184 ();
 sg13g2_decap_4 FILLER_54_1232 ();
 sg13g2_fill_1 FILLER_54_1236 ();
 sg13g2_fill_2 FILLER_54_1246 ();
 sg13g2_fill_1 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1254 ();
 sg13g2_fill_2 FILLER_54_1261 ();
 sg13g2_fill_1 FILLER_54_1263 ();
 sg13g2_fill_2 FILLER_54_1282 ();
 sg13g2_fill_1 FILLER_54_1284 ();
 sg13g2_fill_1 FILLER_54_1315 ();
 sg13g2_fill_1 FILLER_54_1339 ();
 sg13g2_fill_2 FILLER_54_1363 ();
 sg13g2_decap_4 FILLER_54_1402 ();
 sg13g2_fill_1 FILLER_54_1406 ();
 sg13g2_fill_1 FILLER_54_1414 ();
 sg13g2_fill_2 FILLER_54_1428 ();
 sg13g2_fill_1 FILLER_54_1430 ();
 sg13g2_fill_2 FILLER_54_1449 ();
 sg13g2_fill_2 FILLER_54_1469 ();
 sg13g2_fill_1 FILLER_54_1471 ();
 sg13g2_fill_2 FILLER_54_1480 ();
 sg13g2_fill_1 FILLER_54_1482 ();
 sg13g2_fill_1 FILLER_54_1493 ();
 sg13g2_fill_2 FILLER_54_1508 ();
 sg13g2_decap_4 FILLER_54_1515 ();
 sg13g2_fill_1 FILLER_54_1519 ();
 sg13g2_fill_2 FILLER_54_1530 ();
 sg13g2_decap_8 FILLER_54_1578 ();
 sg13g2_decap_8 FILLER_54_1585 ();
 sg13g2_fill_1 FILLER_54_1592 ();
 sg13g2_fill_2 FILLER_54_1598 ();
 sg13g2_fill_1 FILLER_54_1600 ();
 sg13g2_fill_1 FILLER_54_1651 ();
 sg13g2_fill_2 FILLER_54_1656 ();
 sg13g2_decap_4 FILLER_54_1678 ();
 sg13g2_fill_2 FILLER_54_1682 ();
 sg13g2_decap_8 FILLER_54_1719 ();
 sg13g2_decap_4 FILLER_54_1726 ();
 sg13g2_fill_2 FILLER_54_1730 ();
 sg13g2_decap_8 FILLER_54_1815 ();
 sg13g2_decap_4 FILLER_54_1849 ();
 sg13g2_fill_1 FILLER_54_1853 ();
 sg13g2_decap_8 FILLER_54_1877 ();
 sg13g2_fill_2 FILLER_54_1921 ();
 sg13g2_decap_8 FILLER_54_1928 ();
 sg13g2_decap_8 FILLER_54_1935 ();
 sg13g2_decap_4 FILLER_54_1942 ();
 sg13g2_fill_2 FILLER_54_1972 ();
 sg13g2_fill_2 FILLER_54_2001 ();
 sg13g2_decap_8 FILLER_54_2040 ();
 sg13g2_fill_1 FILLER_54_2047 ();
 sg13g2_decap_4 FILLER_54_2114 ();
 sg13g2_fill_2 FILLER_54_2118 ();
 sg13g2_decap_4 FILLER_54_2139 ();
 sg13g2_fill_1 FILLER_54_2143 ();
 sg13g2_decap_8 FILLER_54_2173 ();
 sg13g2_decap_8 FILLER_54_2190 ();
 sg13g2_decap_4 FILLER_54_2243 ();
 sg13g2_fill_2 FILLER_54_2247 ();
 sg13g2_decap_4 FILLER_54_2314 ();
 sg13g2_fill_1 FILLER_54_2318 ();
 sg13g2_decap_4 FILLER_54_2345 ();
 sg13g2_fill_2 FILLER_54_2349 ();
 sg13g2_fill_2 FILLER_54_2378 ();
 sg13g2_fill_1 FILLER_54_2380 ();
 sg13g2_fill_2 FILLER_54_2408 ();
 sg13g2_decap_4 FILLER_54_2437 ();
 sg13g2_fill_1 FILLER_54_2441 ();
 sg13g2_decap_4 FILLER_54_2479 ();
 sg13g2_fill_1 FILLER_54_2483 ();
 sg13g2_decap_4 FILLER_54_2494 ();
 sg13g2_fill_2 FILLER_54_2498 ();
 sg13g2_decap_4 FILLER_54_2553 ();
 sg13g2_fill_1 FILLER_54_2557 ();
 sg13g2_decap_8 FILLER_54_2598 ();
 sg13g2_fill_2 FILLER_54_2605 ();
 sg13g2_fill_1 FILLER_54_2607 ();
 sg13g2_decap_4 FILLER_54_2631 ();
 sg13g2_fill_1 FILLER_54_2635 ();
 sg13g2_fill_1 FILLER_54_2646 ();
 sg13g2_decap_4 FILLER_54_2675 ();
 sg13g2_fill_2 FILLER_54_2679 ();
 sg13g2_fill_1 FILLER_54_2721 ();
 sg13g2_decap_8 FILLER_54_2758 ();
 sg13g2_decap_4 FILLER_54_2765 ();
 sg13g2_fill_1 FILLER_54_2769 ();
 sg13g2_fill_1 FILLER_54_2805 ();
 sg13g2_fill_2 FILLER_54_2843 ();
 sg13g2_fill_1 FILLER_54_2921 ();
 sg13g2_fill_1 FILLER_54_2926 ();
 sg13g2_decap_4 FILLER_54_2945 ();
 sg13g2_fill_2 FILLER_54_2949 ();
 sg13g2_fill_1 FILLER_54_2969 ();
 sg13g2_fill_1 FILLER_54_3022 ();
 sg13g2_decap_8 FILLER_54_3050 ();
 sg13g2_fill_2 FILLER_54_3057 ();
 sg13g2_decap_8 FILLER_54_3069 ();
 sg13g2_fill_2 FILLER_54_3076 ();
 sg13g2_decap_8 FILLER_54_3087 ();
 sg13g2_fill_2 FILLER_54_3107 ();
 sg13g2_fill_1 FILLER_54_3109 ();
 sg13g2_fill_1 FILLER_54_3124 ();
 sg13g2_fill_2 FILLER_54_3148 ();
 sg13g2_fill_1 FILLER_54_3159 ();
 sg13g2_fill_1 FILLER_54_3192 ();
 sg13g2_fill_1 FILLER_54_3198 ();
 sg13g2_fill_2 FILLER_54_3207 ();
 sg13g2_decap_8 FILLER_54_3222 ();
 sg13g2_fill_2 FILLER_54_3243 ();
 sg13g2_fill_1 FILLER_54_3245 ();
 sg13g2_fill_2 FILLER_54_3267 ();
 sg13g2_decap_4 FILLER_54_3280 ();
 sg13g2_fill_1 FILLER_54_3284 ();
 sg13g2_decap_8 FILLER_54_3294 ();
 sg13g2_decap_4 FILLER_54_3301 ();
 sg13g2_fill_1 FILLER_54_3305 ();
 sg13g2_fill_2 FILLER_54_3311 ();
 sg13g2_fill_1 FILLER_54_3313 ();
 sg13g2_decap_8 FILLER_54_3319 ();
 sg13g2_decap_8 FILLER_54_3326 ();
 sg13g2_decap_4 FILLER_54_3333 ();
 sg13g2_decap_8 FILLER_54_3350 ();
 sg13g2_fill_2 FILLER_54_3357 ();
 sg13g2_fill_1 FILLER_54_3376 ();
 sg13g2_fill_2 FILLER_54_3398 ();
 sg13g2_decap_8 FILLER_54_3445 ();
 sg13g2_decap_8 FILLER_54_3452 ();
 sg13g2_decap_8 FILLER_54_3459 ();
 sg13g2_decap_8 FILLER_54_3466 ();
 sg13g2_decap_8 FILLER_54_3473 ();
 sg13g2_decap_8 FILLER_54_3480 ();
 sg13g2_decap_8 FILLER_54_3487 ();
 sg13g2_decap_8 FILLER_54_3494 ();
 sg13g2_decap_8 FILLER_54_3501 ();
 sg13g2_decap_8 FILLER_54_3508 ();
 sg13g2_decap_8 FILLER_54_3515 ();
 sg13g2_decap_8 FILLER_54_3522 ();
 sg13g2_decap_8 FILLER_54_3529 ();
 sg13g2_decap_8 FILLER_54_3536 ();
 sg13g2_decap_8 FILLER_54_3543 ();
 sg13g2_decap_8 FILLER_54_3550 ();
 sg13g2_decap_8 FILLER_54_3557 ();
 sg13g2_decap_8 FILLER_54_3564 ();
 sg13g2_decap_8 FILLER_54_3571 ();
 sg13g2_fill_2 FILLER_54_3578 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_116 ();
 sg13g2_decap_8 FILLER_55_121 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_decap_4 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_142 ();
 sg13g2_decap_8 FILLER_55_180 ();
 sg13g2_decap_8 FILLER_55_187 ();
 sg13g2_fill_1 FILLER_55_194 ();
 sg13g2_decap_4 FILLER_55_211 ();
 sg13g2_fill_2 FILLER_55_215 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_decap_4 FILLER_55_264 ();
 sg13g2_fill_2 FILLER_55_268 ();
 sg13g2_fill_2 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_348 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_447 ();
 sg13g2_decap_8 FILLER_55_454 ();
 sg13g2_fill_2 FILLER_55_466 ();
 sg13g2_fill_1 FILLER_55_468 ();
 sg13g2_fill_2 FILLER_55_506 ();
 sg13g2_fill_1 FILLER_55_517 ();
 sg13g2_decap_4 FILLER_55_551 ();
 sg13g2_fill_1 FILLER_55_555 ();
 sg13g2_decap_8 FILLER_55_584 ();
 sg13g2_fill_2 FILLER_55_591 ();
 sg13g2_fill_1 FILLER_55_593 ();
 sg13g2_fill_1 FILLER_55_599 ();
 sg13g2_decap_8 FILLER_55_604 ();
 sg13g2_decap_4 FILLER_55_611 ();
 sg13g2_fill_2 FILLER_55_615 ();
 sg13g2_decap_8 FILLER_55_636 ();
 sg13g2_fill_2 FILLER_55_643 ();
 sg13g2_fill_1 FILLER_55_645 ();
 sg13g2_decap_8 FILLER_55_660 ();
 sg13g2_decap_8 FILLER_55_667 ();
 sg13g2_fill_1 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_690 ();
 sg13g2_decap_4 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_719 ();
 sg13g2_fill_2 FILLER_55_755 ();
 sg13g2_decap_4 FILLER_55_785 ();
 sg13g2_fill_1 FILLER_55_789 ();
 sg13g2_fill_1 FILLER_55_797 ();
 sg13g2_fill_2 FILLER_55_820 ();
 sg13g2_fill_1 FILLER_55_822 ();
 sg13g2_fill_2 FILLER_55_833 ();
 sg13g2_fill_1 FILLER_55_835 ();
 sg13g2_fill_2 FILLER_55_849 ();
 sg13g2_fill_1 FILLER_55_856 ();
 sg13g2_fill_2 FILLER_55_879 ();
 sg13g2_fill_1 FILLER_55_881 ();
 sg13g2_fill_1 FILLER_55_900 ();
 sg13g2_fill_1 FILLER_55_908 ();
 sg13g2_fill_2 FILLER_55_918 ();
 sg13g2_fill_2 FILLER_55_969 ();
 sg13g2_fill_2 FILLER_55_976 ();
 sg13g2_fill_1 FILLER_55_978 ();
 sg13g2_decap_8 FILLER_55_1002 ();
 sg13g2_fill_2 FILLER_55_1009 ();
 sg13g2_fill_1 FILLER_55_1016 ();
 sg13g2_decap_8 FILLER_55_1027 ();
 sg13g2_decap_4 FILLER_55_1039 ();
 sg13g2_fill_1 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1114 ();
 sg13g2_fill_1 FILLER_55_1121 ();
 sg13g2_fill_2 FILLER_55_1131 ();
 sg13g2_fill_1 FILLER_55_1133 ();
 sg13g2_decap_8 FILLER_55_1153 ();
 sg13g2_decap_4 FILLER_55_1160 ();
 sg13g2_decap_8 FILLER_55_1196 ();
 sg13g2_decap_4 FILLER_55_1203 ();
 sg13g2_fill_1 FILLER_55_1223 ();
 sg13g2_decap_4 FILLER_55_1229 ();
 sg13g2_fill_2 FILLER_55_1233 ();
 sg13g2_fill_2 FILLER_55_1250 ();
 sg13g2_decap_4 FILLER_55_1265 ();
 sg13g2_fill_1 FILLER_55_1269 ();
 sg13g2_fill_2 FILLER_55_1275 ();
 sg13g2_fill_1 FILLER_55_1277 ();
 sg13g2_fill_2 FILLER_55_1307 ();
 sg13g2_fill_1 FILLER_55_1309 ();
 sg13g2_fill_2 FILLER_55_1370 ();
 sg13g2_fill_1 FILLER_55_1372 ();
 sg13g2_fill_1 FILLER_55_1378 ();
 sg13g2_decap_4 FILLER_55_1387 ();
 sg13g2_fill_1 FILLER_55_1404 ();
 sg13g2_decap_8 FILLER_55_1453 ();
 sg13g2_fill_1 FILLER_55_1468 ();
 sg13g2_decap_8 FILLER_55_1482 ();
 sg13g2_decap_8 FILLER_55_1489 ();
 sg13g2_fill_1 FILLER_55_1496 ();
 sg13g2_fill_2 FILLER_55_1509 ();
 sg13g2_fill_1 FILLER_55_1511 ();
 sg13g2_decap_4 FILLER_55_1517 ();
 sg13g2_fill_2 FILLER_55_1521 ();
 sg13g2_fill_2 FILLER_55_1529 ();
 sg13g2_decap_4 FILLER_55_1559 ();
 sg13g2_fill_2 FILLER_55_1583 ();
 sg13g2_decap_4 FILLER_55_1608 ();
 sg13g2_decap_8 FILLER_55_1617 ();
 sg13g2_fill_2 FILLER_55_1624 ();
 sg13g2_fill_1 FILLER_55_1626 ();
 sg13g2_decap_8 FILLER_55_1648 ();
 sg13g2_decap_8 FILLER_55_1655 ();
 sg13g2_decap_4 FILLER_55_1662 ();
 sg13g2_decap_8 FILLER_55_1676 ();
 sg13g2_decap_4 FILLER_55_1683 ();
 sg13g2_fill_2 FILLER_55_1713 ();
 sg13g2_decap_8 FILLER_55_1719 ();
 sg13g2_fill_1 FILLER_55_1726 ();
 sg13g2_fill_2 FILLER_55_1737 ();
 sg13g2_fill_1 FILLER_55_1739 ();
 sg13g2_fill_1 FILLER_55_1744 ();
 sg13g2_decap_4 FILLER_55_1749 ();
 sg13g2_fill_1 FILLER_55_1753 ();
 sg13g2_decap_8 FILLER_55_1773 ();
 sg13g2_decap_4 FILLER_55_1780 ();
 sg13g2_fill_1 FILLER_55_1784 ();
 sg13g2_decap_8 FILLER_55_1790 ();
 sg13g2_decap_8 FILLER_55_1797 ();
 sg13g2_fill_1 FILLER_55_1804 ();
 sg13g2_decap_8 FILLER_55_1834 ();
 sg13g2_decap_4 FILLER_55_1841 ();
 sg13g2_fill_1 FILLER_55_1845 ();
 sg13g2_decap_8 FILLER_55_1908 ();
 sg13g2_decap_4 FILLER_55_1942 ();
 sg13g2_fill_2 FILLER_55_1946 ();
 sg13g2_fill_2 FILLER_55_1970 ();
 sg13g2_fill_1 FILLER_55_1972 ();
 sg13g2_fill_2 FILLER_55_2005 ();
 sg13g2_fill_1 FILLER_55_2007 ();
 sg13g2_fill_1 FILLER_55_2027 ();
 sg13g2_fill_2 FILLER_55_2041 ();
 sg13g2_decap_8 FILLER_55_2053 ();
 sg13g2_fill_1 FILLER_55_2060 ();
 sg13g2_fill_2 FILLER_55_2074 ();
 sg13g2_decap_8 FILLER_55_2103 ();
 sg13g2_fill_2 FILLER_55_2110 ();
 sg13g2_decap_4 FILLER_55_2135 ();
 sg13g2_fill_2 FILLER_55_2139 ();
 sg13g2_fill_1 FILLER_55_2151 ();
 sg13g2_decap_4 FILLER_55_2179 ();
 sg13g2_decap_4 FILLER_55_2210 ();
 sg13g2_decap_8 FILLER_55_2227 ();
 sg13g2_fill_1 FILLER_55_2234 ();
 sg13g2_decap_8 FILLER_55_2272 ();
 sg13g2_decap_4 FILLER_55_2302 ();
 sg13g2_fill_1 FILLER_55_2306 ();
 sg13g2_fill_2 FILLER_55_2428 ();
 sg13g2_fill_2 FILLER_55_2440 ();
 sg13g2_fill_1 FILLER_55_2442 ();
 sg13g2_fill_2 FILLER_55_2501 ();
 sg13g2_fill_1 FILLER_55_2503 ();
 sg13g2_decap_8 FILLER_55_2571 ();
 sg13g2_fill_1 FILLER_55_2578 ();
 sg13g2_fill_2 FILLER_55_2616 ();
 sg13g2_fill_1 FILLER_55_2618 ();
 sg13g2_decap_4 FILLER_55_2673 ();
 sg13g2_fill_2 FILLER_55_2677 ();
 sg13g2_decap_8 FILLER_55_2689 ();
 sg13g2_fill_1 FILLER_55_2722 ();
 sg13g2_decap_8 FILLER_55_2813 ();
 sg13g2_decap_4 FILLER_55_2820 ();
 sg13g2_fill_2 FILLER_55_2824 ();
 sg13g2_decap_4 FILLER_55_2835 ();
 sg13g2_fill_1 FILLER_55_2839 ();
 sg13g2_fill_2 FILLER_55_2849 ();
 sg13g2_fill_1 FILLER_55_2851 ();
 sg13g2_decap_8 FILLER_55_2871 ();
 sg13g2_decap_8 FILLER_55_2878 ();
 sg13g2_decap_4 FILLER_55_2885 ();
 sg13g2_fill_1 FILLER_55_2889 ();
 sg13g2_decap_4 FILLER_55_2917 ();
 sg13g2_fill_1 FILLER_55_2948 ();
 sg13g2_fill_2 FILLER_55_2986 ();
 sg13g2_decap_4 FILLER_55_3001 ();
 sg13g2_decap_8 FILLER_55_3015 ();
 sg13g2_fill_2 FILLER_55_3022 ();
 sg13g2_fill_1 FILLER_55_3037 ();
 sg13g2_decap_8 FILLER_55_3052 ();
 sg13g2_decap_8 FILLER_55_3059 ();
 sg13g2_decap_4 FILLER_55_3094 ();
 sg13g2_fill_2 FILLER_55_3111 ();
 sg13g2_decap_8 FILLER_55_3141 ();
 sg13g2_fill_2 FILLER_55_3148 ();
 sg13g2_decap_4 FILLER_55_3153 ();
 sg13g2_fill_2 FILLER_55_3169 ();
 sg13g2_decap_8 FILLER_55_3189 ();
 sg13g2_decap_4 FILLER_55_3196 ();
 sg13g2_fill_2 FILLER_55_3207 ();
 sg13g2_decap_8 FILLER_55_3218 ();
 sg13g2_fill_2 FILLER_55_3225 ();
 sg13g2_decap_4 FILLER_55_3240 ();
 sg13g2_fill_1 FILLER_55_3244 ();
 sg13g2_decap_8 FILLER_55_3249 ();
 sg13g2_fill_2 FILLER_55_3256 ();
 sg13g2_fill_2 FILLER_55_3324 ();
 sg13g2_fill_1 FILLER_55_3326 ();
 sg13g2_fill_1 FILLER_55_3341 ();
 sg13g2_decap_4 FILLER_55_3355 ();
 sg13g2_fill_2 FILLER_55_3359 ();
 sg13g2_fill_1 FILLER_55_3386 ();
 sg13g2_fill_2 FILLER_55_3396 ();
 sg13g2_decap_4 FILLER_55_3402 ();
 sg13g2_fill_1 FILLER_55_3406 ();
 sg13g2_decap_8 FILLER_55_3435 ();
 sg13g2_decap_8 FILLER_55_3442 ();
 sg13g2_decap_8 FILLER_55_3449 ();
 sg13g2_decap_8 FILLER_55_3456 ();
 sg13g2_decap_8 FILLER_55_3463 ();
 sg13g2_decap_8 FILLER_55_3470 ();
 sg13g2_decap_8 FILLER_55_3477 ();
 sg13g2_decap_8 FILLER_55_3484 ();
 sg13g2_decap_8 FILLER_55_3491 ();
 sg13g2_decap_8 FILLER_55_3498 ();
 sg13g2_decap_8 FILLER_55_3505 ();
 sg13g2_decap_8 FILLER_55_3512 ();
 sg13g2_decap_8 FILLER_55_3519 ();
 sg13g2_decap_8 FILLER_55_3526 ();
 sg13g2_decap_8 FILLER_55_3533 ();
 sg13g2_decap_8 FILLER_55_3540 ();
 sg13g2_decap_8 FILLER_55_3547 ();
 sg13g2_decap_8 FILLER_55_3554 ();
 sg13g2_decap_8 FILLER_55_3561 ();
 sg13g2_decap_8 FILLER_55_3568 ();
 sg13g2_decap_4 FILLER_55_3575 ();
 sg13g2_fill_1 FILLER_55_3579 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_4 FILLER_56_63 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_72 ();
 sg13g2_decap_8 FILLER_56_79 ();
 sg13g2_decap_4 FILLER_56_86 ();
 sg13g2_decap_8 FILLER_56_142 ();
 sg13g2_fill_1 FILLER_56_157 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_2 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_2 FILLER_56_219 ();
 sg13g2_fill_1 FILLER_56_221 ();
 sg13g2_decap_4 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_273 ();
 sg13g2_decap_4 FILLER_56_289 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_367 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_397 ();
 sg13g2_fill_2 FILLER_56_425 ();
 sg13g2_fill_1 FILLER_56_427 ();
 sg13g2_fill_1 FILLER_56_507 ();
 sg13g2_decap_8 FILLER_56_513 ();
 sg13g2_fill_2 FILLER_56_520 ();
 sg13g2_fill_1 FILLER_56_522 ();
 sg13g2_decap_4 FILLER_56_532 ();
 sg13g2_decap_4 FILLER_56_540 ();
 sg13g2_fill_1 FILLER_56_553 ();
 sg13g2_fill_2 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_573 ();
 sg13g2_fill_2 FILLER_56_588 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_decap_8 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_612 ();
 sg13g2_decap_4 FILLER_56_637 ();
 sg13g2_fill_1 FILLER_56_641 ();
 sg13g2_decap_4 FILLER_56_666 ();
 sg13g2_fill_1 FILLER_56_670 ();
 sg13g2_decap_4 FILLER_56_697 ();
 sg13g2_fill_2 FILLER_56_709 ();
 sg13g2_decap_8 FILLER_56_720 ();
 sg13g2_fill_1 FILLER_56_727 ();
 sg13g2_decap_8 FILLER_56_737 ();
 sg13g2_decap_8 FILLER_56_744 ();
 sg13g2_fill_2 FILLER_56_764 ();
 sg13g2_decap_4 FILLER_56_775 ();
 sg13g2_fill_1 FILLER_56_779 ();
 sg13g2_fill_1 FILLER_56_824 ();
 sg13g2_fill_1 FILLER_56_847 ();
 sg13g2_fill_1 FILLER_56_876 ();
 sg13g2_fill_1 FILLER_56_885 ();
 sg13g2_decap_4 FILLER_56_912 ();
 sg13g2_fill_1 FILLER_56_916 ();
 sg13g2_fill_2 FILLER_56_935 ();
 sg13g2_fill_1 FILLER_56_937 ();
 sg13g2_decap_4 FILLER_56_947 ();
 sg13g2_fill_2 FILLER_56_968 ();
 sg13g2_decap_8 FILLER_56_974 ();
 sg13g2_fill_2 FILLER_56_981 ();
 sg13g2_fill_1 FILLER_56_983 ();
 sg13g2_decap_8 FILLER_56_1001 ();
 sg13g2_fill_1 FILLER_56_1021 ();
 sg13g2_fill_2 FILLER_56_1027 ();
 sg13g2_fill_1 FILLER_56_1029 ();
 sg13g2_decap_8 FILLER_56_1035 ();
 sg13g2_decap_8 FILLER_56_1042 ();
 sg13g2_fill_2 FILLER_56_1049 ();
 sg13g2_fill_2 FILLER_56_1062 ();
 sg13g2_fill_1 FILLER_56_1064 ();
 sg13g2_decap_8 FILLER_56_1092 ();
 sg13g2_fill_1 FILLER_56_1116 ();
 sg13g2_fill_1 FILLER_56_1152 ();
 sg13g2_fill_2 FILLER_56_1175 ();
 sg13g2_fill_1 FILLER_56_1177 ();
 sg13g2_decap_4 FILLER_56_1191 ();
 sg13g2_decap_8 FILLER_56_1208 ();
 sg13g2_decap_4 FILLER_56_1236 ();
 sg13g2_decap_8 FILLER_56_1245 ();
 sg13g2_decap_4 FILLER_56_1252 ();
 sg13g2_fill_2 FILLER_56_1256 ();
 sg13g2_decap_8 FILLER_56_1263 ();
 sg13g2_decap_8 FILLER_56_1277 ();
 sg13g2_fill_2 FILLER_56_1284 ();
 sg13g2_fill_1 FILLER_56_1286 ();
 sg13g2_fill_1 FILLER_56_1297 ();
 sg13g2_fill_2 FILLER_56_1316 ();
 sg13g2_fill_1 FILLER_56_1318 ();
 sg13g2_decap_8 FILLER_56_1347 ();
 sg13g2_fill_2 FILLER_56_1359 ();
 sg13g2_fill_2 FILLER_56_1366 ();
 sg13g2_fill_1 FILLER_56_1368 ();
 sg13g2_decap_8 FILLER_56_1379 ();
 sg13g2_decap_4 FILLER_56_1386 ();
 sg13g2_fill_1 FILLER_56_1390 ();
 sg13g2_fill_1 FILLER_56_1441 ();
 sg13g2_decap_4 FILLER_56_1452 ();
 sg13g2_fill_2 FILLER_56_1456 ();
 sg13g2_fill_1 FILLER_56_1463 ();
 sg13g2_decap_8 FILLER_56_1468 ();
 sg13g2_decap_4 FILLER_56_1475 ();
 sg13g2_fill_1 FILLER_56_1485 ();
 sg13g2_decap_8 FILLER_56_1491 ();
 sg13g2_decap_8 FILLER_56_1498 ();
 sg13g2_fill_1 FILLER_56_1505 ();
 sg13g2_decap_4 FILLER_56_1526 ();
 sg13g2_fill_2 FILLER_56_1541 ();
 sg13g2_fill_2 FILLER_56_1556 ();
 sg13g2_fill_1 FILLER_56_1558 ();
 sg13g2_fill_2 FILLER_56_1584 ();
 sg13g2_fill_1 FILLER_56_1595 ();
 sg13g2_fill_1 FILLER_56_1605 ();
 sg13g2_decap_4 FILLER_56_1614 ();
 sg13g2_fill_2 FILLER_56_1623 ();
 sg13g2_fill_1 FILLER_56_1625 ();
 sg13g2_fill_1 FILLER_56_1635 ();
 sg13g2_fill_2 FILLER_56_1651 ();
 sg13g2_fill_1 FILLER_56_1653 ();
 sg13g2_decap_4 FILLER_56_1684 ();
 sg13g2_fill_2 FILLER_56_1688 ();
 sg13g2_fill_2 FILLER_56_1722 ();
 sg13g2_fill_1 FILLER_56_1724 ();
 sg13g2_decap_8 FILLER_56_1875 ();
 sg13g2_decap_4 FILLER_56_1882 ();
 sg13g2_fill_2 FILLER_56_1913 ();
 sg13g2_fill_1 FILLER_56_1915 ();
 sg13g2_decap_4 FILLER_56_1926 ();
 sg13g2_fill_1 FILLER_56_1930 ();
 sg13g2_fill_1 FILLER_56_1940 ();
 sg13g2_decap_4 FILLER_56_1968 ();
 sg13g2_decap_4 FILLER_56_1995 ();
 sg13g2_fill_1 FILLER_56_1999 ();
 sg13g2_decap_4 FILLER_56_2046 ();
 sg13g2_fill_1 FILLER_56_2050 ();
 sg13g2_fill_2 FILLER_56_2078 ();
 sg13g2_fill_1 FILLER_56_2080 ();
 sg13g2_decap_4 FILLER_56_2103 ();
 sg13g2_fill_2 FILLER_56_2170 ();
 sg13g2_fill_2 FILLER_56_2181 ();
 sg13g2_fill_1 FILLER_56_2183 ();
 sg13g2_fill_2 FILLER_56_2207 ();
 sg13g2_decap_8 FILLER_56_2238 ();
 sg13g2_decap_4 FILLER_56_2245 ();
 sg13g2_fill_1 FILLER_56_2258 ();
 sg13g2_fill_1 FILLER_56_2268 ();
 sg13g2_fill_1 FILLER_56_2309 ();
 sg13g2_fill_2 FILLER_56_2364 ();
 sg13g2_fill_1 FILLER_56_2366 ();
 sg13g2_decap_4 FILLER_56_2380 ();
 sg13g2_fill_2 FILLER_56_2384 ();
 sg13g2_fill_2 FILLER_56_2422 ();
 sg13g2_decap_4 FILLER_56_2434 ();
 sg13g2_fill_1 FILLER_56_2438 ();
 sg13g2_decap_8 FILLER_56_2466 ();
 sg13g2_decap_8 FILLER_56_2473 ();
 sg13g2_fill_2 FILLER_56_2480 ();
 sg13g2_fill_2 FILLER_56_2511 ();
 sg13g2_fill_1 FILLER_56_2513 ();
 sg13g2_fill_2 FILLER_56_2527 ();
 sg13g2_decap_4 FILLER_56_2539 ();
 sg13g2_fill_1 FILLER_56_2552 ();
 sg13g2_decap_4 FILLER_56_2590 ();
 sg13g2_decap_8 FILLER_56_2626 ();
 sg13g2_fill_2 FILLER_56_2633 ();
 sg13g2_fill_1 FILLER_56_2635 ();
 sg13g2_fill_2 FILLER_56_2645 ();
 sg13g2_decap_8 FILLER_56_2651 ();
 sg13g2_decap_4 FILLER_56_2703 ();
 sg13g2_fill_1 FILLER_56_2707 ();
 sg13g2_fill_2 FILLER_56_2713 ();
 sg13g2_fill_1 FILLER_56_2715 ();
 sg13g2_decap_8 FILLER_56_2738 ();
 sg13g2_fill_2 FILLER_56_2745 ();
 sg13g2_fill_1 FILLER_56_2747 ();
 sg13g2_fill_2 FILLER_56_2767 ();
 sg13g2_fill_1 FILLER_56_2769 ();
 sg13g2_decap_4 FILLER_56_2790 ();
 sg13g2_fill_2 FILLER_56_2794 ();
 sg13g2_fill_1 FILLER_56_2819 ();
 sg13g2_decap_4 FILLER_56_2857 ();
 sg13g2_decap_4 FILLER_56_2888 ();
 sg13g2_decap_4 FILLER_56_2909 ();
 sg13g2_decap_8 FILLER_56_2972 ();
 sg13g2_decap_4 FILLER_56_3043 ();
 sg13g2_fill_1 FILLER_56_3047 ();
 sg13g2_fill_1 FILLER_56_3068 ();
 sg13g2_fill_1 FILLER_56_3122 ();
 sg13g2_fill_2 FILLER_56_3151 ();
 sg13g2_fill_1 FILLER_56_3157 ();
 sg13g2_fill_1 FILLER_56_3176 ();
 sg13g2_fill_2 FILLER_56_3181 ();
 sg13g2_fill_2 FILLER_56_3193 ();
 sg13g2_fill_2 FILLER_56_3209 ();
 sg13g2_fill_2 FILLER_56_3220 ();
 sg13g2_fill_1 FILLER_56_3222 ();
 sg13g2_decap_4 FILLER_56_3251 ();
 sg13g2_fill_2 FILLER_56_3255 ();
 sg13g2_fill_2 FILLER_56_3274 ();
 sg13g2_fill_1 FILLER_56_3276 ();
 sg13g2_decap_8 FILLER_56_3282 ();
 sg13g2_decap_8 FILLER_56_3289 ();
 sg13g2_decap_4 FILLER_56_3300 ();
 sg13g2_fill_2 FILLER_56_3313 ();
 sg13g2_fill_1 FILLER_56_3315 ();
 sg13g2_fill_1 FILLER_56_3330 ();
 sg13g2_decap_4 FILLER_56_3335 ();
 sg13g2_decap_8 FILLER_56_3361 ();
 sg13g2_fill_2 FILLER_56_3368 ();
 sg13g2_fill_1 FILLER_56_3370 ();
 sg13g2_fill_2 FILLER_56_3381 ();
 sg13g2_decap_8 FILLER_56_3405 ();
 sg13g2_decap_8 FILLER_56_3416 ();
 sg13g2_decap_8 FILLER_56_3423 ();
 sg13g2_decap_8 FILLER_56_3430 ();
 sg13g2_decap_8 FILLER_56_3437 ();
 sg13g2_decap_8 FILLER_56_3444 ();
 sg13g2_decap_8 FILLER_56_3451 ();
 sg13g2_decap_8 FILLER_56_3458 ();
 sg13g2_decap_8 FILLER_56_3465 ();
 sg13g2_decap_8 FILLER_56_3472 ();
 sg13g2_decap_8 FILLER_56_3479 ();
 sg13g2_decap_8 FILLER_56_3486 ();
 sg13g2_decap_8 FILLER_56_3493 ();
 sg13g2_decap_8 FILLER_56_3500 ();
 sg13g2_decap_8 FILLER_56_3507 ();
 sg13g2_decap_8 FILLER_56_3514 ();
 sg13g2_decap_8 FILLER_56_3521 ();
 sg13g2_decap_8 FILLER_56_3528 ();
 sg13g2_decap_8 FILLER_56_3535 ();
 sg13g2_decap_8 FILLER_56_3542 ();
 sg13g2_decap_8 FILLER_56_3549 ();
 sg13g2_decap_8 FILLER_56_3556 ();
 sg13g2_decap_8 FILLER_56_3563 ();
 sg13g2_decap_8 FILLER_56_3570 ();
 sg13g2_fill_2 FILLER_56_3577 ();
 sg13g2_fill_1 FILLER_56_3579 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_4 FILLER_57_56 ();
 sg13g2_fill_2 FILLER_57_60 ();
 sg13g2_fill_1 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_116 ();
 sg13g2_fill_2 FILLER_57_123 ();
 sg13g2_fill_1 FILLER_57_137 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_fill_1 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_176 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_217 ();
 sg13g2_fill_1 FILLER_57_219 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_264 ();
 sg13g2_fill_2 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_303 ();
 sg13g2_decap_4 FILLER_57_349 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_4 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_395 ();
 sg13g2_fill_1 FILLER_57_411 ();
 sg13g2_decap_4 FILLER_57_448 ();
 sg13g2_fill_2 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_536 ();
 sg13g2_decap_4 FILLER_57_542 ();
 sg13g2_fill_1 FILLER_57_573 ();
 sg13g2_fill_1 FILLER_57_597 ();
 sg13g2_fill_2 FILLER_57_613 ();
 sg13g2_decap_8 FILLER_57_627 ();
 sg13g2_decap_8 FILLER_57_634 ();
 sg13g2_decap_8 FILLER_57_641 ();
 sg13g2_decap_4 FILLER_57_672 ();
 sg13g2_fill_2 FILLER_57_676 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_fill_2 FILLER_57_700 ();
 sg13g2_fill_2 FILLER_57_715 ();
 sg13g2_fill_1 FILLER_57_717 ();
 sg13g2_decap_8 FILLER_57_723 ();
 sg13g2_fill_2 FILLER_57_743 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_decap_4 FILLER_57_800 ();
 sg13g2_fill_1 FILLER_57_804 ();
 sg13g2_decap_8 FILLER_57_822 ();
 sg13g2_fill_2 FILLER_57_829 ();
 sg13g2_fill_1 FILLER_57_831 ();
 sg13g2_decap_8 FILLER_57_836 ();
 sg13g2_decap_4 FILLER_57_843 ();
 sg13g2_fill_1 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_874 ();
 sg13g2_fill_2 FILLER_57_894 ();
 sg13g2_decap_4 FILLER_57_909 ();
 sg13g2_fill_1 FILLER_57_926 ();
 sg13g2_fill_2 FILLER_57_931 ();
 sg13g2_fill_1 FILLER_57_933 ();
 sg13g2_fill_2 FILLER_57_954 ();
 sg13g2_fill_1 FILLER_57_969 ();
 sg13g2_fill_2 FILLER_57_978 ();
 sg13g2_fill_2 FILLER_57_1000 ();
 sg13g2_decap_4 FILLER_57_1010 ();
 sg13g2_fill_2 FILLER_57_1014 ();
 sg13g2_decap_8 FILLER_57_1024 ();
 sg13g2_fill_2 FILLER_57_1031 ();
 sg13g2_fill_1 FILLER_57_1033 ();
 sg13g2_decap_4 FILLER_57_1051 ();
 sg13g2_fill_1 FILLER_57_1055 ();
 sg13g2_decap_8 FILLER_57_1060 ();
 sg13g2_decap_4 FILLER_57_1067 ();
 sg13g2_decap_8 FILLER_57_1076 ();
 sg13g2_decap_8 FILLER_57_1083 ();
 sg13g2_decap_4 FILLER_57_1090 ();
 sg13g2_fill_1 FILLER_57_1094 ();
 sg13g2_fill_1 FILLER_57_1108 ();
 sg13g2_decap_8 FILLER_57_1118 ();
 sg13g2_decap_8 FILLER_57_1125 ();
 sg13g2_fill_2 FILLER_57_1132 ();
 sg13g2_fill_1 FILLER_57_1187 ();
 sg13g2_decap_4 FILLER_57_1205 ();
 sg13g2_fill_2 FILLER_57_1209 ();
 sg13g2_fill_2 FILLER_57_1225 ();
 sg13g2_decap_4 FILLER_57_1230 ();
 sg13g2_fill_2 FILLER_57_1234 ();
 sg13g2_decap_4 FILLER_57_1241 ();
 sg13g2_fill_2 FILLER_57_1245 ();
 sg13g2_fill_2 FILLER_57_1265 ();
 sg13g2_fill_1 FILLER_57_1267 ();
 sg13g2_decap_8 FILLER_57_1273 ();
 sg13g2_decap_8 FILLER_57_1280 ();
 sg13g2_fill_1 FILLER_57_1287 ();
 sg13g2_decap_4 FILLER_57_1295 ();
 sg13g2_fill_1 FILLER_57_1299 ();
 sg13g2_decap_8 FILLER_57_1308 ();
 sg13g2_decap_8 FILLER_57_1315 ();
 sg13g2_fill_2 FILLER_57_1322 ();
 sg13g2_fill_2 FILLER_57_1328 ();
 sg13g2_fill_1 FILLER_57_1330 ();
 sg13g2_fill_1 FILLER_57_1344 ();
 sg13g2_decap_8 FILLER_57_1361 ();
 sg13g2_fill_1 FILLER_57_1368 ();
 sg13g2_decap_8 FILLER_57_1385 ();
 sg13g2_decap_8 FILLER_57_1392 ();
 sg13g2_fill_1 FILLER_57_1412 ();
 sg13g2_fill_2 FILLER_57_1420 ();
 sg13g2_fill_1 FILLER_57_1422 ();
 sg13g2_fill_1 FILLER_57_1428 ();
 sg13g2_fill_1 FILLER_57_1442 ();
 sg13g2_decap_4 FILLER_57_1459 ();
 sg13g2_fill_2 FILLER_57_1486 ();
 sg13g2_fill_1 FILLER_57_1488 ();
 sg13g2_decap_4 FILLER_57_1498 ();
 sg13g2_fill_1 FILLER_57_1502 ();
 sg13g2_fill_2 FILLER_57_1507 ();
 sg13g2_fill_1 FILLER_57_1509 ();
 sg13g2_decap_4 FILLER_57_1518 ();
 sg13g2_fill_1 FILLER_57_1522 ();
 sg13g2_fill_1 FILLER_57_1559 ();
 sg13g2_fill_2 FILLER_57_1581 ();
 sg13g2_fill_1 FILLER_57_1583 ();
 sg13g2_fill_1 FILLER_57_1593 ();
 sg13g2_decap_4 FILLER_57_1602 ();
 sg13g2_fill_2 FILLER_57_1606 ();
 sg13g2_fill_1 FILLER_57_1651 ();
 sg13g2_fill_1 FILLER_57_1657 ();
 sg13g2_fill_1 FILLER_57_1671 ();
 sg13g2_decap_4 FILLER_57_1691 ();
 sg13g2_fill_2 FILLER_57_1695 ();
 sg13g2_fill_2 FILLER_57_1707 ();
 sg13g2_decap_8 FILLER_57_1714 ();
 sg13g2_decap_8 FILLER_57_1721 ();
 sg13g2_fill_1 FILLER_57_1728 ();
 sg13g2_fill_2 FILLER_57_1738 ();
 sg13g2_fill_1 FILLER_57_1740 ();
 sg13g2_decap_8 FILLER_57_1746 ();
 sg13g2_fill_1 FILLER_57_1753 ();
 sg13g2_decap_4 FILLER_57_1770 ();
 sg13g2_fill_1 FILLER_57_1797 ();
 sg13g2_fill_1 FILLER_57_1807 ();
 sg13g2_decap_4 FILLER_57_1820 ();
 sg13g2_fill_1 FILLER_57_1824 ();
 sg13g2_fill_1 FILLER_57_1838 ();
 sg13g2_decap_8 FILLER_57_1848 ();
 sg13g2_fill_1 FILLER_57_1855 ();
 sg13g2_decap_4 FILLER_57_1879 ();
 sg13g2_fill_1 FILLER_57_1883 ();
 sg13g2_decap_8 FILLER_57_1894 ();
 sg13g2_fill_2 FILLER_57_1947 ();
 sg13g2_fill_2 FILLER_57_1982 ();
 sg13g2_fill_1 FILLER_57_1984 ();
 sg13g2_fill_2 FILLER_57_2021 ();
 sg13g2_fill_1 FILLER_57_2023 ();
 sg13g2_decap_4 FILLER_57_2033 ();
 sg13g2_fill_2 FILLER_57_2037 ();
 sg13g2_decap_4 FILLER_57_2079 ();
 sg13g2_fill_1 FILLER_57_2083 ();
 sg13g2_decap_4 FILLER_57_2111 ();
 sg13g2_fill_1 FILLER_57_2152 ();
 sg13g2_fill_2 FILLER_57_2167 ();
 sg13g2_fill_1 FILLER_57_2169 ();
 sg13g2_fill_2 FILLER_57_2180 ();
 sg13g2_decap_4 FILLER_57_2191 ();
 sg13g2_fill_1 FILLER_57_2195 ();
 sg13g2_decap_8 FILLER_57_2239 ();
 sg13g2_fill_1 FILLER_57_2278 ();
 sg13g2_fill_1 FILLER_57_2292 ();
 sg13g2_fill_2 FILLER_57_2315 ();
 sg13g2_decap_4 FILLER_57_2330 ();
 sg13g2_fill_1 FILLER_57_2334 ();
 sg13g2_fill_2 FILLER_57_2390 ();
 sg13g2_fill_1 FILLER_57_2411 ();
 sg13g2_decap_4 FILLER_57_2428 ();
 sg13g2_decap_8 FILLER_57_2459 ();
 sg13g2_decap_4 FILLER_57_2466 ();
 sg13g2_fill_1 FILLER_57_2470 ();
 sg13g2_fill_1 FILLER_57_2484 ();
 sg13g2_fill_2 FILLER_57_2503 ();
 sg13g2_fill_1 FILLER_57_2505 ();
 sg13g2_fill_1 FILLER_57_2533 ();
 sg13g2_decap_8 FILLER_57_2566 ();
 sg13g2_decap_8 FILLER_57_2582 ();
 sg13g2_decap_8 FILLER_57_2589 ();
 sg13g2_fill_1 FILLER_57_2596 ();
 sg13g2_decap_4 FILLER_57_2602 ();
 sg13g2_decap_4 FILLER_57_2639 ();
 sg13g2_decap_8 FILLER_57_2666 ();
 sg13g2_fill_2 FILLER_57_2673 ();
 sg13g2_fill_1 FILLER_57_2675 ();
 sg13g2_fill_1 FILLER_57_2680 ();
 sg13g2_fill_1 FILLER_57_2693 ();
 sg13g2_fill_1 FILLER_57_2703 ();
 sg13g2_fill_1 FILLER_57_2713 ();
 sg13g2_decap_4 FILLER_57_2736 ();
 sg13g2_fill_1 FILLER_57_2740 ();
 sg13g2_decap_4 FILLER_57_2777 ();
 sg13g2_fill_2 FILLER_57_2808 ();
 sg13g2_fill_1 FILLER_57_2810 ();
 sg13g2_decap_4 FILLER_57_2838 ();
 sg13g2_fill_2 FILLER_57_2847 ();
 sg13g2_fill_2 FILLER_57_2854 ();
 sg13g2_fill_1 FILLER_57_2861 ();
 sg13g2_fill_2 FILLER_57_2877 ();
 sg13g2_fill_1 FILLER_57_2879 ();
 sg13g2_decap_4 FILLER_57_2889 ();
 sg13g2_fill_2 FILLER_57_2916 ();
 sg13g2_fill_1 FILLER_57_2946 ();
 sg13g2_decap_8 FILLER_57_3003 ();
 sg13g2_decap_8 FILLER_57_3010 ();
 sg13g2_decap_8 FILLER_57_3036 ();
 sg13g2_fill_2 FILLER_57_3043 ();
 sg13g2_fill_2 FILLER_57_3054 ();
 sg13g2_fill_1 FILLER_57_3056 ();
 sg13g2_fill_2 FILLER_57_3094 ();
 sg13g2_fill_1 FILLER_57_3096 ();
 sg13g2_fill_1 FILLER_57_3236 ();
 sg13g2_decap_8 FILLER_57_3277 ();
 sg13g2_decap_4 FILLER_57_3284 ();
 sg13g2_fill_2 FILLER_57_3288 ();
 sg13g2_fill_1 FILLER_57_3300 ();
 sg13g2_decap_4 FILLER_57_3309 ();
 sg13g2_fill_1 FILLER_57_3313 ();
 sg13g2_decap_8 FILLER_57_3341 ();
 sg13g2_fill_1 FILLER_57_3348 ();
 sg13g2_decap_4 FILLER_57_3357 ();
 sg13g2_fill_1 FILLER_57_3361 ();
 sg13g2_fill_2 FILLER_57_3382 ();
 sg13g2_decap_8 FILLER_57_3412 ();
 sg13g2_decap_8 FILLER_57_3419 ();
 sg13g2_decap_8 FILLER_57_3426 ();
 sg13g2_decap_8 FILLER_57_3433 ();
 sg13g2_decap_8 FILLER_57_3440 ();
 sg13g2_decap_8 FILLER_57_3447 ();
 sg13g2_decap_8 FILLER_57_3454 ();
 sg13g2_decap_8 FILLER_57_3461 ();
 sg13g2_decap_8 FILLER_57_3468 ();
 sg13g2_decap_8 FILLER_57_3475 ();
 sg13g2_decap_8 FILLER_57_3482 ();
 sg13g2_decap_8 FILLER_57_3489 ();
 sg13g2_decap_8 FILLER_57_3496 ();
 sg13g2_decap_8 FILLER_57_3503 ();
 sg13g2_decap_8 FILLER_57_3510 ();
 sg13g2_decap_8 FILLER_57_3517 ();
 sg13g2_decap_8 FILLER_57_3524 ();
 sg13g2_decap_8 FILLER_57_3531 ();
 sg13g2_decap_8 FILLER_57_3538 ();
 sg13g2_decap_8 FILLER_57_3545 ();
 sg13g2_decap_8 FILLER_57_3552 ();
 sg13g2_decap_8 FILLER_57_3559 ();
 sg13g2_decap_8 FILLER_57_3566 ();
 sg13g2_decap_8 FILLER_57_3573 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_4 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_fill_2 FILLER_58_92 ();
 sg13g2_fill_2 FILLER_58_111 ();
 sg13g2_fill_1 FILLER_58_113 ();
 sg13g2_fill_2 FILLER_58_119 ();
 sg13g2_decap_4 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_174 ();
 sg13g2_fill_2 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_188 ();
 sg13g2_fill_1 FILLER_58_286 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_332 ();
 sg13g2_fill_1 FILLER_58_334 ();
 sg13g2_decap_8 FILLER_58_348 ();
 sg13g2_decap_4 FILLER_58_364 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_485 ();
 sg13g2_decap_8 FILLER_58_496 ();
 sg13g2_fill_2 FILLER_58_558 ();
 sg13g2_fill_1 FILLER_58_560 ();
 sg13g2_fill_2 FILLER_58_574 ();
 sg13g2_fill_1 FILLER_58_576 ();
 sg13g2_fill_2 FILLER_58_597 ();
 sg13g2_fill_1 FILLER_58_612 ();
 sg13g2_decap_8 FILLER_58_634 ();
 sg13g2_decap_4 FILLER_58_641 ();
 sg13g2_fill_1 FILLER_58_645 ();
 sg13g2_decap_8 FILLER_58_650 ();
 sg13g2_decap_8 FILLER_58_657 ();
 sg13g2_decap_8 FILLER_58_664 ();
 sg13g2_fill_2 FILLER_58_671 ();
 sg13g2_decap_4 FILLER_58_691 ();
 sg13g2_fill_1 FILLER_58_695 ();
 sg13g2_decap_8 FILLER_58_700 ();
 sg13g2_fill_2 FILLER_58_716 ();
 sg13g2_decap_8 FILLER_58_728 ();
 sg13g2_fill_1 FILLER_58_767 ();
 sg13g2_fill_1 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_813 ();
 sg13g2_fill_1 FILLER_58_824 ();
 sg13g2_fill_1 FILLER_58_838 ();
 sg13g2_decap_8 FILLER_58_843 ();
 sg13g2_decap_8 FILLER_58_850 ();
 sg13g2_fill_1 FILLER_58_885 ();
 sg13g2_fill_1 FILLER_58_890 ();
 sg13g2_fill_2 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_949 ();
 sg13g2_fill_1 FILLER_58_951 ();
 sg13g2_decap_8 FILLER_58_1029 ();
 sg13g2_fill_1 FILLER_58_1151 ();
 sg13g2_fill_2 FILLER_58_1198 ();
 sg13g2_fill_2 FILLER_58_1225 ();
 sg13g2_fill_1 FILLER_58_1260 ();
 sg13g2_decap_4 FILLER_58_1265 ();
 sg13g2_fill_2 FILLER_58_1286 ();
 sg13g2_fill_1 FILLER_58_1288 ();
 sg13g2_decap_8 FILLER_58_1297 ();
 sg13g2_decap_8 FILLER_58_1304 ();
 sg13g2_decap_4 FILLER_58_1329 ();
 sg13g2_fill_2 FILLER_58_1333 ();
 sg13g2_decap_8 FILLER_58_1356 ();
 sg13g2_decap_4 FILLER_58_1388 ();
 sg13g2_fill_2 FILLER_58_1414 ();
 sg13g2_fill_2 FILLER_58_1421 ();
 sg13g2_fill_1 FILLER_58_1423 ();
 sg13g2_fill_2 FILLER_58_1429 ();
 sg13g2_fill_1 FILLER_58_1431 ();
 sg13g2_decap_4 FILLER_58_1449 ();
 sg13g2_fill_1 FILLER_58_1453 ();
 sg13g2_fill_1 FILLER_58_1492 ();
 sg13g2_fill_2 FILLER_58_1497 ();
 sg13g2_decap_4 FILLER_58_1578 ();
 sg13g2_fill_2 FILLER_58_1582 ();
 sg13g2_decap_8 FILLER_58_1601 ();
 sg13g2_fill_1 FILLER_58_1608 ();
 sg13g2_decap_8 FILLER_58_1618 ();
 sg13g2_fill_1 FILLER_58_1625 ();
 sg13g2_decap_8 FILLER_58_1644 ();
 sg13g2_fill_1 FILLER_58_1651 ();
 sg13g2_decap_4 FILLER_58_1656 ();
 sg13g2_fill_2 FILLER_58_1660 ();
 sg13g2_decap_8 FILLER_58_1692 ();
 sg13g2_decap_4 FILLER_58_1699 ();
 sg13g2_fill_1 FILLER_58_1703 ();
 sg13g2_decap_4 FILLER_58_1722 ();
 sg13g2_fill_2 FILLER_58_1752 ();
 sg13g2_fill_1 FILLER_58_1784 ();
 sg13g2_decap_8 FILLER_58_1797 ();
 sg13g2_fill_2 FILLER_58_1804 ();
 sg13g2_fill_1 FILLER_58_1806 ();
 sg13g2_decap_4 FILLER_58_1815 ();
 sg13g2_fill_2 FILLER_58_1828 ();
 sg13g2_decap_4 FILLER_58_1895 ();
 sg13g2_fill_2 FILLER_58_1899 ();
 sg13g2_fill_2 FILLER_58_1938 ();
 sg13g2_fill_1 FILLER_58_1956 ();
 sg13g2_decap_8 FILLER_58_1997 ();
 sg13g2_fill_1 FILLER_58_2017 ();
 sg13g2_fill_2 FILLER_58_2073 ();
 sg13g2_fill_1 FILLER_58_2075 ();
 sg13g2_decap_4 FILLER_58_2089 ();
 sg13g2_fill_2 FILLER_58_2122 ();
 sg13g2_fill_1 FILLER_58_2124 ();
 sg13g2_fill_1 FILLER_58_2134 ();
 sg13g2_decap_4 FILLER_58_2157 ();
 sg13g2_fill_2 FILLER_58_2174 ();
 sg13g2_decap_8 FILLER_58_2204 ();
 sg13g2_fill_1 FILLER_58_2211 ();
 sg13g2_decap_8 FILLER_58_2219 ();
 sg13g2_fill_2 FILLER_58_2235 ();
 sg13g2_fill_2 FILLER_58_2255 ();
 sg13g2_fill_1 FILLER_58_2257 ();
 sg13g2_fill_1 FILLER_58_2304 ();
 sg13g2_decap_4 FILLER_58_2331 ();
 sg13g2_fill_1 FILLER_58_2335 ();
 sg13g2_decap_4 FILLER_58_2349 ();
 sg13g2_decap_4 FILLER_58_2385 ();
 sg13g2_fill_2 FILLER_58_2412 ();
 sg13g2_decap_4 FILLER_58_2419 ();
 sg13g2_fill_1 FILLER_58_2423 ();
 sg13g2_decap_8 FILLER_58_2428 ();
 sg13g2_decap_4 FILLER_58_2435 ();
 sg13g2_fill_2 FILLER_58_2452 ();
 sg13g2_fill_1 FILLER_58_2454 ();
 sg13g2_fill_2 FILLER_58_2464 ();
 sg13g2_fill_2 FILLER_58_2492 ();
 sg13g2_fill_1 FILLER_58_2494 ();
 sg13g2_decap_4 FILLER_58_2514 ();
 sg13g2_fill_2 FILLER_58_2527 ();
 sg13g2_fill_2 FILLER_58_2547 ();
 sg13g2_decap_8 FILLER_58_2562 ();
 sg13g2_fill_2 FILLER_58_2583 ();
 sg13g2_fill_2 FILLER_58_2613 ();
 sg13g2_decap_4 FILLER_58_2631 ();
 sg13g2_fill_1 FILLER_58_2635 ();
 sg13g2_decap_8 FILLER_58_2664 ();
 sg13g2_fill_2 FILLER_58_2671 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_decap_8 FILLER_58_2722 ();
 sg13g2_fill_1 FILLER_58_2742 ();
 sg13g2_decap_4 FILLER_58_2747 ();
 sg13g2_fill_1 FILLER_58_2751 ();
 sg13g2_decap_8 FILLER_58_2757 ();
 sg13g2_fill_2 FILLER_58_2764 ();
 sg13g2_fill_2 FILLER_58_2775 ();
 sg13g2_fill_1 FILLER_58_2777 ();
 sg13g2_fill_1 FILLER_58_2822 ();
 sg13g2_fill_2 FILLER_58_2850 ();
 sg13g2_fill_1 FILLER_58_2852 ();
 sg13g2_fill_2 FILLER_58_2893 ();
 sg13g2_fill_1 FILLER_58_2895 ();
 sg13g2_decap_4 FILLER_58_2951 ();
 sg13g2_fill_2 FILLER_58_2985 ();
 sg13g2_fill_2 FILLER_58_3014 ();
 sg13g2_fill_1 FILLER_58_3016 ();
 sg13g2_decap_8 FILLER_58_3026 ();
 sg13g2_fill_2 FILLER_58_3060 ();
 sg13g2_fill_1 FILLER_58_3062 ();
 sg13g2_fill_2 FILLER_58_3077 ();
 sg13g2_decap_4 FILLER_58_3097 ();
 sg13g2_decap_8 FILLER_58_3160 ();
 sg13g2_fill_1 FILLER_58_3167 ();
 sg13g2_decap_8 FILLER_58_3172 ();
 sg13g2_fill_2 FILLER_58_3179 ();
 sg13g2_decap_8 FILLER_58_3185 ();
 sg13g2_fill_1 FILLER_58_3192 ();
 sg13g2_decap_4 FILLER_58_3233 ();
 sg13g2_fill_1 FILLER_58_3246 ();
 sg13g2_decap_4 FILLER_58_3256 ();
 sg13g2_fill_2 FILLER_58_3260 ();
 sg13g2_fill_2 FILLER_58_3272 ();
 sg13g2_fill_2 FILLER_58_3277 ();
 sg13g2_fill_2 FILLER_58_3292 ();
 sg13g2_fill_2 FILLER_58_3298 ();
 sg13g2_fill_1 FILLER_58_3300 ();
 sg13g2_decap_8 FILLER_58_3310 ();
 sg13g2_decap_4 FILLER_58_3317 ();
 sg13g2_fill_1 FILLER_58_3321 ();
 sg13g2_decap_8 FILLER_58_3331 ();
 sg13g2_fill_2 FILLER_58_3402 ();
 sg13g2_decap_8 FILLER_58_3432 ();
 sg13g2_decap_8 FILLER_58_3439 ();
 sg13g2_decap_8 FILLER_58_3446 ();
 sg13g2_decap_8 FILLER_58_3453 ();
 sg13g2_decap_8 FILLER_58_3460 ();
 sg13g2_decap_8 FILLER_58_3467 ();
 sg13g2_decap_8 FILLER_58_3474 ();
 sg13g2_decap_8 FILLER_58_3481 ();
 sg13g2_decap_8 FILLER_58_3488 ();
 sg13g2_decap_8 FILLER_58_3495 ();
 sg13g2_decap_8 FILLER_58_3502 ();
 sg13g2_decap_8 FILLER_58_3509 ();
 sg13g2_decap_8 FILLER_58_3516 ();
 sg13g2_decap_8 FILLER_58_3523 ();
 sg13g2_decap_8 FILLER_58_3530 ();
 sg13g2_decap_8 FILLER_58_3537 ();
 sg13g2_decap_8 FILLER_58_3544 ();
 sg13g2_decap_8 FILLER_58_3551 ();
 sg13g2_decap_8 FILLER_58_3558 ();
 sg13g2_decap_8 FILLER_58_3565 ();
 sg13g2_decap_8 FILLER_58_3572 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_4 FILLER_59_63 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_fill_2 FILLER_59_97 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_114 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_fill_1 FILLER_59_182 ();
 sg13g2_fill_2 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_190 ();
 sg13g2_fill_1 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_decap_4 FILLER_59_230 ();
 sg13g2_fill_1 FILLER_59_234 ();
 sg13g2_decap_4 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_293 ();
 sg13g2_fill_1 FILLER_59_317 ();
 sg13g2_fill_2 FILLER_59_344 ();
 sg13g2_fill_1 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_362 ();
 sg13g2_fill_1 FILLER_59_376 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_402 ();
 sg13g2_fill_1 FILLER_59_404 ();
 sg13g2_decap_4 FILLER_59_440 ();
 sg13g2_fill_1 FILLER_59_444 ();
 sg13g2_fill_2 FILLER_59_509 ();
 sg13g2_fill_1 FILLER_59_529 ();
 sg13g2_decap_4 FILLER_59_535 ();
 sg13g2_fill_2 FILLER_59_539 ();
 sg13g2_fill_1 FILLER_59_550 ();
 sg13g2_decap_8 FILLER_59_555 ();
 sg13g2_decap_4 FILLER_59_562 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_fill_1 FILLER_59_581 ();
 sg13g2_fill_2 FILLER_59_613 ();
 sg13g2_fill_1 FILLER_59_615 ();
 sg13g2_fill_1 FILLER_59_620 ();
 sg13g2_decap_8 FILLER_59_626 ();
 sg13g2_fill_2 FILLER_59_633 ();
 sg13g2_fill_1 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_640 ();
 sg13g2_fill_2 FILLER_59_677 ();
 sg13g2_fill_2 FILLER_59_696 ();
 sg13g2_fill_1 FILLER_59_698 ();
 sg13g2_fill_2 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_714 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_fill_1 FILLER_59_735 ();
 sg13g2_decap_8 FILLER_59_847 ();
 sg13g2_fill_1 FILLER_59_854 ();
 sg13g2_decap_4 FILLER_59_872 ();
 sg13g2_decap_4 FILLER_59_889 ();
 sg13g2_fill_2 FILLER_59_893 ();
 sg13g2_decap_8 FILLER_59_908 ();
 sg13g2_fill_2 FILLER_59_915 ();
 sg13g2_decap_8 FILLER_59_921 ();
 sg13g2_decap_4 FILLER_59_928 ();
 sg13g2_fill_1 FILLER_59_997 ();
 sg13g2_decap_4 FILLER_59_1007 ();
 sg13g2_fill_1 FILLER_59_1056 ();
 sg13g2_fill_2 FILLER_59_1083 ();
 sg13g2_decap_4 FILLER_59_1089 ();
 sg13g2_decap_8 FILLER_59_1107 ();
 sg13g2_fill_2 FILLER_59_1118 ();
 sg13g2_fill_1 FILLER_59_1120 ();
 sg13g2_fill_1 FILLER_59_1140 ();
 sg13g2_decap_4 FILLER_59_1154 ();
 sg13g2_fill_1 FILLER_59_1158 ();
 sg13g2_fill_1 FILLER_59_1184 ();
 sg13g2_fill_1 FILLER_59_1190 ();
 sg13g2_fill_2 FILLER_59_1196 ();
 sg13g2_fill_1 FILLER_59_1198 ();
 sg13g2_fill_2 FILLER_59_1212 ();
 sg13g2_decap_4 FILLER_59_1233 ();
 sg13g2_fill_2 FILLER_59_1237 ();
 sg13g2_decap_4 FILLER_59_1284 ();
 sg13g2_fill_1 FILLER_59_1288 ();
 sg13g2_fill_2 FILLER_59_1307 ();
 sg13g2_decap_8 FILLER_59_1320 ();
 sg13g2_decap_8 FILLER_59_1327 ();
 sg13g2_decap_8 FILLER_59_1352 ();
 sg13g2_fill_2 FILLER_59_1359 ();
 sg13g2_fill_1 FILLER_59_1361 ();
 sg13g2_fill_2 FILLER_59_1384 ();
 sg13g2_fill_2 FILLER_59_1420 ();
 sg13g2_fill_1 FILLER_59_1422 ();
 sg13g2_decap_8 FILLER_59_1434 ();
 sg13g2_decap_8 FILLER_59_1441 ();
 sg13g2_decap_4 FILLER_59_1448 ();
 sg13g2_decap_8 FILLER_59_1466 ();
 sg13g2_decap_4 FILLER_59_1473 ();
 sg13g2_fill_1 FILLER_59_1477 ();
 sg13g2_fill_2 FILLER_59_1491 ();
 sg13g2_fill_1 FILLER_59_1493 ();
 sg13g2_fill_2 FILLER_59_1511 ();
 sg13g2_fill_2 FILLER_59_1526 ();
 sg13g2_fill_1 FILLER_59_1528 ();
 sg13g2_fill_1 FILLER_59_1539 ();
 sg13g2_decap_4 FILLER_59_1582 ();
 sg13g2_fill_1 FILLER_59_1586 ();
 sg13g2_decap_8 FILLER_59_1618 ();
 sg13g2_fill_2 FILLER_59_1625 ();
 sg13g2_fill_2 FILLER_59_1650 ();
 sg13g2_fill_1 FILLER_59_1652 ();
 sg13g2_decap_8 FILLER_59_1689 ();
 sg13g2_fill_2 FILLER_59_1696 ();
 sg13g2_fill_1 FILLER_59_1698 ();
 sg13g2_decap_4 FILLER_59_1717 ();
 sg13g2_decap_8 FILLER_59_1744 ();
 sg13g2_decap_8 FILLER_59_1751 ();
 sg13g2_decap_4 FILLER_59_1770 ();
 sg13g2_decap_4 FILLER_59_1802 ();
 sg13g2_fill_1 FILLER_59_1814 ();
 sg13g2_fill_2 FILLER_59_1828 ();
 sg13g2_fill_2 FILLER_59_1846 ();
 sg13g2_fill_1 FILLER_59_1848 ();
 sg13g2_fill_2 FILLER_59_1867 ();
 sg13g2_fill_1 FILLER_59_1869 ();
 sg13g2_fill_2 FILLER_59_1892 ();
 sg13g2_fill_1 FILLER_59_1894 ();
 sg13g2_fill_2 FILLER_59_1914 ();
 sg13g2_fill_1 FILLER_59_1970 ();
 sg13g2_fill_1 FILLER_59_2018 ();
 sg13g2_fill_2 FILLER_59_2042 ();
 sg13g2_fill_1 FILLER_59_2062 ();
 sg13g2_fill_2 FILLER_59_2076 ();
 sg13g2_fill_1 FILLER_59_2078 ();
 sg13g2_fill_2 FILLER_59_2116 ();
 sg13g2_fill_1 FILLER_59_2118 ();
 sg13g2_fill_2 FILLER_59_2161 ();
 sg13g2_fill_1 FILLER_59_2163 ();
 sg13g2_fill_2 FILLER_59_2178 ();
 sg13g2_fill_1 FILLER_59_2189 ();
 sg13g2_fill_1 FILLER_59_2195 ();
 sg13g2_decap_8 FILLER_59_2201 ();
 sg13g2_fill_1 FILLER_59_2216 ();
 sg13g2_fill_2 FILLER_59_2229 ();
 sg13g2_fill_2 FILLER_59_2279 ();
 sg13g2_fill_1 FILLER_59_2281 ();
 sg13g2_decap_8 FILLER_59_2291 ();
 sg13g2_decap_4 FILLER_59_2316 ();
 sg13g2_decap_4 FILLER_59_2347 ();
 sg13g2_fill_2 FILLER_59_2356 ();
 sg13g2_fill_1 FILLER_59_2358 ();
 sg13g2_fill_2 FILLER_59_2396 ();
 sg13g2_fill_2 FILLER_59_2411 ();
 sg13g2_fill_1 FILLER_59_2413 ();
 sg13g2_decap_4 FILLER_59_2431 ();
 sg13g2_fill_2 FILLER_59_2468 ();
 sg13g2_fill_2 FILLER_59_2498 ();
 sg13g2_fill_2 FILLER_59_2541 ();
 sg13g2_fill_1 FILLER_59_2543 ();
 sg13g2_fill_1 FILLER_59_2595 ();
 sg13g2_fill_2 FILLER_59_2616 ();
 sg13g2_fill_1 FILLER_59_2618 ();
 sg13g2_decap_4 FILLER_59_2665 ();
 sg13g2_fill_1 FILLER_59_2687 ();
 sg13g2_fill_2 FILLER_59_2693 ();
 sg13g2_fill_2 FILLER_59_2699 ();
 sg13g2_fill_1 FILLER_59_2701 ();
 sg13g2_decap_4 FILLER_59_2707 ();
 sg13g2_fill_1 FILLER_59_2711 ();
 sg13g2_decap_4 FILLER_59_2717 ();
 sg13g2_fill_2 FILLER_59_2721 ();
 sg13g2_fill_2 FILLER_59_2736 ();
 sg13g2_decap_8 FILLER_59_2765 ();
 sg13g2_decap_4 FILLER_59_2772 ();
 sg13g2_fill_1 FILLER_59_2776 ();
 sg13g2_decap_4 FILLER_59_2790 ();
 sg13g2_fill_1 FILLER_59_2825 ();
 sg13g2_fill_2 FILLER_59_2856 ();
 sg13g2_decap_8 FILLER_59_2863 ();
 sg13g2_decap_8 FILLER_59_2870 ();
 sg13g2_decap_8 FILLER_59_2877 ();
 sg13g2_fill_1 FILLER_59_2898 ();
 sg13g2_decap_8 FILLER_59_2913 ();
 sg13g2_fill_2 FILLER_59_2920 ();
 sg13g2_fill_1 FILLER_59_2922 ();
 sg13g2_decap_4 FILLER_59_2936 ();
 sg13g2_fill_2 FILLER_59_2940 ();
 sg13g2_decap_8 FILLER_59_2974 ();
 sg13g2_fill_1 FILLER_59_2981 ();
 sg13g2_fill_2 FILLER_59_2985 ();
 sg13g2_decap_4 FILLER_59_2996 ();
 sg13g2_fill_1 FILLER_59_3000 ();
 sg13g2_decap_8 FILLER_59_3050 ();
 sg13g2_fill_2 FILLER_59_3057 ();
 sg13g2_decap_4 FILLER_59_3067 ();
 sg13g2_fill_1 FILLER_59_3071 ();
 sg13g2_fill_2 FILLER_59_3077 ();
 sg13g2_fill_1 FILLER_59_3079 ();
 sg13g2_decap_4 FILLER_59_3106 ();
 sg13g2_fill_2 FILLER_59_3110 ();
 sg13g2_fill_1 FILLER_59_3125 ();
 sg13g2_decap_4 FILLER_59_3204 ();
 sg13g2_fill_2 FILLER_59_3208 ();
 sg13g2_decap_4 FILLER_59_3243 ();
 sg13g2_fill_2 FILLER_59_3247 ();
 sg13g2_fill_1 FILLER_59_3253 ();
 sg13g2_decap_8 FILLER_59_3281 ();
 sg13g2_fill_1 FILLER_59_3288 ();
 sg13g2_fill_1 FILLER_59_3302 ();
 sg13g2_decap_4 FILLER_59_3326 ();
 sg13g2_fill_1 FILLER_59_3330 ();
 sg13g2_fill_1 FILLER_59_3348 ();
 sg13g2_decap_8 FILLER_59_3375 ();
 sg13g2_fill_1 FILLER_59_3382 ();
 sg13g2_decap_8 FILLER_59_3411 ();
 sg13g2_decap_8 FILLER_59_3418 ();
 sg13g2_decap_8 FILLER_59_3425 ();
 sg13g2_decap_8 FILLER_59_3432 ();
 sg13g2_decap_8 FILLER_59_3439 ();
 sg13g2_decap_8 FILLER_59_3446 ();
 sg13g2_decap_8 FILLER_59_3453 ();
 sg13g2_decap_8 FILLER_59_3460 ();
 sg13g2_decap_8 FILLER_59_3467 ();
 sg13g2_decap_8 FILLER_59_3474 ();
 sg13g2_decap_8 FILLER_59_3481 ();
 sg13g2_decap_8 FILLER_59_3488 ();
 sg13g2_decap_8 FILLER_59_3495 ();
 sg13g2_decap_8 FILLER_59_3502 ();
 sg13g2_decap_8 FILLER_59_3509 ();
 sg13g2_decap_8 FILLER_59_3516 ();
 sg13g2_decap_8 FILLER_59_3523 ();
 sg13g2_decap_8 FILLER_59_3530 ();
 sg13g2_decap_8 FILLER_59_3537 ();
 sg13g2_decap_8 FILLER_59_3544 ();
 sg13g2_decap_8 FILLER_59_3551 ();
 sg13g2_decap_8 FILLER_59_3558 ();
 sg13g2_decap_8 FILLER_59_3565 ();
 sg13g2_decap_8 FILLER_59_3572 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_fill_2 FILLER_60_126 ();
 sg13g2_decap_4 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_decap_4 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_174 ();
 sg13g2_decap_8 FILLER_60_181 ();
 sg13g2_fill_2 FILLER_60_188 ();
 sg13g2_fill_2 FILLER_60_259 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_fill_2 FILLER_60_324 ();
 sg13g2_fill_1 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_decap_4 FILLER_60_445 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_fill_2 FILLER_60_471 ();
 sg13g2_fill_2 FILLER_60_562 ();
 sg13g2_fill_2 FILLER_60_592 ();
 sg13g2_fill_1 FILLER_60_603 ();
 sg13g2_fill_1 FILLER_60_630 ();
 sg13g2_decap_4 FILLER_60_658 ();
 sg13g2_fill_2 FILLER_60_662 ();
 sg13g2_decap_8 FILLER_60_695 ();
 sg13g2_decap_8 FILLER_60_702 ();
 sg13g2_fill_2 FILLER_60_709 ();
 sg13g2_fill_2 FILLER_60_720 ();
 sg13g2_fill_2 FILLER_60_727 ();
 sg13g2_fill_1 FILLER_60_737 ();
 sg13g2_fill_2 FILLER_60_741 ();
 sg13g2_fill_1 FILLER_60_743 ();
 sg13g2_decap_4 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_60_770 ();
 sg13g2_decap_8 FILLER_60_777 ();
 sg13g2_decap_4 FILLER_60_787 ();
 sg13g2_fill_2 FILLER_60_791 ();
 sg13g2_fill_1 FILLER_60_819 ();
 sg13g2_fill_1 FILLER_60_864 ();
 sg13g2_fill_2 FILLER_60_870 ();
 sg13g2_fill_1 FILLER_60_872 ();
 sg13g2_decap_4 FILLER_60_901 ();
 sg13g2_decap_4 FILLER_60_931 ();
 sg13g2_fill_2 FILLER_60_948 ();
 sg13g2_decap_8 FILLER_60_979 ();
 sg13g2_fill_1 FILLER_60_986 ();
 sg13g2_fill_1 FILLER_60_1015 ();
 sg13g2_fill_2 FILLER_60_1025 ();
 sg13g2_fill_1 FILLER_60_1027 ();
 sg13g2_fill_1 FILLER_60_1065 ();
 sg13g2_fill_2 FILLER_60_1143 ();
 sg13g2_fill_1 FILLER_60_1145 ();
 sg13g2_fill_1 FILLER_60_1172 ();
 sg13g2_fill_2 FILLER_60_1238 ();
 sg13g2_fill_1 FILLER_60_1240 ();
 sg13g2_decap_4 FILLER_60_1266 ();
 sg13g2_fill_1 FILLER_60_1301 ();
 sg13g2_decap_8 FILLER_60_1320 ();
 sg13g2_fill_2 FILLER_60_1399 ();
 sg13g2_fill_1 FILLER_60_1401 ();
 sg13g2_decap_4 FILLER_60_1413 ();
 sg13g2_fill_1 FILLER_60_1440 ();
 sg13g2_decap_8 FILLER_60_1466 ();
 sg13g2_fill_2 FILLER_60_1473 ();
 sg13g2_fill_1 FILLER_60_1514 ();
 sg13g2_fill_1 FILLER_60_1560 ();
 sg13g2_fill_2 FILLER_60_1596 ();
 sg13g2_decap_8 FILLER_60_1616 ();
 sg13g2_decap_4 FILLER_60_1623 ();
 sg13g2_fill_2 FILLER_60_1653 ();
 sg13g2_fill_1 FILLER_60_1655 ();
 sg13g2_decap_4 FILLER_60_1670 ();
 sg13g2_fill_1 FILLER_60_1674 ();
 sg13g2_decap_8 FILLER_60_1694 ();
 sg13g2_fill_2 FILLER_60_1701 ();
 sg13g2_fill_1 FILLER_60_1703 ();
 sg13g2_decap_8 FILLER_60_1709 ();
 sg13g2_decap_8 FILLER_60_1716 ();
 sg13g2_fill_2 FILLER_60_1723 ();
 sg13g2_fill_1 FILLER_60_1725 ();
 sg13g2_decap_8 FILLER_60_1736 ();
 sg13g2_fill_1 FILLER_60_1760 ();
 sg13g2_decap_8 FILLER_60_1769 ();
 sg13g2_fill_2 FILLER_60_1776 ();
 sg13g2_fill_1 FILLER_60_1778 ();
 sg13g2_decap_4 FILLER_60_1785 ();
 sg13g2_decap_8 FILLER_60_1799 ();
 sg13g2_fill_2 FILLER_60_1806 ();
 sg13g2_fill_1 FILLER_60_1808 ();
 sg13g2_fill_2 FILLER_60_1818 ();
 sg13g2_fill_1 FILLER_60_1820 ();
 sg13g2_fill_1 FILLER_60_1838 ();
 sg13g2_fill_2 FILLER_60_1845 ();
 sg13g2_fill_2 FILLER_60_1875 ();
 sg13g2_fill_1 FILLER_60_1877 ();
 sg13g2_fill_1 FILLER_60_1900 ();
 sg13g2_decap_8 FILLER_60_1910 ();
 sg13g2_fill_2 FILLER_60_1917 ();
 sg13g2_decap_4 FILLER_60_1945 ();
 sg13g2_fill_2 FILLER_60_1949 ();
 sg13g2_fill_1 FILLER_60_1984 ();
 sg13g2_fill_2 FILLER_60_1997 ();
 sg13g2_fill_1 FILLER_60_1999 ();
 sg13g2_decap_8 FILLER_60_2045 ();
 sg13g2_decap_8 FILLER_60_2052 ();
 sg13g2_fill_2 FILLER_60_2064 ();
 sg13g2_fill_1 FILLER_60_2105 ();
 sg13g2_fill_2 FILLER_60_2133 ();
 sg13g2_fill_2 FILLER_60_2190 ();
 sg13g2_fill_1 FILLER_60_2192 ();
 sg13g2_decap_8 FILLER_60_2206 ();
 sg13g2_fill_2 FILLER_60_2213 ();
 sg13g2_fill_2 FILLER_60_2220 ();
 sg13g2_fill_1 FILLER_60_2243 ();
 sg13g2_fill_1 FILLER_60_2315 ();
 sg13g2_decap_4 FILLER_60_2320 ();
 sg13g2_fill_1 FILLER_60_2324 ();
 sg13g2_decap_8 FILLER_60_2351 ();
 sg13g2_decap_4 FILLER_60_2358 ();
 sg13g2_fill_2 FILLER_60_2362 ();
 sg13g2_decap_8 FILLER_60_2400 ();
 sg13g2_decap_8 FILLER_60_2457 ();
 sg13g2_fill_2 FILLER_60_2464 ();
 sg13g2_fill_1 FILLER_60_2492 ();
 sg13g2_fill_2 FILLER_60_2515 ();
 sg13g2_fill_1 FILLER_60_2517 ();
 sg13g2_fill_2 FILLER_60_2541 ();
 sg13g2_decap_8 FILLER_60_2547 ();
 sg13g2_fill_2 FILLER_60_2554 ();
 sg13g2_decap_4 FILLER_60_2592 ();
 sg13g2_fill_2 FILLER_60_2596 ();
 sg13g2_fill_2 FILLER_60_2611 ();
 sg13g2_fill_1 FILLER_60_2619 ();
 sg13g2_decap_4 FILLER_60_2629 ();
 sg13g2_fill_1 FILLER_60_2633 ();
 sg13g2_decap_4 FILLER_60_2639 ();
 sg13g2_fill_1 FILLER_60_2682 ();
 sg13g2_fill_1 FILLER_60_2705 ();
 sg13g2_fill_2 FILLER_60_2724 ();
 sg13g2_fill_1 FILLER_60_2726 ();
 sg13g2_fill_2 FILLER_60_2743 ();
 sg13g2_fill_2 FILLER_60_2773 ();
 sg13g2_fill_2 FILLER_60_2802 ();
 sg13g2_fill_1 FILLER_60_2817 ();
 sg13g2_fill_1 FILLER_60_2827 ();
 sg13g2_fill_2 FILLER_60_2931 ();
 sg13g2_fill_1 FILLER_60_2933 ();
 sg13g2_fill_2 FILLER_60_2939 ();
 sg13g2_fill_1 FILLER_60_2941 ();
 sg13g2_decap_8 FILLER_60_2952 ();
 sg13g2_fill_2 FILLER_60_2959 ();
 sg13g2_decap_8 FILLER_60_2965 ();
 sg13g2_fill_1 FILLER_60_2972 ();
 sg13g2_decap_4 FILLER_60_2995 ();
 sg13g2_fill_2 FILLER_60_2999 ();
 sg13g2_decap_8 FILLER_60_3019 ();
 sg13g2_decap_8 FILLER_60_3026 ();
 sg13g2_fill_2 FILLER_60_3038 ();
 sg13g2_decap_8 FILLER_60_3044 ();
 sg13g2_fill_2 FILLER_60_3051 ();
 sg13g2_fill_1 FILLER_60_3067 ();
 sg13g2_fill_2 FILLER_60_3078 ();
 sg13g2_fill_1 FILLER_60_3080 ();
 sg13g2_fill_2 FILLER_60_3094 ();
 sg13g2_fill_1 FILLER_60_3177 ();
 sg13g2_fill_2 FILLER_60_3204 ();
 sg13g2_fill_2 FILLER_60_3219 ();
 sg13g2_fill_1 FILLER_60_3221 ();
 sg13g2_fill_2 FILLER_60_3272 ();
 sg13g2_fill_1 FILLER_60_3274 ();
 sg13g2_decap_8 FILLER_60_3297 ();
 sg13g2_decap_8 FILLER_60_3304 ();
 sg13g2_fill_2 FILLER_60_3311 ();
 sg13g2_fill_1 FILLER_60_3313 ();
 sg13g2_fill_2 FILLER_60_3324 ();
 sg13g2_fill_1 FILLER_60_3326 ();
 sg13g2_decap_8 FILLER_60_3355 ();
 sg13g2_fill_1 FILLER_60_3362 ();
 sg13g2_fill_2 FILLER_60_3368 ();
 sg13g2_fill_1 FILLER_60_3370 ();
 sg13g2_decap_8 FILLER_60_3375 ();
 sg13g2_fill_1 FILLER_60_3382 ();
 sg13g2_decap_4 FILLER_60_3396 ();
 sg13g2_decap_8 FILLER_60_3409 ();
 sg13g2_decap_8 FILLER_60_3416 ();
 sg13g2_decap_8 FILLER_60_3423 ();
 sg13g2_decap_8 FILLER_60_3430 ();
 sg13g2_decap_8 FILLER_60_3437 ();
 sg13g2_decap_8 FILLER_60_3444 ();
 sg13g2_decap_8 FILLER_60_3451 ();
 sg13g2_decap_8 FILLER_60_3458 ();
 sg13g2_decap_8 FILLER_60_3465 ();
 sg13g2_decap_8 FILLER_60_3472 ();
 sg13g2_decap_8 FILLER_60_3479 ();
 sg13g2_decap_8 FILLER_60_3486 ();
 sg13g2_decap_8 FILLER_60_3493 ();
 sg13g2_decap_8 FILLER_60_3500 ();
 sg13g2_decap_8 FILLER_60_3507 ();
 sg13g2_decap_8 FILLER_60_3514 ();
 sg13g2_decap_8 FILLER_60_3521 ();
 sg13g2_decap_8 FILLER_60_3528 ();
 sg13g2_decap_8 FILLER_60_3535 ();
 sg13g2_decap_8 FILLER_60_3542 ();
 sg13g2_decap_8 FILLER_60_3549 ();
 sg13g2_decap_8 FILLER_60_3556 ();
 sg13g2_decap_8 FILLER_60_3563 ();
 sg13g2_decap_8 FILLER_60_3570 ();
 sg13g2_fill_2 FILLER_60_3577 ();
 sg13g2_fill_1 FILLER_60_3579 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_88 ();
 sg13g2_fill_2 FILLER_61_95 ();
 sg13g2_fill_1 FILLER_61_97 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_decap_8 FILLER_61_173 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_fill_2 FILLER_61_204 ();
 sg13g2_fill_1 FILLER_61_206 ();
 sg13g2_fill_2 FILLER_61_216 ();
 sg13g2_decap_8 FILLER_61_237 ();
 sg13g2_fill_1 FILLER_61_244 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_275 ();
 sg13g2_fill_2 FILLER_61_318 ();
 sg13g2_fill_2 FILLER_61_347 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_fill_2 FILLER_61_370 ();
 sg13g2_decap_4 FILLER_61_392 ();
 sg13g2_fill_1 FILLER_61_495 ();
 sg13g2_fill_1 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_620 ();
 sg13g2_decap_4 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_631 ();
 sg13g2_decap_4 FILLER_61_645 ();
 sg13g2_fill_2 FILLER_61_649 ();
 sg13g2_decap_4 FILLER_61_702 ();
 sg13g2_fill_2 FILLER_61_744 ();
 sg13g2_decap_8 FILLER_61_771 ();
 sg13g2_decap_8 FILLER_61_778 ();
 sg13g2_fill_1 FILLER_61_785 ();
 sg13g2_fill_2 FILLER_61_813 ();
 sg13g2_fill_1 FILLER_61_815 ();
 sg13g2_fill_2 FILLER_61_852 ();
 sg13g2_fill_1 FILLER_61_854 ();
 sg13g2_fill_2 FILLER_61_864 ();
 sg13g2_fill_1 FILLER_61_871 ();
 sg13g2_fill_2 FILLER_61_900 ();
 sg13g2_decap_4 FILLER_61_943 ();
 sg13g2_fill_1 FILLER_61_947 ();
 sg13g2_fill_1 FILLER_61_961 ();
 sg13g2_fill_1 FILLER_61_975 ();
 sg13g2_decap_4 FILLER_61_984 ();
 sg13g2_fill_2 FILLER_61_996 ();
 sg13g2_decap_4 FILLER_61_1002 ();
 sg13g2_fill_1 FILLER_61_1006 ();
 sg13g2_decap_4 FILLER_61_1034 ();
 sg13g2_fill_2 FILLER_61_1038 ();
 sg13g2_fill_2 FILLER_61_1044 ();
 sg13g2_fill_1 FILLER_61_1046 ();
 sg13g2_fill_2 FILLER_61_1092 ();
 sg13g2_fill_1 FILLER_61_1098 ();
 sg13g2_decap_8 FILLER_61_1104 ();
 sg13g2_fill_2 FILLER_61_1111 ();
 sg13g2_fill_1 FILLER_61_1113 ();
 sg13g2_fill_2 FILLER_61_1127 ();
 sg13g2_fill_1 FILLER_61_1129 ();
 sg13g2_fill_2 FILLER_61_1157 ();
 sg13g2_fill_1 FILLER_61_1159 ();
 sg13g2_fill_2 FILLER_61_1173 ();
 sg13g2_fill_2 FILLER_61_1185 ();
 sg13g2_fill_1 FILLER_61_1192 ();
 sg13g2_decap_8 FILLER_61_1205 ();
 sg13g2_decap_8 FILLER_61_1216 ();
 sg13g2_decap_4 FILLER_61_1223 ();
 sg13g2_fill_2 FILLER_61_1232 ();
 sg13g2_decap_4 FILLER_61_1239 ();
 sg13g2_fill_2 FILLER_61_1306 ();
 sg13g2_decap_8 FILLER_61_1336 ();
 sg13g2_decap_4 FILLER_61_1356 ();
 sg13g2_fill_2 FILLER_61_1386 ();
 sg13g2_fill_1 FILLER_61_1388 ();
 sg13g2_fill_2 FILLER_61_1394 ();
 sg13g2_decap_8 FILLER_61_1410 ();
 sg13g2_decap_4 FILLER_61_1417 ();
 sg13g2_fill_1 FILLER_61_1421 ();
 sg13g2_fill_2 FILLER_61_1439 ();
 sg13g2_decap_8 FILLER_61_1459 ();
 sg13g2_fill_2 FILLER_61_1466 ();
 sg13g2_fill_2 FILLER_61_1516 ();
 sg13g2_fill_1 FILLER_61_1518 ();
 sg13g2_fill_2 FILLER_61_1532 ();
 sg13g2_fill_1 FILLER_61_1543 ();
 sg13g2_fill_1 FILLER_61_1556 ();
 sg13g2_fill_1 FILLER_61_1594 ();
 sg13g2_fill_1 FILLER_61_1632 ();
 sg13g2_decap_4 FILLER_61_1643 ();
 sg13g2_fill_2 FILLER_61_1721 ();
 sg13g2_fill_1 FILLER_61_1723 ();
 sg13g2_fill_2 FILLER_61_1752 ();
 sg13g2_fill_2 FILLER_61_1787 ();
 sg13g2_fill_1 FILLER_61_1789 ();
 sg13g2_decap_8 FILLER_61_1848 ();
 sg13g2_decap_4 FILLER_61_1855 ();
 sg13g2_fill_1 FILLER_61_1859 ();
 sg13g2_fill_2 FILLER_61_1873 ();
 sg13g2_fill_2 FILLER_61_1926 ();
 sg13g2_fill_1 FILLER_61_1928 ();
 sg13g2_fill_1 FILLER_61_1970 ();
 sg13g2_fill_1 FILLER_61_1989 ();
 sg13g2_decap_4 FILLER_61_2016 ();
 sg13g2_fill_1 FILLER_61_2033 ();
 sg13g2_fill_2 FILLER_61_2062 ();
 sg13g2_fill_1 FILLER_61_2064 ();
 sg13g2_fill_2 FILLER_61_2106 ();
 sg13g2_fill_1 FILLER_61_2108 ();
 sg13g2_fill_2 FILLER_61_2118 ();
 sg13g2_fill_1 FILLER_61_2120 ();
 sg13g2_decap_8 FILLER_61_2138 ();
 sg13g2_decap_4 FILLER_61_2145 ();
 sg13g2_decap_4 FILLER_61_2153 ();
 sg13g2_fill_2 FILLER_61_2157 ();
 sg13g2_decap_8 FILLER_61_2163 ();
 sg13g2_decap_8 FILLER_61_2170 ();
 sg13g2_decap_4 FILLER_61_2177 ();
 sg13g2_fill_1 FILLER_61_2185 ();
 sg13g2_fill_2 FILLER_61_2199 ();
 sg13g2_fill_1 FILLER_61_2201 ();
 sg13g2_fill_2 FILLER_61_2224 ();
 sg13g2_fill_1 FILLER_61_2226 ();
 sg13g2_decap_4 FILLER_61_2236 ();
 sg13g2_fill_2 FILLER_61_2240 ();
 sg13g2_fill_2 FILLER_61_2258 ();
 sg13g2_fill_2 FILLER_61_2269 ();
 sg13g2_fill_2 FILLER_61_2284 ();
 sg13g2_fill_1 FILLER_61_2286 ();
 sg13g2_decap_4 FILLER_61_2296 ();
 sg13g2_fill_1 FILLER_61_2305 ();
 sg13g2_fill_2 FILLER_61_2374 ();
 sg13g2_fill_1 FILLER_61_2376 ();
 sg13g2_fill_2 FILLER_61_2409 ();
 sg13g2_fill_1 FILLER_61_2411 ();
 sg13g2_fill_1 FILLER_61_2425 ();
 sg13g2_fill_2 FILLER_61_2435 ();
 sg13g2_fill_1 FILLER_61_2437 ();
 sg13g2_decap_8 FILLER_61_2451 ();
 sg13g2_fill_1 FILLER_61_2499 ();
 sg13g2_fill_1 FILLER_61_2509 ();
 sg13g2_fill_2 FILLER_61_2581 ();
 sg13g2_decap_4 FILLER_61_2591 ();
 sg13g2_fill_2 FILLER_61_2595 ();
 sg13g2_fill_1 FILLER_61_2610 ();
 sg13g2_decap_4 FILLER_61_2621 ();
 sg13g2_decap_8 FILLER_61_2640 ();
 sg13g2_decap_8 FILLER_61_2647 ();
 sg13g2_decap_8 FILLER_61_2676 ();
 sg13g2_decap_8 FILLER_61_2683 ();
 sg13g2_fill_2 FILLER_61_2690 ();
 sg13g2_decap_8 FILLER_61_2713 ();
 sg13g2_decap_4 FILLER_61_2720 ();
 sg13g2_fill_1 FILLER_61_2737 ();
 sg13g2_fill_2 FILLER_61_2746 ();
 sg13g2_fill_1 FILLER_61_2748 ();
 sg13g2_decap_4 FILLER_61_2762 ();
 sg13g2_fill_2 FILLER_61_2766 ();
 sg13g2_fill_1 FILLER_61_2774 ();
 sg13g2_fill_1 FILLER_61_2806 ();
 sg13g2_fill_2 FILLER_61_2829 ();
 sg13g2_fill_2 FILLER_61_2835 ();
 sg13g2_fill_1 FILLER_61_2837 ();
 sg13g2_decap_8 FILLER_61_2842 ();
 sg13g2_decap_8 FILLER_61_2849 ();
 sg13g2_decap_4 FILLER_61_2856 ();
 sg13g2_fill_1 FILLER_61_2860 ();
 sg13g2_fill_2 FILLER_61_2865 ();
 sg13g2_fill_2 FILLER_61_2871 ();
 sg13g2_fill_1 FILLER_61_2895 ();
 sg13g2_fill_2 FILLER_61_2909 ();
 sg13g2_decap_8 FILLER_61_2920 ();
 sg13g2_fill_2 FILLER_61_2927 ();
 sg13g2_fill_1 FILLER_61_2929 ();
 sg13g2_fill_1 FILLER_61_2942 ();
 sg13g2_fill_1 FILLER_61_2985 ();
 sg13g2_fill_2 FILLER_61_2991 ();
 sg13g2_fill_1 FILLER_61_2993 ();
 sg13g2_fill_1 FILLER_61_3007 ();
 sg13g2_decap_8 FILLER_61_3018 ();
 sg13g2_decap_4 FILLER_61_3025 ();
 sg13g2_fill_2 FILLER_61_3029 ();
 sg13g2_decap_8 FILLER_61_3064 ();
 sg13g2_fill_2 FILLER_61_3071 ();
 sg13g2_fill_2 FILLER_61_3086 ();
 sg13g2_fill_2 FILLER_61_3116 ();
 sg13g2_fill_1 FILLER_61_3148 ();
 sg13g2_fill_1 FILLER_61_3208 ();
 sg13g2_fill_1 FILLER_61_3217 ();
 sg13g2_fill_1 FILLER_61_3224 ();
 sg13g2_decap_8 FILLER_61_3249 ();
 sg13g2_fill_2 FILLER_61_3256 ();
 sg13g2_fill_1 FILLER_61_3258 ();
 sg13g2_decap_8 FILLER_61_3267 ();
 sg13g2_decap_4 FILLER_61_3274 ();
 sg13g2_fill_2 FILLER_61_3278 ();
 sg13g2_decap_4 FILLER_61_3284 ();
 sg13g2_fill_1 FILLER_61_3288 ();
 sg13g2_fill_2 FILLER_61_3298 ();
 sg13g2_fill_1 FILLER_61_3300 ();
 sg13g2_fill_2 FILLER_61_3305 ();
 sg13g2_fill_1 FILLER_61_3307 ();
 sg13g2_decap_8 FILLER_61_3331 ();
 sg13g2_fill_2 FILLER_61_3338 ();
 sg13g2_fill_2 FILLER_61_3363 ();
 sg13g2_fill_1 FILLER_61_3365 ();
 sg13g2_decap_8 FILLER_61_3394 ();
 sg13g2_decap_8 FILLER_61_3401 ();
 sg13g2_decap_8 FILLER_61_3408 ();
 sg13g2_decap_8 FILLER_61_3415 ();
 sg13g2_decap_8 FILLER_61_3422 ();
 sg13g2_decap_8 FILLER_61_3429 ();
 sg13g2_decap_8 FILLER_61_3436 ();
 sg13g2_decap_8 FILLER_61_3443 ();
 sg13g2_decap_8 FILLER_61_3450 ();
 sg13g2_decap_8 FILLER_61_3457 ();
 sg13g2_decap_8 FILLER_61_3464 ();
 sg13g2_decap_8 FILLER_61_3471 ();
 sg13g2_decap_8 FILLER_61_3478 ();
 sg13g2_decap_8 FILLER_61_3485 ();
 sg13g2_decap_8 FILLER_61_3492 ();
 sg13g2_decap_8 FILLER_61_3499 ();
 sg13g2_decap_8 FILLER_61_3506 ();
 sg13g2_decap_8 FILLER_61_3513 ();
 sg13g2_decap_8 FILLER_61_3520 ();
 sg13g2_decap_8 FILLER_61_3527 ();
 sg13g2_decap_8 FILLER_61_3534 ();
 sg13g2_decap_8 FILLER_61_3541 ();
 sg13g2_decap_8 FILLER_61_3548 ();
 sg13g2_decap_8 FILLER_61_3555 ();
 sg13g2_decap_8 FILLER_61_3562 ();
 sg13g2_decap_8 FILLER_61_3569 ();
 sg13g2_decap_4 FILLER_61_3576 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_131 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_decap_4 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_173 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_189 ();
 sg13g2_fill_2 FILLER_62_194 ();
 sg13g2_fill_2 FILLER_62_223 ();
 sg13g2_decap_4 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_283 ();
 sg13g2_decap_4 FILLER_62_304 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_decap_4 FILLER_62_396 ();
 sg13g2_decap_4 FILLER_62_408 ();
 sg13g2_fill_1 FILLER_62_448 ();
 sg13g2_decap_4 FILLER_62_453 ();
 sg13g2_fill_2 FILLER_62_457 ();
 sg13g2_fill_2 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_506 ();
 sg13g2_fill_2 FILLER_62_562 ();
 sg13g2_fill_1 FILLER_62_564 ();
 sg13g2_decap_4 FILLER_62_583 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_fill_1 FILLER_62_658 ();
 sg13g2_fill_2 FILLER_62_675 ();
 sg13g2_decap_8 FILLER_62_687 ();
 sg13g2_decap_8 FILLER_62_694 ();
 sg13g2_decap_8 FILLER_62_701 ();
 sg13g2_decap_4 FILLER_62_708 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_fill_1 FILLER_62_717 ();
 sg13g2_fill_2 FILLER_62_723 ();
 sg13g2_fill_1 FILLER_62_725 ();
 sg13g2_fill_1 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_791 ();
 sg13g2_fill_1 FILLER_62_822 ();
 sg13g2_fill_1 FILLER_62_832 ();
 sg13g2_fill_1 FILLER_62_856 ();
 sg13g2_fill_2 FILLER_62_874 ();
 sg13g2_fill_1 FILLER_62_876 ();
 sg13g2_fill_2 FILLER_62_882 ();
 sg13g2_fill_1 FILLER_62_884 ();
 sg13g2_fill_1 FILLER_62_900 ();
 sg13g2_fill_1 FILLER_62_906 ();
 sg13g2_fill_1 FILLER_62_929 ();
 sg13g2_fill_1 FILLER_62_962 ();
 sg13g2_fill_2 FILLER_62_999 ();
 sg13g2_fill_1 FILLER_62_1001 ();
 sg13g2_decap_4 FILLER_62_1007 ();
 sg13g2_fill_1 FILLER_62_1011 ();
 sg13g2_fill_2 FILLER_62_1025 ();
 sg13g2_decap_4 FILLER_62_1032 ();
 sg13g2_fill_1 FILLER_62_1036 ();
 sg13g2_fill_1 FILLER_62_1047 ();
 sg13g2_fill_1 FILLER_62_1052 ();
 sg13g2_decap_4 FILLER_62_1057 ();
 sg13g2_fill_2 FILLER_62_1061 ();
 sg13g2_fill_1 FILLER_62_1072 ();
 sg13g2_decap_8 FILLER_62_1114 ();
 sg13g2_decap_4 FILLER_62_1121 ();
 sg13g2_fill_1 FILLER_62_1125 ();
 sg13g2_fill_2 FILLER_62_1135 ();
 sg13g2_fill_1 FILLER_62_1137 ();
 sg13g2_decap_8 FILLER_62_1148 ();
 sg13g2_fill_1 FILLER_62_1155 ();
 sg13g2_fill_2 FILLER_62_1160 ();
 sg13g2_fill_1 FILLER_62_1162 ();
 sg13g2_decap_4 FILLER_62_1212 ();
 sg13g2_fill_1 FILLER_62_1221 ();
 sg13g2_decap_4 FILLER_62_1261 ();
 sg13g2_decap_4 FILLER_62_1270 ();
 sg13g2_decap_4 FILLER_62_1305 ();
 sg13g2_fill_2 FILLER_62_1317 ();
 sg13g2_fill_1 FILLER_62_1319 ();
 sg13g2_decap_4 FILLER_62_1329 ();
 sg13g2_fill_2 FILLER_62_1374 ();
 sg13g2_fill_1 FILLER_62_1376 ();
 sg13g2_fill_2 FILLER_62_1382 ();
 sg13g2_fill_1 FILLER_62_1384 ();
 sg13g2_decap_4 FILLER_62_1389 ();
 sg13g2_fill_1 FILLER_62_1393 ();
 sg13g2_decap_8 FILLER_62_1399 ();
 sg13g2_decap_8 FILLER_62_1406 ();
 sg13g2_fill_1 FILLER_62_1413 ();
 sg13g2_fill_2 FILLER_62_1428 ();
 sg13g2_fill_1 FILLER_62_1430 ();
 sg13g2_fill_2 FILLER_62_1443 ();
 sg13g2_fill_1 FILLER_62_1445 ();
 sg13g2_fill_1 FILLER_62_1469 ();
 sg13g2_fill_2 FILLER_62_1488 ();
 sg13g2_decap_8 FILLER_62_1558 ();
 sg13g2_fill_1 FILLER_62_1565 ();
 sg13g2_fill_2 FILLER_62_1605 ();
 sg13g2_fill_1 FILLER_62_1607 ();
 sg13g2_fill_1 FILLER_62_1631 ();
 sg13g2_fill_1 FILLER_62_1669 ();
 sg13g2_decap_4 FILLER_62_1697 ();
 sg13g2_fill_1 FILLER_62_1701 ();
 sg13g2_decap_4 FILLER_62_1724 ();
 sg13g2_fill_1 FILLER_62_1728 ();
 sg13g2_decap_8 FILLER_62_1733 ();
 sg13g2_fill_2 FILLER_62_1740 ();
 sg13g2_decap_8 FILLER_62_1746 ();
 sg13g2_fill_2 FILLER_62_1753 ();
 sg13g2_fill_1 FILLER_62_1755 ();
 sg13g2_decap_8 FILLER_62_1785 ();
 sg13g2_decap_8 FILLER_62_1792 ();
 sg13g2_decap_4 FILLER_62_1799 ();
 sg13g2_decap_8 FILLER_62_1808 ();
 sg13g2_fill_2 FILLER_62_1827 ();
 sg13g2_fill_1 FILLER_62_1829 ();
 sg13g2_decap_8 FILLER_62_1848 ();
 sg13g2_fill_2 FILLER_62_1918 ();
 sg13g2_fill_1 FILLER_62_1933 ();
 sg13g2_fill_2 FILLER_62_1943 ();
 sg13g2_decap_8 FILLER_62_1954 ();
 sg13g2_decap_8 FILLER_62_1961 ();
 sg13g2_fill_2 FILLER_62_1968 ();
 sg13g2_fill_1 FILLER_62_2004 ();
 sg13g2_fill_2 FILLER_62_2018 ();
 sg13g2_fill_1 FILLER_62_2033 ();
 sg13g2_decap_8 FILLER_62_2045 ();
 sg13g2_fill_2 FILLER_62_2080 ();
 sg13g2_fill_1 FILLER_62_2082 ();
 sg13g2_fill_2 FILLER_62_2087 ();
 sg13g2_fill_1 FILLER_62_2089 ();
 sg13g2_fill_2 FILLER_62_2108 ();
 sg13g2_fill_2 FILLER_62_2132 ();
 sg13g2_decap_4 FILLER_62_2139 ();
 sg13g2_fill_1 FILLER_62_2143 ();
 sg13g2_decap_4 FILLER_62_2171 ();
 sg13g2_fill_2 FILLER_62_2196 ();
 sg13g2_decap_4 FILLER_62_2217 ();
 sg13g2_fill_1 FILLER_62_2221 ();
 sg13g2_fill_2 FILLER_62_2242 ();
 sg13g2_fill_1 FILLER_62_2244 ();
 sg13g2_fill_1 FILLER_62_2261 ();
 sg13g2_fill_2 FILLER_62_2270 ();
 sg13g2_fill_2 FILLER_62_2282 ();
 sg13g2_fill_1 FILLER_62_2284 ();
 sg13g2_fill_2 FILLER_62_2325 ();
 sg13g2_fill_1 FILLER_62_2327 ();
 sg13g2_fill_2 FILLER_62_2365 ();
 sg13g2_fill_1 FILLER_62_2376 ();
 sg13g2_fill_2 FILLER_62_2391 ();
 sg13g2_fill_1 FILLER_62_2393 ();
 sg13g2_decap_8 FILLER_62_2411 ();
 sg13g2_fill_2 FILLER_62_2418 ();
 sg13g2_fill_1 FILLER_62_2420 ();
 sg13g2_decap_8 FILLER_62_2462 ();
 sg13g2_decap_8 FILLER_62_2469 ();
 sg13g2_fill_2 FILLER_62_2480 ();
 sg13g2_fill_1 FILLER_62_2482 ();
 sg13g2_fill_2 FILLER_62_2492 ();
 sg13g2_fill_1 FILLER_62_2512 ();
 sg13g2_decap_8 FILLER_62_2535 ();
 sg13g2_fill_2 FILLER_62_2547 ();
 sg13g2_fill_2 FILLER_62_2571 ();
 sg13g2_fill_1 FILLER_62_2593 ();
 sg13g2_fill_1 FILLER_62_2605 ();
 sg13g2_decap_8 FILLER_62_2610 ();
 sg13g2_fill_2 FILLER_62_2617 ();
 sg13g2_fill_1 FILLER_62_2619 ();
 sg13g2_decap_8 FILLER_62_2624 ();
 sg13g2_fill_1 FILLER_62_2631 ();
 sg13g2_fill_2 FILLER_62_2636 ();
 sg13g2_fill_1 FILLER_62_2638 ();
 sg13g2_decap_8 FILLER_62_2647 ();
 sg13g2_decap_4 FILLER_62_2654 ();
 sg13g2_fill_2 FILLER_62_2658 ();
 sg13g2_decap_8 FILLER_62_2665 ();
 sg13g2_decap_4 FILLER_62_2672 ();
 sg13g2_fill_2 FILLER_62_2676 ();
 sg13g2_decap_8 FILLER_62_2692 ();
 sg13g2_fill_2 FILLER_62_2699 ();
 sg13g2_decap_8 FILLER_62_2709 ();
 sg13g2_decap_4 FILLER_62_2716 ();
 sg13g2_fill_2 FILLER_62_2720 ();
 sg13g2_decap_8 FILLER_62_2747 ();
 sg13g2_fill_2 FILLER_62_2754 ();
 sg13g2_decap_8 FILLER_62_2784 ();
 sg13g2_fill_2 FILLER_62_2799 ();
 sg13g2_fill_1 FILLER_62_2812 ();
 sg13g2_fill_2 FILLER_62_2827 ();
 sg13g2_fill_1 FILLER_62_2844 ();
 sg13g2_fill_2 FILLER_62_2859 ();
 sg13g2_fill_1 FILLER_62_2861 ();
 sg13g2_decap_8 FILLER_62_2866 ();
 sg13g2_decap_8 FILLER_62_2873 ();
 sg13g2_decap_4 FILLER_62_2880 ();
 sg13g2_fill_1 FILLER_62_2897 ();
 sg13g2_fill_1 FILLER_62_2919 ();
 sg13g2_decap_4 FILLER_62_2949 ();
 sg13g2_fill_2 FILLER_62_2953 ();
 sg13g2_fill_2 FILLER_62_3004 ();
 sg13g2_fill_1 FILLER_62_3006 ();
 sg13g2_fill_1 FILLER_62_3011 ();
 sg13g2_decap_8 FILLER_62_3057 ();
 sg13g2_decap_4 FILLER_62_3064 ();
 sg13g2_fill_1 FILLER_62_3068 ();
 sg13g2_decap_8 FILLER_62_3074 ();
 sg13g2_fill_1 FILLER_62_3081 ();
 sg13g2_decap_8 FILLER_62_3119 ();
 sg13g2_fill_1 FILLER_62_3126 ();
 sg13g2_fill_2 FILLER_62_3149 ();
 sg13g2_decap_8 FILLER_62_3156 ();
 sg13g2_fill_1 FILLER_62_3163 ();
 sg13g2_decap_4 FILLER_62_3171 ();
 sg13g2_fill_2 FILLER_62_3178 ();
 sg13g2_fill_1 FILLER_62_3180 ();
 sg13g2_fill_2 FILLER_62_3207 ();
 sg13g2_decap_4 FILLER_62_3227 ();
 sg13g2_fill_1 FILLER_62_3239 ();
 sg13g2_decap_8 FILLER_62_3245 ();
 sg13g2_decap_4 FILLER_62_3252 ();
 sg13g2_decap_8 FILLER_62_3268 ();
 sg13g2_decap_8 FILLER_62_3275 ();
 sg13g2_fill_1 FILLER_62_3282 ();
 sg13g2_decap_4 FILLER_62_3310 ();
 sg13g2_fill_1 FILLER_62_3314 ();
 sg13g2_fill_1 FILLER_62_3338 ();
 sg13g2_fill_2 FILLER_62_3360 ();
 sg13g2_fill_1 FILLER_62_3362 ();
 sg13g2_decap_8 FILLER_62_3376 ();
 sg13g2_decap_8 FILLER_62_3383 ();
 sg13g2_decap_8 FILLER_62_3390 ();
 sg13g2_decap_8 FILLER_62_3397 ();
 sg13g2_decap_8 FILLER_62_3404 ();
 sg13g2_decap_8 FILLER_62_3411 ();
 sg13g2_decap_8 FILLER_62_3418 ();
 sg13g2_decap_8 FILLER_62_3425 ();
 sg13g2_decap_8 FILLER_62_3432 ();
 sg13g2_decap_8 FILLER_62_3439 ();
 sg13g2_decap_8 FILLER_62_3446 ();
 sg13g2_decap_8 FILLER_62_3453 ();
 sg13g2_decap_8 FILLER_62_3460 ();
 sg13g2_decap_8 FILLER_62_3467 ();
 sg13g2_decap_8 FILLER_62_3474 ();
 sg13g2_decap_8 FILLER_62_3481 ();
 sg13g2_decap_8 FILLER_62_3488 ();
 sg13g2_decap_8 FILLER_62_3495 ();
 sg13g2_decap_8 FILLER_62_3502 ();
 sg13g2_decap_8 FILLER_62_3509 ();
 sg13g2_decap_8 FILLER_62_3516 ();
 sg13g2_decap_8 FILLER_62_3523 ();
 sg13g2_decap_8 FILLER_62_3530 ();
 sg13g2_decap_8 FILLER_62_3537 ();
 sg13g2_decap_8 FILLER_62_3544 ();
 sg13g2_decap_8 FILLER_62_3551 ();
 sg13g2_decap_8 FILLER_62_3558 ();
 sg13g2_decap_8 FILLER_62_3565 ();
 sg13g2_decap_8 FILLER_62_3572 ();
 sg13g2_fill_1 FILLER_62_3579 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_107 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_4 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_decap_4 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_174 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_decap_8 FILLER_63_235 ();
 sg13g2_fill_2 FILLER_63_242 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_decap_8 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_267 ();
 sg13g2_fill_2 FILLER_63_297 ();
 sg13g2_fill_1 FILLER_63_299 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_4 FILLER_63_349 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_fill_2 FILLER_63_448 ();
 sg13g2_fill_1 FILLER_63_450 ();
 sg13g2_fill_1 FILLER_63_459 ();
 sg13g2_fill_2 FILLER_63_473 ();
 sg13g2_decap_4 FILLER_63_493 ();
 sg13g2_fill_1 FILLER_63_497 ();
 sg13g2_decap_8 FILLER_63_507 ();
 sg13g2_decap_8 FILLER_63_514 ();
 sg13g2_decap_8 FILLER_63_521 ();
 sg13g2_fill_2 FILLER_63_528 ();
 sg13g2_fill_1 FILLER_63_530 ();
 sg13g2_decap_8 FILLER_63_604 ();
 sg13g2_fill_2 FILLER_63_611 ();
 sg13g2_fill_1 FILLER_63_613 ();
 sg13g2_fill_1 FILLER_63_653 ();
 sg13g2_fill_2 FILLER_63_686 ();
 sg13g2_fill_2 FILLER_63_749 ();
 sg13g2_fill_1 FILLER_63_751 ();
 sg13g2_fill_1 FILLER_63_765 ();
 sg13g2_fill_2 FILLER_63_875 ();
 sg13g2_fill_2 FILLER_63_886 ();
 sg13g2_decap_4 FILLER_63_902 ();
 sg13g2_decap_8 FILLER_63_952 ();
 sg13g2_fill_2 FILLER_63_959 ();
 sg13g2_fill_1 FILLER_63_961 ();
 sg13g2_fill_2 FILLER_63_996 ();
 sg13g2_decap_4 FILLER_63_1020 ();
 sg13g2_fill_2 FILLER_63_1037 ();
 sg13g2_fill_2 FILLER_63_1118 ();
 sg13g2_fill_1 FILLER_63_1120 ();
 sg13g2_fill_2 FILLER_63_1144 ();
 sg13g2_fill_2 FILLER_63_1186 ();
 sg13g2_fill_1 FILLER_63_1188 ();
 sg13g2_decap_4 FILLER_63_1214 ();
 sg13g2_decap_8 FILLER_63_1223 ();
 sg13g2_decap_4 FILLER_63_1230 ();
 sg13g2_fill_1 FILLER_63_1234 ();
 sg13g2_decap_4 FILLER_63_1239 ();
 sg13g2_fill_2 FILLER_63_1243 ();
 sg13g2_fill_2 FILLER_63_1250 ();
 sg13g2_fill_1 FILLER_63_1252 ();
 sg13g2_fill_2 FILLER_63_1263 ();
 sg13g2_fill_2 FILLER_63_1288 ();
 sg13g2_decap_4 FILLER_63_1358 ();
 sg13g2_fill_1 FILLER_63_1362 ();
 sg13g2_fill_2 FILLER_63_1403 ();
 sg13g2_fill_2 FILLER_63_1422 ();
 sg13g2_fill_2 FILLER_63_1433 ();
 sg13g2_fill_1 FILLER_63_1435 ();
 sg13g2_decap_8 FILLER_63_1453 ();
 sg13g2_decap_4 FILLER_63_1460 ();
 sg13g2_fill_2 FILLER_63_1464 ();
 sg13g2_fill_1 FILLER_63_1530 ();
 sg13g2_decap_8 FILLER_63_1581 ();
 sg13g2_decap_4 FILLER_63_1588 ();
 sg13g2_fill_1 FILLER_63_1631 ();
 sg13g2_decap_4 FILLER_63_1672 ();
 sg13g2_fill_1 FILLER_63_1676 ();
 sg13g2_fill_2 FILLER_63_1709 ();
 sg13g2_fill_1 FILLER_63_1711 ();
 sg13g2_fill_2 FILLER_63_1771 ();
 sg13g2_fill_2 FILLER_63_1777 ();
 sg13g2_fill_2 FILLER_63_1783 ();
 sg13g2_fill_1 FILLER_63_1785 ();
 sg13g2_decap_4 FILLER_63_1791 ();
 sg13g2_fill_2 FILLER_63_1795 ();
 sg13g2_fill_1 FILLER_63_1802 ();
 sg13g2_fill_2 FILLER_63_1816 ();
 sg13g2_decap_4 FILLER_63_1823 ();
 sg13g2_fill_2 FILLER_63_1827 ();
 sg13g2_decap_8 FILLER_63_1851 ();
 sg13g2_decap_4 FILLER_63_1858 ();
 sg13g2_fill_2 FILLER_63_1862 ();
 sg13g2_decap_4 FILLER_63_1868 ();
 sg13g2_fill_1 FILLER_63_1872 ();
 sg13g2_decap_4 FILLER_63_1901 ();
 sg13g2_fill_2 FILLER_63_1905 ();
 sg13g2_decap_8 FILLER_63_1935 ();
 sg13g2_fill_2 FILLER_63_1942 ();
 sg13g2_fill_1 FILLER_63_1944 ();
 sg13g2_fill_2 FILLER_63_1950 ();
 sg13g2_decap_8 FILLER_63_2026 ();
 sg13g2_decap_8 FILLER_63_2033 ();
 sg13g2_decap_4 FILLER_63_2040 ();
 sg13g2_fill_2 FILLER_63_2067 ();
 sg13g2_decap_4 FILLER_63_2110 ();
 sg13g2_decap_4 FILLER_63_2119 ();
 sg13g2_fill_2 FILLER_63_2123 ();
 sg13g2_decap_8 FILLER_63_2129 ();
 sg13g2_decap_8 FILLER_63_2136 ();
 sg13g2_decap_8 FILLER_63_2143 ();
 sg13g2_fill_2 FILLER_63_2150 ();
 sg13g2_decap_8 FILLER_63_2156 ();
 sg13g2_decap_8 FILLER_63_2163 ();
 sg13g2_fill_2 FILLER_63_2170 ();
 sg13g2_fill_1 FILLER_63_2172 ();
 sg13g2_fill_1 FILLER_63_2209 ();
 sg13g2_decap_4 FILLER_63_2217 ();
 sg13g2_fill_1 FILLER_63_2221 ();
 sg13g2_decap_8 FILLER_63_2237 ();
 sg13g2_decap_8 FILLER_63_2244 ();
 sg13g2_decap_4 FILLER_63_2251 ();
 sg13g2_fill_1 FILLER_63_2255 ();
 sg13g2_fill_1 FILLER_63_2271 ();
 sg13g2_fill_1 FILLER_63_2289 ();
 sg13g2_fill_2 FILLER_63_2294 ();
 sg13g2_fill_1 FILLER_63_2296 ();
 sg13g2_decap_4 FILLER_63_2306 ();
 sg13g2_fill_1 FILLER_63_2350 ();
 sg13g2_fill_2 FILLER_63_2366 ();
 sg13g2_fill_1 FILLER_63_2392 ();
 sg13g2_decap_4 FILLER_63_2401 ();
 sg13g2_fill_1 FILLER_63_2440 ();
 sg13g2_decap_8 FILLER_63_2476 ();
 sg13g2_fill_2 FILLER_63_2483 ();
 sg13g2_decap_4 FILLER_63_2532 ();
 sg13g2_fill_1 FILLER_63_2536 ();
 sg13g2_fill_2 FILLER_63_2637 ();
 sg13g2_fill_2 FILLER_63_2655 ();
 sg13g2_fill_1 FILLER_63_2657 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_fill_1 FILLER_63_2675 ();
 sg13g2_fill_2 FILLER_63_2688 ();
 sg13g2_fill_1 FILLER_63_2690 ();
 sg13g2_fill_2 FILLER_63_2705 ();
 sg13g2_fill_1 FILLER_63_2707 ();
 sg13g2_decap_4 FILLER_63_2719 ();
 sg13g2_decap_4 FILLER_63_2733 ();
 sg13g2_fill_2 FILLER_63_2743 ();
 sg13g2_fill_1 FILLER_63_2754 ();
 sg13g2_fill_1 FILLER_63_2764 ();
 sg13g2_decap_8 FILLER_63_2796 ();
 sg13g2_decap_4 FILLER_63_2803 ();
 sg13g2_fill_1 FILLER_63_2807 ();
 sg13g2_fill_2 FILLER_63_2811 ();
 sg13g2_fill_1 FILLER_63_2813 ();
 sg13g2_fill_1 FILLER_63_2823 ();
 sg13g2_decap_8 FILLER_63_2834 ();
 sg13g2_decap_4 FILLER_63_2841 ();
 sg13g2_fill_2 FILLER_63_2855 ();
 sg13g2_fill_2 FILLER_63_2898 ();
 sg13g2_fill_1 FILLER_63_2900 ();
 sg13g2_fill_2 FILLER_63_2906 ();
 sg13g2_fill_2 FILLER_63_2936 ();
 sg13g2_fill_1 FILLER_63_2955 ();
 sg13g2_fill_2 FILLER_63_2964 ();
 sg13g2_fill_2 FILLER_63_2982 ();
 sg13g2_fill_2 FILLER_63_2994 ();
 sg13g2_fill_1 FILLER_63_3005 ();
 sg13g2_fill_2 FILLER_63_3024 ();
 sg13g2_fill_2 FILLER_63_3030 ();
 sg13g2_fill_1 FILLER_63_3032 ();
 sg13g2_fill_2 FILLER_63_3082 ();
 sg13g2_fill_1 FILLER_63_3097 ();
 sg13g2_fill_1 FILLER_63_3103 ();
 sg13g2_decap_8 FILLER_63_3174 ();
 sg13g2_fill_1 FILLER_63_3181 ();
 sg13g2_decap_8 FILLER_63_3200 ();
 sg13g2_decap_4 FILLER_63_3207 ();
 sg13g2_fill_2 FILLER_63_3211 ();
 sg13g2_decap_4 FILLER_63_3226 ();
 sg13g2_fill_1 FILLER_63_3254 ();
 sg13g2_decap_8 FILLER_63_3273 ();
 sg13g2_decap_4 FILLER_63_3280 ();
 sg13g2_fill_1 FILLER_63_3284 ();
 sg13g2_decap_8 FILLER_63_3306 ();
 sg13g2_decap_4 FILLER_63_3313 ();
 sg13g2_fill_2 FILLER_63_3317 ();
 sg13g2_decap_8 FILLER_63_3328 ();
 sg13g2_decap_4 FILLER_63_3335 ();
 sg13g2_fill_1 FILLER_63_3339 ();
 sg13g2_fill_2 FILLER_63_3370 ();
 sg13g2_fill_1 FILLER_63_3372 ();
 sg13g2_decap_8 FILLER_63_3400 ();
 sg13g2_decap_8 FILLER_63_3407 ();
 sg13g2_decap_8 FILLER_63_3414 ();
 sg13g2_decap_8 FILLER_63_3421 ();
 sg13g2_decap_8 FILLER_63_3428 ();
 sg13g2_decap_8 FILLER_63_3435 ();
 sg13g2_decap_8 FILLER_63_3442 ();
 sg13g2_decap_8 FILLER_63_3449 ();
 sg13g2_decap_8 FILLER_63_3456 ();
 sg13g2_decap_8 FILLER_63_3463 ();
 sg13g2_decap_8 FILLER_63_3470 ();
 sg13g2_decap_8 FILLER_63_3477 ();
 sg13g2_decap_8 FILLER_63_3484 ();
 sg13g2_decap_8 FILLER_63_3491 ();
 sg13g2_decap_8 FILLER_63_3498 ();
 sg13g2_decap_8 FILLER_63_3505 ();
 sg13g2_decap_8 FILLER_63_3512 ();
 sg13g2_decap_8 FILLER_63_3519 ();
 sg13g2_decap_8 FILLER_63_3526 ();
 sg13g2_decap_8 FILLER_63_3533 ();
 sg13g2_decap_8 FILLER_63_3540 ();
 sg13g2_decap_8 FILLER_63_3547 ();
 sg13g2_decap_8 FILLER_63_3554 ();
 sg13g2_decap_8 FILLER_63_3561 ();
 sg13g2_decap_8 FILLER_63_3568 ();
 sg13g2_decap_4 FILLER_63_3575 ();
 sg13g2_fill_1 FILLER_63_3579 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_279 ();
 sg13g2_decap_4 FILLER_64_289 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_fill_1 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_405 ();
 sg13g2_fill_1 FILLER_64_412 ();
 sg13g2_fill_2 FILLER_64_441 ();
 sg13g2_fill_2 FILLER_64_456 ();
 sg13g2_fill_1 FILLER_64_458 ();
 sg13g2_decap_8 FILLER_64_472 ();
 sg13g2_decap_8 FILLER_64_479 ();
 sg13g2_fill_2 FILLER_64_486 ();
 sg13g2_fill_1 FILLER_64_488 ();
 sg13g2_decap_4 FILLER_64_517 ();
 sg13g2_fill_1 FILLER_64_547 ();
 sg13g2_fill_2 FILLER_64_558 ();
 sg13g2_fill_1 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_570 ();
 sg13g2_decap_8 FILLER_64_582 ();
 sg13g2_decap_8 FILLER_64_601 ();
 sg13g2_decap_4 FILLER_64_608 ();
 sg13g2_fill_1 FILLER_64_667 ();
 sg13g2_fill_2 FILLER_64_684 ();
 sg13g2_decap_4 FILLER_64_707 ();
 sg13g2_fill_1 FILLER_64_711 ();
 sg13g2_fill_2 FILLER_64_723 ();
 sg13g2_decap_8 FILLER_64_729 ();
 sg13g2_fill_2 FILLER_64_773 ();
 sg13g2_fill_2 FILLER_64_812 ();
 sg13g2_fill_2 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_decap_4 FILLER_64_900 ();
 sg13g2_decap_4 FILLER_64_950 ();
 sg13g2_decap_4 FILLER_64_990 ();
 sg13g2_fill_2 FILLER_64_1026 ();
 sg13g2_fill_2 FILLER_64_1041 ();
 sg13g2_fill_1 FILLER_64_1043 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_fill_1 FILLER_64_1055 ();
 sg13g2_fill_1 FILLER_64_1071 ();
 sg13g2_fill_1 FILLER_64_1090 ();
 sg13g2_fill_2 FILLER_64_1141 ();
 sg13g2_fill_1 FILLER_64_1143 ();
 sg13g2_fill_2 FILLER_64_1153 ();
 sg13g2_fill_1 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1187 ();
 sg13g2_fill_2 FILLER_64_1197 ();
 sg13g2_fill_1 FILLER_64_1199 ();
 sg13g2_fill_1 FILLER_64_1205 ();
 sg13g2_fill_1 FILLER_64_1283 ();
 sg13g2_fill_2 FILLER_64_1321 ();
 sg13g2_decap_4 FILLER_64_1346 ();
 sg13g2_fill_1 FILLER_64_1350 ();
 sg13g2_decap_4 FILLER_64_1360 ();
 sg13g2_fill_1 FILLER_64_1364 ();
 sg13g2_decap_8 FILLER_64_1378 ();
 sg13g2_decap_8 FILLER_64_1385 ();
 sg13g2_decap_8 FILLER_64_1461 ();
 sg13g2_decap_4 FILLER_64_1468 ();
 sg13g2_decap_4 FILLER_64_1481 ();
 sg13g2_decap_4 FILLER_64_1495 ();
 sg13g2_fill_2 FILLER_64_1499 ();
 sg13g2_fill_1 FILLER_64_1518 ();
 sg13g2_decap_4 FILLER_64_1560 ();
 sg13g2_decap_4 FILLER_64_1577 ();
 sg13g2_fill_2 FILLER_64_1591 ();
 sg13g2_fill_2 FILLER_64_1620 ();
 sg13g2_fill_2 FILLER_64_1664 ();
 sg13g2_fill_1 FILLER_64_1666 ();
 sg13g2_fill_1 FILLER_64_1694 ();
 sg13g2_decap_4 FILLER_64_1704 ();
 sg13g2_fill_1 FILLER_64_1708 ();
 sg13g2_fill_2 FILLER_64_1729 ();
 sg13g2_fill_2 FILLER_64_1771 ();
 sg13g2_fill_2 FILLER_64_1781 ();
 sg13g2_fill_1 FILLER_64_1796 ();
 sg13g2_fill_1 FILLER_64_1802 ();
 sg13g2_fill_2 FILLER_64_1808 ();
 sg13g2_fill_1 FILLER_64_1810 ();
 sg13g2_decap_8 FILLER_64_1826 ();
 sg13g2_fill_2 FILLER_64_1843 ();
 sg13g2_fill_1 FILLER_64_1845 ();
 sg13g2_fill_2 FILLER_64_1859 ();
 sg13g2_fill_1 FILLER_64_1861 ();
 sg13g2_decap_8 FILLER_64_1889 ();
 sg13g2_fill_1 FILLER_64_1896 ();
 sg13g2_fill_2 FILLER_64_1916 ();
 sg13g2_fill_1 FILLER_64_1921 ();
 sg13g2_decap_4 FILLER_64_1943 ();
 sg13g2_fill_2 FILLER_64_1956 ();
 sg13g2_fill_1 FILLER_64_1962 ();
 sg13g2_fill_1 FILLER_64_1972 ();
 sg13g2_fill_1 FILLER_64_2011 ();
 sg13g2_decap_8 FILLER_64_2034 ();
 sg13g2_fill_1 FILLER_64_2041 ();
 sg13g2_fill_2 FILLER_64_2080 ();
 sg13g2_decap_8 FILLER_64_2095 ();
 sg13g2_decap_8 FILLER_64_2102 ();
 sg13g2_decap_4 FILLER_64_2109 ();
 sg13g2_fill_1 FILLER_64_2113 ();
 sg13g2_fill_2 FILLER_64_2145 ();
 sg13g2_decap_4 FILLER_64_2214 ();
 sg13g2_fill_2 FILLER_64_2218 ();
 sg13g2_fill_2 FILLER_64_2224 ();
 sg13g2_fill_1 FILLER_64_2226 ();
 sg13g2_decap_8 FILLER_64_2235 ();
 sg13g2_fill_1 FILLER_64_2242 ();
 sg13g2_decap_4 FILLER_64_2248 ();
 sg13g2_fill_1 FILLER_64_2252 ();
 sg13g2_fill_2 FILLER_64_2261 ();
 sg13g2_fill_1 FILLER_64_2263 ();
 sg13g2_fill_2 FILLER_64_2274 ();
 sg13g2_decap_8 FILLER_64_2290 ();
 sg13g2_decap_4 FILLER_64_2297 ();
 sg13g2_fill_1 FILLER_64_2301 ();
 sg13g2_decap_8 FILLER_64_2334 ();
 sg13g2_decap_4 FILLER_64_2341 ();
 sg13g2_fill_1 FILLER_64_2345 ();
 sg13g2_fill_1 FILLER_64_2374 ();
 sg13g2_fill_2 FILLER_64_2396 ();
 sg13g2_decap_8 FILLER_64_2403 ();
 sg13g2_fill_1 FILLER_64_2410 ();
 sg13g2_decap_8 FILLER_64_2415 ();
 sg13g2_fill_1 FILLER_64_2431 ();
 sg13g2_fill_2 FILLER_64_2473 ();
 sg13g2_fill_1 FILLER_64_2475 ();
 sg13g2_fill_1 FILLER_64_2489 ();
 sg13g2_fill_2 FILLER_64_2516 ();
 sg13g2_fill_1 FILLER_64_2518 ();
 sg13g2_decap_4 FILLER_64_2531 ();
 sg13g2_fill_2 FILLER_64_2535 ();
 sg13g2_decap_4 FILLER_64_2563 ();
 sg13g2_fill_1 FILLER_64_2567 ();
 sg13g2_decap_8 FILLER_64_2572 ();
 sg13g2_decap_8 FILLER_64_2579 ();
 sg13g2_fill_2 FILLER_64_2586 ();
 sg13g2_fill_1 FILLER_64_2588 ();
 sg13g2_fill_1 FILLER_64_2593 ();
 sg13g2_fill_2 FILLER_64_2608 ();
 sg13g2_fill_2 FILLER_64_2632 ();
 sg13g2_fill_1 FILLER_64_2634 ();
 sg13g2_fill_2 FILLER_64_2639 ();
 sg13g2_fill_1 FILLER_64_2641 ();
 sg13g2_decap_4 FILLER_64_2647 ();
 sg13g2_decap_8 FILLER_64_2672 ();
 sg13g2_decap_4 FILLER_64_2682 ();
 sg13g2_fill_1 FILLER_64_2686 ();
 sg13g2_decap_8 FILLER_64_2691 ();
 sg13g2_fill_2 FILLER_64_2698 ();
 sg13g2_fill_1 FILLER_64_2700 ();
 sg13g2_fill_2 FILLER_64_2712 ();
 sg13g2_fill_2 FILLER_64_2723 ();
 sg13g2_decap_8 FILLER_64_2751 ();
 sg13g2_fill_2 FILLER_64_2758 ();
 sg13g2_fill_1 FILLER_64_2769 ();
 sg13g2_fill_2 FILLER_64_2783 ();
 sg13g2_fill_1 FILLER_64_2785 ();
 sg13g2_fill_2 FILLER_64_2807 ();
 sg13g2_decap_4 FILLER_64_2821 ();
 sg13g2_decap_4 FILLER_64_2844 ();
 sg13g2_fill_1 FILLER_64_2848 ();
 sg13g2_fill_1 FILLER_64_2867 ();
 sg13g2_decap_8 FILLER_64_2877 ();
 sg13g2_decap_4 FILLER_64_2910 ();
 sg13g2_fill_1 FILLER_64_2914 ();
 sg13g2_fill_2 FILLER_64_2932 ();
 sg13g2_fill_1 FILLER_64_2934 ();
 sg13g2_fill_2 FILLER_64_2955 ();
 sg13g2_fill_1 FILLER_64_2957 ();
 sg13g2_fill_2 FILLER_64_2963 ();
 sg13g2_fill_1 FILLER_64_2965 ();
 sg13g2_decap_4 FILLER_64_2978 ();
 sg13g2_decap_4 FILLER_64_3013 ();
 sg13g2_fill_2 FILLER_64_3017 ();
 sg13g2_fill_2 FILLER_64_3024 ();
 sg13g2_fill_1 FILLER_64_3026 ();
 sg13g2_decap_4 FILLER_64_3042 ();
 sg13g2_fill_1 FILLER_64_3046 ();
 sg13g2_fill_1 FILLER_64_3072 ();
 sg13g2_decap_4 FILLER_64_3088 ();
 sg13g2_fill_1 FILLER_64_3092 ();
 sg13g2_fill_2 FILLER_64_3113 ();
 sg13g2_fill_1 FILLER_64_3115 ();
 sg13g2_decap_8 FILLER_64_3137 ();
 sg13g2_decap_8 FILLER_64_3152 ();
 sg13g2_decap_8 FILLER_64_3159 ();
 sg13g2_decap_8 FILLER_64_3197 ();
 sg13g2_fill_2 FILLER_64_3204 ();
 sg13g2_fill_1 FILLER_64_3217 ();
 sg13g2_fill_2 FILLER_64_3245 ();
 sg13g2_fill_1 FILLER_64_3247 ();
 sg13g2_decap_4 FILLER_64_3251 ();
 sg13g2_fill_2 FILLER_64_3255 ();
 sg13g2_fill_2 FILLER_64_3282 ();
 sg13g2_fill_2 FILLER_64_3312 ();
 sg13g2_fill_1 FILLER_64_3314 ();
 sg13g2_fill_2 FILLER_64_3356 ();
 sg13g2_fill_1 FILLER_64_3358 ();
 sg13g2_decap_8 FILLER_64_3396 ();
 sg13g2_decap_8 FILLER_64_3403 ();
 sg13g2_decap_8 FILLER_64_3410 ();
 sg13g2_decap_8 FILLER_64_3417 ();
 sg13g2_decap_8 FILLER_64_3424 ();
 sg13g2_decap_8 FILLER_64_3431 ();
 sg13g2_decap_8 FILLER_64_3438 ();
 sg13g2_decap_8 FILLER_64_3445 ();
 sg13g2_decap_8 FILLER_64_3452 ();
 sg13g2_decap_8 FILLER_64_3459 ();
 sg13g2_decap_8 FILLER_64_3466 ();
 sg13g2_decap_8 FILLER_64_3473 ();
 sg13g2_decap_8 FILLER_64_3480 ();
 sg13g2_decap_8 FILLER_64_3487 ();
 sg13g2_decap_8 FILLER_64_3494 ();
 sg13g2_decap_8 FILLER_64_3501 ();
 sg13g2_decap_8 FILLER_64_3508 ();
 sg13g2_decap_8 FILLER_64_3515 ();
 sg13g2_decap_8 FILLER_64_3522 ();
 sg13g2_decap_8 FILLER_64_3529 ();
 sg13g2_decap_8 FILLER_64_3536 ();
 sg13g2_decap_8 FILLER_64_3543 ();
 sg13g2_decap_8 FILLER_64_3550 ();
 sg13g2_decap_8 FILLER_64_3557 ();
 sg13g2_decap_8 FILLER_64_3564 ();
 sg13g2_decap_8 FILLER_64_3571 ();
 sg13g2_fill_2 FILLER_64_3578 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_fill_2 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_182 ();
 sg13g2_fill_1 FILLER_65_192 ();
 sg13g2_decap_4 FILLER_65_220 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_fill_1 FILLER_65_287 ();
 sg13g2_fill_2 FILLER_65_321 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_fill_1 FILLER_65_436 ();
 sg13g2_fill_1 FILLER_65_446 ();
 sg13g2_decap_4 FILLER_65_482 ();
 sg13g2_decap_8 FILLER_65_506 ();
 sg13g2_decap_8 FILLER_65_513 ();
 sg13g2_decap_8 FILLER_65_520 ();
 sg13g2_fill_2 FILLER_65_527 ();
 sg13g2_fill_1 FILLER_65_533 ();
 sg13g2_fill_2 FILLER_65_547 ();
 sg13g2_fill_2 FILLER_65_639 ();
 sg13g2_fill_1 FILLER_65_650 ();
 sg13g2_fill_2 FILLER_65_691 ();
 sg13g2_fill_2 FILLER_65_704 ();
 sg13g2_decap_4 FILLER_65_712 ();
 sg13g2_fill_1 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_754 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_fill_2 FILLER_65_783 ();
 sg13g2_fill_1 FILLER_65_785 ();
 sg13g2_decap_4 FILLER_65_878 ();
 sg13g2_decap_4 FILLER_65_892 ();
 sg13g2_fill_1 FILLER_65_896 ();
 sg13g2_decap_4 FILLER_65_907 ();
 sg13g2_fill_1 FILLER_65_911 ();
 sg13g2_decap_8 FILLER_65_916 ();
 sg13g2_decap_8 FILLER_65_923 ();
 sg13g2_fill_2 FILLER_65_930 ();
 sg13g2_fill_2 FILLER_65_946 ();
 sg13g2_fill_1 FILLER_65_948 ();
 sg13g2_decap_4 FILLER_65_963 ();
 sg13g2_fill_1 FILLER_65_967 ();
 sg13g2_fill_2 FILLER_65_977 ();
 sg13g2_fill_2 FILLER_65_1006 ();
 sg13g2_fill_2 FILLER_65_1022 ();
 sg13g2_fill_1 FILLER_65_1024 ();
 sg13g2_fill_2 FILLER_65_1070 ();
 sg13g2_fill_1 FILLER_65_1081 ();
 sg13g2_fill_2 FILLER_65_1119 ();
 sg13g2_fill_1 FILLER_65_1121 ();
 sg13g2_decap_4 FILLER_65_1127 ();
 sg13g2_fill_1 FILLER_65_1204 ();
 sg13g2_decap_8 FILLER_65_1218 ();
 sg13g2_decap_8 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1232 ();
 sg13g2_fill_1 FILLER_65_1239 ();
 sg13g2_fill_2 FILLER_65_1249 ();
 sg13g2_decap_8 FILLER_65_1264 ();
 sg13g2_decap_8 FILLER_65_1271 ();
 sg13g2_decap_4 FILLER_65_1283 ();
 sg13g2_fill_2 FILLER_65_1311 ();
 sg13g2_decap_4 FILLER_65_1362 ();
 sg13g2_fill_1 FILLER_65_1421 ();
 sg13g2_fill_1 FILLER_65_1435 ();
 sg13g2_fill_2 FILLER_65_1449 ();
 sg13g2_fill_1 FILLER_65_1460 ();
 sg13g2_fill_2 FILLER_65_1488 ();
 sg13g2_decap_4 FILLER_65_1502 ();
 sg13g2_fill_2 FILLER_65_1506 ();
 sg13g2_decap_4 FILLER_65_1535 ();
 sg13g2_fill_1 FILLER_65_1552 ();
 sg13g2_decap_4 FILLER_65_1602 ();
 sg13g2_fill_1 FILLER_65_1606 ();
 sg13g2_fill_2 FILLER_65_1630 ();
 sg13g2_fill_2 FILLER_65_1645 ();
 sg13g2_fill_1 FILLER_65_1659 ();
 sg13g2_fill_1 FILLER_65_1686 ();
 sg13g2_fill_2 FILLER_65_1692 ();
 sg13g2_fill_2 FILLER_65_1730 ();
 sg13g2_fill_1 FILLER_65_1751 ();
 sg13g2_fill_2 FILLER_65_1765 ();
 sg13g2_fill_1 FILLER_65_1767 ();
 sg13g2_fill_2 FILLER_65_1780 ();
 sg13g2_decap_8 FILLER_65_1795 ();
 sg13g2_decap_4 FILLER_65_1802 ();
 sg13g2_fill_1 FILLER_65_1806 ();
 sg13g2_decap_8 FILLER_65_1824 ();
 sg13g2_decap_4 FILLER_65_1831 ();
 sg13g2_fill_1 FILLER_65_1835 ();
 sg13g2_decap_4 FILLER_65_1878 ();
 sg13g2_fill_2 FILLER_65_1882 ();
 sg13g2_decap_4 FILLER_65_1925 ();
 sg13g2_fill_1 FILLER_65_1929 ();
 sg13g2_fill_1 FILLER_65_1965 ();
 sg13g2_fill_1 FILLER_65_1985 ();
 sg13g2_fill_1 FILLER_65_2003 ();
 sg13g2_fill_1 FILLER_65_2025 ();
 sg13g2_decap_8 FILLER_65_2034 ();
 sg13g2_decap_8 FILLER_65_2041 ();
 sg13g2_fill_2 FILLER_65_2048 ();
 sg13g2_fill_1 FILLER_65_2050 ();
 sg13g2_fill_2 FILLER_65_2068 ();
 sg13g2_fill_1 FILLER_65_2076 ();
 sg13g2_fill_1 FILLER_65_2114 ();
 sg13g2_decap_8 FILLER_65_2152 ();
 sg13g2_fill_1 FILLER_65_2159 ();
 sg13g2_decap_8 FILLER_65_2221 ();
 sg13g2_decap_4 FILLER_65_2228 ();
 sg13g2_decap_8 FILLER_65_2254 ();
 sg13g2_fill_2 FILLER_65_2261 ();
 sg13g2_fill_1 FILLER_65_2263 ();
 sg13g2_fill_2 FILLER_65_2279 ();
 sg13g2_fill_1 FILLER_65_2281 ();
 sg13g2_fill_1 FILLER_65_2288 ();
 sg13g2_fill_2 FILLER_65_2301 ();
 sg13g2_decap_8 FILLER_65_2316 ();
 sg13g2_decap_8 FILLER_65_2336 ();
 sg13g2_fill_2 FILLER_65_2343 ();
 sg13g2_decap_4 FILLER_65_2353 ();
 sg13g2_fill_1 FILLER_65_2357 ();
 sg13g2_fill_2 FILLER_65_2369 ();
 sg13g2_fill_1 FILLER_65_2389 ();
 sg13g2_decap_4 FILLER_65_2400 ();
 sg13g2_fill_1 FILLER_65_2404 ();
 sg13g2_decap_8 FILLER_65_2409 ();
 sg13g2_decap_8 FILLER_65_2416 ();
 sg13g2_fill_1 FILLER_65_2423 ();
 sg13g2_fill_2 FILLER_65_2432 ();
 sg13g2_fill_2 FILLER_65_2438 ();
 sg13g2_fill_1 FILLER_65_2440 ();
 sg13g2_fill_1 FILLER_65_2446 ();
 sg13g2_decap_8 FILLER_65_2458 ();
 sg13g2_fill_2 FILLER_65_2465 ();
 sg13g2_decap_8 FILLER_65_2476 ();
 sg13g2_decap_4 FILLER_65_2483 ();
 sg13g2_fill_1 FILLER_65_2487 ();
 sg13g2_fill_2 FILLER_65_2498 ();
 sg13g2_fill_1 FILLER_65_2500 ();
 sg13g2_fill_2 FILLER_65_2510 ();
 sg13g2_fill_1 FILLER_65_2512 ();
 sg13g2_fill_2 FILLER_65_2518 ();
 sg13g2_fill_1 FILLER_65_2535 ();
 sg13g2_decap_8 FILLER_65_2552 ();
 sg13g2_decap_8 FILLER_65_2559 ();
 sg13g2_decap_8 FILLER_65_2566 ();
 sg13g2_fill_2 FILLER_65_2573 ();
 sg13g2_fill_2 FILLER_65_2581 ();
 sg13g2_fill_1 FILLER_65_2583 ();
 sg13g2_fill_1 FILLER_65_2639 ();
 sg13g2_fill_2 FILLER_65_2653 ();
 sg13g2_fill_2 FILLER_65_2664 ();
 sg13g2_fill_1 FILLER_65_2666 ();
 sg13g2_decap_8 FILLER_65_2671 ();
 sg13g2_decap_4 FILLER_65_2678 ();
 sg13g2_fill_2 FILLER_65_2710 ();
 sg13g2_decap_4 FILLER_65_2730 ();
 sg13g2_fill_2 FILLER_65_2734 ();
 sg13g2_fill_2 FILLER_65_2740 ();
 sg13g2_fill_1 FILLER_65_2742 ();
 sg13g2_decap_8 FILLER_65_2747 ();
 sg13g2_fill_2 FILLER_65_2778 ();
 sg13g2_decap_8 FILLER_65_2784 ();
 sg13g2_decap_4 FILLER_65_2791 ();
 sg13g2_fill_2 FILLER_65_2795 ();
 sg13g2_fill_2 FILLER_65_2802 ();
 sg13g2_fill_1 FILLER_65_2816 ();
 sg13g2_decap_4 FILLER_65_2822 ();
 sg13g2_fill_2 FILLER_65_2836 ();
 sg13g2_fill_1 FILLER_65_2849 ();
 sg13g2_decap_4 FILLER_65_2881 ();
 sg13g2_fill_2 FILLER_65_2890 ();
 sg13g2_fill_2 FILLER_65_2928 ();
 sg13g2_fill_1 FILLER_65_2930 ();
 sg13g2_fill_2 FILLER_65_2959 ();
 sg13g2_fill_1 FILLER_65_2961 ();
 sg13g2_fill_1 FILLER_65_2970 ();
 sg13g2_decap_8 FILLER_65_2975 ();
 sg13g2_decap_8 FILLER_65_2982 ();
 sg13g2_fill_1 FILLER_65_2989 ();
 sg13g2_decap_8 FILLER_65_2995 ();
 sg13g2_decap_8 FILLER_65_3002 ();
 sg13g2_fill_2 FILLER_65_3009 ();
 sg13g2_fill_1 FILLER_65_3011 ();
 sg13g2_decap_8 FILLER_65_3024 ();
 sg13g2_fill_1 FILLER_65_3039 ();
 sg13g2_decap_4 FILLER_65_3057 ();
 sg13g2_fill_1 FILLER_65_3061 ();
 sg13g2_fill_2 FILLER_65_3071 ();
 sg13g2_fill_1 FILLER_65_3073 ();
 sg13g2_fill_1 FILLER_65_3110 ();
 sg13g2_decap_8 FILLER_65_3132 ();
 sg13g2_fill_2 FILLER_65_3139 ();
 sg13g2_decap_4 FILLER_65_3186 ();
 sg13g2_decap_8 FILLER_65_3238 ();
 sg13g2_decap_4 FILLER_65_3245 ();
 sg13g2_fill_1 FILLER_65_3249 ();
 sg13g2_fill_2 FILLER_65_3271 ();
 sg13g2_fill_2 FILLER_65_3285 ();
 sg13g2_fill_2 FILLER_65_3313 ();
 sg13g2_fill_2 FILLER_65_3336 ();
 sg13g2_fill_1 FILLER_65_3338 ();
 sg13g2_decap_4 FILLER_65_3358 ();
 sg13g2_fill_2 FILLER_65_3362 ();
 sg13g2_decap_8 FILLER_65_3368 ();
 sg13g2_fill_2 FILLER_65_3375 ();
 sg13g2_fill_1 FILLER_65_3377 ();
 sg13g2_decap_8 FILLER_65_3382 ();
 sg13g2_decap_8 FILLER_65_3389 ();
 sg13g2_decap_8 FILLER_65_3396 ();
 sg13g2_decap_8 FILLER_65_3403 ();
 sg13g2_decap_8 FILLER_65_3410 ();
 sg13g2_decap_8 FILLER_65_3417 ();
 sg13g2_decap_8 FILLER_65_3424 ();
 sg13g2_decap_8 FILLER_65_3431 ();
 sg13g2_decap_8 FILLER_65_3438 ();
 sg13g2_decap_8 FILLER_65_3445 ();
 sg13g2_decap_8 FILLER_65_3452 ();
 sg13g2_decap_8 FILLER_65_3459 ();
 sg13g2_decap_8 FILLER_65_3466 ();
 sg13g2_decap_8 FILLER_65_3473 ();
 sg13g2_decap_8 FILLER_65_3480 ();
 sg13g2_decap_8 FILLER_65_3487 ();
 sg13g2_decap_8 FILLER_65_3494 ();
 sg13g2_decap_8 FILLER_65_3501 ();
 sg13g2_decap_8 FILLER_65_3508 ();
 sg13g2_decap_8 FILLER_65_3515 ();
 sg13g2_decap_8 FILLER_65_3522 ();
 sg13g2_decap_8 FILLER_65_3529 ();
 sg13g2_decap_8 FILLER_65_3536 ();
 sg13g2_decap_8 FILLER_65_3543 ();
 sg13g2_decap_8 FILLER_65_3550 ();
 sg13g2_decap_8 FILLER_65_3557 ();
 sg13g2_decap_8 FILLER_65_3564 ();
 sg13g2_decap_8 FILLER_65_3571 ();
 sg13g2_fill_2 FILLER_65_3578 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_4 FILLER_66_147 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_216 ();
 sg13g2_fill_1 FILLER_66_218 ();
 sg13g2_fill_2 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_267 ();
 sg13g2_decap_8 FILLER_66_290 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_fill_1 FILLER_66_299 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_339 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_359 ();
 sg13g2_fill_2 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_407 ();
 sg13g2_decap_4 FILLER_66_414 ();
 sg13g2_fill_1 FILLER_66_418 ();
 sg13g2_decap_8 FILLER_66_472 ();
 sg13g2_decap_4 FILLER_66_479 ();
 sg13g2_decap_8 FILLER_66_488 ();
 sg13g2_decap_4 FILLER_66_495 ();
 sg13g2_fill_1 FILLER_66_499 ();
 sg13g2_decap_4 FILLER_66_513 ();
 sg13g2_decap_4 FILLER_66_560 ();
 sg13g2_fill_2 FILLER_66_573 ();
 sg13g2_fill_1 FILLER_66_584 ();
 sg13g2_fill_2 FILLER_66_599 ();
 sg13g2_fill_2 FILLER_66_624 ();
 sg13g2_fill_1 FILLER_66_635 ();
 sg13g2_fill_2 FILLER_66_646 ();
 sg13g2_fill_1 FILLER_66_648 ();
 sg13g2_fill_1 FILLER_66_663 ();
 sg13g2_fill_2 FILLER_66_677 ();
 sg13g2_decap_8 FILLER_66_683 ();
 sg13g2_fill_2 FILLER_66_690 ();
 sg13g2_fill_1 FILLER_66_720 ();
 sg13g2_fill_2 FILLER_66_734 ();
 sg13g2_fill_1 FILLER_66_736 ();
 sg13g2_fill_1 FILLER_66_774 ();
 sg13g2_fill_1 FILLER_66_816 ();
 sg13g2_fill_2 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_868 ();
 sg13g2_fill_2 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_950 ();
 sg13g2_decap_4 FILLER_66_988 ();
 sg13g2_fill_1 FILLER_66_992 ();
 sg13g2_fill_2 FILLER_66_1030 ();
 sg13g2_fill_2 FILLER_66_1041 ();
 sg13g2_fill_1 FILLER_66_1043 ();
 sg13g2_fill_2 FILLER_66_1108 ();
 sg13g2_decap_8 FILLER_66_1119 ();
 sg13g2_decap_8 FILLER_66_1126 ();
 sg13g2_fill_2 FILLER_66_1133 ();
 sg13g2_fill_1 FILLER_66_1135 ();
 sg13g2_fill_2 FILLER_66_1212 ();
 sg13g2_fill_1 FILLER_66_1214 ();
 sg13g2_fill_2 FILLER_66_1253 ();
 sg13g2_decap_8 FILLER_66_1309 ();
 sg13g2_fill_1 FILLER_66_1316 ();
 sg13g2_fill_1 FILLER_66_1320 ();
 sg13g2_decap_8 FILLER_66_1363 ();
 sg13g2_fill_1 FILLER_66_1370 ();
 sg13g2_decap_4 FILLER_66_1379 ();
 sg13g2_fill_1 FILLER_66_1383 ();
 sg13g2_fill_1 FILLER_66_1393 ();
 sg13g2_fill_1 FILLER_66_1452 ();
 sg13g2_fill_2 FILLER_66_1503 ();
 sg13g2_fill_1 FILLER_66_1505 ();
 sg13g2_fill_2 FILLER_66_1516 ();
 sg13g2_fill_1 FILLER_66_1532 ();
 sg13g2_decap_4 FILLER_66_1570 ();
 sg13g2_decap_8 FILLER_66_1583 ();
 sg13g2_fill_2 FILLER_66_1590 ();
 sg13g2_fill_1 FILLER_66_1592 ();
 sg13g2_fill_1 FILLER_66_1645 ();
 sg13g2_decap_4 FILLER_66_1673 ();
 sg13g2_fill_1 FILLER_66_1677 ();
 sg13g2_decap_4 FILLER_66_1715 ();
 sg13g2_fill_1 FILLER_66_1719 ();
 sg13g2_decap_8 FILLER_66_1777 ();
 sg13g2_fill_2 FILLER_66_1784 ();
 sg13g2_fill_1 FILLER_66_1786 ();
 sg13g2_fill_1 FILLER_66_1800 ();
 sg13g2_fill_2 FILLER_66_1846 ();
 sg13g2_decap_8 FILLER_66_1861 ();
 sg13g2_fill_2 FILLER_66_1868 ();
 sg13g2_fill_1 FILLER_66_1870 ();
 sg13g2_decap_8 FILLER_66_1884 ();
 sg13g2_decap_8 FILLER_66_1891 ();
 sg13g2_fill_1 FILLER_66_1898 ();
 sg13g2_fill_2 FILLER_66_1903 ();
 sg13g2_decap_4 FILLER_66_1915 ();
 sg13g2_fill_1 FILLER_66_1919 ();
 sg13g2_fill_2 FILLER_66_1930 ();
 sg13g2_decap_4 FILLER_66_1940 ();
 sg13g2_fill_2 FILLER_66_1944 ();
 sg13g2_decap_4 FILLER_66_1956 ();
 sg13g2_fill_1 FILLER_66_1960 ();
 sg13g2_fill_1 FILLER_66_2005 ();
 sg13g2_fill_1 FILLER_66_2015 ();
 sg13g2_fill_1 FILLER_66_2026 ();
 sg13g2_decap_8 FILLER_66_2035 ();
 sg13g2_decap_4 FILLER_66_2063 ();
 sg13g2_fill_1 FILLER_66_2067 ();
 sg13g2_fill_1 FILLER_66_2092 ();
 sg13g2_fill_2 FILLER_66_2127 ();
 sg13g2_fill_1 FILLER_66_2129 ();
 sg13g2_decap_4 FILLER_66_2160 ();
 sg13g2_fill_1 FILLER_66_2164 ();
 sg13g2_decap_8 FILLER_66_2169 ();
 sg13g2_decap_8 FILLER_66_2176 ();
 sg13g2_decap_4 FILLER_66_2183 ();
 sg13g2_fill_2 FILLER_66_2187 ();
 sg13g2_fill_2 FILLER_66_2192 ();
 sg13g2_fill_1 FILLER_66_2199 ();
 sg13g2_decap_8 FILLER_66_2220 ();
 sg13g2_fill_2 FILLER_66_2227 ();
 sg13g2_fill_2 FILLER_66_2237 ();
 sg13g2_fill_1 FILLER_66_2239 ();
 sg13g2_fill_1 FILLER_66_2255 ();
 sg13g2_fill_2 FILLER_66_2265 ();
 sg13g2_fill_2 FILLER_66_2283 ();
 sg13g2_decap_8 FILLER_66_2310 ();
 sg13g2_fill_2 FILLER_66_2317 ();
 sg13g2_fill_1 FILLER_66_2319 ();
 sg13g2_decap_8 FILLER_66_2324 ();
 sg13g2_fill_1 FILLER_66_2331 ();
 sg13g2_fill_2 FILLER_66_2342 ();
 sg13g2_fill_2 FILLER_66_2367 ();
 sg13g2_fill_1 FILLER_66_2369 ();
 sg13g2_fill_1 FILLER_66_2375 ();
 sg13g2_fill_1 FILLER_66_2388 ();
 sg13g2_fill_2 FILLER_66_2394 ();
 sg13g2_fill_2 FILLER_66_2400 ();
 sg13g2_fill_1 FILLER_66_2402 ();
 sg13g2_fill_2 FILLER_66_2420 ();
 sg13g2_fill_2 FILLER_66_2444 ();
 sg13g2_decap_8 FILLER_66_2451 ();
 sg13g2_decap_8 FILLER_66_2458 ();
 sg13g2_fill_2 FILLER_66_2465 ();
 sg13g2_fill_1 FILLER_66_2467 ();
 sg13g2_fill_2 FILLER_66_2481 ();
 sg13g2_fill_1 FILLER_66_2483 ();
 sg13g2_fill_2 FILLER_66_2534 ();
 sg13g2_fill_2 FILLER_66_2540 ();
 sg13g2_fill_1 FILLER_66_2542 ();
 sg13g2_fill_1 FILLER_66_2547 ();
 sg13g2_decap_4 FILLER_66_2557 ();
 sg13g2_decap_8 FILLER_66_2587 ();
 sg13g2_fill_2 FILLER_66_2594 ();
 sg13g2_decap_4 FILLER_66_2609 ();
 sg13g2_fill_1 FILLER_66_2613 ();
 sg13g2_fill_1 FILLER_66_2627 ();
 sg13g2_fill_2 FILLER_66_2641 ();
 sg13g2_fill_1 FILLER_66_2643 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_4 FILLER_66_2656 ();
 sg13g2_fill_2 FILLER_66_2660 ();
 sg13g2_fill_2 FILLER_66_2667 ();
 sg13g2_decap_8 FILLER_66_2674 ();
 sg13g2_fill_1 FILLER_66_2681 ();
 sg13g2_decap_8 FILLER_66_2688 ();
 sg13g2_fill_2 FILLER_66_2695 ();
 sg13g2_decap_8 FILLER_66_2726 ();
 sg13g2_fill_1 FILLER_66_2733 ();
 sg13g2_fill_1 FILLER_66_2738 ();
 sg13g2_decap_8 FILLER_66_2748 ();
 sg13g2_fill_2 FILLER_66_2755 ();
 sg13g2_fill_1 FILLER_66_2757 ();
 sg13g2_decap_8 FILLER_66_2780 ();
 sg13g2_fill_1 FILLER_66_2787 ();
 sg13g2_fill_2 FILLER_66_2793 ();
 sg13g2_fill_2 FILLER_66_2800 ();
 sg13g2_fill_1 FILLER_66_2802 ();
 sg13g2_decap_8 FILLER_66_2819 ();
 sg13g2_fill_1 FILLER_66_2839 ();
 sg13g2_decap_4 FILLER_66_2844 ();
 sg13g2_fill_1 FILLER_66_2848 ();
 sg13g2_fill_2 FILLER_66_2863 ();
 sg13g2_fill_2 FILLER_66_2878 ();
 sg13g2_fill_1 FILLER_66_2880 ();
 sg13g2_fill_2 FILLER_66_2894 ();
 sg13g2_decap_4 FILLER_66_2907 ();
 sg13g2_fill_1 FILLER_66_2920 ();
 sg13g2_fill_1 FILLER_66_2934 ();
 sg13g2_decap_8 FILLER_66_2956 ();
 sg13g2_fill_2 FILLER_66_2963 ();
 sg13g2_fill_1 FILLER_66_2965 ();
 sg13g2_fill_2 FILLER_66_2974 ();
 sg13g2_decap_4 FILLER_66_2980 ();
 sg13g2_fill_1 FILLER_66_2984 ();
 sg13g2_fill_2 FILLER_66_2990 ();
 sg13g2_fill_2 FILLER_66_3027 ();
 sg13g2_decap_4 FILLER_66_3047 ();
 sg13g2_fill_2 FILLER_66_3051 ();
 sg13g2_decap_4 FILLER_66_3074 ();
 sg13g2_fill_1 FILLER_66_3078 ();
 sg13g2_fill_2 FILLER_66_3083 ();
 sg13g2_decap_8 FILLER_66_3090 ();
 sg13g2_decap_4 FILLER_66_3122 ();
 sg13g2_fill_2 FILLER_66_3126 ();
 sg13g2_decap_4 FILLER_66_3153 ();
 sg13g2_fill_1 FILLER_66_3157 ();
 sg13g2_fill_1 FILLER_66_3162 ();
 sg13g2_decap_8 FILLER_66_3179 ();
 sg13g2_decap_8 FILLER_66_3186 ();
 sg13g2_fill_2 FILLER_66_3193 ();
 sg13g2_decap_8 FILLER_66_3199 ();
 sg13g2_fill_2 FILLER_66_3206 ();
 sg13g2_fill_1 FILLER_66_3208 ();
 sg13g2_fill_1 FILLER_66_3236 ();
 sg13g2_decap_4 FILLER_66_3246 ();
 sg13g2_fill_2 FILLER_66_3250 ();
 sg13g2_decap_8 FILLER_66_3261 ();
 sg13g2_decap_4 FILLER_66_3268 ();
 sg13g2_fill_1 FILLER_66_3277 ();
 sg13g2_fill_2 FILLER_66_3287 ();
 sg13g2_decap_8 FILLER_66_3310 ();
 sg13g2_decap_8 FILLER_66_3317 ();
 sg13g2_fill_1 FILLER_66_3345 ();
 sg13g2_decap_8 FILLER_66_3373 ();
 sg13g2_decap_8 FILLER_66_3380 ();
 sg13g2_decap_8 FILLER_66_3387 ();
 sg13g2_decap_8 FILLER_66_3394 ();
 sg13g2_decap_8 FILLER_66_3401 ();
 sg13g2_decap_8 FILLER_66_3408 ();
 sg13g2_decap_8 FILLER_66_3415 ();
 sg13g2_decap_8 FILLER_66_3422 ();
 sg13g2_decap_8 FILLER_66_3429 ();
 sg13g2_decap_8 FILLER_66_3436 ();
 sg13g2_decap_8 FILLER_66_3443 ();
 sg13g2_decap_8 FILLER_66_3450 ();
 sg13g2_decap_8 FILLER_66_3457 ();
 sg13g2_decap_8 FILLER_66_3464 ();
 sg13g2_decap_8 FILLER_66_3471 ();
 sg13g2_decap_8 FILLER_66_3478 ();
 sg13g2_decap_8 FILLER_66_3485 ();
 sg13g2_decap_8 FILLER_66_3492 ();
 sg13g2_decap_8 FILLER_66_3499 ();
 sg13g2_decap_8 FILLER_66_3506 ();
 sg13g2_decap_8 FILLER_66_3513 ();
 sg13g2_decap_8 FILLER_66_3520 ();
 sg13g2_decap_8 FILLER_66_3527 ();
 sg13g2_decap_8 FILLER_66_3534 ();
 sg13g2_decap_8 FILLER_66_3541 ();
 sg13g2_decap_8 FILLER_66_3548 ();
 sg13g2_decap_8 FILLER_66_3555 ();
 sg13g2_decap_8 FILLER_66_3562 ();
 sg13g2_decap_8 FILLER_66_3569 ();
 sg13g2_decap_4 FILLER_66_3576 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_221 ();
 sg13g2_decap_4 FILLER_67_237 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_decap_4 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_309 ();
 sg13g2_decap_8 FILLER_67_348 ();
 sg13g2_decap_8 FILLER_67_355 ();
 sg13g2_fill_2 FILLER_67_362 ();
 sg13g2_decap_4 FILLER_67_368 ();
 sg13g2_fill_1 FILLER_67_372 ();
 sg13g2_fill_1 FILLER_67_392 ();
 sg13g2_fill_1 FILLER_67_397 ();
 sg13g2_fill_2 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_fill_2 FILLER_67_417 ();
 sg13g2_fill_1 FILLER_67_419 ();
 sg13g2_fill_1 FILLER_67_433 ();
 sg13g2_fill_2 FILLER_67_469 ();
 sg13g2_fill_2 FILLER_67_484 ();
 sg13g2_decap_4 FILLER_67_491 ();
 sg13g2_decap_4 FILLER_67_515 ();
 sg13g2_fill_1 FILLER_67_519 ();
 sg13g2_decap_4 FILLER_67_541 ();
 sg13g2_fill_2 FILLER_67_545 ();
 sg13g2_decap_4 FILLER_67_584 ();
 sg13g2_decap_4 FILLER_67_651 ();
 sg13g2_fill_2 FILLER_67_695 ();
 sg13g2_fill_1 FILLER_67_714 ();
 sg13g2_fill_2 FILLER_67_724 ();
 sg13g2_fill_1 FILLER_67_726 ();
 sg13g2_fill_1 FILLER_67_740 ();
 sg13g2_decap_8 FILLER_67_758 ();
 sg13g2_decap_8 FILLER_67_765 ();
 sg13g2_decap_8 FILLER_67_772 ();
 sg13g2_fill_1 FILLER_67_789 ();
 sg13g2_fill_1 FILLER_67_832 ();
 sg13g2_fill_2 FILLER_67_842 ();
 sg13g2_fill_2 FILLER_67_884 ();
 sg13g2_fill_1 FILLER_67_886 ();
 sg13g2_fill_2 FILLER_67_906 ();
 sg13g2_decap_8 FILLER_67_948 ();
 sg13g2_fill_2 FILLER_67_955 ();
 sg13g2_decap_4 FILLER_67_960 ();
 sg13g2_fill_2 FILLER_67_964 ();
 sg13g2_fill_2 FILLER_67_989 ();
 sg13g2_fill_1 FILLER_67_991 ();
 sg13g2_fill_2 FILLER_67_1042 ();
 sg13g2_fill_2 FILLER_67_1062 ();
 sg13g2_decap_8 FILLER_67_1101 ();
 sg13g2_decap_8 FILLER_67_1108 ();
 sg13g2_decap_4 FILLER_67_1115 ();
 sg13g2_fill_2 FILLER_67_1119 ();
 sg13g2_decap_8 FILLER_67_1131 ();
 sg13g2_fill_2 FILLER_67_1138 ();
 sg13g2_fill_1 FILLER_67_1140 ();
 sg13g2_fill_1 FILLER_67_1182 ();
 sg13g2_fill_1 FILLER_67_1211 ();
 sg13g2_decap_8 FILLER_67_1239 ();
 sg13g2_fill_1 FILLER_67_1246 ();
 sg13g2_fill_1 FILLER_67_1283 ();
 sg13g2_decap_4 FILLER_67_1297 ();
 sg13g2_decap_8 FILLER_67_1333 ();
 sg13g2_fill_1 FILLER_67_1340 ();
 sg13g2_fill_2 FILLER_67_1353 ();
 sg13g2_fill_1 FILLER_67_1355 ();
 sg13g2_decap_4 FILLER_67_1397 ();
 sg13g2_fill_2 FILLER_67_1401 ();
 sg13g2_decap_4 FILLER_67_1424 ();
 sg13g2_fill_1 FILLER_67_1428 ();
 sg13g2_decap_8 FILLER_67_1433 ();
 sg13g2_decap_8 FILLER_67_1440 ();
 sg13g2_decap_4 FILLER_67_1447 ();
 sg13g2_fill_2 FILLER_67_1455 ();
 sg13g2_decap_4 FILLER_67_1462 ();
 sg13g2_fill_1 FILLER_67_1466 ();
 sg13g2_fill_2 FILLER_67_1499 ();
 sg13g2_fill_2 FILLER_67_1545 ();
 sg13g2_decap_8 FILLER_67_1569 ();
 sg13g2_decap_8 FILLER_67_1603 ();
 sg13g2_fill_1 FILLER_67_1610 ();
 sg13g2_fill_2 FILLER_67_1616 ();
 sg13g2_fill_1 FILLER_67_1618 ();
 sg13g2_fill_2 FILLER_67_1637 ();
 sg13g2_fill_1 FILLER_67_1639 ();
 sg13g2_decap_4 FILLER_67_1662 ();
 sg13g2_decap_4 FILLER_67_1686 ();
 sg13g2_decap_4 FILLER_67_1722 ();
 sg13g2_fill_1 FILLER_67_1726 ();
 sg13g2_decap_8 FILLER_67_1732 ();
 sg13g2_fill_2 FILLER_67_1739 ();
 sg13g2_fill_1 FILLER_67_1741 ();
 sg13g2_fill_2 FILLER_67_1756 ();
 sg13g2_decap_4 FILLER_67_1808 ();
 sg13g2_fill_2 FILLER_67_1829 ();
 sg13g2_fill_1 FILLER_67_1831 ();
 sg13g2_decap_4 FILLER_67_1840 ();
 sg13g2_fill_2 FILLER_67_1844 ();
 sg13g2_decap_4 FILLER_67_1849 ();
 sg13g2_fill_1 FILLER_67_1853 ();
 sg13g2_decap_4 FILLER_67_1882 ();
 sg13g2_fill_2 FILLER_67_1901 ();
 sg13g2_fill_1 FILLER_67_1903 ();
 sg13g2_fill_2 FILLER_67_1914 ();
 sg13g2_decap_8 FILLER_67_1926 ();
 sg13g2_fill_2 FILLER_67_1933 ();
 sg13g2_fill_1 FILLER_67_1935 ();
 sg13g2_decap_8 FILLER_67_1954 ();
 sg13g2_decap_4 FILLER_67_1961 ();
 sg13g2_fill_1 FILLER_67_1965 ();
 sg13g2_decap_8 FILLER_67_1970 ();
 sg13g2_fill_1 FILLER_67_1977 ();
 sg13g2_fill_1 FILLER_67_2018 ();
 sg13g2_decap_8 FILLER_67_2041 ();
 sg13g2_decap_8 FILLER_67_2048 ();
 sg13g2_fill_1 FILLER_67_2055 ();
 sg13g2_decap_4 FILLER_67_2073 ();
 sg13g2_fill_2 FILLER_67_2083 ();
 sg13g2_fill_1 FILLER_67_2085 ();
 sg13g2_fill_2 FILLER_67_2094 ();
 sg13g2_fill_1 FILLER_67_2096 ();
 sg13g2_fill_1 FILLER_67_2102 ();
 sg13g2_fill_1 FILLER_67_2143 ();
 sg13g2_decap_8 FILLER_67_2181 ();
 sg13g2_decap_8 FILLER_67_2188 ();
 sg13g2_decap_4 FILLER_67_2195 ();
 sg13g2_fill_2 FILLER_67_2199 ();
 sg13g2_decap_8 FILLER_67_2215 ();
 sg13g2_fill_1 FILLER_67_2222 ();
 sg13g2_fill_2 FILLER_67_2249 ();
 sg13g2_fill_1 FILLER_67_2251 ();
 sg13g2_decap_8 FILLER_67_2256 ();
 sg13g2_decap_4 FILLER_67_2263 ();
 sg13g2_decap_8 FILLER_67_2276 ();
 sg13g2_decap_8 FILLER_67_2283 ();
 sg13g2_fill_2 FILLER_67_2290 ();
 sg13g2_decap_8 FILLER_67_2305 ();
 sg13g2_fill_2 FILLER_67_2312 ();
 sg13g2_fill_1 FILLER_67_2314 ();
 sg13g2_fill_2 FILLER_67_2343 ();
 sg13g2_decap_8 FILLER_67_2366 ();
 sg13g2_fill_2 FILLER_67_2373 ();
 sg13g2_decap_8 FILLER_67_2380 ();
 sg13g2_fill_2 FILLER_67_2387 ();
 sg13g2_decap_8 FILLER_67_2393 ();
 sg13g2_decap_4 FILLER_67_2400 ();
 sg13g2_fill_2 FILLER_67_2404 ();
 sg13g2_decap_8 FILLER_67_2412 ();
 sg13g2_decap_8 FILLER_67_2419 ();
 sg13g2_fill_2 FILLER_67_2435 ();
 sg13g2_fill_1 FILLER_67_2437 ();
 sg13g2_decap_8 FILLER_67_2442 ();
 sg13g2_decap_4 FILLER_67_2467 ();
 sg13g2_fill_2 FILLER_67_2471 ();
 sg13g2_fill_2 FILLER_67_2478 ();
 sg13g2_decap_8 FILLER_67_2499 ();
 sg13g2_fill_2 FILLER_67_2506 ();
 sg13g2_fill_1 FILLER_67_2508 ();
 sg13g2_decap_8 FILLER_67_2523 ();
 sg13g2_fill_1 FILLER_67_2530 ();
 sg13g2_fill_2 FILLER_67_2559 ();
 sg13g2_fill_1 FILLER_67_2561 ();
 sg13g2_fill_2 FILLER_67_2568 ();
 sg13g2_fill_2 FILLER_67_2587 ();
 sg13g2_fill_1 FILLER_67_2589 ();
 sg13g2_fill_2 FILLER_67_2597 ();
 sg13g2_fill_1 FILLER_67_2599 ();
 sg13g2_fill_2 FILLER_67_2613 ();
 sg13g2_fill_1 FILLER_67_2677 ();
 sg13g2_fill_2 FILLER_67_2694 ();
 sg13g2_fill_1 FILLER_67_2696 ();
 sg13g2_decap_8 FILLER_67_2772 ();
 sg13g2_decap_4 FILLER_67_2779 ();
 sg13g2_fill_2 FILLER_67_2787 ();
 sg13g2_fill_2 FILLER_67_2797 ();
 sg13g2_fill_1 FILLER_67_2799 ();
 sg13g2_decap_4 FILLER_67_2823 ();
 sg13g2_fill_2 FILLER_67_2841 ();
 sg13g2_fill_1 FILLER_67_2843 ();
 sg13g2_decap_4 FILLER_67_2886 ();
 sg13g2_fill_1 FILLER_67_2909 ();
 sg13g2_fill_2 FILLER_67_2932 ();
 sg13g2_fill_1 FILLER_67_2934 ();
 sg13g2_decap_8 FILLER_67_2951 ();
 sg13g2_fill_2 FILLER_67_2958 ();
 sg13g2_fill_1 FILLER_67_2960 ();
 sg13g2_decap_8 FILLER_67_2979 ();
 sg13g2_fill_2 FILLER_67_2986 ();
 sg13g2_fill_1 FILLER_67_2988 ();
 sg13g2_decap_8 FILLER_67_3000 ();
 sg13g2_fill_2 FILLER_67_3007 ();
 sg13g2_fill_1 FILLER_67_3009 ();
 sg13g2_decap_8 FILLER_67_3036 ();
 sg13g2_decap_8 FILLER_67_3043 ();
 sg13g2_decap_4 FILLER_67_3050 ();
 sg13g2_fill_1 FILLER_67_3064 ();
 sg13g2_fill_2 FILLER_67_3071 ();
 sg13g2_fill_1 FILLER_67_3073 ();
 sg13g2_fill_2 FILLER_67_3095 ();
 sg13g2_fill_1 FILLER_67_3102 ();
 sg13g2_fill_2 FILLER_67_3119 ();
 sg13g2_decap_8 FILLER_67_3136 ();
 sg13g2_decap_4 FILLER_67_3143 ();
 sg13g2_fill_1 FILLER_67_3147 ();
 sg13g2_fill_1 FILLER_67_3180 ();
 sg13g2_fill_2 FILLER_67_3209 ();
 sg13g2_decap_8 FILLER_67_3224 ();
 sg13g2_fill_2 FILLER_67_3231 ();
 sg13g2_decap_8 FILLER_67_3330 ();
 sg13g2_fill_1 FILLER_67_3337 ();
 sg13g2_decap_8 FILLER_67_3351 ();
 sg13g2_decap_8 FILLER_67_3358 ();
 sg13g2_decap_8 FILLER_67_3365 ();
 sg13g2_decap_8 FILLER_67_3372 ();
 sg13g2_decap_8 FILLER_67_3379 ();
 sg13g2_decap_8 FILLER_67_3386 ();
 sg13g2_decap_8 FILLER_67_3393 ();
 sg13g2_decap_8 FILLER_67_3400 ();
 sg13g2_decap_8 FILLER_67_3407 ();
 sg13g2_decap_8 FILLER_67_3414 ();
 sg13g2_decap_8 FILLER_67_3421 ();
 sg13g2_decap_8 FILLER_67_3428 ();
 sg13g2_decap_8 FILLER_67_3435 ();
 sg13g2_decap_8 FILLER_67_3442 ();
 sg13g2_decap_8 FILLER_67_3449 ();
 sg13g2_decap_8 FILLER_67_3456 ();
 sg13g2_decap_8 FILLER_67_3463 ();
 sg13g2_decap_8 FILLER_67_3470 ();
 sg13g2_decap_8 FILLER_67_3477 ();
 sg13g2_decap_8 FILLER_67_3484 ();
 sg13g2_decap_8 FILLER_67_3491 ();
 sg13g2_decap_8 FILLER_67_3498 ();
 sg13g2_decap_8 FILLER_67_3505 ();
 sg13g2_decap_8 FILLER_67_3512 ();
 sg13g2_decap_8 FILLER_67_3519 ();
 sg13g2_decap_8 FILLER_67_3526 ();
 sg13g2_decap_8 FILLER_67_3533 ();
 sg13g2_decap_8 FILLER_67_3540 ();
 sg13g2_decap_8 FILLER_67_3547 ();
 sg13g2_decap_8 FILLER_67_3554 ();
 sg13g2_decap_8 FILLER_67_3561 ();
 sg13g2_decap_8 FILLER_67_3568 ();
 sg13g2_decap_4 FILLER_67_3575 ();
 sg13g2_fill_1 FILLER_67_3579 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_176 ();
 sg13g2_fill_2 FILLER_68_191 ();
 sg13g2_decap_8 FILLER_68_232 ();
 sg13g2_decap_4 FILLER_68_239 ();
 sg13g2_decap_8 FILLER_68_247 ();
 sg13g2_decap_8 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_293 ();
 sg13g2_fill_2 FILLER_68_322 ();
 sg13g2_fill_1 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_415 ();
 sg13g2_decap_8 FILLER_68_471 ();
 sg13g2_fill_1 FILLER_68_488 ();
 sg13g2_decap_4 FILLER_68_495 ();
 sg13g2_fill_2 FILLER_68_499 ();
 sg13g2_decap_8 FILLER_68_521 ();
 sg13g2_fill_1 FILLER_68_528 ();
 sg13g2_decap_8 FILLER_68_533 ();
 sg13g2_decap_8 FILLER_68_540 ();
 sg13g2_decap_4 FILLER_68_547 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_fill_2 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_629 ();
 sg13g2_fill_1 FILLER_68_640 ();
 sg13g2_decap_4 FILLER_68_664 ();
 sg13g2_fill_2 FILLER_68_668 ();
 sg13g2_decap_4 FILLER_68_684 ();
 sg13g2_fill_2 FILLER_68_688 ();
 sg13g2_fill_2 FILLER_68_752 ();
 sg13g2_decap_4 FILLER_68_781 ();
 sg13g2_fill_1 FILLER_68_798 ();
 sg13g2_fill_1 FILLER_68_812 ();
 sg13g2_decap_4 FILLER_68_822 ();
 sg13g2_fill_1 FILLER_68_853 ();
 sg13g2_decap_8 FILLER_68_863 ();
 sg13g2_fill_2 FILLER_68_870 ();
 sg13g2_fill_1 FILLER_68_872 ();
 sg13g2_decap_4 FILLER_68_942 ();
 sg13g2_fill_2 FILLER_68_946 ();
 sg13g2_decap_8 FILLER_68_953 ();
 sg13g2_fill_2 FILLER_68_960 ();
 sg13g2_fill_2 FILLER_68_989 ();
 sg13g2_fill_1 FILLER_68_991 ();
 sg13g2_decap_8 FILLER_68_1019 ();
 sg13g2_decap_4 FILLER_68_1026 ();
 sg13g2_fill_2 FILLER_68_1030 ();
 sg13g2_fill_1 FILLER_68_1059 ();
 sg13g2_decap_4 FILLER_68_1070 ();
 sg13g2_fill_2 FILLER_68_1074 ();
 sg13g2_fill_1 FILLER_68_1143 ();
 sg13g2_fill_2 FILLER_68_1163 ();
 sg13g2_fill_2 FILLER_68_1192 ();
 sg13g2_fill_1 FILLER_68_1194 ();
 sg13g2_fill_1 FILLER_68_1223 ();
 sg13g2_decap_4 FILLER_68_1246 ();
 sg13g2_decap_4 FILLER_68_1282 ();
 sg13g2_fill_2 FILLER_68_1286 ();
 sg13g2_fill_1 FILLER_68_1305 ();
 sg13g2_fill_1 FILLER_68_1330 ();
 sg13g2_fill_2 FILLER_68_1344 ();
 sg13g2_fill_1 FILLER_68_1351 ();
 sg13g2_fill_1 FILLER_68_1369 ();
 sg13g2_fill_1 FILLER_68_1383 ();
 sg13g2_fill_2 FILLER_68_1410 ();
 sg13g2_fill_1 FILLER_68_1412 ();
 sg13g2_decap_4 FILLER_68_1440 ();
 sg13g2_fill_2 FILLER_68_1444 ();
 sg13g2_fill_2 FILLER_68_1506 ();
 sg13g2_fill_1 FILLER_68_1508 ();
 sg13g2_decap_8 FILLER_68_1551 ();
 sg13g2_decap_8 FILLER_68_1562 ();
 sg13g2_decap_8 FILLER_68_1569 ();
 sg13g2_fill_2 FILLER_68_1576 ();
 sg13g2_decap_8 FILLER_68_1594 ();
 sg13g2_fill_1 FILLER_68_1601 ();
 sg13g2_fill_2 FILLER_68_1630 ();
 sg13g2_decap_4 FILLER_68_1645 ();
 sg13g2_fill_1 FILLER_68_1649 ();
 sg13g2_fill_2 FILLER_68_1682 ();
 sg13g2_fill_1 FILLER_68_1684 ();
 sg13g2_fill_2 FILLER_68_1711 ();
 sg13g2_fill_2 FILLER_68_1740 ();
 sg13g2_fill_1 FILLER_68_1742 ();
 sg13g2_fill_2 FILLER_68_1776 ();
 sg13g2_decap_8 FILLER_68_1791 ();
 sg13g2_decap_8 FILLER_68_1798 ();
 sg13g2_fill_2 FILLER_68_1805 ();
 sg13g2_decap_8 FILLER_68_1835 ();
 sg13g2_fill_2 FILLER_68_1842 ();
 sg13g2_decap_8 FILLER_68_1848 ();
 sg13g2_decap_4 FILLER_68_1855 ();
 sg13g2_decap_8 FILLER_68_1863 ();
 sg13g2_fill_1 FILLER_68_1895 ();
 sg13g2_decap_8 FILLER_68_1912 ();
 sg13g2_fill_2 FILLER_68_1919 ();
 sg13g2_decap_8 FILLER_68_1939 ();
 sg13g2_decap_8 FILLER_68_1946 ();
 sg13g2_decap_8 FILLER_68_1953 ();
 sg13g2_fill_1 FILLER_68_1960 ();
 sg13g2_decap_8 FILLER_68_1974 ();
 sg13g2_fill_2 FILLER_68_1981 ();
 sg13g2_decap_4 FILLER_68_1987 ();
 sg13g2_fill_1 FILLER_68_1991 ();
 sg13g2_fill_1 FILLER_68_2045 ();
 sg13g2_fill_1 FILLER_68_2060 ();
 sg13g2_decap_8 FILLER_68_2073 ();
 sg13g2_decap_4 FILLER_68_2080 ();
 sg13g2_decap_8 FILLER_68_2099 ();
 sg13g2_decap_4 FILLER_68_2106 ();
 sg13g2_fill_1 FILLER_68_2110 ();
 sg13g2_fill_2 FILLER_68_2134 ();
 sg13g2_fill_2 FILLER_68_2191 ();
 sg13g2_decap_4 FILLER_68_2230 ();
 sg13g2_fill_2 FILLER_68_2242 ();
 sg13g2_fill_1 FILLER_68_2244 ();
 sg13g2_decap_8 FILLER_68_2250 ();
 sg13g2_decap_8 FILLER_68_2284 ();
 sg13g2_fill_1 FILLER_68_2291 ();
 sg13g2_fill_2 FILLER_68_2305 ();
 sg13g2_decap_8 FILLER_68_2312 ();
 sg13g2_fill_2 FILLER_68_2328 ();
 sg13g2_fill_1 FILLER_68_2330 ();
 sg13g2_decap_8 FILLER_68_2347 ();
 sg13g2_fill_1 FILLER_68_2354 ();
 sg13g2_fill_2 FILLER_68_2360 ();
 sg13g2_fill_2 FILLER_68_2373 ();
 sg13g2_decap_8 FILLER_68_2446 ();
 sg13g2_decap_4 FILLER_68_2453 ();
 sg13g2_fill_1 FILLER_68_2457 ();
 sg13g2_decap_4 FILLER_68_2462 ();
 sg13g2_fill_2 FILLER_68_2466 ();
 sg13g2_decap_8 FILLER_68_2473 ();
 sg13g2_decap_8 FILLER_68_2480 ();
 sg13g2_fill_2 FILLER_68_2487 ();
 sg13g2_fill_2 FILLER_68_2492 ();
 sg13g2_decap_8 FILLER_68_2504 ();
 sg13g2_fill_2 FILLER_68_2511 ();
 sg13g2_fill_2 FILLER_68_2525 ();
 sg13g2_fill_1 FILLER_68_2527 ();
 sg13g2_decap_8 FILLER_68_2532 ();
 sg13g2_decap_8 FILLER_68_2539 ();
 sg13g2_decap_8 FILLER_68_2546 ();
 sg13g2_fill_1 FILLER_68_2559 ();
 sg13g2_fill_2 FILLER_68_2565 ();
 sg13g2_decap_4 FILLER_68_2595 ();
 sg13g2_fill_1 FILLER_68_2599 ();
 sg13g2_fill_2 FILLER_68_2637 ();
 sg13g2_fill_1 FILLER_68_2639 ();
 sg13g2_decap_8 FILLER_68_2658 ();
 sg13g2_decap_4 FILLER_68_2665 ();
 sg13g2_fill_2 FILLER_68_2669 ();
 sg13g2_decap_4 FILLER_68_2689 ();
 sg13g2_decap_8 FILLER_68_2697 ();
 sg13g2_fill_2 FILLER_68_2704 ();
 sg13g2_decap_4 FILLER_68_2715 ();
 sg13g2_fill_1 FILLER_68_2719 ();
 sg13g2_decap_8 FILLER_68_2733 ();
 sg13g2_decap_4 FILLER_68_2740 ();
 sg13g2_decap_8 FILLER_68_2757 ();
 sg13g2_fill_2 FILLER_68_2764 ();
 sg13g2_fill_1 FILLER_68_2766 ();
 sg13g2_fill_2 FILLER_68_2771 ();
 sg13g2_fill_1 FILLER_68_2773 ();
 sg13g2_fill_2 FILLER_68_2806 ();
 sg13g2_decap_8 FILLER_68_2820 ();
 sg13g2_fill_1 FILLER_68_2827 ();
 sg13g2_decap_8 FILLER_68_2860 ();
 sg13g2_decap_8 FILLER_68_2867 ();
 sg13g2_decap_8 FILLER_68_2874 ();
 sg13g2_decap_8 FILLER_68_2881 ();
 sg13g2_fill_1 FILLER_68_2892 ();
 sg13g2_decap_8 FILLER_68_2898 ();
 sg13g2_decap_8 FILLER_68_2905 ();
 sg13g2_decap_4 FILLER_68_2921 ();
 sg13g2_fill_1 FILLER_68_2933 ();
 sg13g2_decap_8 FILLER_68_2942 ();
 sg13g2_decap_4 FILLER_68_2949 ();
 sg13g2_fill_2 FILLER_68_2953 ();
 sg13g2_decap_8 FILLER_68_2972 ();
 sg13g2_fill_2 FILLER_68_2979 ();
 sg13g2_fill_1 FILLER_68_2981 ();
 sg13g2_decap_4 FILLER_68_3005 ();
 sg13g2_decap_8 FILLER_68_3050 ();
 sg13g2_decap_4 FILLER_68_3063 ();
 sg13g2_fill_1 FILLER_68_3067 ();
 sg13g2_decap_8 FILLER_68_3073 ();
 sg13g2_decap_4 FILLER_68_3080 ();
 sg13g2_fill_2 FILLER_68_3084 ();
 sg13g2_fill_2 FILLER_68_3090 ();
 sg13g2_fill_1 FILLER_68_3092 ();
 sg13g2_decap_4 FILLER_68_3100 ();
 sg13g2_fill_1 FILLER_68_3104 ();
 sg13g2_decap_8 FILLER_68_3114 ();
 sg13g2_fill_1 FILLER_68_3121 ();
 sg13g2_fill_2 FILLER_68_3142 ();
 sg13g2_decap_4 FILLER_68_3154 ();
 sg13g2_decap_8 FILLER_68_3166 ();
 sg13g2_fill_1 FILLER_68_3173 ();
 sg13g2_decap_8 FILLER_68_3193 ();
 sg13g2_decap_8 FILLER_68_3200 ();
 sg13g2_decap_8 FILLER_68_3207 ();
 sg13g2_decap_8 FILLER_68_3214 ();
 sg13g2_decap_8 FILLER_68_3221 ();
 sg13g2_decap_8 FILLER_68_3228 ();
 sg13g2_fill_2 FILLER_68_3235 ();
 sg13g2_fill_1 FILLER_68_3237 ();
 sg13g2_decap_8 FILLER_68_3242 ();
 sg13g2_decap_8 FILLER_68_3249 ();
 sg13g2_decap_4 FILLER_68_3256 ();
 sg13g2_decap_8 FILLER_68_3264 ();
 sg13g2_decap_8 FILLER_68_3271 ();
 sg13g2_fill_2 FILLER_68_3278 ();
 sg13g2_decap_8 FILLER_68_3312 ();
 sg13g2_decap_8 FILLER_68_3319 ();
 sg13g2_decap_8 FILLER_68_3326 ();
 sg13g2_decap_4 FILLER_68_3333 ();
 sg13g2_fill_1 FILLER_68_3337 ();
 sg13g2_decap_8 FILLER_68_3351 ();
 sg13g2_decap_8 FILLER_68_3358 ();
 sg13g2_decap_8 FILLER_68_3365 ();
 sg13g2_decap_8 FILLER_68_3372 ();
 sg13g2_decap_8 FILLER_68_3379 ();
 sg13g2_decap_8 FILLER_68_3386 ();
 sg13g2_decap_8 FILLER_68_3393 ();
 sg13g2_decap_8 FILLER_68_3400 ();
 sg13g2_decap_8 FILLER_68_3407 ();
 sg13g2_decap_8 FILLER_68_3414 ();
 sg13g2_decap_8 FILLER_68_3421 ();
 sg13g2_decap_8 FILLER_68_3428 ();
 sg13g2_decap_8 FILLER_68_3435 ();
 sg13g2_decap_8 FILLER_68_3442 ();
 sg13g2_decap_8 FILLER_68_3449 ();
 sg13g2_decap_8 FILLER_68_3456 ();
 sg13g2_decap_8 FILLER_68_3463 ();
 sg13g2_decap_8 FILLER_68_3470 ();
 sg13g2_decap_8 FILLER_68_3477 ();
 sg13g2_decap_8 FILLER_68_3484 ();
 sg13g2_decap_8 FILLER_68_3491 ();
 sg13g2_decap_8 FILLER_68_3498 ();
 sg13g2_decap_8 FILLER_68_3505 ();
 sg13g2_decap_8 FILLER_68_3512 ();
 sg13g2_decap_8 FILLER_68_3519 ();
 sg13g2_decap_8 FILLER_68_3526 ();
 sg13g2_decap_8 FILLER_68_3533 ();
 sg13g2_decap_8 FILLER_68_3540 ();
 sg13g2_decap_8 FILLER_68_3547 ();
 sg13g2_decap_8 FILLER_68_3554 ();
 sg13g2_decap_8 FILLER_68_3561 ();
 sg13g2_decap_8 FILLER_68_3568 ();
 sg13g2_decap_4 FILLER_68_3575 ();
 sg13g2_fill_1 FILLER_68_3579 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_decap_4 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_decap_4 FILLER_69_295 ();
 sg13g2_fill_2 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_337 ();
 sg13g2_decap_4 FILLER_69_351 ();
 sg13g2_fill_1 FILLER_69_355 ();
 sg13g2_fill_1 FILLER_69_384 ();
 sg13g2_fill_1 FILLER_69_394 ();
 sg13g2_fill_2 FILLER_69_400 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_69_439 ();
 sg13g2_decap_8 FILLER_69_466 ();
 sg13g2_decap_4 FILLER_69_473 ();
 sg13g2_fill_2 FILLER_69_477 ();
 sg13g2_decap_8 FILLER_69_488 ();
 sg13g2_decap_4 FILLER_69_495 ();
 sg13g2_fill_1 FILLER_69_499 ();
 sg13g2_decap_4 FILLER_69_551 ();
 sg13g2_fill_2 FILLER_69_555 ();
 sg13g2_decap_4 FILLER_69_561 ();
 sg13g2_fill_2 FILLER_69_565 ();
 sg13g2_decap_4 FILLER_69_570 ();
 sg13g2_fill_1 FILLER_69_574 ();
 sg13g2_fill_1 FILLER_69_589 ();
 sg13g2_fill_2 FILLER_69_650 ();
 sg13g2_fill_1 FILLER_69_652 ();
 sg13g2_fill_1 FILLER_69_670 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_fill_1 FILLER_69_732 ();
 sg13g2_fill_2 FILLER_69_743 ();
 sg13g2_fill_1 FILLER_69_745 ();
 sg13g2_decap_8 FILLER_69_759 ();
 sg13g2_fill_2 FILLER_69_766 ();
 sg13g2_fill_1 FILLER_69_768 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_fill_2 FILLER_69_830 ();
 sg13g2_fill_1 FILLER_69_832 ();
 sg13g2_decap_8 FILLER_69_857 ();
 sg13g2_decap_8 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_69_884 ();
 sg13g2_fill_1 FILLER_69_891 ();
 sg13g2_decap_8 FILLER_69_897 ();
 sg13g2_fill_1 FILLER_69_904 ();
 sg13g2_decap_8 FILLER_69_943 ();
 sg13g2_fill_2 FILLER_69_950 ();
 sg13g2_fill_2 FILLER_69_978 ();
 sg13g2_fill_1 FILLER_69_993 ();
 sg13g2_decap_4 FILLER_69_997 ();
 sg13g2_decap_4 FILLER_69_1006 ();
 sg13g2_decap_4 FILLER_69_1038 ();
 sg13g2_decap_4 FILLER_69_1074 ();
 sg13g2_fill_2 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_fill_2 FILLER_69_1124 ();
 sg13g2_fill_1 FILLER_69_1126 ();
 sg13g2_fill_1 FILLER_69_1154 ();
 sg13g2_decap_4 FILLER_69_1234 ();
 sg13g2_fill_2 FILLER_69_1242 ();
 sg13g2_fill_2 FILLER_69_1249 ();
 sg13g2_decap_8 FILLER_69_1272 ();
 sg13g2_decap_8 FILLER_69_1279 ();
 sg13g2_fill_2 FILLER_69_1286 ();
 sg13g2_fill_2 FILLER_69_1356 ();
 sg13g2_fill_2 FILLER_69_1425 ();
 sg13g2_fill_1 FILLER_69_1427 ();
 sg13g2_decap_4 FILLER_69_1431 ();
 sg13g2_fill_2 FILLER_69_1444 ();
 sg13g2_fill_1 FILLER_69_1452 ();
 sg13g2_fill_2 FILLER_69_1459 ();
 sg13g2_fill_2 FILLER_69_1477 ();
 sg13g2_fill_2 FILLER_69_1488 ();
 sg13g2_fill_1 FILLER_69_1490 ();
 sg13g2_decap_8 FILLER_69_1500 ();
 sg13g2_decap_4 FILLER_69_1507 ();
 sg13g2_fill_2 FILLER_69_1511 ();
 sg13g2_fill_2 FILLER_69_1518 ();
 sg13g2_fill_2 FILLER_69_1551 ();
 sg13g2_fill_2 FILLER_69_1580 ();
 sg13g2_fill_2 FILLER_69_1591 ();
 sg13g2_fill_1 FILLER_69_1615 ();
 sg13g2_fill_1 FILLER_69_1629 ();
 sg13g2_decap_4 FILLER_69_1665 ();
 sg13g2_fill_2 FILLER_69_1669 ();
 sg13g2_fill_2 FILLER_69_1702 ();
 sg13g2_decap_8 FILLER_69_1730 ();
 sg13g2_fill_2 FILLER_69_1751 ();
 sg13g2_decap_4 FILLER_69_1757 ();
 sg13g2_decap_4 FILLER_69_1774 ();
 sg13g2_decap_4 FILLER_69_1801 ();
 sg13g2_fill_2 FILLER_69_1805 ();
 sg13g2_fill_2 FILLER_69_1811 ();
 sg13g2_fill_1 FILLER_69_1813 ();
 sg13g2_decap_8 FILLER_69_1828 ();
 sg13g2_fill_2 FILLER_69_1835 ();
 sg13g2_fill_1 FILLER_69_1837 ();
 sg13g2_decap_4 FILLER_69_1881 ();
 sg13g2_decap_8 FILLER_69_1908 ();
 sg13g2_fill_1 FILLER_69_1915 ();
 sg13g2_fill_2 FILLER_69_1933 ();
 sg13g2_decap_4 FILLER_69_1944 ();
 sg13g2_decap_8 FILLER_69_2040 ();
 sg13g2_decap_8 FILLER_69_2065 ();
 sg13g2_decap_8 FILLER_69_2072 ();
 sg13g2_decap_4 FILLER_69_2079 ();
 sg13g2_fill_1 FILLER_69_2083 ();
 sg13g2_decap_8 FILLER_69_2094 ();
 sg13g2_decap_8 FILLER_69_2101 ();
 sg13g2_fill_1 FILLER_69_2108 ();
 sg13g2_fill_2 FILLER_69_2114 ();
 sg13g2_fill_2 FILLER_69_2162 ();
 sg13g2_decap_8 FILLER_69_2177 ();
 sg13g2_decap_8 FILLER_69_2184 ();
 sg13g2_decap_4 FILLER_69_2191 ();
 sg13g2_decap_4 FILLER_69_2203 ();
 sg13g2_fill_1 FILLER_69_2207 ();
 sg13g2_decap_8 FILLER_69_2213 ();
 sg13g2_fill_2 FILLER_69_2220 ();
 sg13g2_fill_2 FILLER_69_2238 ();
 sg13g2_decap_8 FILLER_69_2277 ();
 sg13g2_decap_4 FILLER_69_2284 ();
 sg13g2_fill_1 FILLER_69_2288 ();
 sg13g2_decap_4 FILLER_69_2314 ();
 sg13g2_fill_2 FILLER_69_2318 ();
 sg13g2_fill_2 FILLER_69_2333 ();
 sg13g2_fill_1 FILLER_69_2335 ();
 sg13g2_fill_1 FILLER_69_2348 ();
 sg13g2_decap_4 FILLER_69_2354 ();
 sg13g2_fill_2 FILLER_69_2358 ();
 sg13g2_fill_2 FILLER_69_2365 ();
 sg13g2_decap_8 FILLER_69_2372 ();
 sg13g2_fill_2 FILLER_69_2379 ();
 sg13g2_fill_1 FILLER_69_2381 ();
 sg13g2_fill_2 FILLER_69_2387 ();
 sg13g2_fill_1 FILLER_69_2389 ();
 sg13g2_decap_4 FILLER_69_2395 ();
 sg13g2_fill_2 FILLER_69_2399 ();
 sg13g2_decap_4 FILLER_69_2411 ();
 sg13g2_fill_2 FILLER_69_2421 ();
 sg13g2_fill_1 FILLER_69_2423 ();
 sg13g2_fill_1 FILLER_69_2437 ();
 sg13g2_fill_2 FILLER_69_2444 ();
 sg13g2_decap_8 FILLER_69_2501 ();
 sg13g2_fill_2 FILLER_69_2508 ();
 sg13g2_fill_1 FILLER_69_2510 ();
 sg13g2_decap_4 FILLER_69_2558 ();
 sg13g2_fill_1 FILLER_69_2571 ();
 sg13g2_decap_8 FILLER_69_2576 ();
 sg13g2_fill_2 FILLER_69_2583 ();
 sg13g2_fill_1 FILLER_69_2585 ();
 sg13g2_decap_4 FILLER_69_2591 ();
 sg13g2_fill_1 FILLER_69_2595 ();
 sg13g2_decap_8 FILLER_69_2613 ();
 sg13g2_fill_2 FILLER_69_2620 ();
 sg13g2_fill_1 FILLER_69_2622 ();
 sg13g2_decap_4 FILLER_69_2670 ();
 sg13g2_fill_2 FILLER_69_2674 ();
 sg13g2_fill_2 FILLER_69_2686 ();
 sg13g2_decap_4 FILLER_69_2716 ();
 sg13g2_fill_2 FILLER_69_2720 ();
 sg13g2_fill_2 FILLER_69_2759 ();
 sg13g2_fill_1 FILLER_69_2761 ();
 sg13g2_decap_8 FILLER_69_2788 ();
 sg13g2_fill_2 FILLER_69_2844 ();
 sg13g2_fill_1 FILLER_69_2859 ();
 sg13g2_fill_1 FILLER_69_2888 ();
 sg13g2_decap_8 FILLER_69_2904 ();
 sg13g2_fill_2 FILLER_69_2911 ();
 sg13g2_decap_4 FILLER_69_2917 ();
 sg13g2_decap_8 FILLER_69_2934 ();
 sg13g2_fill_2 FILLER_69_2941 ();
 sg13g2_decap_4 FILLER_69_2956 ();
 sg13g2_fill_2 FILLER_69_2960 ();
 sg13g2_decap_8 FILLER_69_2973 ();
 sg13g2_fill_2 FILLER_69_2980 ();
 sg13g2_fill_2 FILLER_69_2987 ();
 sg13g2_decap_4 FILLER_69_2994 ();
 sg13g2_fill_2 FILLER_69_2998 ();
 sg13g2_decap_8 FILLER_69_3019 ();
 sg13g2_decap_8 FILLER_69_3026 ();
 sg13g2_fill_2 FILLER_69_3033 ();
 sg13g2_decap_8 FILLER_69_3039 ();
 sg13g2_decap_4 FILLER_69_3071 ();
 sg13g2_fill_2 FILLER_69_3075 ();
 sg13g2_decap_4 FILLER_69_3081 ();
 sg13g2_decap_8 FILLER_69_3105 ();
 sg13g2_fill_1 FILLER_69_3112 ();
 sg13g2_fill_2 FILLER_69_3117 ();
 sg13g2_decap_4 FILLER_69_3147 ();
 sg13g2_fill_2 FILLER_69_3151 ();
 sg13g2_fill_1 FILLER_69_3165 ();
 sg13g2_decap_8 FILLER_69_3201 ();
 sg13g2_decap_8 FILLER_69_3208 ();
 sg13g2_decap_8 FILLER_69_3215 ();
 sg13g2_decap_8 FILLER_69_3222 ();
 sg13g2_decap_8 FILLER_69_3229 ();
 sg13g2_decap_8 FILLER_69_3236 ();
 sg13g2_decap_8 FILLER_69_3243 ();
 sg13g2_decap_8 FILLER_69_3250 ();
 sg13g2_decap_8 FILLER_69_3257 ();
 sg13g2_decap_8 FILLER_69_3264 ();
 sg13g2_decap_8 FILLER_69_3271 ();
 sg13g2_decap_8 FILLER_69_3278 ();
 sg13g2_decap_8 FILLER_69_3292 ();
 sg13g2_decap_8 FILLER_69_3308 ();
 sg13g2_decap_8 FILLER_69_3315 ();
 sg13g2_decap_8 FILLER_69_3322 ();
 sg13g2_decap_8 FILLER_69_3329 ();
 sg13g2_decap_8 FILLER_69_3336 ();
 sg13g2_decap_8 FILLER_69_3343 ();
 sg13g2_decap_8 FILLER_69_3350 ();
 sg13g2_decap_8 FILLER_69_3357 ();
 sg13g2_decap_8 FILLER_69_3364 ();
 sg13g2_decap_8 FILLER_69_3371 ();
 sg13g2_decap_8 FILLER_69_3378 ();
 sg13g2_decap_8 FILLER_69_3385 ();
 sg13g2_decap_8 FILLER_69_3392 ();
 sg13g2_decap_8 FILLER_69_3399 ();
 sg13g2_decap_8 FILLER_69_3406 ();
 sg13g2_decap_8 FILLER_69_3413 ();
 sg13g2_decap_8 FILLER_69_3420 ();
 sg13g2_decap_8 FILLER_69_3427 ();
 sg13g2_decap_8 FILLER_69_3434 ();
 sg13g2_decap_8 FILLER_69_3441 ();
 sg13g2_decap_8 FILLER_69_3448 ();
 sg13g2_decap_8 FILLER_69_3455 ();
 sg13g2_decap_8 FILLER_69_3462 ();
 sg13g2_decap_8 FILLER_69_3469 ();
 sg13g2_decap_8 FILLER_69_3476 ();
 sg13g2_decap_8 FILLER_69_3483 ();
 sg13g2_decap_8 FILLER_69_3490 ();
 sg13g2_decap_8 FILLER_69_3497 ();
 sg13g2_decap_8 FILLER_69_3504 ();
 sg13g2_decap_8 FILLER_69_3511 ();
 sg13g2_decap_8 FILLER_69_3518 ();
 sg13g2_decap_8 FILLER_69_3525 ();
 sg13g2_decap_8 FILLER_69_3532 ();
 sg13g2_decap_8 FILLER_69_3539 ();
 sg13g2_decap_8 FILLER_69_3546 ();
 sg13g2_decap_8 FILLER_69_3553 ();
 sg13g2_decap_8 FILLER_69_3560 ();
 sg13g2_decap_8 FILLER_69_3567 ();
 sg13g2_decap_4 FILLER_69_3574 ();
 sg13g2_fill_2 FILLER_69_3578 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_2 FILLER_70_227 ();
 sg13g2_decap_8 FILLER_70_242 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_251 ();
 sg13g2_decap_8 FILLER_70_261 ();
 sg13g2_decap_8 FILLER_70_268 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_decap_4 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_424 ();
 sg13g2_fill_1 FILLER_70_431 ();
 sg13g2_fill_2 FILLER_70_437 ();
 sg13g2_decap_8 FILLER_70_463 ();
 sg13g2_fill_1 FILLER_70_470 ();
 sg13g2_fill_2 FILLER_70_503 ();
 sg13g2_decap_8 FILLER_70_527 ();
 sg13g2_decap_8 FILLER_70_534 ();
 sg13g2_fill_2 FILLER_70_541 ();
 sg13g2_decap_4 FILLER_70_547 ();
 sg13g2_fill_1 FILLER_70_551 ();
 sg13g2_fill_1 FILLER_70_580 ();
 sg13g2_fill_1 FILLER_70_597 ();
 sg13g2_fill_2 FILLER_70_626 ();
 sg13g2_fill_2 FILLER_70_633 ();
 sg13g2_decap_4 FILLER_70_644 ();
 sg13g2_fill_1 FILLER_70_648 ();
 sg13g2_decap_4 FILLER_70_682 ();
 sg13g2_decap_8 FILLER_70_692 ();
 sg13g2_fill_2 FILLER_70_699 ();
 sg13g2_fill_1 FILLER_70_701 ();
 sg13g2_fill_2 FILLER_70_706 ();
 sg13g2_fill_2 FILLER_70_738 ();
 sg13g2_fill_1 FILLER_70_740 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_784 ();
 sg13g2_decap_4 FILLER_70_830 ();
 sg13g2_decap_4 FILLER_70_867 ();
 sg13g2_fill_1 FILLER_70_902 ();
 sg13g2_decap_4 FILLER_70_906 ();
 sg13g2_fill_2 FILLER_70_910 ();
 sg13g2_fill_2 FILLER_70_916 ();
 sg13g2_fill_1 FILLER_70_918 ();
 sg13g2_fill_2 FILLER_70_932 ();
 sg13g2_decap_4 FILLER_70_968 ();
 sg13g2_fill_2 FILLER_70_1011 ();
 sg13g2_fill_1 FILLER_70_1013 ();
 sg13g2_fill_2 FILLER_70_1032 ();
 sg13g2_fill_2 FILLER_70_1043 ();
 sg13g2_fill_1 FILLER_70_1045 ();
 sg13g2_fill_2 FILLER_70_1054 ();
 sg13g2_fill_1 FILLER_70_1056 ();
 sg13g2_decap_4 FILLER_70_1063 ();
 sg13g2_decap_4 FILLER_70_1100 ();
 sg13g2_fill_2 FILLER_70_1104 ();
 sg13g2_decap_8 FILLER_70_1110 ();
 sg13g2_decap_4 FILLER_70_1117 ();
 sg13g2_fill_1 FILLER_70_1121 ();
 sg13g2_decap_8 FILLER_70_1127 ();
 sg13g2_decap_8 FILLER_70_1134 ();
 sg13g2_fill_1 FILLER_70_1141 ();
 sg13g2_decap_8 FILLER_70_1167 ();
 sg13g2_decap_4 FILLER_70_1174 ();
 sg13g2_fill_2 FILLER_70_1178 ();
 sg13g2_fill_2 FILLER_70_1188 ();
 sg13g2_fill_1 FILLER_70_1220 ();
 sg13g2_fill_1 FILLER_70_1244 ();
 sg13g2_fill_1 FILLER_70_1251 ();
 sg13g2_decap_8 FILLER_70_1289 ();
 sg13g2_decap_4 FILLER_70_1296 ();
 sg13g2_fill_1 FILLER_70_1322 ();
 sg13g2_decap_4 FILLER_70_1337 ();
 sg13g2_fill_2 FILLER_70_1341 ();
 sg13g2_decap_8 FILLER_70_1348 ();
 sg13g2_decap_8 FILLER_70_1355 ();
 sg13g2_decap_8 FILLER_70_1362 ();
 sg13g2_decap_8 FILLER_70_1369 ();
 sg13g2_fill_2 FILLER_70_1380 ();
 sg13g2_fill_1 FILLER_70_1410 ();
 sg13g2_fill_2 FILLER_70_1424 ();
 sg13g2_fill_2 FILLER_70_1435 ();
 sg13g2_fill_2 FILLER_70_1450 ();
 sg13g2_fill_1 FILLER_70_1460 ();
 sg13g2_fill_1 FILLER_70_1495 ();
 sg13g2_fill_2 FILLER_70_1513 ();
 sg13g2_decap_8 FILLER_70_1550 ();
 sg13g2_fill_2 FILLER_70_1557 ();
 sg13g2_fill_1 FILLER_70_1559 ();
 sg13g2_fill_1 FILLER_70_1566 ();
 sg13g2_decap_4 FILLER_70_1623 ();
 sg13g2_fill_1 FILLER_70_1627 ();
 sg13g2_fill_2 FILLER_70_1666 ();
 sg13g2_fill_1 FILLER_70_1673 ();
 sg13g2_fill_1 FILLER_70_1711 ();
 sg13g2_fill_1 FILLER_70_1740 ();
 sg13g2_fill_1 FILLER_70_1750 ();
 sg13g2_fill_2 FILLER_70_1762 ();
 sg13g2_fill_1 FILLER_70_1764 ();
 sg13g2_fill_2 FILLER_70_1778 ();
 sg13g2_fill_1 FILLER_70_1780 ();
 sg13g2_decap_4 FILLER_70_1791 ();
 sg13g2_fill_2 FILLER_70_1795 ();
 sg13g2_fill_1 FILLER_70_1801 ();
 sg13g2_decap_8 FILLER_70_1830 ();
 sg13g2_decap_8 FILLER_70_1837 ();
 sg13g2_decap_4 FILLER_70_1893 ();
 sg13g2_fill_1 FILLER_70_1897 ();
 sg13g2_decap_4 FILLER_70_1914 ();
 sg13g2_fill_2 FILLER_70_1918 ();
 sg13g2_fill_2 FILLER_70_1945 ();
 sg13g2_fill_2 FILLER_70_1994 ();
 sg13g2_fill_1 FILLER_70_1996 ();
 sg13g2_fill_1 FILLER_70_2006 ();
 sg13g2_fill_1 FILLER_70_2030 ();
 sg13g2_fill_2 FILLER_70_2034 ();
 sg13g2_fill_1 FILLER_70_2044 ();
 sg13g2_fill_1 FILLER_70_2055 ();
 sg13g2_decap_8 FILLER_70_2066 ();
 sg13g2_fill_2 FILLER_70_2073 ();
 sg13g2_decap_4 FILLER_70_2107 ();
 sg13g2_fill_2 FILLER_70_2124 ();
 sg13g2_fill_1 FILLER_70_2139 ();
 sg13g2_decap_8 FILLER_70_2144 ();
 sg13g2_fill_2 FILLER_70_2151 ();
 sg13g2_fill_1 FILLER_70_2153 ();
 sg13g2_fill_1 FILLER_70_2208 ();
 sg13g2_fill_2 FILLER_70_2215 ();
 sg13g2_fill_1 FILLER_70_2217 ();
 sg13g2_fill_2 FILLER_70_2228 ();
 sg13g2_decap_4 FILLER_70_2233 ();
 sg13g2_fill_1 FILLER_70_2237 ();
 sg13g2_fill_2 FILLER_70_2270 ();
 sg13g2_fill_1 FILLER_70_2272 ();
 sg13g2_decap_8 FILLER_70_2283 ();
 sg13g2_decap_8 FILLER_70_2290 ();
 sg13g2_fill_1 FILLER_70_2297 ();
 sg13g2_fill_2 FILLER_70_2311 ();
 sg13g2_decap_4 FILLER_70_2325 ();
 sg13g2_fill_2 FILLER_70_2329 ();
 sg13g2_fill_1 FILLER_70_2346 ();
 sg13g2_decap_4 FILLER_70_2356 ();
 sg13g2_decap_8 FILLER_70_2365 ();
 sg13g2_fill_2 FILLER_70_2385 ();
 sg13g2_fill_2 FILLER_70_2398 ();
 sg13g2_fill_1 FILLER_70_2400 ();
 sg13g2_fill_2 FILLER_70_2423 ();
 sg13g2_decap_4 FILLER_70_2467 ();
 sg13g2_fill_2 FILLER_70_2471 ();
 sg13g2_fill_2 FILLER_70_2482 ();
 sg13g2_decap_8 FILLER_70_2509 ();
 sg13g2_fill_2 FILLER_70_2516 ();
 sg13g2_decap_4 FILLER_70_2524 ();
 sg13g2_fill_1 FILLER_70_2538 ();
 sg13g2_fill_1 FILLER_70_2549 ();
 sg13g2_fill_2 FILLER_70_2555 ();
 sg13g2_fill_2 FILLER_70_2565 ();
 sg13g2_fill_1 FILLER_70_2567 ();
 sg13g2_fill_2 FILLER_70_2577 ();
 sg13g2_fill_1 FILLER_70_2579 ();
 sg13g2_decap_4 FILLER_70_2589 ();
 sg13g2_fill_2 FILLER_70_2593 ();
 sg13g2_decap_8 FILLER_70_2599 ();
 sg13g2_decap_4 FILLER_70_2606 ();
 sg13g2_fill_1 FILLER_70_2610 ();
 sg13g2_decap_4 FILLER_70_2616 ();
 sg13g2_fill_1 FILLER_70_2620 ();
 sg13g2_fill_1 FILLER_70_2626 ();
 sg13g2_decap_4 FILLER_70_2642 ();
 sg13g2_fill_2 FILLER_70_2646 ();
 sg13g2_fill_1 FILLER_70_2657 ();
 sg13g2_fill_2 FILLER_70_2684 ();
 sg13g2_fill_1 FILLER_70_2686 ();
 sg13g2_fill_1 FILLER_70_2696 ();
 sg13g2_fill_2 FILLER_70_2725 ();
 sg13g2_fill_2 FILLER_70_2745 ();
 sg13g2_fill_1 FILLER_70_2747 ();
 sg13g2_fill_1 FILLER_70_2769 ();
 sg13g2_fill_1 FILLER_70_2776 ();
 sg13g2_decap_4 FILLER_70_2803 ();
 sg13g2_fill_2 FILLER_70_2825 ();
 sg13g2_fill_2 FILLER_70_2832 ();
 sg13g2_decap_4 FILLER_70_2848 ();
 sg13g2_decap_8 FILLER_70_2869 ();
 sg13g2_decap_8 FILLER_70_2876 ();
 sg13g2_decap_4 FILLER_70_2912 ();
 sg13g2_fill_2 FILLER_70_2943 ();
 sg13g2_fill_1 FILLER_70_2945 ();
 sg13g2_fill_1 FILLER_70_2959 ();
 sg13g2_decap_4 FILLER_70_2969 ();
 sg13g2_fill_2 FILLER_70_2973 ();
 sg13g2_fill_2 FILLER_70_2987 ();
 sg13g2_decap_8 FILLER_70_3013 ();
 sg13g2_decap_8 FILLER_70_3020 ();
 sg13g2_decap_4 FILLER_70_3027 ();
 sg13g2_decap_4 FILLER_70_3047 ();
 sg13g2_fill_2 FILLER_70_3051 ();
 sg13g2_decap_4 FILLER_70_3063 ();
 sg13g2_decap_4 FILLER_70_3072 ();
 sg13g2_fill_1 FILLER_70_3076 ();
 sg13g2_decap_8 FILLER_70_3086 ();
 sg13g2_fill_2 FILLER_70_3093 ();
 sg13g2_fill_1 FILLER_70_3095 ();
 sg13g2_fill_2 FILLER_70_3117 ();
 sg13g2_fill_2 FILLER_70_3128 ();
 sg13g2_fill_1 FILLER_70_3130 ();
 sg13g2_decap_8 FILLER_70_3135 ();
 sg13g2_fill_2 FILLER_70_3142 ();
 sg13g2_decap_8 FILLER_70_3148 ();
 sg13g2_decap_8 FILLER_70_3155 ();
 sg13g2_decap_8 FILLER_70_3162 ();
 sg13g2_decap_4 FILLER_70_3169 ();
 sg13g2_fill_1 FILLER_70_3173 ();
 sg13g2_decap_8 FILLER_70_3205 ();
 sg13g2_decap_8 FILLER_70_3212 ();
 sg13g2_decap_8 FILLER_70_3219 ();
 sg13g2_decap_8 FILLER_70_3226 ();
 sg13g2_decap_8 FILLER_70_3233 ();
 sg13g2_decap_8 FILLER_70_3240 ();
 sg13g2_decap_8 FILLER_70_3247 ();
 sg13g2_decap_8 FILLER_70_3254 ();
 sg13g2_decap_8 FILLER_70_3261 ();
 sg13g2_decap_8 FILLER_70_3268 ();
 sg13g2_decap_8 FILLER_70_3275 ();
 sg13g2_decap_8 FILLER_70_3282 ();
 sg13g2_decap_8 FILLER_70_3289 ();
 sg13g2_decap_8 FILLER_70_3296 ();
 sg13g2_decap_8 FILLER_70_3303 ();
 sg13g2_decap_8 FILLER_70_3310 ();
 sg13g2_decap_8 FILLER_70_3317 ();
 sg13g2_decap_8 FILLER_70_3324 ();
 sg13g2_decap_8 FILLER_70_3331 ();
 sg13g2_decap_8 FILLER_70_3338 ();
 sg13g2_decap_8 FILLER_70_3345 ();
 sg13g2_decap_8 FILLER_70_3352 ();
 sg13g2_decap_8 FILLER_70_3359 ();
 sg13g2_decap_8 FILLER_70_3366 ();
 sg13g2_decap_8 FILLER_70_3373 ();
 sg13g2_decap_8 FILLER_70_3380 ();
 sg13g2_decap_8 FILLER_70_3387 ();
 sg13g2_decap_8 FILLER_70_3394 ();
 sg13g2_decap_8 FILLER_70_3401 ();
 sg13g2_decap_8 FILLER_70_3408 ();
 sg13g2_decap_8 FILLER_70_3415 ();
 sg13g2_decap_8 FILLER_70_3422 ();
 sg13g2_decap_8 FILLER_70_3429 ();
 sg13g2_decap_8 FILLER_70_3436 ();
 sg13g2_decap_8 FILLER_70_3443 ();
 sg13g2_decap_8 FILLER_70_3450 ();
 sg13g2_decap_8 FILLER_70_3457 ();
 sg13g2_decap_8 FILLER_70_3464 ();
 sg13g2_decap_8 FILLER_70_3471 ();
 sg13g2_decap_8 FILLER_70_3478 ();
 sg13g2_decap_8 FILLER_70_3485 ();
 sg13g2_decap_8 FILLER_70_3492 ();
 sg13g2_decap_8 FILLER_70_3499 ();
 sg13g2_decap_8 FILLER_70_3506 ();
 sg13g2_decap_8 FILLER_70_3513 ();
 sg13g2_decap_8 FILLER_70_3520 ();
 sg13g2_decap_8 FILLER_70_3527 ();
 sg13g2_decap_8 FILLER_70_3534 ();
 sg13g2_decap_8 FILLER_70_3541 ();
 sg13g2_decap_8 FILLER_70_3548 ();
 sg13g2_decap_8 FILLER_70_3555 ();
 sg13g2_decap_8 FILLER_70_3562 ();
 sg13g2_decap_8 FILLER_70_3569 ();
 sg13g2_decap_4 FILLER_70_3576 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_fill_2 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_265 ();
 sg13g2_decap_8 FILLER_71_272 ();
 sg13g2_decap_8 FILLER_71_279 ();
 sg13g2_fill_2 FILLER_71_286 ();
 sg13g2_fill_1 FILLER_71_301 ();
 sg13g2_fill_2 FILLER_71_310 ();
 sg13g2_fill_2 FILLER_71_338 ();
 sg13g2_decap_4 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_371 ();
 sg13g2_decap_4 FILLER_71_380 ();
 sg13g2_fill_1 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_419 ();
 sg13g2_fill_1 FILLER_71_421 ();
 sg13g2_fill_2 FILLER_71_438 ();
 sg13g2_decap_8 FILLER_71_459 ();
 sg13g2_decap_8 FILLER_71_466 ();
 sg13g2_fill_2 FILLER_71_473 ();
 sg13g2_fill_1 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_481 ();
 sg13g2_fill_1 FILLER_71_493 ();
 sg13g2_decap_4 FILLER_71_498 ();
 sg13g2_decap_8 FILLER_71_526 ();
 sg13g2_decap_4 FILLER_71_533 ();
 sg13g2_fill_1 FILLER_71_537 ();
 sg13g2_fill_1 FILLER_71_616 ();
 sg13g2_decap_8 FILLER_71_657 ();
 sg13g2_fill_2 FILLER_71_664 ();
 sg13g2_fill_2 FILLER_71_703 ();
 sg13g2_fill_1 FILLER_71_705 ();
 sg13g2_fill_1 FILLER_71_714 ();
 sg13g2_fill_2 FILLER_71_821 ();
 sg13g2_fill_1 FILLER_71_823 ();
 sg13g2_fill_1 FILLER_71_829 ();
 sg13g2_fill_2 FILLER_71_852 ();
 sg13g2_decap_8 FILLER_71_863 ();
 sg13g2_fill_1 FILLER_71_892 ();
 sg13g2_fill_2 FILLER_71_918 ();
 sg13g2_fill_2 FILLER_71_924 ();
 sg13g2_fill_1 FILLER_71_931 ();
 sg13g2_decap_4 FILLER_71_935 ();
 sg13g2_decap_8 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_959 ();
 sg13g2_decap_8 FILLER_71_966 ();
 sg13g2_decap_4 FILLER_71_973 ();
 sg13g2_fill_1 FILLER_71_981 ();
 sg13g2_fill_1 FILLER_71_996 ();
 sg13g2_fill_2 FILLER_71_1024 ();
 sg13g2_decap_4 FILLER_71_1055 ();
 sg13g2_decap_4 FILLER_71_1072 ();
 sg13g2_fill_1 FILLER_71_1076 ();
 sg13g2_decap_4 FILLER_71_1081 ();
 sg13g2_fill_2 FILLER_71_1094 ();
 sg13g2_fill_1 FILLER_71_1096 ();
 sg13g2_decap_4 FILLER_71_1129 ();
 sg13g2_fill_2 FILLER_71_1133 ();
 sg13g2_decap_8 FILLER_71_1169 ();
 sg13g2_fill_1 FILLER_71_1176 ();
 sg13g2_fill_1 FILLER_71_1236 ();
 sg13g2_fill_2 FILLER_71_1243 ();
 sg13g2_fill_1 FILLER_71_1245 ();
 sg13g2_fill_2 FILLER_71_1251 ();
 sg13g2_decap_4 FILLER_71_1264 ();
 sg13g2_fill_2 FILLER_71_1294 ();
 sg13g2_fill_1 FILLER_71_1296 ();
 sg13g2_fill_1 FILLER_71_1321 ();
 sg13g2_fill_1 FILLER_71_1326 ();
 sg13g2_decap_8 FILLER_71_1353 ();
 sg13g2_decap_4 FILLER_71_1360 ();
 sg13g2_fill_2 FILLER_71_1364 ();
 sg13g2_decap_4 FILLER_71_1390 ();
 sg13g2_fill_1 FILLER_71_1394 ();
 sg13g2_fill_1 FILLER_71_1415 ();
 sg13g2_fill_2 FILLER_71_1423 ();
 sg13g2_fill_1 FILLER_71_1438 ();
 sg13g2_decap_8 FILLER_71_1454 ();
 sg13g2_decap_8 FILLER_71_1464 ();
 sg13g2_fill_2 FILLER_71_1471 ();
 sg13g2_fill_1 FILLER_71_1473 ();
 sg13g2_decap_8 FILLER_71_1501 ();
 sg13g2_decap_4 FILLER_71_1508 ();
 sg13g2_decap_8 FILLER_71_1524 ();
 sg13g2_fill_2 FILLER_71_1531 ();
 sg13g2_decap_8 FILLER_71_1544 ();
 sg13g2_decap_8 FILLER_71_1551 ();
 sg13g2_fill_2 FILLER_71_1558 ();
 sg13g2_fill_1 FILLER_71_1560 ();
 sg13g2_fill_2 FILLER_71_1566 ();
 sg13g2_fill_2 FILLER_71_1577 ();
 sg13g2_fill_2 FILLER_71_1583 ();
 sg13g2_fill_1 FILLER_71_1600 ();
 sg13g2_fill_2 FILLER_71_1605 ();
 sg13g2_decap_8 FILLER_71_1625 ();
 sg13g2_decap_4 FILLER_71_1632 ();
 sg13g2_decap_4 FILLER_71_1673 ();
 sg13g2_fill_1 FILLER_71_1682 ();
 sg13g2_fill_1 FILLER_71_1692 ();
 sg13g2_decap_4 FILLER_71_1702 ();
 sg13g2_decap_8 FILLER_71_1714 ();
 sg13g2_decap_4 FILLER_71_1721 ();
 sg13g2_fill_1 FILLER_71_1725 ();
 sg13g2_decap_4 FILLER_71_1753 ();
 sg13g2_fill_1 FILLER_71_1757 ();
 sg13g2_fill_2 FILLER_71_1768 ();
 sg13g2_fill_1 FILLER_71_1770 ();
 sg13g2_fill_2 FILLER_71_1779 ();
 sg13g2_decap_8 FILLER_71_1797 ();
 sg13g2_decap_4 FILLER_71_1804 ();
 sg13g2_fill_2 FILLER_71_1808 ();
 sg13g2_fill_2 FILLER_71_1829 ();
 sg13g2_fill_1 FILLER_71_1831 ();
 sg13g2_fill_1 FILLER_71_1841 ();
 sg13g2_fill_2 FILLER_71_1847 ();
 sg13g2_fill_1 FILLER_71_1849 ();
 sg13g2_decap_4 FILLER_71_1854 ();
 sg13g2_fill_1 FILLER_71_1858 ();
 sg13g2_fill_2 FILLER_71_1887 ();
 sg13g2_decap_8 FILLER_71_1906 ();
 sg13g2_fill_2 FILLER_71_1913 ();
 sg13g2_fill_1 FILLER_71_1915 ();
 sg13g2_decap_8 FILLER_71_1939 ();
 sg13g2_fill_2 FILLER_71_1946 ();
 sg13g2_fill_1 FILLER_71_1948 ();
 sg13g2_fill_2 FILLER_71_1956 ();
 sg13g2_fill_1 FILLER_71_1958 ();
 sg13g2_decap_8 FILLER_71_1992 ();
 sg13g2_decap_8 FILLER_71_1999 ();
 sg13g2_fill_1 FILLER_71_2006 ();
 sg13g2_fill_2 FILLER_71_2015 ();
 sg13g2_fill_1 FILLER_71_2023 ();
 sg13g2_fill_1 FILLER_71_2029 ();
 sg13g2_fill_1 FILLER_71_2049 ();
 sg13g2_decap_8 FILLER_71_2062 ();
 sg13g2_decap_8 FILLER_71_2069 ();
 sg13g2_decap_8 FILLER_71_2076 ();
 sg13g2_fill_2 FILLER_71_2083 ();
 sg13g2_decap_8 FILLER_71_2121 ();
 sg13g2_fill_2 FILLER_71_2128 ();
 sg13g2_fill_1 FILLER_71_2130 ();
 sg13g2_decap_4 FILLER_71_2136 ();
 sg13g2_fill_1 FILLER_71_2148 ();
 sg13g2_decap_4 FILLER_71_2157 ();
 sg13g2_fill_1 FILLER_71_2161 ();
 sg13g2_fill_2 FILLER_71_2171 ();
 sg13g2_fill_2 FILLER_71_2190 ();
 sg13g2_decap_8 FILLER_71_2204 ();
 sg13g2_fill_2 FILLER_71_2211 ();
 sg13g2_decap_8 FILLER_71_2279 ();
 sg13g2_fill_1 FILLER_71_2286 ();
 sg13g2_fill_2 FILLER_71_2304 ();
 sg13g2_fill_2 FILLER_71_2311 ();
 sg13g2_fill_2 FILLER_71_2328 ();
 sg13g2_fill_1 FILLER_71_2330 ();
 sg13g2_decap_4 FILLER_71_2358 ();
 sg13g2_fill_2 FILLER_71_2362 ();
 sg13g2_decap_8 FILLER_71_2398 ();
 sg13g2_decap_4 FILLER_71_2405 ();
 sg13g2_decap_4 FILLER_71_2413 ();
 sg13g2_decap_8 FILLER_71_2458 ();
 sg13g2_fill_2 FILLER_71_2490 ();
 sg13g2_fill_1 FILLER_71_2492 ();
 sg13g2_decap_8 FILLER_71_2507 ();
 sg13g2_decap_8 FILLER_71_2514 ();
 sg13g2_decap_4 FILLER_71_2521 ();
 sg13g2_fill_2 FILLER_71_2525 ();
 sg13g2_decap_4 FILLER_71_2560 ();
 sg13g2_fill_2 FILLER_71_2564 ();
 sg13g2_fill_1 FILLER_71_2595 ();
 sg13g2_fill_1 FILLER_71_2606 ();
 sg13g2_decap_4 FILLER_71_2633 ();
 sg13g2_fill_1 FILLER_71_2637 ();
 sg13g2_decap_8 FILLER_71_2643 ();
 sg13g2_decap_8 FILLER_71_2666 ();
 sg13g2_fill_2 FILLER_71_2673 ();
 sg13g2_decap_8 FILLER_71_2689 ();
 sg13g2_decap_8 FILLER_71_2710 ();
 sg13g2_decap_8 FILLER_71_2717 ();
 sg13g2_decap_8 FILLER_71_2747 ();
 sg13g2_fill_2 FILLER_71_2754 ();
 sg13g2_fill_1 FILLER_71_2768 ();
 sg13g2_fill_2 FILLER_71_2800 ();
 sg13g2_fill_1 FILLER_71_2802 ();
 sg13g2_fill_2 FILLER_71_2822 ();
 sg13g2_fill_2 FILLER_71_2829 ();
 sg13g2_fill_1 FILLER_71_2831 ();
 sg13g2_decap_8 FILLER_71_2850 ();
 sg13g2_decap_8 FILLER_71_2861 ();
 sg13g2_decap_4 FILLER_71_2916 ();
 sg13g2_fill_2 FILLER_71_2944 ();
 sg13g2_fill_1 FILLER_71_2946 ();
 sg13g2_fill_1 FILLER_71_2951 ();
 sg13g2_fill_1 FILLER_71_2961 ();
 sg13g2_decap_4 FILLER_71_2971 ();
 sg13g2_fill_1 FILLER_71_2997 ();
 sg13g2_fill_1 FILLER_71_3023 ();
 sg13g2_fill_2 FILLER_71_3032 ();
 sg13g2_fill_2 FILLER_71_3050 ();
 sg13g2_fill_2 FILLER_71_3057 ();
 sg13g2_fill_1 FILLER_71_3059 ();
 sg13g2_fill_1 FILLER_71_3076 ();
 sg13g2_decap_4 FILLER_71_3090 ();
 sg13g2_fill_2 FILLER_71_3094 ();
 sg13g2_decap_8 FILLER_71_3100 ();
 sg13g2_fill_1 FILLER_71_3107 ();
 sg13g2_fill_2 FILLER_71_3136 ();
 sg13g2_fill_1 FILLER_71_3138 ();
 sg13g2_decap_4 FILLER_71_3176 ();
 sg13g2_fill_2 FILLER_71_3180 ();
 sg13g2_fill_2 FILLER_71_3186 ();
 sg13g2_fill_1 FILLER_71_3188 ();
 sg13g2_decap_8 FILLER_71_3202 ();
 sg13g2_decap_8 FILLER_71_3209 ();
 sg13g2_decap_8 FILLER_71_3216 ();
 sg13g2_decap_8 FILLER_71_3223 ();
 sg13g2_decap_8 FILLER_71_3230 ();
 sg13g2_decap_8 FILLER_71_3237 ();
 sg13g2_decap_8 FILLER_71_3244 ();
 sg13g2_decap_8 FILLER_71_3251 ();
 sg13g2_decap_8 FILLER_71_3258 ();
 sg13g2_decap_8 FILLER_71_3265 ();
 sg13g2_decap_8 FILLER_71_3272 ();
 sg13g2_decap_8 FILLER_71_3279 ();
 sg13g2_decap_8 FILLER_71_3286 ();
 sg13g2_decap_8 FILLER_71_3293 ();
 sg13g2_decap_8 FILLER_71_3300 ();
 sg13g2_decap_8 FILLER_71_3307 ();
 sg13g2_decap_8 FILLER_71_3314 ();
 sg13g2_decap_8 FILLER_71_3321 ();
 sg13g2_decap_8 FILLER_71_3328 ();
 sg13g2_decap_8 FILLER_71_3335 ();
 sg13g2_decap_8 FILLER_71_3342 ();
 sg13g2_decap_8 FILLER_71_3349 ();
 sg13g2_decap_8 FILLER_71_3356 ();
 sg13g2_decap_8 FILLER_71_3363 ();
 sg13g2_decap_8 FILLER_71_3370 ();
 sg13g2_decap_8 FILLER_71_3377 ();
 sg13g2_decap_8 FILLER_71_3384 ();
 sg13g2_decap_8 FILLER_71_3391 ();
 sg13g2_decap_8 FILLER_71_3398 ();
 sg13g2_decap_8 FILLER_71_3405 ();
 sg13g2_decap_8 FILLER_71_3412 ();
 sg13g2_decap_8 FILLER_71_3419 ();
 sg13g2_decap_8 FILLER_71_3426 ();
 sg13g2_decap_8 FILLER_71_3433 ();
 sg13g2_decap_8 FILLER_71_3440 ();
 sg13g2_decap_8 FILLER_71_3447 ();
 sg13g2_decap_8 FILLER_71_3454 ();
 sg13g2_decap_8 FILLER_71_3461 ();
 sg13g2_decap_8 FILLER_71_3468 ();
 sg13g2_decap_8 FILLER_71_3475 ();
 sg13g2_decap_8 FILLER_71_3482 ();
 sg13g2_decap_8 FILLER_71_3489 ();
 sg13g2_decap_8 FILLER_71_3496 ();
 sg13g2_decap_8 FILLER_71_3503 ();
 sg13g2_decap_8 FILLER_71_3510 ();
 sg13g2_decap_8 FILLER_71_3517 ();
 sg13g2_decap_8 FILLER_71_3524 ();
 sg13g2_decap_8 FILLER_71_3531 ();
 sg13g2_decap_8 FILLER_71_3538 ();
 sg13g2_decap_8 FILLER_71_3545 ();
 sg13g2_decap_8 FILLER_71_3552 ();
 sg13g2_decap_8 FILLER_71_3559 ();
 sg13g2_decap_8 FILLER_71_3566 ();
 sg13g2_decap_8 FILLER_71_3573 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_4 FILLER_72_182 ();
 sg13g2_fill_2 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_246 ();
 sg13g2_fill_1 FILLER_72_248 ();
 sg13g2_decap_8 FILLER_72_258 ();
 sg13g2_decap_8 FILLER_72_265 ();
 sg13g2_decap_8 FILLER_72_272 ();
 sg13g2_decap_8 FILLER_72_279 ();
 sg13g2_fill_2 FILLER_72_286 ();
 sg13g2_fill_1 FILLER_72_288 ();
 sg13g2_fill_2 FILLER_72_321 ();
 sg13g2_decap_4 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_fill_1 FILLER_72_434 ();
 sg13g2_decap_4 FILLER_72_450 ();
 sg13g2_decap_4 FILLER_72_458 ();
 sg13g2_fill_2 FILLER_72_462 ();
 sg13g2_fill_1 FILLER_72_490 ();
 sg13g2_decap_8 FILLER_72_496 ();
 sg13g2_fill_2 FILLER_72_507 ();
 sg13g2_fill_1 FILLER_72_509 ();
 sg13g2_fill_2 FILLER_72_518 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_fill_1 FILLER_72_538 ();
 sg13g2_decap_4 FILLER_72_576 ();
 sg13g2_fill_2 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_590 ();
 sg13g2_fill_2 FILLER_72_606 ();
 sg13g2_fill_1 FILLER_72_635 ();
 sg13g2_fill_2 FILLER_72_646 ();
 sg13g2_fill_1 FILLER_72_648 ();
 sg13g2_decap_4 FILLER_72_659 ();
 sg13g2_fill_1 FILLER_72_695 ();
 sg13g2_fill_1 FILLER_72_705 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_4 FILLER_72_725 ();
 sg13g2_fill_2 FILLER_72_729 ();
 sg13g2_fill_2 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_4 FILLER_72_780 ();
 sg13g2_fill_2 FILLER_72_784 ();
 sg13g2_fill_2 FILLER_72_802 ();
 sg13g2_fill_1 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_830 ();
 sg13g2_decap_4 FILLER_72_837 ();
 sg13g2_fill_1 FILLER_72_854 ();
 sg13g2_fill_2 FILLER_72_881 ();
 sg13g2_fill_1 FILLER_72_883 ();
 sg13g2_fill_1 FILLER_72_900 ();
 sg13g2_fill_2 FILLER_72_913 ();
 sg13g2_fill_1 FILLER_72_915 ();
 sg13g2_fill_2 FILLER_72_937 ();
 sg13g2_decap_8 FILLER_72_1019 ();
 sg13g2_decap_4 FILLER_72_1026 ();
 sg13g2_fill_2 FILLER_72_1049 ();
 sg13g2_decap_4 FILLER_72_1057 ();
 sg13g2_fill_2 FILLER_72_1061 ();
 sg13g2_decap_8 FILLER_72_1067 ();
 sg13g2_decap_8 FILLER_72_1074 ();
 sg13g2_decap_4 FILLER_72_1081 ();
 sg13g2_decap_8 FILLER_72_1162 ();
 sg13g2_decap_8 FILLER_72_1169 ();
 sg13g2_fill_2 FILLER_72_1176 ();
 sg13g2_fill_2 FILLER_72_1186 ();
 sg13g2_fill_2 FILLER_72_1202 ();
 sg13g2_fill_1 FILLER_72_1222 ();
 sg13g2_fill_2 FILLER_72_1238 ();
 sg13g2_fill_1 FILLER_72_1240 ();
 sg13g2_decap_8 FILLER_72_1245 ();
 sg13g2_decap_8 FILLER_72_1257 ();
 sg13g2_decap_4 FILLER_72_1264 ();
 sg13g2_decap_8 FILLER_72_1287 ();
 sg13g2_decap_8 FILLER_72_1294 ();
 sg13g2_fill_2 FILLER_72_1301 ();
 sg13g2_decap_4 FILLER_72_1330 ();
 sg13g2_fill_1 FILLER_72_1334 ();
 sg13g2_decap_8 FILLER_72_1356 ();
 sg13g2_fill_2 FILLER_72_1404 ();
 sg13g2_fill_2 FILLER_72_1429 ();
 sg13g2_fill_2 FILLER_72_1446 ();
 sg13g2_decap_4 FILLER_72_1466 ();
 sg13g2_fill_1 FILLER_72_1470 ();
 sg13g2_fill_1 FILLER_72_1480 ();
 sg13g2_fill_1 FILLER_72_1499 ();
 sg13g2_decap_8 FILLER_72_1504 ();
 sg13g2_fill_2 FILLER_72_1524 ();
 sg13g2_fill_2 FILLER_72_1530 ();
 sg13g2_fill_1 FILLER_72_1532 ();
 sg13g2_fill_1 FILLER_72_1557 ();
 sg13g2_fill_1 FILLER_72_1564 ();
 sg13g2_decap_8 FILLER_72_1579 ();
 sg13g2_decap_4 FILLER_72_1586 ();
 sg13g2_fill_1 FILLER_72_1590 ();
 sg13g2_fill_1 FILLER_72_1599 ();
 sg13g2_decap_8 FILLER_72_1604 ();
 sg13g2_fill_1 FILLER_72_1611 ();
 sg13g2_decap_8 FILLER_72_1621 ();
 sg13g2_decap_8 FILLER_72_1628 ();
 sg13g2_decap_4 FILLER_72_1635 ();
 sg13g2_fill_2 FILLER_72_1639 ();
 sg13g2_fill_1 FILLER_72_1672 ();
 sg13g2_fill_1 FILLER_72_1696 ();
 sg13g2_fill_1 FILLER_72_1700 ();
 sg13g2_decap_4 FILLER_72_1707 ();
 sg13g2_fill_2 FILLER_72_1711 ();
 sg13g2_decap_8 FILLER_72_1722 ();
 sg13g2_fill_1 FILLER_72_1729 ();
 sg13g2_decap_8 FILLER_72_1735 ();
 sg13g2_decap_4 FILLER_72_1742 ();
 sg13g2_fill_1 FILLER_72_1746 ();
 sg13g2_fill_2 FILLER_72_1759 ();
 sg13g2_decap_8 FILLER_72_1766 ();
 sg13g2_decap_4 FILLER_72_1773 ();
 sg13g2_fill_2 FILLER_72_1781 ();
 sg13g2_fill_1 FILLER_72_1783 ();
 sg13g2_decap_4 FILLER_72_1788 ();
 sg13g2_fill_1 FILLER_72_1792 ();
 sg13g2_decap_8 FILLER_72_1802 ();
 sg13g2_decap_8 FILLER_72_1827 ();
 sg13g2_fill_2 FILLER_72_1834 ();
 sg13g2_fill_2 FILLER_72_1853 ();
 sg13g2_fill_1 FILLER_72_1892 ();
 sg13g2_decap_8 FILLER_72_1908 ();
 sg13g2_decap_4 FILLER_72_1915 ();
 sg13g2_fill_1 FILLER_72_1919 ();
 sg13g2_fill_1 FILLER_72_1935 ();
 sg13g2_decap_8 FILLER_72_1944 ();
 sg13g2_fill_2 FILLER_72_1951 ();
 sg13g2_fill_1 FILLER_72_1953 ();
 sg13g2_fill_2 FILLER_72_1987 ();
 sg13g2_fill_1 FILLER_72_1994 ();
 sg13g2_decap_8 FILLER_72_2010 ();
 sg13g2_decap_8 FILLER_72_2022 ();
 sg13g2_decap_8 FILLER_72_2029 ();
 sg13g2_decap_8 FILLER_72_2046 ();
 sg13g2_decap_8 FILLER_72_2053 ();
 sg13g2_fill_1 FILLER_72_2093 ();
 sg13g2_fill_2 FILLER_72_2124 ();
 sg13g2_decap_4 FILLER_72_2148 ();
 sg13g2_fill_1 FILLER_72_2152 ();
 sg13g2_fill_1 FILLER_72_2165 ();
 sg13g2_decap_8 FILLER_72_2181 ();
 sg13g2_decap_8 FILLER_72_2203 ();
 sg13g2_decap_8 FILLER_72_2210 ();
 sg13g2_fill_2 FILLER_72_2217 ();
 sg13g2_decap_8 FILLER_72_2223 ();
 sg13g2_decap_8 FILLER_72_2230 ();
 sg13g2_decap_4 FILLER_72_2237 ();
 sg13g2_fill_1 FILLER_72_2297 ();
 sg13g2_fill_1 FILLER_72_2314 ();
 sg13g2_decap_4 FILLER_72_2324 ();
 sg13g2_fill_1 FILLER_72_2328 ();
 sg13g2_decap_8 FILLER_72_2334 ();
 sg13g2_decap_8 FILLER_72_2358 ();
 sg13g2_fill_1 FILLER_72_2377 ();
 sg13g2_decap_8 FILLER_72_2386 ();
 sg13g2_decap_8 FILLER_72_2393 ();
 sg13g2_decap_4 FILLER_72_2400 ();
 sg13g2_decap_8 FILLER_72_2460 ();
 sg13g2_fill_2 FILLER_72_2467 ();
 sg13g2_fill_1 FILLER_72_2469 ();
 sg13g2_fill_1 FILLER_72_2502 ();
 sg13g2_decap_8 FILLER_72_2553 ();
 sg13g2_decap_8 FILLER_72_2560 ();
 sg13g2_fill_2 FILLER_72_2567 ();
 sg13g2_fill_1 FILLER_72_2569 ();
 sg13g2_fill_2 FILLER_72_2573 ();
 sg13g2_fill_1 FILLER_72_2575 ();
 sg13g2_fill_2 FILLER_72_2581 ();
 sg13g2_fill_1 FILLER_72_2583 ();
 sg13g2_decap_8 FILLER_72_2602 ();
 sg13g2_decap_8 FILLER_72_2609 ();
 sg13g2_decap_4 FILLER_72_2616 ();
 sg13g2_fill_1 FILLER_72_2620 ();
 sg13g2_decap_4 FILLER_72_2630 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_fill_2 FILLER_72_2673 ();
 sg13g2_fill_1 FILLER_72_2685 ();
 sg13g2_fill_2 FILLER_72_2693 ();
 sg13g2_fill_1 FILLER_72_2695 ();
 sg13g2_decap_4 FILLER_72_2714 ();
 sg13g2_fill_1 FILLER_72_2718 ();
 sg13g2_fill_2 FILLER_72_2740 ();
 sg13g2_fill_1 FILLER_72_2742 ();
 sg13g2_decap_8 FILLER_72_2750 ();
 sg13g2_decap_8 FILLER_72_2757 ();
 sg13g2_decap_4 FILLER_72_2764 ();
 sg13g2_fill_1 FILLER_72_2768 ();
 sg13g2_fill_1 FILLER_72_2778 ();
 sg13g2_decap_4 FILLER_72_2794 ();
 sg13g2_fill_1 FILLER_72_2854 ();
 sg13g2_decap_8 FILLER_72_2879 ();
 sg13g2_decap_8 FILLER_72_2886 ();
 sg13g2_decap_4 FILLER_72_2893 ();
 sg13g2_fill_1 FILLER_72_2903 ();
 sg13g2_fill_1 FILLER_72_2916 ();
 sg13g2_fill_2 FILLER_72_2928 ();
 sg13g2_fill_1 FILLER_72_2930 ();
 sg13g2_decap_4 FILLER_72_2935 ();
 sg13g2_decap_8 FILLER_72_2942 ();
 sg13g2_decap_8 FILLER_72_2949 ();
 sg13g2_decap_8 FILLER_72_2956 ();
 sg13g2_fill_1 FILLER_72_2979 ();
 sg13g2_decap_8 FILLER_72_3004 ();
 sg13g2_decap_4 FILLER_72_3011 ();
 sg13g2_fill_2 FILLER_72_3015 ();
 sg13g2_fill_2 FILLER_72_3022 ();
 sg13g2_decap_8 FILLER_72_3028 ();
 sg13g2_fill_2 FILLER_72_3035 ();
 sg13g2_fill_1 FILLER_72_3037 ();
 sg13g2_decap_8 FILLER_72_3050 ();
 sg13g2_fill_2 FILLER_72_3057 ();
 sg13g2_decap_4 FILLER_72_3073 ();
 sg13g2_fill_1 FILLER_72_3077 ();
 sg13g2_fill_2 FILLER_72_3082 ();
 sg13g2_fill_1 FILLER_72_3090 ();
 sg13g2_decap_8 FILLER_72_3119 ();
 sg13g2_decap_8 FILLER_72_3126 ();
 sg13g2_decap_8 FILLER_72_3133 ();
 sg13g2_decap_8 FILLER_72_3140 ();
 sg13g2_decap_8 FILLER_72_3147 ();
 sg13g2_decap_8 FILLER_72_3154 ();
 sg13g2_decap_8 FILLER_72_3161 ();
 sg13g2_decap_8 FILLER_72_3168 ();
 sg13g2_decap_8 FILLER_72_3175 ();
 sg13g2_decap_8 FILLER_72_3182 ();
 sg13g2_decap_8 FILLER_72_3198 ();
 sg13g2_decap_8 FILLER_72_3205 ();
 sg13g2_decap_8 FILLER_72_3212 ();
 sg13g2_decap_8 FILLER_72_3219 ();
 sg13g2_decap_8 FILLER_72_3226 ();
 sg13g2_decap_8 FILLER_72_3233 ();
 sg13g2_decap_8 FILLER_72_3240 ();
 sg13g2_decap_8 FILLER_72_3247 ();
 sg13g2_decap_8 FILLER_72_3254 ();
 sg13g2_decap_8 FILLER_72_3261 ();
 sg13g2_decap_8 FILLER_72_3268 ();
 sg13g2_decap_8 FILLER_72_3275 ();
 sg13g2_decap_8 FILLER_72_3282 ();
 sg13g2_decap_8 FILLER_72_3289 ();
 sg13g2_decap_8 FILLER_72_3296 ();
 sg13g2_decap_8 FILLER_72_3303 ();
 sg13g2_decap_8 FILLER_72_3310 ();
 sg13g2_decap_8 FILLER_72_3317 ();
 sg13g2_decap_8 FILLER_72_3324 ();
 sg13g2_decap_8 FILLER_72_3331 ();
 sg13g2_decap_8 FILLER_72_3338 ();
 sg13g2_decap_8 FILLER_72_3345 ();
 sg13g2_decap_8 FILLER_72_3352 ();
 sg13g2_decap_8 FILLER_72_3359 ();
 sg13g2_decap_8 FILLER_72_3366 ();
 sg13g2_decap_8 FILLER_72_3373 ();
 sg13g2_decap_8 FILLER_72_3380 ();
 sg13g2_decap_8 FILLER_72_3387 ();
 sg13g2_decap_8 FILLER_72_3394 ();
 sg13g2_decap_8 FILLER_72_3401 ();
 sg13g2_decap_8 FILLER_72_3408 ();
 sg13g2_decap_8 FILLER_72_3415 ();
 sg13g2_decap_8 FILLER_72_3422 ();
 sg13g2_decap_8 FILLER_72_3429 ();
 sg13g2_decap_8 FILLER_72_3436 ();
 sg13g2_decap_8 FILLER_72_3443 ();
 sg13g2_decap_8 FILLER_72_3450 ();
 sg13g2_decap_8 FILLER_72_3457 ();
 sg13g2_decap_8 FILLER_72_3464 ();
 sg13g2_decap_8 FILLER_72_3471 ();
 sg13g2_decap_8 FILLER_72_3478 ();
 sg13g2_decap_8 FILLER_72_3485 ();
 sg13g2_decap_8 FILLER_72_3492 ();
 sg13g2_decap_8 FILLER_72_3499 ();
 sg13g2_decap_8 FILLER_72_3506 ();
 sg13g2_decap_8 FILLER_72_3513 ();
 sg13g2_decap_8 FILLER_72_3520 ();
 sg13g2_decap_8 FILLER_72_3527 ();
 sg13g2_decap_8 FILLER_72_3534 ();
 sg13g2_decap_8 FILLER_72_3541 ();
 sg13g2_decap_8 FILLER_72_3548 ();
 sg13g2_decap_8 FILLER_72_3555 ();
 sg13g2_decap_8 FILLER_72_3562 ();
 sg13g2_decap_8 FILLER_72_3569 ();
 sg13g2_decap_4 FILLER_72_3576 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_4 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_214 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_2 FILLER_73_229 ();
 sg13g2_decap_8 FILLER_73_240 ();
 sg13g2_decap_8 FILLER_73_247 ();
 sg13g2_decap_8 FILLER_73_254 ();
 sg13g2_decap_8 FILLER_73_261 ();
 sg13g2_decap_8 FILLER_73_268 ();
 sg13g2_decap_8 FILLER_73_275 ();
 sg13g2_decap_8 FILLER_73_282 ();
 sg13g2_decap_8 FILLER_73_289 ();
 sg13g2_fill_2 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_319 ();
 sg13g2_fill_1 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_fill_2 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_379 ();
 sg13g2_fill_2 FILLER_73_386 ();
 sg13g2_fill_1 FILLER_73_388 ();
 sg13g2_decap_4 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_73_431 ();
 sg13g2_decap_4 FILLER_73_444 ();
 sg13g2_fill_1 FILLER_73_448 ();
 sg13g2_fill_1 FILLER_73_506 ();
 sg13g2_fill_1 FILLER_73_522 ();
 sg13g2_decap_8 FILLER_73_528 ();
 sg13g2_decap_8 FILLER_73_535 ();
 sg13g2_fill_2 FILLER_73_574 ();
 sg13g2_fill_1 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_fill_2 FILLER_73_616 ();
 sg13g2_fill_1 FILLER_73_618 ();
 sg13g2_decap_4 FILLER_73_623 ();
 sg13g2_fill_2 FILLER_73_636 ();
 sg13g2_decap_8 FILLER_73_660 ();
 sg13g2_decap_8 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_674 ();
 sg13g2_fill_2 FILLER_73_691 ();
 sg13g2_decap_4 FILLER_73_697 ();
 sg13g2_fill_2 FILLER_73_701 ();
 sg13g2_fill_1 FILLER_73_717 ();
 sg13g2_decap_4 FILLER_73_722 ();
 sg13g2_fill_1 FILLER_73_726 ();
 sg13g2_decap_4 FILLER_73_749 ();
 sg13g2_fill_2 FILLER_73_758 ();
 sg13g2_fill_1 FILLER_73_808 ();
 sg13g2_fill_2 FILLER_73_814 ();
 sg13g2_decap_4 FILLER_73_825 ();
 sg13g2_fill_2 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_856 ();
 sg13g2_decap_8 FILLER_73_863 ();
 sg13g2_fill_1 FILLER_73_900 ();
 sg13g2_decap_8 FILLER_73_906 ();
 sg13g2_fill_2 FILLER_73_913 ();
 sg13g2_fill_1 FILLER_73_915 ();
 sg13g2_fill_2 FILLER_73_924 ();
 sg13g2_fill_1 FILLER_73_926 ();
 sg13g2_decap_4 FILLER_73_931 ();
 sg13g2_fill_2 FILLER_73_940 ();
 sg13g2_decap_8 FILLER_73_960 ();
 sg13g2_fill_1 FILLER_73_967 ();
 sg13g2_decap_4 FILLER_73_972 ();
 sg13g2_decap_8 FILLER_73_980 ();
 sg13g2_decap_4 FILLER_73_987 ();
 sg13g2_decap_4 FILLER_73_1005 ();
 sg13g2_decap_8 FILLER_73_1024 ();
 sg13g2_fill_2 FILLER_73_1117 ();
 sg13g2_fill_1 FILLER_73_1119 ();
 sg13g2_fill_2 FILLER_73_1191 ();
 sg13g2_fill_1 FILLER_73_1202 ();
 sg13g2_fill_1 FILLER_73_1219 ();
 sg13g2_decap_8 FILLER_73_1235 ();
 sg13g2_decap_4 FILLER_73_1242 ();
 sg13g2_fill_2 FILLER_73_1246 ();
 sg13g2_fill_1 FILLER_73_1267 ();
 sg13g2_fill_1 FILLER_73_1276 ();
 sg13g2_fill_1 FILLER_73_1282 ();
 sg13g2_fill_1 FILLER_73_1289 ();
 sg13g2_fill_1 FILLER_73_1307 ();
 sg13g2_decap_8 FILLER_73_1317 ();
 sg13g2_fill_1 FILLER_73_1345 ();
 sg13g2_fill_1 FILLER_73_1358 ();
 sg13g2_decap_8 FILLER_73_1381 ();
 sg13g2_fill_2 FILLER_73_1388 ();
 sg13g2_fill_1 FILLER_73_1399 ();
 sg13g2_decap_8 FILLER_73_1413 ();
 sg13g2_decap_4 FILLER_73_1420 ();
 sg13g2_fill_1 FILLER_73_1424 ();
 sg13g2_decap_8 FILLER_73_1514 ();
 sg13g2_fill_2 FILLER_73_1564 ();
 sg13g2_fill_1 FILLER_73_1566 ();
 sg13g2_decap_4 FILLER_73_1581 ();
 sg13g2_fill_2 FILLER_73_1585 ();
 sg13g2_fill_1 FILLER_73_1608 ();
 sg13g2_decap_8 FILLER_73_1632 ();
 sg13g2_decap_4 FILLER_73_1639 ();
 sg13g2_decap_8 FILLER_73_1660 ();
 sg13g2_decap_8 FILLER_73_1685 ();
 sg13g2_decap_8 FILLER_73_1692 ();
 sg13g2_fill_1 FILLER_73_1699 ();
 sg13g2_fill_2 FILLER_73_1735 ();
 sg13g2_fill_2 FILLER_73_1774 ();
 sg13g2_fill_1 FILLER_73_1776 ();
 sg13g2_decap_4 FILLER_73_1794 ();
 sg13g2_fill_2 FILLER_73_1802 ();
 sg13g2_decap_8 FILLER_73_1831 ();
 sg13g2_decap_4 FILLER_73_1838 ();
 sg13g2_fill_1 FILLER_73_1842 ();
 sg13g2_decap_4 FILLER_73_1846 ();
 sg13g2_decap_4 FILLER_73_1854 ();
 sg13g2_fill_2 FILLER_73_1858 ();
 sg13g2_decap_8 FILLER_73_1864 ();
 sg13g2_decap_8 FILLER_73_1871 ();
 sg13g2_decap_8 FILLER_73_1878 ();
 sg13g2_decap_8 FILLER_73_1921 ();
 sg13g2_fill_2 FILLER_73_1928 ();
 sg13g2_decap_4 FILLER_73_1940 ();
 sg13g2_decap_4 FILLER_73_1949 ();
 sg13g2_fill_1 FILLER_73_1953 ();
 sg13g2_fill_1 FILLER_73_1957 ();
 sg13g2_fill_1 FILLER_73_2002 ();
 sg13g2_fill_2 FILLER_73_2006 ();
 sg13g2_fill_1 FILLER_73_2012 ();
 sg13g2_decap_8 FILLER_73_2028 ();
 sg13g2_decap_8 FILLER_73_2044 ();
 sg13g2_decap_4 FILLER_73_2051 ();
 sg13g2_fill_1 FILLER_73_2055 ();
 sg13g2_decap_4 FILLER_73_2061 ();
 sg13g2_decap_8 FILLER_73_2069 ();
 sg13g2_fill_2 FILLER_73_2091 ();
 sg13g2_fill_2 FILLER_73_2100 ();
 sg13g2_fill_2 FILLER_73_2123 ();
 sg13g2_decap_8 FILLER_73_2147 ();
 sg13g2_fill_1 FILLER_73_2154 ();
 sg13g2_fill_2 FILLER_73_2160 ();
 sg13g2_fill_1 FILLER_73_2162 ();
 sg13g2_decap_4 FILLER_73_2183 ();
 sg13g2_fill_1 FILLER_73_2187 ();
 sg13g2_decap_4 FILLER_73_2210 ();
 sg13g2_fill_2 FILLER_73_2242 ();
 sg13g2_fill_1 FILLER_73_2244 ();
 sg13g2_decap_8 FILLER_73_2254 ();
 sg13g2_decap_8 FILLER_73_2261 ();
 sg13g2_fill_1 FILLER_73_2268 ();
 sg13g2_fill_1 FILLER_73_2278 ();
 sg13g2_decap_8 FILLER_73_2283 ();
 sg13g2_decap_4 FILLER_73_2290 ();
 sg13g2_fill_2 FILLER_73_2294 ();
 sg13g2_fill_2 FILLER_73_2310 ();
 sg13g2_fill_1 FILLER_73_2312 ();
 sg13g2_fill_2 FILLER_73_2343 ();
 sg13g2_fill_1 FILLER_73_2345 ();
 sg13g2_fill_2 FILLER_73_2367 ();
 sg13g2_fill_1 FILLER_73_2369 ();
 sg13g2_decap_4 FILLER_73_2389 ();
 sg13g2_decap_4 FILLER_73_2404 ();
 sg13g2_decap_4 FILLER_73_2421 ();
 sg13g2_fill_2 FILLER_73_2425 ();
 sg13g2_decap_4 FILLER_73_2449 ();
 sg13g2_decap_4 FILLER_73_2501 ();
 sg13g2_fill_1 FILLER_73_2505 ();
 sg13g2_fill_1 FILLER_73_2519 ();
 sg13g2_fill_2 FILLER_73_2541 ();
 sg13g2_decap_8 FILLER_73_2550 ();
 sg13g2_fill_2 FILLER_73_2576 ();
 sg13g2_fill_1 FILLER_73_2583 ();
 sg13g2_fill_2 FILLER_73_2588 ();
 sg13g2_fill_1 FILLER_73_2594 ();
 sg13g2_fill_2 FILLER_73_2610 ();
 sg13g2_fill_1 FILLER_73_2612 ();
 sg13g2_fill_2 FILLER_73_2622 ();
 sg13g2_fill_1 FILLER_73_2624 ();
 sg13g2_decap_8 FILLER_73_2630 ();
 sg13g2_fill_2 FILLER_73_2637 ();
 sg13g2_fill_2 FILLER_73_2644 ();
 sg13g2_fill_1 FILLER_73_2646 ();
 sg13g2_decap_8 FILLER_73_2656 ();
 sg13g2_fill_2 FILLER_73_2663 ();
 sg13g2_fill_1 FILLER_73_2665 ();
 sg13g2_decap_8 FILLER_73_2682 ();
 sg13g2_fill_2 FILLER_73_2694 ();
 sg13g2_decap_8 FILLER_73_2710 ();
 sg13g2_decap_8 FILLER_73_2717 ();
 sg13g2_decap_8 FILLER_73_2724 ();
 sg13g2_decap_4 FILLER_73_2731 ();
 sg13g2_decap_8 FILLER_73_2755 ();
 sg13g2_decap_4 FILLER_73_2762 ();
 sg13g2_fill_1 FILLER_73_2790 ();
 sg13g2_decap_8 FILLER_73_2796 ();
 sg13g2_fill_2 FILLER_73_2803 ();
 sg13g2_fill_2 FILLER_73_2813 ();
 sg13g2_fill_1 FILLER_73_2815 ();
 sg13g2_fill_1 FILLER_73_2822 ();
 sg13g2_decap_4 FILLER_73_2827 ();
 sg13g2_fill_2 FILLER_73_2831 ();
 sg13g2_decap_4 FILLER_73_2837 ();
 sg13g2_decap_4 FILLER_73_2849 ();
 sg13g2_fill_2 FILLER_73_2853 ();
 sg13g2_decap_4 FILLER_73_2923 ();
 sg13g2_fill_2 FILLER_73_2927 ();
 sg13g2_fill_1 FILLER_73_2978 ();
 sg13g2_fill_2 FILLER_73_2992 ();
 sg13g2_fill_2 FILLER_73_3003 ();
 sg13g2_fill_1 FILLER_73_3035 ();
 sg13g2_fill_1 FILLER_73_3077 ();
 sg13g2_fill_2 FILLER_73_3093 ();
 sg13g2_fill_2 FILLER_73_3099 ();
 sg13g2_decap_8 FILLER_73_3110 ();
 sg13g2_decap_8 FILLER_73_3117 ();
 sg13g2_decap_8 FILLER_73_3124 ();
 sg13g2_decap_8 FILLER_73_3131 ();
 sg13g2_decap_8 FILLER_73_3138 ();
 sg13g2_decap_8 FILLER_73_3145 ();
 sg13g2_decap_8 FILLER_73_3152 ();
 sg13g2_decap_8 FILLER_73_3159 ();
 sg13g2_decap_8 FILLER_73_3166 ();
 sg13g2_decap_8 FILLER_73_3173 ();
 sg13g2_decap_8 FILLER_73_3180 ();
 sg13g2_decap_8 FILLER_73_3187 ();
 sg13g2_decap_8 FILLER_73_3194 ();
 sg13g2_decap_8 FILLER_73_3201 ();
 sg13g2_decap_8 FILLER_73_3208 ();
 sg13g2_decap_8 FILLER_73_3215 ();
 sg13g2_decap_8 FILLER_73_3222 ();
 sg13g2_decap_8 FILLER_73_3229 ();
 sg13g2_decap_8 FILLER_73_3236 ();
 sg13g2_decap_8 FILLER_73_3243 ();
 sg13g2_decap_8 FILLER_73_3250 ();
 sg13g2_decap_8 FILLER_73_3257 ();
 sg13g2_decap_8 FILLER_73_3264 ();
 sg13g2_decap_8 FILLER_73_3271 ();
 sg13g2_decap_8 FILLER_73_3278 ();
 sg13g2_decap_8 FILLER_73_3285 ();
 sg13g2_decap_8 FILLER_73_3292 ();
 sg13g2_decap_8 FILLER_73_3299 ();
 sg13g2_decap_8 FILLER_73_3306 ();
 sg13g2_decap_8 FILLER_73_3313 ();
 sg13g2_decap_8 FILLER_73_3320 ();
 sg13g2_decap_8 FILLER_73_3327 ();
 sg13g2_decap_8 FILLER_73_3334 ();
 sg13g2_decap_8 FILLER_73_3341 ();
 sg13g2_decap_8 FILLER_73_3348 ();
 sg13g2_decap_8 FILLER_73_3355 ();
 sg13g2_decap_8 FILLER_73_3362 ();
 sg13g2_decap_8 FILLER_73_3369 ();
 sg13g2_decap_8 FILLER_73_3376 ();
 sg13g2_decap_8 FILLER_73_3383 ();
 sg13g2_decap_8 FILLER_73_3390 ();
 sg13g2_decap_8 FILLER_73_3397 ();
 sg13g2_decap_8 FILLER_73_3404 ();
 sg13g2_decap_8 FILLER_73_3411 ();
 sg13g2_decap_8 FILLER_73_3418 ();
 sg13g2_decap_8 FILLER_73_3425 ();
 sg13g2_decap_8 FILLER_73_3432 ();
 sg13g2_decap_8 FILLER_73_3439 ();
 sg13g2_decap_8 FILLER_73_3446 ();
 sg13g2_decap_8 FILLER_73_3453 ();
 sg13g2_decap_8 FILLER_73_3460 ();
 sg13g2_decap_8 FILLER_73_3467 ();
 sg13g2_decap_8 FILLER_73_3474 ();
 sg13g2_decap_8 FILLER_73_3481 ();
 sg13g2_decap_8 FILLER_73_3488 ();
 sg13g2_decap_8 FILLER_73_3495 ();
 sg13g2_decap_8 FILLER_73_3502 ();
 sg13g2_decap_8 FILLER_73_3509 ();
 sg13g2_decap_8 FILLER_73_3516 ();
 sg13g2_decap_8 FILLER_73_3523 ();
 sg13g2_decap_8 FILLER_73_3530 ();
 sg13g2_decap_8 FILLER_73_3537 ();
 sg13g2_decap_8 FILLER_73_3544 ();
 sg13g2_decap_8 FILLER_73_3551 ();
 sg13g2_decap_8 FILLER_73_3558 ();
 sg13g2_decap_8 FILLER_73_3565 ();
 sg13g2_decap_8 FILLER_73_3572 ();
 sg13g2_fill_1 FILLER_73_3579 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_fill_2 FILLER_74_294 ();
 sg13g2_fill_1 FILLER_74_296 ();
 sg13g2_fill_2 FILLER_74_420 ();
 sg13g2_fill_2 FILLER_74_459 ();
 sg13g2_decap_8 FILLER_74_465 ();
 sg13g2_fill_2 FILLER_74_490 ();
 sg13g2_fill_2 FILLER_74_508 ();
 sg13g2_fill_1 FILLER_74_510 ();
 sg13g2_fill_2 FILLER_74_535 ();
 sg13g2_fill_1 FILLER_74_537 ();
 sg13g2_decap_4 FILLER_74_553 ();
 sg13g2_decap_4 FILLER_74_583 ();
 sg13g2_fill_1 FILLER_74_587 ();
 sg13g2_fill_1 FILLER_74_606 ();
 sg13g2_decap_4 FILLER_74_612 ();
 sg13g2_fill_1 FILLER_74_639 ();
 sg13g2_decap_4 FILLER_74_645 ();
 sg13g2_fill_2 FILLER_74_649 ();
 sg13g2_fill_2 FILLER_74_656 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_fill_2 FILLER_74_695 ();
 sg13g2_decap_4 FILLER_74_704 ();
 sg13g2_fill_1 FILLER_74_708 ();
 sg13g2_fill_1 FILLER_74_730 ();
 sg13g2_fill_2 FILLER_74_744 ();
 sg13g2_fill_2 FILLER_74_761 ();
 sg13g2_fill_1 FILLER_74_776 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_fill_1 FILLER_74_797 ();
 sg13g2_decap_4 FILLER_74_804 ();
 sg13g2_fill_1 FILLER_74_808 ();
 sg13g2_fill_1 FILLER_74_818 ();
 sg13g2_fill_2 FILLER_74_829 ();
 sg13g2_fill_1 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_855 ();
 sg13g2_decap_4 FILLER_74_862 ();
 sg13g2_fill_2 FILLER_74_866 ();
 sg13g2_fill_1 FILLER_74_882 ();
 sg13g2_decap_4 FILLER_74_909 ();
 sg13g2_fill_2 FILLER_74_913 ();
 sg13g2_decap_8 FILLER_74_936 ();
 sg13g2_decap_8 FILLER_74_943 ();
 sg13g2_fill_2 FILLER_74_950 ();
 sg13g2_fill_1 FILLER_74_958 ();
 sg13g2_fill_2 FILLER_74_977 ();
 sg13g2_fill_1 FILLER_74_979 ();
 sg13g2_fill_1 FILLER_74_1049 ();
 sg13g2_decap_8 FILLER_74_1060 ();
 sg13g2_decap_8 FILLER_74_1067 ();
 sg13g2_decap_4 FILLER_74_1074 ();
 sg13g2_fill_1 FILLER_74_1078 ();
 sg13g2_fill_2 FILLER_74_1114 ();
 sg13g2_fill_2 FILLER_74_1120 ();
 sg13g2_fill_1 FILLER_74_1122 ();
 sg13g2_fill_1 FILLER_74_1136 ();
 sg13g2_fill_2 FILLER_74_1151 ();
 sg13g2_fill_1 FILLER_74_1153 ();
 sg13g2_fill_1 FILLER_74_1168 ();
 sg13g2_fill_2 FILLER_74_1209 ();
 sg13g2_decap_4 FILLER_74_1239 ();
 sg13g2_fill_1 FILLER_74_1243 ();
 sg13g2_fill_2 FILLER_74_1262 ();
 sg13g2_fill_1 FILLER_74_1271 ();
 sg13g2_decap_8 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_fill_1 FILLER_74_1302 ();
 sg13g2_fill_1 FILLER_74_1308 ();
 sg13g2_fill_1 FILLER_74_1312 ();
 sg13g2_fill_1 FILLER_74_1319 ();
 sg13g2_decap_8 FILLER_74_1324 ();
 sg13g2_decap_8 FILLER_74_1331 ();
 sg13g2_fill_1 FILLER_74_1338 ();
 sg13g2_fill_2 FILLER_74_1347 ();
 sg13g2_decap_8 FILLER_74_1377 ();
 sg13g2_decap_8 FILLER_74_1384 ();
 sg13g2_fill_2 FILLER_74_1396 ();
 sg13g2_fill_1 FILLER_74_1398 ();
 sg13g2_decap_4 FILLER_74_1416 ();
 sg13g2_decap_4 FILLER_74_1425 ();
 sg13g2_fill_2 FILLER_74_1429 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_decap_8 FILLER_74_1456 ();
 sg13g2_decap_4 FILLER_74_1463 ();
 sg13g2_fill_2 FILLER_74_1467 ();
 sg13g2_fill_1 FILLER_74_1485 ();
 sg13g2_fill_1 FILLER_74_1491 ();
 sg13g2_fill_2 FILLER_74_1497 ();
 sg13g2_fill_1 FILLER_74_1499 ();
 sg13g2_fill_2 FILLER_74_1505 ();
 sg13g2_fill_1 FILLER_74_1507 ();
 sg13g2_decap_8 FILLER_74_1521 ();
 sg13g2_fill_2 FILLER_74_1528 ();
 sg13g2_decap_8 FILLER_74_1534 ();
 sg13g2_decap_8 FILLER_74_1541 ();
 sg13g2_decap_4 FILLER_74_1588 ();
 sg13g2_decap_8 FILLER_74_1607 ();
 sg13g2_decap_4 FILLER_74_1614 ();
 sg13g2_fill_1 FILLER_74_1618 ();
 sg13g2_decap_8 FILLER_74_1624 ();
 sg13g2_decap_4 FILLER_74_1631 ();
 sg13g2_decap_8 FILLER_74_1657 ();
 sg13g2_fill_1 FILLER_74_1688 ();
 sg13g2_decap_8 FILLER_74_1715 ();
 sg13g2_decap_4 FILLER_74_1722 ();
 sg13g2_fill_1 FILLER_74_1726 ();
 sg13g2_fill_1 FILLER_74_1745 ();
 sg13g2_fill_1 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1769 ();
 sg13g2_decap_4 FILLER_74_1782 ();
 sg13g2_fill_2 FILLER_74_1790 ();
 sg13g2_decap_8 FILLER_74_1829 ();
 sg13g2_decap_8 FILLER_74_1836 ();
 sg13g2_fill_2 FILLER_74_1843 ();
 sg13g2_fill_2 FILLER_74_1893 ();
 sg13g2_decap_8 FILLER_74_1918 ();
 sg13g2_fill_2 FILLER_74_1946 ();
 sg13g2_fill_1 FILLER_74_1948 ();
 sg13g2_decap_4 FILLER_74_1959 ();
 sg13g2_decap_8 FILLER_74_1967 ();
 sg13g2_decap_4 FILLER_74_1974 ();
 sg13g2_fill_1 FILLER_74_1984 ();
 sg13g2_fill_1 FILLER_74_1997 ();
 sg13g2_fill_2 FILLER_74_2015 ();
 sg13g2_fill_1 FILLER_74_2017 ();
 sg13g2_decap_4 FILLER_74_2026 ();
 sg13g2_fill_1 FILLER_74_2030 ();
 sg13g2_fill_1 FILLER_74_2051 ();
 sg13g2_fill_2 FILLER_74_2061 ();
 sg13g2_fill_1 FILLER_74_2063 ();
 sg13g2_decap_8 FILLER_74_2125 ();
 sg13g2_decap_4 FILLER_74_2132 ();
 sg13g2_fill_1 FILLER_74_2136 ();
 sg13g2_decap_4 FILLER_74_2154 ();
 sg13g2_fill_1 FILLER_74_2158 ();
 sg13g2_decap_8 FILLER_74_2172 ();
 sg13g2_decap_8 FILLER_74_2179 ();
 sg13g2_fill_1 FILLER_74_2186 ();
 sg13g2_fill_1 FILLER_74_2205 ();
 sg13g2_decap_4 FILLER_74_2242 ();
 sg13g2_decap_8 FILLER_74_2254 ();
 sg13g2_decap_4 FILLER_74_2261 ();
 sg13g2_decap_4 FILLER_74_2311 ();
 sg13g2_decap_4 FILLER_74_2320 ();
 sg13g2_fill_1 FILLER_74_2324 ();
 sg13g2_fill_1 FILLER_74_2330 ();
 sg13g2_fill_2 FILLER_74_2335 ();
 sg13g2_fill_2 FILLER_74_2341 ();
 sg13g2_fill_2 FILLER_74_2358 ();
 sg13g2_decap_4 FILLER_74_2423 ();
 sg13g2_fill_1 FILLER_74_2427 ();
 sg13g2_fill_1 FILLER_74_2456 ();
 sg13g2_decap_4 FILLER_74_2552 ();
 sg13g2_fill_1 FILLER_74_2556 ();
 sg13g2_decap_4 FILLER_74_2591 ();
 sg13g2_decap_4 FILLER_74_2607 ();
 sg13g2_fill_2 FILLER_74_2611 ();
 sg13g2_fill_1 FILLER_74_2641 ();
 sg13g2_decap_8 FILLER_74_2671 ();
 sg13g2_decap_4 FILLER_74_2678 ();
 sg13g2_fill_1 FILLER_74_2682 ();
 sg13g2_decap_4 FILLER_74_2707 ();
 sg13g2_decap_4 FILLER_74_2786 ();
 sg13g2_fill_2 FILLER_74_2790 ();
 sg13g2_fill_1 FILLER_74_2797 ();
 sg13g2_fill_2 FILLER_74_2811 ();
 sg13g2_fill_2 FILLER_74_2843 ();
 sg13g2_decap_8 FILLER_74_2849 ();
 sg13g2_fill_2 FILLER_74_2856 ();
 sg13g2_fill_1 FILLER_74_2858 ();
 sg13g2_decap_4 FILLER_74_2887 ();
 sg13g2_decap_4 FILLER_74_2895 ();
 sg13g2_fill_2 FILLER_74_2899 ();
 sg13g2_decap_4 FILLER_74_2929 ();
 sg13g2_fill_2 FILLER_74_2939 ();
 sg13g2_decap_8 FILLER_74_2944 ();
 sg13g2_decap_4 FILLER_74_2951 ();
 sg13g2_decap_8 FILLER_74_2959 ();
 sg13g2_decap_4 FILLER_74_2966 ();
 sg13g2_fill_1 FILLER_74_2998 ();
 sg13g2_decap_8 FILLER_74_3012 ();
 sg13g2_fill_2 FILLER_74_3019 ();
 sg13g2_decap_8 FILLER_74_3026 ();
 sg13g2_decap_8 FILLER_74_3033 ();
 sg13g2_fill_1 FILLER_74_3040 ();
 sg13g2_decap_8 FILLER_74_3054 ();
 sg13g2_decap_4 FILLER_74_3061 ();
 sg13g2_fill_1 FILLER_74_3065 ();
 sg13g2_decap_8 FILLER_74_3122 ();
 sg13g2_decap_8 FILLER_74_3129 ();
 sg13g2_decap_8 FILLER_74_3136 ();
 sg13g2_decap_8 FILLER_74_3143 ();
 sg13g2_decap_8 FILLER_74_3150 ();
 sg13g2_decap_8 FILLER_74_3157 ();
 sg13g2_decap_8 FILLER_74_3164 ();
 sg13g2_decap_8 FILLER_74_3171 ();
 sg13g2_decap_8 FILLER_74_3178 ();
 sg13g2_decap_8 FILLER_74_3185 ();
 sg13g2_decap_8 FILLER_74_3192 ();
 sg13g2_decap_8 FILLER_74_3199 ();
 sg13g2_decap_8 FILLER_74_3206 ();
 sg13g2_decap_8 FILLER_74_3213 ();
 sg13g2_decap_8 FILLER_74_3220 ();
 sg13g2_decap_8 FILLER_74_3227 ();
 sg13g2_decap_8 FILLER_74_3234 ();
 sg13g2_decap_8 FILLER_74_3241 ();
 sg13g2_decap_8 FILLER_74_3248 ();
 sg13g2_decap_8 FILLER_74_3255 ();
 sg13g2_decap_8 FILLER_74_3262 ();
 sg13g2_decap_8 FILLER_74_3269 ();
 sg13g2_decap_8 FILLER_74_3276 ();
 sg13g2_decap_8 FILLER_74_3283 ();
 sg13g2_decap_8 FILLER_74_3290 ();
 sg13g2_decap_8 FILLER_74_3297 ();
 sg13g2_decap_8 FILLER_74_3304 ();
 sg13g2_decap_8 FILLER_74_3311 ();
 sg13g2_decap_8 FILLER_74_3318 ();
 sg13g2_decap_8 FILLER_74_3325 ();
 sg13g2_decap_8 FILLER_74_3332 ();
 sg13g2_decap_8 FILLER_74_3339 ();
 sg13g2_decap_8 FILLER_74_3346 ();
 sg13g2_decap_8 FILLER_74_3353 ();
 sg13g2_decap_8 FILLER_74_3360 ();
 sg13g2_decap_8 FILLER_74_3367 ();
 sg13g2_decap_8 FILLER_74_3374 ();
 sg13g2_decap_8 FILLER_74_3381 ();
 sg13g2_decap_8 FILLER_74_3388 ();
 sg13g2_decap_8 FILLER_74_3395 ();
 sg13g2_decap_8 FILLER_74_3402 ();
 sg13g2_decap_8 FILLER_74_3409 ();
 sg13g2_decap_8 FILLER_74_3416 ();
 sg13g2_decap_8 FILLER_74_3423 ();
 sg13g2_decap_8 FILLER_74_3430 ();
 sg13g2_decap_8 FILLER_74_3437 ();
 sg13g2_decap_8 FILLER_74_3444 ();
 sg13g2_decap_8 FILLER_74_3451 ();
 sg13g2_decap_8 FILLER_74_3458 ();
 sg13g2_decap_8 FILLER_74_3465 ();
 sg13g2_decap_8 FILLER_74_3472 ();
 sg13g2_decap_8 FILLER_74_3479 ();
 sg13g2_decap_8 FILLER_74_3486 ();
 sg13g2_decap_8 FILLER_74_3493 ();
 sg13g2_decap_8 FILLER_74_3500 ();
 sg13g2_decap_8 FILLER_74_3507 ();
 sg13g2_decap_8 FILLER_74_3514 ();
 sg13g2_decap_8 FILLER_74_3521 ();
 sg13g2_decap_8 FILLER_74_3528 ();
 sg13g2_decap_8 FILLER_74_3535 ();
 sg13g2_decap_8 FILLER_74_3542 ();
 sg13g2_decap_8 FILLER_74_3549 ();
 sg13g2_decap_8 FILLER_74_3556 ();
 sg13g2_decap_8 FILLER_74_3563 ();
 sg13g2_decap_8 FILLER_74_3570 ();
 sg13g2_fill_2 FILLER_74_3577 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_4 FILLER_75_308 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_fill_2 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_4 FILLER_75_388 ();
 sg13g2_fill_2 FILLER_75_392 ();
 sg13g2_fill_1 FILLER_75_413 ();
 sg13g2_fill_2 FILLER_75_423 ();
 sg13g2_fill_2 FILLER_75_505 ();
 sg13g2_fill_1 FILLER_75_507 ();
 sg13g2_decap_4 FILLER_75_524 ();
 sg13g2_fill_2 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_535 ();
 sg13g2_fill_2 FILLER_75_542 ();
 sg13g2_fill_2 FILLER_75_552 ();
 sg13g2_decap_8 FILLER_75_559 ();
 sg13g2_decap_8 FILLER_75_581 ();
 sg13g2_decap_4 FILLER_75_596 ();
 sg13g2_decap_8 FILLER_75_610 ();
 sg13g2_decap_4 FILLER_75_617 ();
 sg13g2_fill_2 FILLER_75_621 ();
 sg13g2_decap_4 FILLER_75_646 ();
 sg13g2_decap_8 FILLER_75_667 ();
 sg13g2_fill_1 FILLER_75_674 ();
 sg13g2_decap_8 FILLER_75_694 ();
 sg13g2_decap_4 FILLER_75_701 ();
 sg13g2_fill_2 FILLER_75_720 ();
 sg13g2_fill_2 FILLER_75_727 ();
 sg13g2_fill_2 FILLER_75_750 ();
 sg13g2_decap_4 FILLER_75_758 ();
 sg13g2_fill_1 FILLER_75_762 ();
 sg13g2_fill_2 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_807 ();
 sg13g2_decap_8 FILLER_75_827 ();
 sg13g2_decap_8 FILLER_75_834 ();
 sg13g2_fill_2 FILLER_75_841 ();
 sg13g2_fill_1 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_fill_1 FILLER_75_855 ();
 sg13g2_decap_4 FILLER_75_882 ();
 sg13g2_fill_1 FILLER_75_895 ();
 sg13g2_decap_8 FILLER_75_905 ();
 sg13g2_decap_4 FILLER_75_912 ();
 sg13g2_fill_2 FILLER_75_916 ();
 sg13g2_decap_4 FILLER_75_930 ();
 sg13g2_decap_4 FILLER_75_941 ();
 sg13g2_decap_4 FILLER_75_963 ();
 sg13g2_fill_1 FILLER_75_970 ();
 sg13g2_decap_8 FILLER_75_976 ();
 sg13g2_decap_4 FILLER_75_986 ();
 sg13g2_decap_8 FILLER_75_995 ();
 sg13g2_decap_4 FILLER_75_1002 ();
 sg13g2_fill_1 FILLER_75_1006 ();
 sg13g2_fill_1 FILLER_75_1035 ();
 sg13g2_fill_1 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1059 ();
 sg13g2_fill_1 FILLER_75_1071 ();
 sg13g2_decap_8 FILLER_75_1101 ();
 sg13g2_decap_8 FILLER_75_1108 ();
 sg13g2_fill_1 FILLER_75_1149 ();
 sg13g2_fill_2 FILLER_75_1172 ();
 sg13g2_decap_8 FILLER_75_1187 ();
 sg13g2_fill_1 FILLER_75_1194 ();
 sg13g2_decap_8 FILLER_75_1199 ();
 sg13g2_fill_1 FILLER_75_1206 ();
 sg13g2_fill_1 FILLER_75_1228 ();
 sg13g2_fill_2 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1257 ();
 sg13g2_decap_4 FILLER_75_1264 ();
 sg13g2_fill_1 FILLER_75_1268 ();
 sg13g2_fill_2 FILLER_75_1272 ();
 sg13g2_fill_2 FILLER_75_1283 ();
 sg13g2_fill_1 FILLER_75_1285 ();
 sg13g2_decap_4 FILLER_75_1291 ();
 sg13g2_fill_2 FILLER_75_1312 ();
 sg13g2_decap_4 FILLER_75_1328 ();
 sg13g2_fill_2 FILLER_75_1332 ();
 sg13g2_decap_8 FILLER_75_1345 ();
 sg13g2_fill_2 FILLER_75_1352 ();
 sg13g2_decap_8 FILLER_75_1358 ();
 sg13g2_fill_1 FILLER_75_1365 ();
 sg13g2_decap_4 FILLER_75_1402 ();
 sg13g2_decap_8 FILLER_75_1426 ();
 sg13g2_fill_1 FILLER_75_1433 ();
 sg13g2_decap_4 FILLER_75_1438 ();
 sg13g2_fill_2 FILLER_75_1442 ();
 sg13g2_fill_1 FILLER_75_1462 ();
 sg13g2_decap_4 FILLER_75_1468 ();
 sg13g2_fill_1 FILLER_75_1472 ();
 sg13g2_fill_1 FILLER_75_1479 ();
 sg13g2_fill_2 FILLER_75_1493 ();
 sg13g2_fill_1 FILLER_75_1495 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_decap_8 FILLER_75_1509 ();
 sg13g2_decap_8 FILLER_75_1516 ();
 sg13g2_fill_1 FILLER_75_1523 ();
 sg13g2_fill_2 FILLER_75_1574 ();
 sg13g2_decap_8 FILLER_75_1590 ();
 sg13g2_fill_1 FILLER_75_1607 ();
 sg13g2_decap_8 FILLER_75_1629 ();
 sg13g2_decap_8 FILLER_75_1652 ();
 sg13g2_decap_8 FILLER_75_1659 ();
 sg13g2_fill_2 FILLER_75_1767 ();
 sg13g2_fill_1 FILLER_75_1769 ();
 sg13g2_fill_2 FILLER_75_1807 ();
 sg13g2_fill_2 FILLER_75_1813 ();
 sg13g2_decap_8 FILLER_75_1843 ();
 sg13g2_decap_8 FILLER_75_1850 ();
 sg13g2_decap_4 FILLER_75_1857 ();
 sg13g2_fill_1 FILLER_75_1861 ();
 sg13g2_fill_2 FILLER_75_1887 ();
 sg13g2_decap_4 FILLER_75_1918 ();
 sg13g2_fill_2 FILLER_75_1922 ();
 sg13g2_decap_8 FILLER_75_1936 ();
 sg13g2_fill_1 FILLER_75_1943 ();
 sg13g2_fill_2 FILLER_75_1959 ();
 sg13g2_decap_4 FILLER_75_1966 ();
 sg13g2_fill_1 FILLER_75_1970 ();
 sg13g2_fill_2 FILLER_75_1978 ();
 sg13g2_fill_1 FILLER_75_1980 ();
 sg13g2_decap_4 FILLER_75_1992 ();
 sg13g2_decap_8 FILLER_75_2012 ();
 sg13g2_decap_8 FILLER_75_2036 ();
 sg13g2_fill_2 FILLER_75_2056 ();
 sg13g2_decap_4 FILLER_75_2076 ();
 sg13g2_fill_2 FILLER_75_2080 ();
 sg13g2_decap_4 FILLER_75_2086 ();
 sg13g2_fill_2 FILLER_75_2106 ();
 sg13g2_fill_1 FILLER_75_2114 ();
 sg13g2_decap_8 FILLER_75_2118 ();
 sg13g2_decap_8 FILLER_75_2130 ();
 sg13g2_decap_8 FILLER_75_2137 ();
 sg13g2_fill_2 FILLER_75_2144 ();
 sg13g2_fill_1 FILLER_75_2169 ();
 sg13g2_fill_2 FILLER_75_2196 ();
 sg13g2_fill_2 FILLER_75_2214 ();
 sg13g2_decap_8 FILLER_75_2233 ();
 sg13g2_fill_2 FILLER_75_2240 ();
 sg13g2_fill_1 FILLER_75_2242 ();
 sg13g2_decap_4 FILLER_75_2303 ();
 sg13g2_fill_2 FILLER_75_2324 ();
 sg13g2_fill_1 FILLER_75_2326 ();
 sg13g2_decap_4 FILLER_75_2360 ();
 sg13g2_fill_2 FILLER_75_2364 ();
 sg13g2_fill_2 FILLER_75_2408 ();
 sg13g2_fill_1 FILLER_75_2419 ();
 sg13g2_decap_8 FILLER_75_2448 ();
 sg13g2_decap_8 FILLER_75_2455 ();
 sg13g2_decap_4 FILLER_75_2462 ();
 sg13g2_decap_8 FILLER_75_2470 ();
 sg13g2_decap_8 FILLER_75_2477 ();
 sg13g2_fill_1 FILLER_75_2484 ();
 sg13g2_decap_8 FILLER_75_2498 ();
 sg13g2_decap_8 FILLER_75_2505 ();
 sg13g2_decap_4 FILLER_75_2512 ();
 sg13g2_fill_2 FILLER_75_2516 ();
 sg13g2_decap_8 FILLER_75_2522 ();
 sg13g2_decap_4 FILLER_75_2529 ();
 sg13g2_fill_2 FILLER_75_2533 ();
 sg13g2_fill_2 FILLER_75_2572 ();
 sg13g2_fill_2 FILLER_75_2599 ();
 sg13g2_fill_2 FILLER_75_2629 ();
 sg13g2_fill_1 FILLER_75_2631 ();
 sg13g2_fill_1 FILLER_75_2641 ();
 sg13g2_fill_2 FILLER_75_2695 ();
 sg13g2_fill_1 FILLER_75_2697 ();
 sg13g2_decap_4 FILLER_75_2707 ();
 sg13g2_fill_1 FILLER_75_2715 ();
 sg13g2_decap_8 FILLER_75_2729 ();
 sg13g2_fill_2 FILLER_75_2753 ();
 sg13g2_decap_8 FILLER_75_2785 ();
 sg13g2_decap_8 FILLER_75_2792 ();
 sg13g2_fill_1 FILLER_75_2799 ();
 sg13g2_decap_8 FILLER_75_2813 ();
 sg13g2_decap_8 FILLER_75_2820 ();
 sg13g2_decap_4 FILLER_75_2827 ();
 sg13g2_fill_1 FILLER_75_2831 ();
 sg13g2_decap_4 FILLER_75_2835 ();
 sg13g2_fill_1 FILLER_75_2839 ();
 sg13g2_decap_8 FILLER_75_2868 ();
 sg13g2_decap_8 FILLER_75_2875 ();
 sg13g2_decap_8 FILLER_75_2882 ();
 sg13g2_decap_8 FILLER_75_2889 ();
 sg13g2_decap_8 FILLER_75_2896 ();
 sg13g2_fill_2 FILLER_75_2903 ();
 sg13g2_fill_1 FILLER_75_2905 ();
 sg13g2_decap_8 FILLER_75_2910 ();
 sg13g2_decap_8 FILLER_75_2917 ();
 sg13g2_fill_1 FILLER_75_2924 ();
 sg13g2_decap_8 FILLER_75_2961 ();
 sg13g2_decap_8 FILLER_75_2968 ();
 sg13g2_fill_1 FILLER_75_2975 ();
 sg13g2_decap_8 FILLER_75_2980 ();
 sg13g2_decap_4 FILLER_75_3015 ();
 sg13g2_fill_1 FILLER_75_3019 ();
 sg13g2_decap_8 FILLER_75_3056 ();
 sg13g2_fill_2 FILLER_75_3063 ();
 sg13g2_decap_8 FILLER_75_3078 ();
 sg13g2_decap_4 FILLER_75_3085 ();
 sg13g2_fill_2 FILLER_75_3089 ();
 sg13g2_fill_2 FILLER_75_3100 ();
 sg13g2_decap_8 FILLER_75_3111 ();
 sg13g2_decap_8 FILLER_75_3118 ();
 sg13g2_decap_8 FILLER_75_3125 ();
 sg13g2_decap_8 FILLER_75_3132 ();
 sg13g2_decap_8 FILLER_75_3139 ();
 sg13g2_decap_8 FILLER_75_3146 ();
 sg13g2_decap_8 FILLER_75_3153 ();
 sg13g2_decap_8 FILLER_75_3160 ();
 sg13g2_decap_8 FILLER_75_3167 ();
 sg13g2_decap_8 FILLER_75_3174 ();
 sg13g2_decap_8 FILLER_75_3181 ();
 sg13g2_decap_8 FILLER_75_3188 ();
 sg13g2_decap_8 FILLER_75_3195 ();
 sg13g2_decap_8 FILLER_75_3202 ();
 sg13g2_decap_8 FILLER_75_3209 ();
 sg13g2_decap_8 FILLER_75_3216 ();
 sg13g2_decap_8 FILLER_75_3223 ();
 sg13g2_decap_8 FILLER_75_3230 ();
 sg13g2_decap_8 FILLER_75_3237 ();
 sg13g2_decap_8 FILLER_75_3244 ();
 sg13g2_decap_8 FILLER_75_3251 ();
 sg13g2_decap_8 FILLER_75_3258 ();
 sg13g2_decap_8 FILLER_75_3265 ();
 sg13g2_decap_8 FILLER_75_3272 ();
 sg13g2_decap_8 FILLER_75_3279 ();
 sg13g2_decap_8 FILLER_75_3286 ();
 sg13g2_decap_8 FILLER_75_3293 ();
 sg13g2_decap_8 FILLER_75_3300 ();
 sg13g2_decap_8 FILLER_75_3307 ();
 sg13g2_decap_8 FILLER_75_3314 ();
 sg13g2_decap_8 FILLER_75_3321 ();
 sg13g2_decap_8 FILLER_75_3328 ();
 sg13g2_decap_8 FILLER_75_3335 ();
 sg13g2_decap_8 FILLER_75_3342 ();
 sg13g2_decap_8 FILLER_75_3349 ();
 sg13g2_decap_8 FILLER_75_3356 ();
 sg13g2_decap_8 FILLER_75_3363 ();
 sg13g2_decap_8 FILLER_75_3370 ();
 sg13g2_decap_8 FILLER_75_3377 ();
 sg13g2_decap_8 FILLER_75_3384 ();
 sg13g2_decap_8 FILLER_75_3391 ();
 sg13g2_decap_8 FILLER_75_3398 ();
 sg13g2_decap_8 FILLER_75_3405 ();
 sg13g2_decap_8 FILLER_75_3412 ();
 sg13g2_decap_8 FILLER_75_3419 ();
 sg13g2_decap_8 FILLER_75_3426 ();
 sg13g2_decap_8 FILLER_75_3433 ();
 sg13g2_decap_8 FILLER_75_3440 ();
 sg13g2_decap_8 FILLER_75_3447 ();
 sg13g2_decap_8 FILLER_75_3454 ();
 sg13g2_decap_8 FILLER_75_3461 ();
 sg13g2_decap_8 FILLER_75_3468 ();
 sg13g2_decap_8 FILLER_75_3475 ();
 sg13g2_decap_8 FILLER_75_3482 ();
 sg13g2_decap_8 FILLER_75_3489 ();
 sg13g2_decap_8 FILLER_75_3496 ();
 sg13g2_decap_8 FILLER_75_3503 ();
 sg13g2_decap_8 FILLER_75_3510 ();
 sg13g2_decap_8 FILLER_75_3517 ();
 sg13g2_decap_8 FILLER_75_3524 ();
 sg13g2_decap_8 FILLER_75_3531 ();
 sg13g2_decap_8 FILLER_75_3538 ();
 sg13g2_decap_8 FILLER_75_3545 ();
 sg13g2_decap_8 FILLER_75_3552 ();
 sg13g2_decap_8 FILLER_75_3559 ();
 sg13g2_decap_8 FILLER_75_3566 ();
 sg13g2_decap_8 FILLER_75_3573 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_315 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_decap_8 FILLER_76_338 ();
 sg13g2_decap_8 FILLER_76_345 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_8 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_4 FILLER_76_401 ();
 sg13g2_fill_2 FILLER_76_405 ();
 sg13g2_decap_8 FILLER_76_410 ();
 sg13g2_decap_8 FILLER_76_417 ();
 sg13g2_decap_4 FILLER_76_424 ();
 sg13g2_fill_2 FILLER_76_428 ();
 sg13g2_decap_8 FILLER_76_443 ();
 sg13g2_decap_8 FILLER_76_450 ();
 sg13g2_decap_4 FILLER_76_457 ();
 sg13g2_fill_1 FILLER_76_461 ();
 sg13g2_decap_8 FILLER_76_498 ();
 sg13g2_decap_4 FILLER_76_505 ();
 sg13g2_fill_1 FILLER_76_509 ();
 sg13g2_decap_8 FILLER_76_555 ();
 sg13g2_fill_2 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_8 FILLER_76_599 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_617 ();
 sg13g2_fill_2 FILLER_76_624 ();
 sg13g2_fill_1 FILLER_76_626 ();
 sg13g2_fill_2 FILLER_76_638 ();
 sg13g2_fill_1 FILLER_76_645 ();
 sg13g2_decap_8 FILLER_76_650 ();
 sg13g2_fill_1 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_674 ();
 sg13g2_fill_1 FILLER_76_681 ();
 sg13g2_fill_1 FILLER_76_705 ();
 sg13g2_fill_1 FILLER_76_714 ();
 sg13g2_fill_2 FILLER_76_727 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_741 ();
 sg13g2_fill_1 FILLER_76_743 ();
 sg13g2_decap_8 FILLER_76_752 ();
 sg13g2_decap_4 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_fill_2 FILLER_76_797 ();
 sg13g2_fill_1 FILLER_76_799 ();
 sg13g2_fill_2 FILLER_76_816 ();
 sg13g2_fill_1 FILLER_76_818 ();
 sg13g2_fill_2 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_fill_2 FILLER_76_865 ();
 sg13g2_fill_1 FILLER_76_867 ();
 sg13g2_decap_8 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_901 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_fill_2 FILLER_76_909 ();
 sg13g2_fill_2 FILLER_76_948 ();
 sg13g2_decap_8 FILLER_76_959 ();
 sg13g2_decap_4 FILLER_76_966 ();
 sg13g2_fill_1 FILLER_76_970 ();
 sg13g2_fill_2 FILLER_76_984 ();
 sg13g2_fill_2 FILLER_76_1004 ();
 sg13g2_decap_8 FILLER_76_1027 ();
 sg13g2_decap_4 FILLER_76_1034 ();
 sg13g2_fill_2 FILLER_76_1038 ();
 sg13g2_fill_1 FILLER_76_1068 ();
 sg13g2_fill_2 FILLER_76_1081 ();
 sg13g2_fill_1 FILLER_76_1083 ();
 sg13g2_decap_4 FILLER_76_1087 ();
 sg13g2_fill_2 FILLER_76_1095 ();
 sg13g2_fill_1 FILLER_76_1097 ();
 sg13g2_decap_8 FILLER_76_1110 ();
 sg13g2_decap_8 FILLER_76_1117 ();
 sg13g2_fill_2 FILLER_76_1141 ();
 sg13g2_fill_1 FILLER_76_1143 ();
 sg13g2_fill_1 FILLER_76_1163 ();
 sg13g2_fill_2 FILLER_76_1191 ();
 sg13g2_decap_8 FILLER_76_1202 ();
 sg13g2_fill_1 FILLER_76_1209 ();
 sg13g2_decap_8 FILLER_76_1213 ();
 sg13g2_fill_1 FILLER_76_1220 ();
 sg13g2_fill_1 FILLER_76_1231 ();
 sg13g2_decap_4 FILLER_76_1249 ();
 sg13g2_decap_8 FILLER_76_1257 ();
 sg13g2_decap_4 FILLER_76_1264 ();
 sg13g2_fill_2 FILLER_76_1268 ();
 sg13g2_decap_4 FILLER_76_1286 ();
 sg13g2_fill_2 FILLER_76_1316 ();
 sg13g2_fill_1 FILLER_76_1318 ();
 sg13g2_fill_1 FILLER_76_1323 ();
 sg13g2_fill_2 FILLER_76_1338 ();
 sg13g2_decap_8 FILLER_76_1359 ();
 sg13g2_decap_4 FILLER_76_1366 ();
 sg13g2_fill_1 FILLER_76_1370 ();
 sg13g2_decap_4 FILLER_76_1375 ();
 sg13g2_fill_2 FILLER_76_1398 ();
 sg13g2_fill_1 FILLER_76_1400 ();
 sg13g2_fill_2 FILLER_76_1409 ();
 sg13g2_fill_2 FILLER_76_1417 ();
 sg13g2_fill_2 FILLER_76_1434 ();
 sg13g2_fill_1 FILLER_76_1436 ();
 sg13g2_decap_4 FILLER_76_1442 ();
 sg13g2_fill_1 FILLER_76_1446 ();
 sg13g2_fill_2 FILLER_76_1453 ();
 sg13g2_fill_2 FILLER_76_1463 ();
 sg13g2_fill_1 FILLER_76_1465 ();
 sg13g2_decap_8 FILLER_76_1471 ();
 sg13g2_decap_4 FILLER_76_1478 ();
 sg13g2_fill_1 FILLER_76_1482 ();
 sg13g2_decap_8 FILLER_76_1493 ();
 sg13g2_fill_2 FILLER_76_1500 ();
 sg13g2_fill_1 FILLER_76_1520 ();
 sg13g2_decap_4 FILLER_76_1530 ();
 sg13g2_fill_1 FILLER_76_1534 ();
 sg13g2_decap_8 FILLER_76_1539 ();
 sg13g2_fill_2 FILLER_76_1546 ();
 sg13g2_fill_1 FILLER_76_1582 ();
 sg13g2_fill_1 FILLER_76_1599 ();
 sg13g2_fill_2 FILLER_76_1612 ();
 sg13g2_fill_1 FILLER_76_1614 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_decap_4 FILLER_76_1634 ();
 sg13g2_fill_1 FILLER_76_1638 ();
 sg13g2_fill_2 FILLER_76_1658 ();
 sg13g2_fill_1 FILLER_76_1660 ();
 sg13g2_fill_1 FILLER_76_1676 ();
 sg13g2_fill_2 FILLER_76_1682 ();
 sg13g2_decap_8 FILLER_76_1692 ();
 sg13g2_decap_8 FILLER_76_1699 ();
 sg13g2_fill_2 FILLER_76_1706 ();
 sg13g2_decap_8 FILLER_76_1712 ();
 sg13g2_decap_8 FILLER_76_1719 ();
 sg13g2_decap_8 FILLER_76_1726 ();
 sg13g2_fill_2 FILLER_76_1733 ();
 sg13g2_decap_8 FILLER_76_1739 ();
 sg13g2_decap_8 FILLER_76_1746 ();
 sg13g2_fill_2 FILLER_76_1753 ();
 sg13g2_fill_2 FILLER_76_1782 ();
 sg13g2_decap_8 FILLER_76_1788 ();
 sg13g2_fill_1 FILLER_76_1795 ();
 sg13g2_decap_4 FILLER_76_1827 ();
 sg13g2_fill_2 FILLER_76_1910 ();
 sg13g2_fill_1 FILLER_76_1912 ();
 sg13g2_fill_1 FILLER_76_1922 ();
 sg13g2_fill_2 FILLER_76_1942 ();
 sg13g2_decap_4 FILLER_76_1956 ();
 sg13g2_decap_4 FILLER_76_1964 ();
 sg13g2_fill_2 FILLER_76_1968 ();
 sg13g2_fill_2 FILLER_76_1992 ();
 sg13g2_fill_1 FILLER_76_2000 ();
 sg13g2_fill_1 FILLER_76_2005 ();
 sg13g2_decap_4 FILLER_76_2010 ();
 sg13g2_fill_2 FILLER_76_2029 ();
 sg13g2_fill_1 FILLER_76_2031 ();
 sg13g2_decap_4 FILLER_76_2037 ();
 sg13g2_fill_1 FILLER_76_2041 ();
 sg13g2_fill_2 FILLER_76_2046 ();
 sg13g2_fill_1 FILLER_76_2048 ();
 sg13g2_fill_2 FILLER_76_2054 ();
 sg13g2_decap_4 FILLER_76_2064 ();
 sg13g2_fill_2 FILLER_76_2068 ();
 sg13g2_decap_4 FILLER_76_2074 ();
 sg13g2_fill_1 FILLER_76_2078 ();
 sg13g2_decap_8 FILLER_76_2082 ();
 sg13g2_decap_4 FILLER_76_2089 ();
 sg13g2_fill_1 FILLER_76_2093 ();
 sg13g2_decap_8 FILLER_76_2101 ();
 sg13g2_fill_1 FILLER_76_2117 ();
 sg13g2_decap_8 FILLER_76_2143 ();
 sg13g2_fill_2 FILLER_76_2167 ();
 sg13g2_fill_1 FILLER_76_2169 ();
 sg13g2_fill_2 FILLER_76_2186 ();
 sg13g2_fill_1 FILLER_76_2188 ();
 sg13g2_fill_2 FILLER_76_2208 ();
 sg13g2_fill_1 FILLER_76_2210 ();
 sg13g2_decap_8 FILLER_76_2239 ();
 sg13g2_decap_8 FILLER_76_2246 ();
 sg13g2_decap_8 FILLER_76_2253 ();
 sg13g2_decap_8 FILLER_76_2260 ();
 sg13g2_fill_2 FILLER_76_2267 ();
 sg13g2_fill_1 FILLER_76_2269 ();
 sg13g2_decap_4 FILLER_76_2287 ();
 sg13g2_fill_2 FILLER_76_2295 ();
 sg13g2_fill_1 FILLER_76_2325 ();
 sg13g2_decap_4 FILLER_76_2331 ();
 sg13g2_fill_1 FILLER_76_2335 ();
 sg13g2_fill_1 FILLER_76_2346 ();
 sg13g2_decap_4 FILLER_76_2388 ();
 sg13g2_fill_2 FILLER_76_2392 ();
 sg13g2_fill_2 FILLER_76_2422 ();
 sg13g2_fill_1 FILLER_76_2424 ();
 sg13g2_decap_8 FILLER_76_2429 ();
 sg13g2_decap_8 FILLER_76_2436 ();
 sg13g2_decap_8 FILLER_76_2443 ();
 sg13g2_decap_8 FILLER_76_2450 ();
 sg13g2_decap_8 FILLER_76_2457 ();
 sg13g2_decap_8 FILLER_76_2464 ();
 sg13g2_decap_8 FILLER_76_2471 ();
 sg13g2_decap_8 FILLER_76_2478 ();
 sg13g2_decap_8 FILLER_76_2485 ();
 sg13g2_decap_8 FILLER_76_2492 ();
 sg13g2_decap_8 FILLER_76_2499 ();
 sg13g2_decap_8 FILLER_76_2506 ();
 sg13g2_decap_8 FILLER_76_2513 ();
 sg13g2_decap_8 FILLER_76_2520 ();
 sg13g2_decap_8 FILLER_76_2527 ();
 sg13g2_decap_8 FILLER_76_2534 ();
 sg13g2_decap_8 FILLER_76_2545 ();
 sg13g2_fill_2 FILLER_76_2552 ();
 sg13g2_decap_4 FILLER_76_2614 ();
 sg13g2_decap_4 FILLER_76_2622 ();
 sg13g2_fill_2 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2684 ();
 sg13g2_decap_8 FILLER_76_2691 ();
 sg13g2_decap_8 FILLER_76_2698 ();
 sg13g2_fill_1 FILLER_76_2705 ();
 sg13g2_decap_8 FILLER_76_2734 ();
 sg13g2_decap_4 FILLER_76_2741 ();
 sg13g2_fill_1 FILLER_76_2745 ();
 sg13g2_fill_1 FILLER_76_2774 ();
 sg13g2_fill_2 FILLER_76_2812 ();
 sg13g2_fill_1 FILLER_76_2814 ();
 sg13g2_decap_8 FILLER_76_2837 ();
 sg13g2_decap_8 FILLER_76_2844 ();
 sg13g2_decap_8 FILLER_76_2851 ();
 sg13g2_decap_8 FILLER_76_2858 ();
 sg13g2_decap_8 FILLER_76_2865 ();
 sg13g2_decap_8 FILLER_76_2872 ();
 sg13g2_decap_8 FILLER_76_2879 ();
 sg13g2_decap_8 FILLER_76_2886 ();
 sg13g2_decap_8 FILLER_76_2893 ();
 sg13g2_decap_8 FILLER_76_2900 ();
 sg13g2_decap_8 FILLER_76_2907 ();
 sg13g2_decap_8 FILLER_76_2914 ();
 sg13g2_decap_8 FILLER_76_2921 ();
 sg13g2_fill_2 FILLER_76_2928 ();
 sg13g2_decap_8 FILLER_76_2934 ();
 sg13g2_decap_8 FILLER_76_2941 ();
 sg13g2_decap_8 FILLER_76_2948 ();
 sg13g2_decap_8 FILLER_76_2955 ();
 sg13g2_decap_8 FILLER_76_2962 ();
 sg13g2_decap_8 FILLER_76_2969 ();
 sg13g2_decap_8 FILLER_76_2976 ();
 sg13g2_decap_8 FILLER_76_2983 ();
 sg13g2_fill_2 FILLER_76_2990 ();
 sg13g2_decap_8 FILLER_76_2996 ();
 sg13g2_decap_4 FILLER_76_3003 ();
 sg13g2_fill_1 FILLER_76_3007 ();
 sg13g2_decap_8 FILLER_76_3017 ();
 sg13g2_fill_1 FILLER_76_3024 ();
 sg13g2_decap_8 FILLER_76_3029 ();
 sg13g2_decap_8 FILLER_76_3036 ();
 sg13g2_decap_8 FILLER_76_3043 ();
 sg13g2_decap_8 FILLER_76_3050 ();
 sg13g2_decap_8 FILLER_76_3057 ();
 sg13g2_decap_8 FILLER_76_3064 ();
 sg13g2_decap_8 FILLER_76_3071 ();
 sg13g2_decap_8 FILLER_76_3078 ();
 sg13g2_decap_8 FILLER_76_3085 ();
 sg13g2_decap_8 FILLER_76_3092 ();
 sg13g2_decap_8 FILLER_76_3099 ();
 sg13g2_decap_8 FILLER_76_3106 ();
 sg13g2_decap_8 FILLER_76_3113 ();
 sg13g2_decap_8 FILLER_76_3120 ();
 sg13g2_decap_8 FILLER_76_3127 ();
 sg13g2_decap_8 FILLER_76_3134 ();
 sg13g2_decap_8 FILLER_76_3141 ();
 sg13g2_decap_8 FILLER_76_3148 ();
 sg13g2_decap_8 FILLER_76_3155 ();
 sg13g2_decap_8 FILLER_76_3162 ();
 sg13g2_decap_8 FILLER_76_3169 ();
 sg13g2_decap_8 FILLER_76_3176 ();
 sg13g2_decap_8 FILLER_76_3183 ();
 sg13g2_decap_8 FILLER_76_3190 ();
 sg13g2_decap_8 FILLER_76_3197 ();
 sg13g2_decap_8 FILLER_76_3204 ();
 sg13g2_decap_8 FILLER_76_3211 ();
 sg13g2_decap_8 FILLER_76_3218 ();
 sg13g2_decap_8 FILLER_76_3225 ();
 sg13g2_decap_8 FILLER_76_3232 ();
 sg13g2_decap_8 FILLER_76_3239 ();
 sg13g2_decap_8 FILLER_76_3246 ();
 sg13g2_decap_8 FILLER_76_3253 ();
 sg13g2_decap_8 FILLER_76_3260 ();
 sg13g2_decap_8 FILLER_76_3267 ();
 sg13g2_decap_8 FILLER_76_3274 ();
 sg13g2_decap_8 FILLER_76_3281 ();
 sg13g2_decap_8 FILLER_76_3288 ();
 sg13g2_decap_8 FILLER_76_3295 ();
 sg13g2_decap_8 FILLER_76_3302 ();
 sg13g2_decap_8 FILLER_76_3309 ();
 sg13g2_decap_8 FILLER_76_3316 ();
 sg13g2_decap_8 FILLER_76_3323 ();
 sg13g2_decap_8 FILLER_76_3330 ();
 sg13g2_decap_8 FILLER_76_3337 ();
 sg13g2_decap_8 FILLER_76_3344 ();
 sg13g2_decap_8 FILLER_76_3351 ();
 sg13g2_decap_8 FILLER_76_3358 ();
 sg13g2_decap_8 FILLER_76_3365 ();
 sg13g2_decap_8 FILLER_76_3372 ();
 sg13g2_decap_8 FILLER_76_3379 ();
 sg13g2_decap_8 FILLER_76_3386 ();
 sg13g2_decap_8 FILLER_76_3393 ();
 sg13g2_decap_8 FILLER_76_3400 ();
 sg13g2_decap_8 FILLER_76_3407 ();
 sg13g2_decap_8 FILLER_76_3414 ();
 sg13g2_decap_8 FILLER_76_3421 ();
 sg13g2_decap_8 FILLER_76_3428 ();
 sg13g2_decap_8 FILLER_76_3435 ();
 sg13g2_decap_8 FILLER_76_3442 ();
 sg13g2_decap_8 FILLER_76_3449 ();
 sg13g2_decap_8 FILLER_76_3456 ();
 sg13g2_decap_8 FILLER_76_3463 ();
 sg13g2_decap_8 FILLER_76_3470 ();
 sg13g2_decap_8 FILLER_76_3477 ();
 sg13g2_decap_8 FILLER_76_3484 ();
 sg13g2_decap_8 FILLER_76_3491 ();
 sg13g2_decap_8 FILLER_76_3498 ();
 sg13g2_decap_8 FILLER_76_3505 ();
 sg13g2_decap_8 FILLER_76_3512 ();
 sg13g2_decap_8 FILLER_76_3519 ();
 sg13g2_decap_8 FILLER_76_3526 ();
 sg13g2_decap_8 FILLER_76_3533 ();
 sg13g2_decap_8 FILLER_76_3540 ();
 sg13g2_decap_8 FILLER_76_3547 ();
 sg13g2_decap_8 FILLER_76_3554 ();
 sg13g2_decap_8 FILLER_76_3561 ();
 sg13g2_decap_8 FILLER_76_3568 ();
 sg13g2_decap_4 FILLER_76_3575 ();
 sg13g2_fill_1 FILLER_76_3579 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_4 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_466 ();
 sg13g2_decap_8 FILLER_77_472 ();
 sg13g2_decap_8 FILLER_77_479 ();
 sg13g2_fill_1 FILLER_77_486 ();
 sg13g2_fill_1 FILLER_77_552 ();
 sg13g2_fill_1 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_fill_2 FILLER_77_659 ();
 sg13g2_fill_1 FILLER_77_668 ();
 sg13g2_decap_4 FILLER_77_711 ();
 sg13g2_fill_1 FILLER_77_715 ();
 sg13g2_fill_2 FILLER_77_740 ();
 sg13g2_fill_1 FILLER_77_836 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_2 FILLER_77_861 ();
 sg13g2_fill_1 FILLER_77_863 ();
 sg13g2_decap_8 FILLER_77_898 ();
 sg13g2_fill_1 FILLER_77_918 ();
 sg13g2_decap_8 FILLER_77_927 ();
 sg13g2_fill_2 FILLER_77_934 ();
 sg13g2_fill_1 FILLER_77_936 ();
 sg13g2_fill_2 FILLER_77_1008 ();
 sg13g2_decap_8 FILLER_77_1019 ();
 sg13g2_decap_8 FILLER_77_1026 ();
 sg13g2_decap_8 FILLER_77_1037 ();
 sg13g2_decap_8 FILLER_77_1044 ();
 sg13g2_decap_8 FILLER_77_1051 ();
 sg13g2_fill_1 FILLER_77_1074 ();
 sg13g2_fill_2 FILLER_77_1089 ();
 sg13g2_fill_1 FILLER_77_1091 ();
 sg13g2_decap_4 FILLER_77_1107 ();
 sg13g2_fill_1 FILLER_77_1130 ();
 sg13g2_fill_1 FILLER_77_1135 ();
 sg13g2_fill_2 FILLER_77_1151 ();
 sg13g2_fill_1 FILLER_77_1153 ();
 sg13g2_decap_8 FILLER_77_1175 ();
 sg13g2_decap_8 FILLER_77_1182 ();
 sg13g2_fill_1 FILLER_77_1189 ();
 sg13g2_fill_1 FILLER_77_1227 ();
 sg13g2_fill_1 FILLER_77_1237 ();
 sg13g2_fill_2 FILLER_77_1252 ();
 sg13g2_fill_1 FILLER_77_1254 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_4 FILLER_77_1271 ();
 sg13g2_decap_4 FILLER_77_1280 ();
 sg13g2_fill_1 FILLER_77_1284 ();
 sg13g2_decap_4 FILLER_77_1290 ();
 sg13g2_fill_1 FILLER_77_1294 ();
 sg13g2_fill_1 FILLER_77_1308 ();
 sg13g2_fill_2 FILLER_77_1321 ();
 sg13g2_fill_1 FILLER_77_1323 ();
 sg13g2_decap_4 FILLER_77_1329 ();
 sg13g2_fill_1 FILLER_77_1333 ();
 sg13g2_fill_1 FILLER_77_1407 ();
 sg13g2_decap_4 FILLER_77_1430 ();
 sg13g2_decap_8 FILLER_77_1443 ();
 sg13g2_fill_2 FILLER_77_1450 ();
 sg13g2_fill_1 FILLER_77_1457 ();
 sg13g2_fill_2 FILLER_77_1477 ();
 sg13g2_fill_2 FILLER_77_1500 ();
 sg13g2_decap_4 FILLER_77_1597 ();
 sg13g2_fill_1 FILLER_77_1610 ();
 sg13g2_fill_1 FILLER_77_1625 ();
 sg13g2_fill_1 FILLER_77_1634 ();
 sg13g2_fill_2 FILLER_77_1643 ();
 sg13g2_decap_4 FILLER_77_1657 ();
 sg13g2_decap_8 FILLER_77_1677 ();
 sg13g2_decap_8 FILLER_77_1684 ();
 sg13g2_fill_1 FILLER_77_1691 ();
 sg13g2_decap_8 FILLER_77_1727 ();
 sg13g2_decap_8 FILLER_77_1734 ();
 sg13g2_decap_8 FILLER_77_1741 ();
 sg13g2_decap_8 FILLER_77_1748 ();
 sg13g2_decap_8 FILLER_77_1755 ();
 sg13g2_decap_8 FILLER_77_1762 ();
 sg13g2_decap_8 FILLER_77_1769 ();
 sg13g2_decap_8 FILLER_77_1776 ();
 sg13g2_decap_8 FILLER_77_1783 ();
 sg13g2_decap_8 FILLER_77_1790 ();
 sg13g2_decap_4 FILLER_77_1797 ();
 sg13g2_decap_4 FILLER_77_1805 ();
 sg13g2_decap_8 FILLER_77_1818 ();
 sg13g2_decap_8 FILLER_77_1825 ();
 sg13g2_decap_4 FILLER_77_1832 ();
 sg13g2_decap_8 FILLER_77_1840 ();
 sg13g2_fill_2 FILLER_77_1847 ();
 sg13g2_fill_1 FILLER_77_1849 ();
 sg13g2_fill_2 FILLER_77_1867 ();
 sg13g2_fill_1 FILLER_77_1869 ();
 sg13g2_decap_8 FILLER_77_1898 ();
 sg13g2_fill_1 FILLER_77_1905 ();
 sg13g2_decap_4 FILLER_77_1915 ();
 sg13g2_fill_1 FILLER_77_1965 ();
 sg13g2_fill_2 FILLER_77_2009 ();
 sg13g2_fill_2 FILLER_77_2029 ();
 sg13g2_fill_1 FILLER_77_2031 ();
 sg13g2_fill_2 FILLER_77_2052 ();
 sg13g2_fill_1 FILLER_77_2054 ();
 sg13g2_fill_2 FILLER_77_2118 ();
 sg13g2_fill_1 FILLER_77_2120 ();
 sg13g2_fill_1 FILLER_77_2139 ();
 sg13g2_fill_2 FILLER_77_2172 ();
 sg13g2_fill_2 FILLER_77_2179 ();
 sg13g2_fill_2 FILLER_77_2194 ();
 sg13g2_fill_1 FILLER_77_2196 ();
 sg13g2_decap_8 FILLER_77_2200 ();
 sg13g2_fill_2 FILLER_77_2207 ();
 sg13g2_fill_1 FILLER_77_2209 ();
 sg13g2_fill_1 FILLER_77_2214 ();
 sg13g2_fill_1 FILLER_77_2224 ();
 sg13g2_decap_8 FILLER_77_2234 ();
 sg13g2_decap_8 FILLER_77_2241 ();
 sg13g2_decap_8 FILLER_77_2248 ();
 sg13g2_decap_8 FILLER_77_2255 ();
 sg13g2_decap_8 FILLER_77_2262 ();
 sg13g2_decap_8 FILLER_77_2269 ();
 sg13g2_decap_8 FILLER_77_2276 ();
 sg13g2_fill_2 FILLER_77_2283 ();
 sg13g2_fill_1 FILLER_77_2285 ();
 sg13g2_fill_2 FILLER_77_2316 ();
 sg13g2_fill_1 FILLER_77_2318 ();
 sg13g2_decap_8 FILLER_77_2360 ();
 sg13g2_fill_1 FILLER_77_2367 ();
 sg13g2_decap_8 FILLER_77_2414 ();
 sg13g2_decap_8 FILLER_77_2421 ();
 sg13g2_decap_8 FILLER_77_2428 ();
 sg13g2_decap_8 FILLER_77_2435 ();
 sg13g2_decap_8 FILLER_77_2442 ();
 sg13g2_decap_8 FILLER_77_2449 ();
 sg13g2_decap_8 FILLER_77_2456 ();
 sg13g2_decap_8 FILLER_77_2463 ();
 sg13g2_decap_8 FILLER_77_2470 ();
 sg13g2_decap_8 FILLER_77_2477 ();
 sg13g2_decap_8 FILLER_77_2484 ();
 sg13g2_decap_8 FILLER_77_2491 ();
 sg13g2_decap_8 FILLER_77_2498 ();
 sg13g2_decap_8 FILLER_77_2505 ();
 sg13g2_decap_8 FILLER_77_2512 ();
 sg13g2_decap_8 FILLER_77_2519 ();
 sg13g2_decap_8 FILLER_77_2526 ();
 sg13g2_decap_8 FILLER_77_2533 ();
 sg13g2_decap_8 FILLER_77_2540 ();
 sg13g2_decap_8 FILLER_77_2547 ();
 sg13g2_decap_4 FILLER_77_2554 ();
 sg13g2_fill_1 FILLER_77_2558 ();
 sg13g2_decap_8 FILLER_77_2563 ();
 sg13g2_decap_8 FILLER_77_2570 ();
 sg13g2_decap_8 FILLER_77_2577 ();
 sg13g2_decap_8 FILLER_77_2584 ();
 sg13g2_decap_8 FILLER_77_2591 ();
 sg13g2_decap_8 FILLER_77_2598 ();
 sg13g2_decap_8 FILLER_77_2605 ();
 sg13g2_decap_8 FILLER_77_2612 ();
 sg13g2_decap_8 FILLER_77_2619 ();
 sg13g2_fill_2 FILLER_77_2626 ();
 sg13g2_fill_2 FILLER_77_2638 ();
 sg13g2_fill_1 FILLER_77_2640 ();
 sg13g2_decap_8 FILLER_77_2648 ();
 sg13g2_decap_8 FILLER_77_2655 ();
 sg13g2_decap_8 FILLER_77_2662 ();
 sg13g2_decap_8 FILLER_77_2669 ();
 sg13g2_fill_2 FILLER_77_2676 ();
 sg13g2_decap_8 FILLER_77_2715 ();
 sg13g2_decap_8 FILLER_77_2722 ();
 sg13g2_decap_8 FILLER_77_2729 ();
 sg13g2_decap_8 FILLER_77_2736 ();
 sg13g2_decap_8 FILLER_77_2743 ();
 sg13g2_decap_8 FILLER_77_2750 ();
 sg13g2_decap_8 FILLER_77_2757 ();
 sg13g2_decap_8 FILLER_77_2764 ();
 sg13g2_decap_8 FILLER_77_2771 ();
 sg13g2_decap_8 FILLER_77_2778 ();
 sg13g2_decap_8 FILLER_77_2785 ();
 sg13g2_fill_2 FILLER_77_2792 ();
 sg13g2_fill_1 FILLER_77_2794 ();
 sg13g2_decap_8 FILLER_77_2822 ();
 sg13g2_decap_8 FILLER_77_2829 ();
 sg13g2_decap_8 FILLER_77_2836 ();
 sg13g2_decap_8 FILLER_77_2843 ();
 sg13g2_decap_8 FILLER_77_2850 ();
 sg13g2_decap_8 FILLER_77_2857 ();
 sg13g2_decap_8 FILLER_77_2864 ();
 sg13g2_decap_8 FILLER_77_2871 ();
 sg13g2_decap_8 FILLER_77_2878 ();
 sg13g2_decap_8 FILLER_77_2885 ();
 sg13g2_decap_8 FILLER_77_2892 ();
 sg13g2_decap_8 FILLER_77_2899 ();
 sg13g2_decap_8 FILLER_77_2906 ();
 sg13g2_decap_8 FILLER_77_2913 ();
 sg13g2_decap_8 FILLER_77_2920 ();
 sg13g2_decap_8 FILLER_77_2927 ();
 sg13g2_decap_8 FILLER_77_2934 ();
 sg13g2_decap_8 FILLER_77_2941 ();
 sg13g2_decap_8 FILLER_77_2948 ();
 sg13g2_decap_8 FILLER_77_2955 ();
 sg13g2_decap_8 FILLER_77_2962 ();
 sg13g2_decap_8 FILLER_77_2969 ();
 sg13g2_decap_8 FILLER_77_2976 ();
 sg13g2_decap_8 FILLER_77_2983 ();
 sg13g2_decap_8 FILLER_77_2990 ();
 sg13g2_decap_8 FILLER_77_2997 ();
 sg13g2_decap_8 FILLER_77_3004 ();
 sg13g2_decap_8 FILLER_77_3011 ();
 sg13g2_decap_8 FILLER_77_3018 ();
 sg13g2_decap_8 FILLER_77_3025 ();
 sg13g2_decap_8 FILLER_77_3032 ();
 sg13g2_decap_8 FILLER_77_3039 ();
 sg13g2_decap_8 FILLER_77_3046 ();
 sg13g2_decap_8 FILLER_77_3053 ();
 sg13g2_decap_8 FILLER_77_3060 ();
 sg13g2_decap_8 FILLER_77_3067 ();
 sg13g2_decap_8 FILLER_77_3074 ();
 sg13g2_decap_8 FILLER_77_3081 ();
 sg13g2_decap_8 FILLER_77_3088 ();
 sg13g2_decap_8 FILLER_77_3095 ();
 sg13g2_decap_8 FILLER_77_3102 ();
 sg13g2_decap_8 FILLER_77_3109 ();
 sg13g2_decap_8 FILLER_77_3116 ();
 sg13g2_decap_8 FILLER_77_3123 ();
 sg13g2_decap_8 FILLER_77_3130 ();
 sg13g2_decap_8 FILLER_77_3137 ();
 sg13g2_decap_8 FILLER_77_3144 ();
 sg13g2_decap_8 FILLER_77_3151 ();
 sg13g2_decap_8 FILLER_77_3158 ();
 sg13g2_decap_8 FILLER_77_3165 ();
 sg13g2_decap_8 FILLER_77_3172 ();
 sg13g2_decap_8 FILLER_77_3179 ();
 sg13g2_decap_8 FILLER_77_3186 ();
 sg13g2_decap_8 FILLER_77_3193 ();
 sg13g2_decap_8 FILLER_77_3200 ();
 sg13g2_decap_8 FILLER_77_3207 ();
 sg13g2_decap_8 FILLER_77_3214 ();
 sg13g2_decap_8 FILLER_77_3221 ();
 sg13g2_decap_8 FILLER_77_3228 ();
 sg13g2_decap_8 FILLER_77_3235 ();
 sg13g2_decap_8 FILLER_77_3242 ();
 sg13g2_decap_8 FILLER_77_3249 ();
 sg13g2_decap_8 FILLER_77_3256 ();
 sg13g2_decap_8 FILLER_77_3263 ();
 sg13g2_decap_8 FILLER_77_3270 ();
 sg13g2_decap_8 FILLER_77_3277 ();
 sg13g2_decap_8 FILLER_77_3284 ();
 sg13g2_decap_8 FILLER_77_3291 ();
 sg13g2_decap_8 FILLER_77_3298 ();
 sg13g2_decap_8 FILLER_77_3305 ();
 sg13g2_decap_8 FILLER_77_3312 ();
 sg13g2_decap_8 FILLER_77_3319 ();
 sg13g2_decap_8 FILLER_77_3326 ();
 sg13g2_decap_8 FILLER_77_3333 ();
 sg13g2_decap_8 FILLER_77_3340 ();
 sg13g2_decap_8 FILLER_77_3347 ();
 sg13g2_decap_8 FILLER_77_3354 ();
 sg13g2_decap_8 FILLER_77_3361 ();
 sg13g2_decap_8 FILLER_77_3368 ();
 sg13g2_decap_8 FILLER_77_3375 ();
 sg13g2_decap_8 FILLER_77_3382 ();
 sg13g2_decap_8 FILLER_77_3389 ();
 sg13g2_decap_8 FILLER_77_3396 ();
 sg13g2_decap_8 FILLER_77_3403 ();
 sg13g2_decap_8 FILLER_77_3410 ();
 sg13g2_decap_8 FILLER_77_3417 ();
 sg13g2_decap_8 FILLER_77_3424 ();
 sg13g2_decap_8 FILLER_77_3431 ();
 sg13g2_decap_8 FILLER_77_3438 ();
 sg13g2_decap_8 FILLER_77_3445 ();
 sg13g2_decap_8 FILLER_77_3452 ();
 sg13g2_decap_8 FILLER_77_3459 ();
 sg13g2_decap_8 FILLER_77_3466 ();
 sg13g2_decap_8 FILLER_77_3473 ();
 sg13g2_decap_8 FILLER_77_3480 ();
 sg13g2_decap_8 FILLER_77_3487 ();
 sg13g2_decap_8 FILLER_77_3494 ();
 sg13g2_decap_8 FILLER_77_3501 ();
 sg13g2_decap_8 FILLER_77_3508 ();
 sg13g2_decap_8 FILLER_77_3515 ();
 sg13g2_decap_8 FILLER_77_3522 ();
 sg13g2_decap_8 FILLER_77_3529 ();
 sg13g2_decap_8 FILLER_77_3536 ();
 sg13g2_decap_8 FILLER_77_3543 ();
 sg13g2_decap_8 FILLER_77_3550 ();
 sg13g2_decap_8 FILLER_77_3557 ();
 sg13g2_decap_8 FILLER_77_3564 ();
 sg13g2_decap_8 FILLER_77_3571 ();
 sg13g2_fill_2 FILLER_77_3578 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_4 FILLER_78_511 ();
 sg13g2_fill_1 FILLER_78_515 ();
 sg13g2_decap_8 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_536 ();
 sg13g2_decap_8 FILLER_78_543 ();
 sg13g2_fill_1 FILLER_78_550 ();
 sg13g2_fill_1 FILLER_78_569 ();
 sg13g2_fill_1 FILLER_78_579 ();
 sg13g2_decap_8 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_610 ();
 sg13g2_decap_4 FILLER_78_617 ();
 sg13g2_fill_1 FILLER_78_621 ();
 sg13g2_decap_8 FILLER_78_647 ();
 sg13g2_fill_2 FILLER_78_654 ();
 sg13g2_fill_1 FILLER_78_656 ();
 sg13g2_decap_4 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_683 ();
 sg13g2_decap_4 FILLER_78_690 ();
 sg13g2_fill_2 FILLER_78_726 ();
 sg13g2_fill_1 FILLER_78_728 ();
 sg13g2_fill_1 FILLER_78_733 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_fill_1 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_750 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_4 FILLER_78_784 ();
 sg13g2_fill_1 FILLER_78_788 ();
 sg13g2_fill_2 FILLER_78_832 ();
 sg13g2_fill_1 FILLER_78_834 ();
 sg13g2_fill_2 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_fill_2 FILLER_78_857 ();
 sg13g2_fill_1 FILLER_78_881 ();
 sg13g2_fill_2 FILLER_78_896 ();
 sg13g2_fill_2 FILLER_78_902 ();
 sg13g2_fill_1 FILLER_78_904 ();
 sg13g2_decap_4 FILLER_78_911 ();
 sg13g2_decap_8 FILLER_78_943 ();
 sg13g2_decap_8 FILLER_78_950 ();
 sg13g2_decap_8 FILLER_78_957 ();
 sg13g2_decap_8 FILLER_78_964 ();
 sg13g2_decap_8 FILLER_78_971 ();
 sg13g2_decap_8 FILLER_78_978 ();
 sg13g2_decap_4 FILLER_78_985 ();
 sg13g2_fill_2 FILLER_78_989 ();
 sg13g2_decap_4 FILLER_78_1022 ();
 sg13g2_fill_2 FILLER_78_1026 ();
 sg13g2_fill_1 FILLER_78_1055 ();
 sg13g2_decap_4 FILLER_78_1084 ();
 sg13g2_fill_1 FILLER_78_1088 ();
 sg13g2_decap_4 FILLER_78_1093 ();
 sg13g2_fill_1 FILLER_78_1097 ();
 sg13g2_fill_2 FILLER_78_1102 ();
 sg13g2_fill_1 FILLER_78_1104 ();
 sg13g2_decap_4 FILLER_78_1114 ();
 sg13g2_decap_4 FILLER_78_1131 ();
 sg13g2_decap_4 FILLER_78_1138 ();
 sg13g2_fill_1 FILLER_78_1142 ();
 sg13g2_decap_8 FILLER_78_1170 ();
 sg13g2_decap_8 FILLER_78_1177 ();
 sg13g2_decap_8 FILLER_78_1184 ();
 sg13g2_decap_4 FILLER_78_1191 ();
 sg13g2_decap_8 FILLER_78_1199 ();
 sg13g2_decap_8 FILLER_78_1206 ();
 sg13g2_decap_4 FILLER_78_1213 ();
 sg13g2_fill_2 FILLER_78_1217 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_4 FILLER_78_1282 ();
 sg13g2_fill_2 FILLER_78_1312 ();
 sg13g2_fill_2 FILLER_78_1320 ();
 sg13g2_fill_1 FILLER_78_1322 ();
 sg13g2_decap_8 FILLER_78_1358 ();
 sg13g2_decap_8 FILLER_78_1365 ();
 sg13g2_decap_4 FILLER_78_1372 ();
 sg13g2_fill_2 FILLER_78_1376 ();
 sg13g2_decap_4 FILLER_78_1391 ();
 sg13g2_fill_2 FILLER_78_1395 ();
 sg13g2_fill_2 FILLER_78_1400 ();
 sg13g2_decap_4 FILLER_78_1406 ();
 sg13g2_decap_4 FILLER_78_1446 ();
 sg13g2_fill_2 FILLER_78_1450 ();
 sg13g2_decap_8 FILLER_78_1473 ();
 sg13g2_decap_8 FILLER_78_1480 ();
 sg13g2_decap_8 FILLER_78_1492 ();
 sg13g2_decap_8 FILLER_78_1499 ();
 sg13g2_decap_4 FILLER_78_1506 ();
 sg13g2_fill_1 FILLER_78_1510 ();
 sg13g2_decap_8 FILLER_78_1515 ();
 sg13g2_decap_8 FILLER_78_1522 ();
 sg13g2_decap_8 FILLER_78_1529 ();
 sg13g2_decap_8 FILLER_78_1536 ();
 sg13g2_fill_1 FILLER_78_1543 ();
 sg13g2_fill_1 FILLER_78_1624 ();
 sg13g2_fill_1 FILLER_78_1634 ();
 sg13g2_decap_4 FILLER_78_1638 ();
 sg13g2_fill_2 FILLER_78_1651 ();
 sg13g2_fill_1 FILLER_78_1703 ();
 sg13g2_fill_2 FILLER_78_1708 ();
 sg13g2_decap_8 FILLER_78_1719 ();
 sg13g2_decap_8 FILLER_78_1726 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_8 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1754 ();
 sg13g2_decap_8 FILLER_78_1761 ();
 sg13g2_decap_8 FILLER_78_1768 ();
 sg13g2_decap_8 FILLER_78_1775 ();
 sg13g2_decap_8 FILLER_78_1782 ();
 sg13g2_decap_8 FILLER_78_1789 ();
 sg13g2_decap_8 FILLER_78_1796 ();
 sg13g2_decap_8 FILLER_78_1803 ();
 sg13g2_decap_8 FILLER_78_1810 ();
 sg13g2_decap_8 FILLER_78_1817 ();
 sg13g2_decap_8 FILLER_78_1824 ();
 sg13g2_decap_8 FILLER_78_1831 ();
 sg13g2_decap_8 FILLER_78_1838 ();
 sg13g2_decap_8 FILLER_78_1845 ();
 sg13g2_decap_8 FILLER_78_1852 ();
 sg13g2_decap_8 FILLER_78_1859 ();
 sg13g2_fill_2 FILLER_78_1866 ();
 sg13g2_fill_1 FILLER_78_1868 ();
 sg13g2_decap_4 FILLER_78_1931 ();
 sg13g2_fill_2 FILLER_78_1935 ();
 sg13g2_decap_4 FILLER_78_1974 ();
 sg13g2_fill_1 FILLER_78_1978 ();
 sg13g2_fill_1 FILLER_78_1988 ();
 sg13g2_decap_8 FILLER_78_2025 ();
 sg13g2_fill_1 FILLER_78_2032 ();
 sg13g2_decap_8 FILLER_78_2053 ();
 sg13g2_decap_8 FILLER_78_2060 ();
 sg13g2_decap_4 FILLER_78_2067 ();
 sg13g2_fill_1 FILLER_78_2071 ();
 sg13g2_decap_4 FILLER_78_2099 ();
 sg13g2_fill_2 FILLER_78_2103 ();
 sg13g2_decap_8 FILLER_78_2109 ();
 sg13g2_fill_2 FILLER_78_2116 ();
 sg13g2_decap_4 FILLER_78_2138 ();
 sg13g2_fill_1 FILLER_78_2151 ();
 sg13g2_decap_4 FILLER_78_2163 ();
 sg13g2_fill_2 FILLER_78_2167 ();
 sg13g2_fill_2 FILLER_78_2181 ();
 sg13g2_fill_2 FILLER_78_2202 ();
 sg13g2_decap_8 FILLER_78_2232 ();
 sg13g2_decap_8 FILLER_78_2239 ();
 sg13g2_decap_8 FILLER_78_2246 ();
 sg13g2_decap_8 FILLER_78_2253 ();
 sg13g2_decap_8 FILLER_78_2260 ();
 sg13g2_decap_8 FILLER_78_2267 ();
 sg13g2_decap_8 FILLER_78_2274 ();
 sg13g2_decap_8 FILLER_78_2281 ();
 sg13g2_decap_8 FILLER_78_2288 ();
 sg13g2_fill_2 FILLER_78_2295 ();
 sg13g2_decap_8 FILLER_78_2306 ();
 sg13g2_decap_8 FILLER_78_2313 ();
 sg13g2_decap_4 FILLER_78_2320 ();
 sg13g2_decap_8 FILLER_78_2328 ();
 sg13g2_decap_8 FILLER_78_2335 ();
 sg13g2_fill_1 FILLER_78_2342 ();
 sg13g2_fill_2 FILLER_78_2371 ();
 sg13g2_fill_1 FILLER_78_2373 ();
 sg13g2_decap_4 FILLER_78_2378 ();
 sg13g2_decap_8 FILLER_78_2395 ();
 sg13g2_decap_8 FILLER_78_2402 ();
 sg13g2_decap_8 FILLER_78_2409 ();
 sg13g2_decap_8 FILLER_78_2416 ();
 sg13g2_decap_8 FILLER_78_2423 ();
 sg13g2_decap_8 FILLER_78_2430 ();
 sg13g2_decap_8 FILLER_78_2437 ();
 sg13g2_decap_8 FILLER_78_2444 ();
 sg13g2_decap_8 FILLER_78_2451 ();
 sg13g2_decap_8 FILLER_78_2458 ();
 sg13g2_decap_8 FILLER_78_2465 ();
 sg13g2_decap_8 FILLER_78_2472 ();
 sg13g2_decap_8 FILLER_78_2479 ();
 sg13g2_decap_8 FILLER_78_2486 ();
 sg13g2_decap_8 FILLER_78_2493 ();
 sg13g2_decap_8 FILLER_78_2500 ();
 sg13g2_decap_8 FILLER_78_2507 ();
 sg13g2_decap_8 FILLER_78_2514 ();
 sg13g2_decap_8 FILLER_78_2521 ();
 sg13g2_decap_8 FILLER_78_2528 ();
 sg13g2_decap_8 FILLER_78_2535 ();
 sg13g2_decap_8 FILLER_78_2542 ();
 sg13g2_decap_8 FILLER_78_2549 ();
 sg13g2_decap_8 FILLER_78_2556 ();
 sg13g2_decap_8 FILLER_78_2563 ();
 sg13g2_decap_8 FILLER_78_2570 ();
 sg13g2_decap_8 FILLER_78_2577 ();
 sg13g2_decap_8 FILLER_78_2584 ();
 sg13g2_decap_8 FILLER_78_2591 ();
 sg13g2_decap_8 FILLER_78_2598 ();
 sg13g2_decap_8 FILLER_78_2605 ();
 sg13g2_decap_8 FILLER_78_2612 ();
 sg13g2_decap_8 FILLER_78_2619 ();
 sg13g2_decap_8 FILLER_78_2626 ();
 sg13g2_decap_8 FILLER_78_2633 ();
 sg13g2_decap_8 FILLER_78_2640 ();
 sg13g2_decap_8 FILLER_78_2647 ();
 sg13g2_decap_8 FILLER_78_2654 ();
 sg13g2_decap_8 FILLER_78_2661 ();
 sg13g2_decap_8 FILLER_78_2668 ();
 sg13g2_decap_8 FILLER_78_2675 ();
 sg13g2_fill_1 FILLER_78_2682 ();
 sg13g2_decap_8 FILLER_78_2687 ();
 sg13g2_decap_8 FILLER_78_2694 ();
 sg13g2_decap_8 FILLER_78_2701 ();
 sg13g2_decap_8 FILLER_78_2708 ();
 sg13g2_decap_8 FILLER_78_2715 ();
 sg13g2_decap_8 FILLER_78_2722 ();
 sg13g2_decap_8 FILLER_78_2729 ();
 sg13g2_decap_8 FILLER_78_2736 ();
 sg13g2_decap_8 FILLER_78_2743 ();
 sg13g2_decap_8 FILLER_78_2750 ();
 sg13g2_decap_8 FILLER_78_2757 ();
 sg13g2_decap_8 FILLER_78_2764 ();
 sg13g2_decap_8 FILLER_78_2771 ();
 sg13g2_decap_8 FILLER_78_2778 ();
 sg13g2_decap_8 FILLER_78_2785 ();
 sg13g2_decap_8 FILLER_78_2792 ();
 sg13g2_fill_1 FILLER_78_2799 ();
 sg13g2_decap_8 FILLER_78_2804 ();
 sg13g2_decap_8 FILLER_78_2811 ();
 sg13g2_decap_8 FILLER_78_2818 ();
 sg13g2_decap_8 FILLER_78_2825 ();
 sg13g2_decap_8 FILLER_78_2832 ();
 sg13g2_decap_8 FILLER_78_2839 ();
 sg13g2_decap_8 FILLER_78_2846 ();
 sg13g2_decap_8 FILLER_78_2853 ();
 sg13g2_decap_8 FILLER_78_2860 ();
 sg13g2_decap_8 FILLER_78_2867 ();
 sg13g2_decap_8 FILLER_78_2874 ();
 sg13g2_decap_8 FILLER_78_2881 ();
 sg13g2_decap_8 FILLER_78_2888 ();
 sg13g2_decap_8 FILLER_78_2895 ();
 sg13g2_decap_8 FILLER_78_2902 ();
 sg13g2_decap_8 FILLER_78_2909 ();
 sg13g2_decap_8 FILLER_78_2916 ();
 sg13g2_decap_8 FILLER_78_2923 ();
 sg13g2_decap_8 FILLER_78_2930 ();
 sg13g2_decap_8 FILLER_78_2937 ();
 sg13g2_decap_8 FILLER_78_2944 ();
 sg13g2_decap_8 FILLER_78_2951 ();
 sg13g2_decap_8 FILLER_78_2958 ();
 sg13g2_decap_8 FILLER_78_2965 ();
 sg13g2_decap_8 FILLER_78_2972 ();
 sg13g2_decap_8 FILLER_78_2979 ();
 sg13g2_decap_8 FILLER_78_2986 ();
 sg13g2_decap_8 FILLER_78_2993 ();
 sg13g2_decap_8 FILLER_78_3000 ();
 sg13g2_decap_8 FILLER_78_3007 ();
 sg13g2_decap_8 FILLER_78_3014 ();
 sg13g2_decap_8 FILLER_78_3021 ();
 sg13g2_decap_8 FILLER_78_3028 ();
 sg13g2_decap_8 FILLER_78_3035 ();
 sg13g2_decap_8 FILLER_78_3042 ();
 sg13g2_decap_8 FILLER_78_3049 ();
 sg13g2_decap_8 FILLER_78_3056 ();
 sg13g2_decap_8 FILLER_78_3063 ();
 sg13g2_decap_8 FILLER_78_3070 ();
 sg13g2_decap_8 FILLER_78_3077 ();
 sg13g2_decap_8 FILLER_78_3084 ();
 sg13g2_decap_8 FILLER_78_3091 ();
 sg13g2_decap_8 FILLER_78_3098 ();
 sg13g2_decap_8 FILLER_78_3105 ();
 sg13g2_decap_8 FILLER_78_3112 ();
 sg13g2_decap_8 FILLER_78_3119 ();
 sg13g2_decap_8 FILLER_78_3126 ();
 sg13g2_decap_8 FILLER_78_3133 ();
 sg13g2_decap_8 FILLER_78_3140 ();
 sg13g2_decap_8 FILLER_78_3147 ();
 sg13g2_decap_8 FILLER_78_3154 ();
 sg13g2_decap_8 FILLER_78_3161 ();
 sg13g2_decap_8 FILLER_78_3168 ();
 sg13g2_decap_8 FILLER_78_3175 ();
 sg13g2_decap_8 FILLER_78_3182 ();
 sg13g2_decap_8 FILLER_78_3189 ();
 sg13g2_decap_8 FILLER_78_3196 ();
 sg13g2_decap_8 FILLER_78_3203 ();
 sg13g2_decap_8 FILLER_78_3210 ();
 sg13g2_decap_8 FILLER_78_3217 ();
 sg13g2_decap_8 FILLER_78_3224 ();
 sg13g2_decap_8 FILLER_78_3231 ();
 sg13g2_decap_8 FILLER_78_3238 ();
 sg13g2_decap_8 FILLER_78_3245 ();
 sg13g2_decap_8 FILLER_78_3252 ();
 sg13g2_decap_8 FILLER_78_3259 ();
 sg13g2_decap_8 FILLER_78_3266 ();
 sg13g2_decap_8 FILLER_78_3273 ();
 sg13g2_decap_8 FILLER_78_3280 ();
 sg13g2_decap_8 FILLER_78_3287 ();
 sg13g2_decap_8 FILLER_78_3294 ();
 sg13g2_decap_8 FILLER_78_3301 ();
 sg13g2_decap_8 FILLER_78_3308 ();
 sg13g2_decap_8 FILLER_78_3315 ();
 sg13g2_decap_8 FILLER_78_3322 ();
 sg13g2_decap_8 FILLER_78_3329 ();
 sg13g2_decap_8 FILLER_78_3336 ();
 sg13g2_decap_8 FILLER_78_3343 ();
 sg13g2_decap_8 FILLER_78_3350 ();
 sg13g2_decap_8 FILLER_78_3357 ();
 sg13g2_decap_8 FILLER_78_3364 ();
 sg13g2_decap_8 FILLER_78_3371 ();
 sg13g2_decap_8 FILLER_78_3378 ();
 sg13g2_decap_8 FILLER_78_3385 ();
 sg13g2_decap_8 FILLER_78_3392 ();
 sg13g2_decap_8 FILLER_78_3399 ();
 sg13g2_decap_8 FILLER_78_3406 ();
 sg13g2_decap_8 FILLER_78_3413 ();
 sg13g2_decap_8 FILLER_78_3420 ();
 sg13g2_decap_8 FILLER_78_3427 ();
 sg13g2_decap_8 FILLER_78_3434 ();
 sg13g2_decap_8 FILLER_78_3441 ();
 sg13g2_decap_8 FILLER_78_3448 ();
 sg13g2_decap_8 FILLER_78_3455 ();
 sg13g2_decap_8 FILLER_78_3462 ();
 sg13g2_decap_8 FILLER_78_3469 ();
 sg13g2_decap_8 FILLER_78_3476 ();
 sg13g2_decap_8 FILLER_78_3483 ();
 sg13g2_decap_8 FILLER_78_3490 ();
 sg13g2_decap_8 FILLER_78_3497 ();
 sg13g2_decap_8 FILLER_78_3504 ();
 sg13g2_decap_8 FILLER_78_3511 ();
 sg13g2_decap_8 FILLER_78_3518 ();
 sg13g2_decap_8 FILLER_78_3525 ();
 sg13g2_decap_8 FILLER_78_3532 ();
 sg13g2_decap_8 FILLER_78_3539 ();
 sg13g2_decap_8 FILLER_78_3546 ();
 sg13g2_decap_8 FILLER_78_3553 ();
 sg13g2_decap_8 FILLER_78_3560 ();
 sg13g2_decap_8 FILLER_78_3567 ();
 sg13g2_decap_4 FILLER_78_3574 ();
 sg13g2_fill_2 FILLER_78_3578 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_fill_2 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_604 ();
 sg13g2_decap_8 FILLER_79_611 ();
 sg13g2_decap_4 FILLER_79_618 ();
 sg13g2_fill_1 FILLER_79_622 ();
 sg13g2_fill_2 FILLER_79_650 ();
 sg13g2_fill_2 FILLER_79_701 ();
 sg13g2_fill_2 FILLER_79_737 ();
 sg13g2_fill_1 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_decap_8 FILLER_79_775 ();
 sg13g2_fill_2 FILLER_79_782 ();
 sg13g2_fill_1 FILLER_79_784 ();
 sg13g2_fill_2 FILLER_79_821 ();
 sg13g2_fill_2 FILLER_79_846 ();
 sg13g2_fill_1 FILLER_79_848 ();
 sg13g2_decap_4 FILLER_79_853 ();
 sg13g2_decap_4 FILLER_79_866 ();
 sg13g2_decap_8 FILLER_79_907 ();
 sg13g2_decap_4 FILLER_79_914 ();
 sg13g2_fill_2 FILLER_79_918 ();
 sg13g2_decap_8 FILLER_79_924 ();
 sg13g2_fill_2 FILLER_79_931 ();
 sg13g2_fill_1 FILLER_79_933 ();
 sg13g2_decap_8 FILLER_79_943 ();
 sg13g2_decap_8 FILLER_79_950 ();
 sg13g2_decap_8 FILLER_79_957 ();
 sg13g2_decap_8 FILLER_79_964 ();
 sg13g2_decap_8 FILLER_79_971 ();
 sg13g2_decap_8 FILLER_79_978 ();
 sg13g2_decap_8 FILLER_79_985 ();
 sg13g2_decap_8 FILLER_79_992 ();
 sg13g2_decap_8 FILLER_79_1003 ();
 sg13g2_decap_8 FILLER_79_1010 ();
 sg13g2_decap_8 FILLER_79_1017 ();
 sg13g2_decap_8 FILLER_79_1024 ();
 sg13g2_decap_8 FILLER_79_1031 ();
 sg13g2_decap_8 FILLER_79_1038 ();
 sg13g2_fill_2 FILLER_79_1045 ();
 sg13g2_decap_8 FILLER_79_1084 ();
 sg13g2_fill_2 FILLER_79_1091 ();
 sg13g2_decap_8 FILLER_79_1152 ();
 sg13g2_decap_8 FILLER_79_1159 ();
 sg13g2_decap_8 FILLER_79_1166 ();
 sg13g2_decap_8 FILLER_79_1173 ();
 sg13g2_decap_8 FILLER_79_1180 ();
 sg13g2_decap_8 FILLER_79_1187 ();
 sg13g2_decap_8 FILLER_79_1194 ();
 sg13g2_decap_8 FILLER_79_1201 ();
 sg13g2_decap_8 FILLER_79_1208 ();
 sg13g2_decap_8 FILLER_79_1215 ();
 sg13g2_decap_8 FILLER_79_1222 ();
 sg13g2_decap_8 FILLER_79_1229 ();
 sg13g2_decap_8 FILLER_79_1243 ();
 sg13g2_decap_8 FILLER_79_1250 ();
 sg13g2_decap_8 FILLER_79_1257 ();
 sg13g2_decap_8 FILLER_79_1264 ();
 sg13g2_decap_8 FILLER_79_1271 ();
 sg13g2_fill_2 FILLER_79_1278 ();
 sg13g2_fill_1 FILLER_79_1280 ();
 sg13g2_fill_2 FILLER_79_1321 ();
 sg13g2_fill_2 FILLER_79_1332 ();
 sg13g2_fill_1 FILLER_79_1334 ();
 sg13g2_decap_8 FILLER_79_1339 ();
 sg13g2_decap_8 FILLER_79_1346 ();
 sg13g2_decap_8 FILLER_79_1353 ();
 sg13g2_decap_8 FILLER_79_1360 ();
 sg13g2_decap_8 FILLER_79_1367 ();
 sg13g2_decap_8 FILLER_79_1374 ();
 sg13g2_decap_8 FILLER_79_1381 ();
 sg13g2_decap_8 FILLER_79_1388 ();
 sg13g2_decap_8 FILLER_79_1395 ();
 sg13g2_fill_2 FILLER_79_1402 ();
 sg13g2_fill_1 FILLER_79_1422 ();
 sg13g2_fill_2 FILLER_79_1427 ();
 sg13g2_decap_8 FILLER_79_1438 ();
 sg13g2_decap_8 FILLER_79_1445 ();
 sg13g2_decap_4 FILLER_79_1452 ();
 sg13g2_fill_1 FILLER_79_1456 ();
 sg13g2_decap_8 FILLER_79_1488 ();
 sg13g2_decap_8 FILLER_79_1495 ();
 sg13g2_decap_8 FILLER_79_1502 ();
 sg13g2_decap_8 FILLER_79_1509 ();
 sg13g2_decap_8 FILLER_79_1516 ();
 sg13g2_decap_8 FILLER_79_1523 ();
 sg13g2_decap_8 FILLER_79_1530 ();
 sg13g2_decap_8 FILLER_79_1537 ();
 sg13g2_decap_4 FILLER_79_1544 ();
 sg13g2_fill_1 FILLER_79_1548 ();
 sg13g2_fill_2 FILLER_79_1562 ();
 sg13g2_fill_1 FILLER_79_1585 ();
 sg13g2_fill_2 FILLER_79_1599 ();
 sg13g2_decap_8 FILLER_79_1609 ();
 sg13g2_fill_2 FILLER_79_1616 ();
 sg13g2_fill_1 FILLER_79_1618 ();
 sg13g2_fill_1 FILLER_79_1632 ();
 sg13g2_fill_1 FILLER_79_1642 ();
 sg13g2_decap_4 FILLER_79_1677 ();
 sg13g2_fill_2 FILLER_79_1685 ();
 sg13g2_decap_8 FILLER_79_1696 ();
 sg13g2_decap_8 FILLER_79_1703 ();
 sg13g2_decap_8 FILLER_79_1710 ();
 sg13g2_decap_8 FILLER_79_1717 ();
 sg13g2_decap_8 FILLER_79_1724 ();
 sg13g2_decap_8 FILLER_79_1731 ();
 sg13g2_decap_8 FILLER_79_1738 ();
 sg13g2_decap_8 FILLER_79_1745 ();
 sg13g2_decap_8 FILLER_79_1752 ();
 sg13g2_decap_8 FILLER_79_1759 ();
 sg13g2_decap_8 FILLER_79_1766 ();
 sg13g2_decap_8 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_79_1780 ();
 sg13g2_decap_8 FILLER_79_1787 ();
 sg13g2_decap_8 FILLER_79_1794 ();
 sg13g2_decap_8 FILLER_79_1801 ();
 sg13g2_decap_8 FILLER_79_1808 ();
 sg13g2_decap_8 FILLER_79_1815 ();
 sg13g2_decap_8 FILLER_79_1822 ();
 sg13g2_decap_8 FILLER_79_1829 ();
 sg13g2_decap_8 FILLER_79_1836 ();
 sg13g2_decap_8 FILLER_79_1843 ();
 sg13g2_decap_8 FILLER_79_1850 ();
 sg13g2_decap_8 FILLER_79_1857 ();
 sg13g2_decap_8 FILLER_79_1864 ();
 sg13g2_decap_8 FILLER_79_1871 ();
 sg13g2_decap_8 FILLER_79_1878 ();
 sg13g2_decap_8 FILLER_79_1885 ();
 sg13g2_decap_8 FILLER_79_1892 ();
 sg13g2_fill_2 FILLER_79_1899 ();
 sg13g2_decap_8 FILLER_79_1905 ();
 sg13g2_decap_8 FILLER_79_1912 ();
 sg13g2_fill_1 FILLER_79_1919 ();
 sg13g2_decap_8 FILLER_79_1948 ();
 sg13g2_decap_4 FILLER_79_1955 ();
 sg13g2_fill_2 FILLER_79_2013 ();
 sg13g2_fill_2 FILLER_79_2071 ();
 sg13g2_fill_1 FILLER_79_2073 ();
 sg13g2_decap_4 FILLER_79_2096 ();
 sg13g2_decap_4 FILLER_79_2155 ();
 sg13g2_fill_2 FILLER_79_2159 ();
 sg13g2_decap_8 FILLER_79_2165 ();
 sg13g2_decap_4 FILLER_79_2172 ();
 sg13g2_fill_2 FILLER_79_2181 ();
 sg13g2_fill_1 FILLER_79_2183 ();
 sg13g2_decap_8 FILLER_79_2211 ();
 sg13g2_decap_8 FILLER_79_2218 ();
 sg13g2_decap_8 FILLER_79_2225 ();
 sg13g2_decap_8 FILLER_79_2232 ();
 sg13g2_decap_8 FILLER_79_2239 ();
 sg13g2_decap_8 FILLER_79_2246 ();
 sg13g2_decap_8 FILLER_79_2253 ();
 sg13g2_decap_8 FILLER_79_2260 ();
 sg13g2_decap_8 FILLER_79_2267 ();
 sg13g2_decap_8 FILLER_79_2274 ();
 sg13g2_decap_8 FILLER_79_2281 ();
 sg13g2_decap_8 FILLER_79_2288 ();
 sg13g2_decap_8 FILLER_79_2295 ();
 sg13g2_decap_8 FILLER_79_2302 ();
 sg13g2_decap_8 FILLER_79_2309 ();
 sg13g2_decap_8 FILLER_79_2316 ();
 sg13g2_decap_8 FILLER_79_2323 ();
 sg13g2_decap_8 FILLER_79_2330 ();
 sg13g2_decap_8 FILLER_79_2337 ();
 sg13g2_decap_8 FILLER_79_2344 ();
 sg13g2_decap_8 FILLER_79_2351 ();
 sg13g2_decap_8 FILLER_79_2358 ();
 sg13g2_decap_8 FILLER_79_2365 ();
 sg13g2_decap_8 FILLER_79_2372 ();
 sg13g2_decap_8 FILLER_79_2379 ();
 sg13g2_decap_8 FILLER_79_2386 ();
 sg13g2_decap_8 FILLER_79_2393 ();
 sg13g2_decap_8 FILLER_79_2400 ();
 sg13g2_decap_8 FILLER_79_2407 ();
 sg13g2_decap_8 FILLER_79_2414 ();
 sg13g2_decap_8 FILLER_79_2421 ();
 sg13g2_decap_8 FILLER_79_2428 ();
 sg13g2_decap_8 FILLER_79_2435 ();
 sg13g2_decap_8 FILLER_79_2442 ();
 sg13g2_decap_8 FILLER_79_2449 ();
 sg13g2_decap_8 FILLER_79_2456 ();
 sg13g2_decap_8 FILLER_79_2463 ();
 sg13g2_decap_8 FILLER_79_2470 ();
 sg13g2_decap_8 FILLER_79_2477 ();
 sg13g2_decap_8 FILLER_79_2484 ();
 sg13g2_decap_8 FILLER_79_2491 ();
 sg13g2_decap_8 FILLER_79_2498 ();
 sg13g2_decap_8 FILLER_79_2505 ();
 sg13g2_decap_8 FILLER_79_2512 ();
 sg13g2_decap_8 FILLER_79_2519 ();
 sg13g2_decap_8 FILLER_79_2526 ();
 sg13g2_decap_8 FILLER_79_2533 ();
 sg13g2_decap_8 FILLER_79_2540 ();
 sg13g2_decap_8 FILLER_79_2547 ();
 sg13g2_decap_8 FILLER_79_2554 ();
 sg13g2_decap_8 FILLER_79_2561 ();
 sg13g2_decap_8 FILLER_79_2568 ();
 sg13g2_decap_8 FILLER_79_2575 ();
 sg13g2_decap_8 FILLER_79_2582 ();
 sg13g2_decap_8 FILLER_79_2589 ();
 sg13g2_decap_8 FILLER_79_2596 ();
 sg13g2_decap_8 FILLER_79_2603 ();
 sg13g2_decap_8 FILLER_79_2610 ();
 sg13g2_decap_8 FILLER_79_2617 ();
 sg13g2_decap_8 FILLER_79_2624 ();
 sg13g2_decap_8 FILLER_79_2631 ();
 sg13g2_decap_8 FILLER_79_2638 ();
 sg13g2_decap_8 FILLER_79_2645 ();
 sg13g2_decap_8 FILLER_79_2652 ();
 sg13g2_decap_8 FILLER_79_2659 ();
 sg13g2_decap_8 FILLER_79_2666 ();
 sg13g2_decap_8 FILLER_79_2673 ();
 sg13g2_decap_8 FILLER_79_2680 ();
 sg13g2_decap_8 FILLER_79_2687 ();
 sg13g2_decap_8 FILLER_79_2694 ();
 sg13g2_decap_8 FILLER_79_2701 ();
 sg13g2_decap_8 FILLER_79_2708 ();
 sg13g2_decap_8 FILLER_79_2715 ();
 sg13g2_decap_8 FILLER_79_2722 ();
 sg13g2_decap_8 FILLER_79_2729 ();
 sg13g2_decap_8 FILLER_79_2736 ();
 sg13g2_decap_8 FILLER_79_2743 ();
 sg13g2_decap_8 FILLER_79_2750 ();
 sg13g2_decap_8 FILLER_79_2757 ();
 sg13g2_decap_8 FILLER_79_2764 ();
 sg13g2_decap_8 FILLER_79_2771 ();
 sg13g2_decap_8 FILLER_79_2778 ();
 sg13g2_decap_8 FILLER_79_2785 ();
 sg13g2_decap_8 FILLER_79_2792 ();
 sg13g2_decap_8 FILLER_79_2799 ();
 sg13g2_decap_8 FILLER_79_2806 ();
 sg13g2_decap_8 FILLER_79_2813 ();
 sg13g2_decap_8 FILLER_79_2820 ();
 sg13g2_decap_8 FILLER_79_2827 ();
 sg13g2_decap_8 FILLER_79_2834 ();
 sg13g2_decap_8 FILLER_79_2841 ();
 sg13g2_decap_8 FILLER_79_2848 ();
 sg13g2_decap_8 FILLER_79_2855 ();
 sg13g2_decap_8 FILLER_79_2862 ();
 sg13g2_decap_8 FILLER_79_2869 ();
 sg13g2_decap_8 FILLER_79_2876 ();
 sg13g2_decap_8 FILLER_79_2883 ();
 sg13g2_decap_8 FILLER_79_2890 ();
 sg13g2_decap_8 FILLER_79_2897 ();
 sg13g2_decap_8 FILLER_79_2904 ();
 sg13g2_decap_8 FILLER_79_2911 ();
 sg13g2_decap_8 FILLER_79_2918 ();
 sg13g2_decap_8 FILLER_79_2925 ();
 sg13g2_decap_8 FILLER_79_2932 ();
 sg13g2_decap_8 FILLER_79_2939 ();
 sg13g2_decap_8 FILLER_79_2946 ();
 sg13g2_decap_8 FILLER_79_2953 ();
 sg13g2_decap_8 FILLER_79_2960 ();
 sg13g2_decap_8 FILLER_79_2967 ();
 sg13g2_decap_8 FILLER_79_2974 ();
 sg13g2_decap_8 FILLER_79_2981 ();
 sg13g2_decap_8 FILLER_79_2988 ();
 sg13g2_decap_8 FILLER_79_2995 ();
 sg13g2_decap_8 FILLER_79_3002 ();
 sg13g2_decap_8 FILLER_79_3009 ();
 sg13g2_decap_8 FILLER_79_3016 ();
 sg13g2_decap_8 FILLER_79_3023 ();
 sg13g2_decap_8 FILLER_79_3030 ();
 sg13g2_decap_8 FILLER_79_3037 ();
 sg13g2_decap_8 FILLER_79_3044 ();
 sg13g2_decap_8 FILLER_79_3051 ();
 sg13g2_decap_8 FILLER_79_3058 ();
 sg13g2_decap_8 FILLER_79_3065 ();
 sg13g2_decap_8 FILLER_79_3072 ();
 sg13g2_decap_8 FILLER_79_3079 ();
 sg13g2_decap_8 FILLER_79_3086 ();
 sg13g2_decap_8 FILLER_79_3093 ();
 sg13g2_decap_8 FILLER_79_3100 ();
 sg13g2_decap_8 FILLER_79_3107 ();
 sg13g2_decap_8 FILLER_79_3114 ();
 sg13g2_decap_8 FILLER_79_3121 ();
 sg13g2_decap_8 FILLER_79_3128 ();
 sg13g2_decap_8 FILLER_79_3135 ();
 sg13g2_decap_8 FILLER_79_3142 ();
 sg13g2_decap_8 FILLER_79_3149 ();
 sg13g2_decap_8 FILLER_79_3156 ();
 sg13g2_decap_8 FILLER_79_3163 ();
 sg13g2_decap_8 FILLER_79_3170 ();
 sg13g2_decap_8 FILLER_79_3177 ();
 sg13g2_decap_8 FILLER_79_3184 ();
 sg13g2_decap_8 FILLER_79_3191 ();
 sg13g2_decap_8 FILLER_79_3198 ();
 sg13g2_decap_8 FILLER_79_3205 ();
 sg13g2_decap_8 FILLER_79_3212 ();
 sg13g2_decap_8 FILLER_79_3219 ();
 sg13g2_decap_8 FILLER_79_3226 ();
 sg13g2_decap_8 FILLER_79_3233 ();
 sg13g2_decap_8 FILLER_79_3240 ();
 sg13g2_decap_8 FILLER_79_3247 ();
 sg13g2_decap_8 FILLER_79_3254 ();
 sg13g2_decap_8 FILLER_79_3261 ();
 sg13g2_decap_8 FILLER_79_3268 ();
 sg13g2_decap_8 FILLER_79_3275 ();
 sg13g2_decap_8 FILLER_79_3282 ();
 sg13g2_decap_8 FILLER_79_3289 ();
 sg13g2_decap_8 FILLER_79_3296 ();
 sg13g2_decap_8 FILLER_79_3303 ();
 sg13g2_decap_8 FILLER_79_3310 ();
 sg13g2_decap_8 FILLER_79_3317 ();
 sg13g2_decap_8 FILLER_79_3324 ();
 sg13g2_decap_8 FILLER_79_3331 ();
 sg13g2_decap_8 FILLER_79_3338 ();
 sg13g2_decap_8 FILLER_79_3345 ();
 sg13g2_decap_8 FILLER_79_3352 ();
 sg13g2_decap_8 FILLER_79_3359 ();
 sg13g2_decap_8 FILLER_79_3366 ();
 sg13g2_decap_8 FILLER_79_3373 ();
 sg13g2_decap_8 FILLER_79_3380 ();
 sg13g2_decap_8 FILLER_79_3387 ();
 sg13g2_decap_8 FILLER_79_3394 ();
 sg13g2_decap_8 FILLER_79_3401 ();
 sg13g2_decap_8 FILLER_79_3408 ();
 sg13g2_decap_8 FILLER_79_3415 ();
 sg13g2_decap_8 FILLER_79_3422 ();
 sg13g2_decap_8 FILLER_79_3429 ();
 sg13g2_decap_8 FILLER_79_3436 ();
 sg13g2_decap_8 FILLER_79_3443 ();
 sg13g2_decap_8 FILLER_79_3450 ();
 sg13g2_decap_8 FILLER_79_3457 ();
 sg13g2_decap_8 FILLER_79_3464 ();
 sg13g2_decap_8 FILLER_79_3471 ();
 sg13g2_decap_8 FILLER_79_3478 ();
 sg13g2_decap_8 FILLER_79_3485 ();
 sg13g2_decap_8 FILLER_79_3492 ();
 sg13g2_decap_8 FILLER_79_3499 ();
 sg13g2_decap_8 FILLER_79_3506 ();
 sg13g2_decap_8 FILLER_79_3513 ();
 sg13g2_decap_8 FILLER_79_3520 ();
 sg13g2_decap_8 FILLER_79_3527 ();
 sg13g2_decap_8 FILLER_79_3534 ();
 sg13g2_decap_8 FILLER_79_3541 ();
 sg13g2_decap_8 FILLER_79_3548 ();
 sg13g2_decap_8 FILLER_79_3555 ();
 sg13g2_decap_8 FILLER_79_3562 ();
 sg13g2_decap_8 FILLER_79_3569 ();
 sg13g2_decap_4 FILLER_79_3576 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_171 ();
 sg13g2_decap_8 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_185 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_213 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_4 FILLER_80_276 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_4 FILLER_80_306 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_decap_4 FILLER_80_316 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_decap_8 FILLER_80_428 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_decap_8 FILLER_80_456 ();
 sg13g2_decap_8 FILLER_80_463 ();
 sg13g2_decap_8 FILLER_80_470 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_4 FILLER_80_554 ();
 sg13g2_fill_2 FILLER_80_558 ();
 sg13g2_decap_4 FILLER_80_564 ();
 sg13g2_fill_2 FILLER_80_568 ();
 sg13g2_fill_1 FILLER_80_586 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_4 FILLER_80_652 ();
 sg13g2_fill_1 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_4 FILLER_80_675 ();
 sg13g2_decap_4 FILLER_80_739 ();
 sg13g2_fill_2 FILLER_80_743 ();
 sg13g2_fill_2 FILLER_80_749 ();
 sg13g2_fill_1 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_fill_1 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_4 FILLER_80_801 ();
 sg13g2_fill_2 FILLER_80_805 ();
 sg13g2_fill_2 FILLER_80_841 ();
 sg13g2_fill_1 FILLER_80_843 ();
 sg13g2_fill_2 FILLER_80_872 ();
 sg13g2_fill_1 FILLER_80_874 ();
 sg13g2_decap_8 FILLER_80_879 ();
 sg13g2_decap_4 FILLER_80_886 ();
 sg13g2_fill_1 FILLER_80_890 ();
 sg13g2_decap_8 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_933 ();
 sg13g2_decap_8 FILLER_80_940 ();
 sg13g2_decap_8 FILLER_80_947 ();
 sg13g2_decap_8 FILLER_80_954 ();
 sg13g2_decap_8 FILLER_80_961 ();
 sg13g2_decap_8 FILLER_80_968 ();
 sg13g2_decap_8 FILLER_80_975 ();
 sg13g2_decap_8 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_decap_8 FILLER_80_1003 ();
 sg13g2_decap_8 FILLER_80_1010 ();
 sg13g2_decap_8 FILLER_80_1017 ();
 sg13g2_decap_8 FILLER_80_1024 ();
 sg13g2_decap_8 FILLER_80_1031 ();
 sg13g2_decap_8 FILLER_80_1038 ();
 sg13g2_decap_8 FILLER_80_1045 ();
 sg13g2_decap_8 FILLER_80_1056 ();
 sg13g2_decap_4 FILLER_80_1063 ();
 sg13g2_fill_1 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1071 ();
 sg13g2_decap_8 FILLER_80_1078 ();
 sg13g2_decap_8 FILLER_80_1085 ();
 sg13g2_decap_8 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1106 ();
 sg13g2_decap_4 FILLER_80_1113 ();
 sg13g2_fill_1 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_fill_2 FILLER_80_1292 ();
 sg13g2_fill_1 FILLER_80_1294 ();
 sg13g2_decap_8 FILLER_80_1336 ();
 sg13g2_decap_8 FILLER_80_1343 ();
 sg13g2_decap_8 FILLER_80_1350 ();
 sg13g2_decap_8 FILLER_80_1357 ();
 sg13g2_decap_8 FILLER_80_1364 ();
 sg13g2_decap_8 FILLER_80_1371 ();
 sg13g2_decap_8 FILLER_80_1378 ();
 sg13g2_decap_8 FILLER_80_1385 ();
 sg13g2_decap_8 FILLER_80_1392 ();
 sg13g2_decap_8 FILLER_80_1399 ();
 sg13g2_fill_1 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1439 ();
 sg13g2_decap_8 FILLER_80_1446 ();
 sg13g2_decap_8 FILLER_80_1453 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_4 FILLER_80_1467 ();
 sg13g2_fill_2 FILLER_80_1471 ();
 sg13g2_decap_8 FILLER_80_1482 ();
 sg13g2_decap_8 FILLER_80_1489 ();
 sg13g2_decap_8 FILLER_80_1496 ();
 sg13g2_decap_8 FILLER_80_1503 ();
 sg13g2_decap_8 FILLER_80_1510 ();
 sg13g2_decap_8 FILLER_80_1517 ();
 sg13g2_decap_8 FILLER_80_1524 ();
 sg13g2_decap_8 FILLER_80_1531 ();
 sg13g2_decap_8 FILLER_80_1538 ();
 sg13g2_decap_8 FILLER_80_1545 ();
 sg13g2_decap_8 FILLER_80_1552 ();
 sg13g2_decap_8 FILLER_80_1559 ();
 sg13g2_fill_2 FILLER_80_1566 ();
 sg13g2_fill_1 FILLER_80_1568 ();
 sg13g2_decap_8 FILLER_80_1603 ();
 sg13g2_decap_4 FILLER_80_1610 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1691 ();
 sg13g2_decap_8 FILLER_80_1698 ();
 sg13g2_decap_8 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1712 ();
 sg13g2_decap_8 FILLER_80_1719 ();
 sg13g2_decap_8 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_80_1768 ();
 sg13g2_decap_8 FILLER_80_1775 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_8 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1803 ();
 sg13g2_decap_8 FILLER_80_1810 ();
 sg13g2_decap_8 FILLER_80_1817 ();
 sg13g2_decap_8 FILLER_80_1824 ();
 sg13g2_decap_8 FILLER_80_1831 ();
 sg13g2_decap_8 FILLER_80_1838 ();
 sg13g2_decap_8 FILLER_80_1845 ();
 sg13g2_decap_8 FILLER_80_1852 ();
 sg13g2_decap_8 FILLER_80_1859 ();
 sg13g2_decap_8 FILLER_80_1866 ();
 sg13g2_decap_8 FILLER_80_1873 ();
 sg13g2_decap_8 FILLER_80_1880 ();
 sg13g2_decap_8 FILLER_80_1887 ();
 sg13g2_decap_8 FILLER_80_1894 ();
 sg13g2_decap_8 FILLER_80_1901 ();
 sg13g2_decap_8 FILLER_80_1908 ();
 sg13g2_decap_8 FILLER_80_1915 ();
 sg13g2_fill_2 FILLER_80_1922 ();
 sg13g2_fill_1 FILLER_80_1924 ();
 sg13g2_decap_8 FILLER_80_1929 ();
 sg13g2_decap_4 FILLER_80_1936 ();
 sg13g2_fill_2 FILLER_80_1940 ();
 sg13g2_decap_8 FILLER_80_1946 ();
 sg13g2_decap_4 FILLER_80_1953 ();
 sg13g2_fill_1 FILLER_80_1957 ();
 sg13g2_decap_8 FILLER_80_1971 ();
 sg13g2_fill_2 FILLER_80_1978 ();
 sg13g2_decap_8 FILLER_80_2012 ();
 sg13g2_fill_1 FILLER_80_2019 ();
 sg13g2_decap_8 FILLER_80_2024 ();
 sg13g2_decap_8 FILLER_80_2031 ();
 sg13g2_decap_8 FILLER_80_2038 ();
 sg13g2_decap_8 FILLER_80_2049 ();
 sg13g2_fill_1 FILLER_80_2056 ();
 sg13g2_decap_8 FILLER_80_2089 ();
 sg13g2_decap_8 FILLER_80_2096 ();
 sg13g2_decap_8 FILLER_80_2103 ();
 sg13g2_decap_8 FILLER_80_2110 ();
 sg13g2_decap_8 FILLER_80_2117 ();
 sg13g2_fill_2 FILLER_80_2124 ();
 sg13g2_fill_1 FILLER_80_2126 ();
 sg13g2_decap_8 FILLER_80_2140 ();
 sg13g2_decap_8 FILLER_80_2147 ();
 sg13g2_fill_2 FILLER_80_2154 ();
 sg13g2_decap_8 FILLER_80_2197 ();
 sg13g2_decap_8 FILLER_80_2204 ();
 sg13g2_decap_8 FILLER_80_2211 ();
 sg13g2_decap_8 FILLER_80_2218 ();
 sg13g2_decap_8 FILLER_80_2225 ();
 sg13g2_decap_8 FILLER_80_2232 ();
 sg13g2_decap_8 FILLER_80_2239 ();
 sg13g2_decap_8 FILLER_80_2246 ();
 sg13g2_decap_8 FILLER_80_2253 ();
 sg13g2_decap_8 FILLER_80_2260 ();
 sg13g2_decap_8 FILLER_80_2267 ();
 sg13g2_decap_8 FILLER_80_2274 ();
 sg13g2_decap_8 FILLER_80_2281 ();
 sg13g2_decap_8 FILLER_80_2288 ();
 sg13g2_decap_8 FILLER_80_2295 ();
 sg13g2_decap_8 FILLER_80_2302 ();
 sg13g2_decap_8 FILLER_80_2309 ();
 sg13g2_decap_8 FILLER_80_2316 ();
 sg13g2_decap_8 FILLER_80_2323 ();
 sg13g2_decap_8 FILLER_80_2330 ();
 sg13g2_decap_8 FILLER_80_2337 ();
 sg13g2_decap_8 FILLER_80_2344 ();
 sg13g2_decap_8 FILLER_80_2351 ();
 sg13g2_decap_8 FILLER_80_2358 ();
 sg13g2_decap_8 FILLER_80_2365 ();
 sg13g2_decap_8 FILLER_80_2372 ();
 sg13g2_decap_8 FILLER_80_2379 ();
 sg13g2_decap_8 FILLER_80_2386 ();
 sg13g2_decap_8 FILLER_80_2393 ();
 sg13g2_decap_8 FILLER_80_2400 ();
 sg13g2_decap_8 FILLER_80_2407 ();
 sg13g2_decap_8 FILLER_80_2414 ();
 sg13g2_decap_8 FILLER_80_2421 ();
 sg13g2_decap_8 FILLER_80_2428 ();
 sg13g2_decap_8 FILLER_80_2435 ();
 sg13g2_decap_8 FILLER_80_2442 ();
 sg13g2_decap_8 FILLER_80_2449 ();
 sg13g2_decap_8 FILLER_80_2456 ();
 sg13g2_decap_8 FILLER_80_2463 ();
 sg13g2_decap_8 FILLER_80_2470 ();
 sg13g2_decap_8 FILLER_80_2477 ();
 sg13g2_decap_8 FILLER_80_2484 ();
 sg13g2_decap_8 FILLER_80_2491 ();
 sg13g2_decap_8 FILLER_80_2498 ();
 sg13g2_decap_8 FILLER_80_2505 ();
 sg13g2_decap_8 FILLER_80_2512 ();
 sg13g2_decap_8 FILLER_80_2519 ();
 sg13g2_decap_8 FILLER_80_2526 ();
 sg13g2_decap_8 FILLER_80_2533 ();
 sg13g2_decap_8 FILLER_80_2540 ();
 sg13g2_decap_8 FILLER_80_2547 ();
 sg13g2_decap_8 FILLER_80_2554 ();
 sg13g2_decap_8 FILLER_80_2561 ();
 sg13g2_decap_8 FILLER_80_2568 ();
 sg13g2_decap_8 FILLER_80_2575 ();
 sg13g2_decap_8 FILLER_80_2582 ();
 sg13g2_decap_8 FILLER_80_2589 ();
 sg13g2_decap_8 FILLER_80_2596 ();
 sg13g2_decap_8 FILLER_80_2603 ();
 sg13g2_decap_8 FILLER_80_2610 ();
 sg13g2_decap_8 FILLER_80_2617 ();
 sg13g2_decap_8 FILLER_80_2624 ();
 sg13g2_decap_8 FILLER_80_2631 ();
 sg13g2_decap_8 FILLER_80_2638 ();
 sg13g2_decap_8 FILLER_80_2645 ();
 sg13g2_decap_8 FILLER_80_2652 ();
 sg13g2_decap_8 FILLER_80_2659 ();
 sg13g2_decap_8 FILLER_80_2666 ();
 sg13g2_decap_8 FILLER_80_2673 ();
 sg13g2_decap_8 FILLER_80_2680 ();
 sg13g2_decap_8 FILLER_80_2687 ();
 sg13g2_decap_8 FILLER_80_2694 ();
 sg13g2_decap_8 FILLER_80_2701 ();
 sg13g2_decap_8 FILLER_80_2708 ();
 sg13g2_decap_8 FILLER_80_2715 ();
 sg13g2_decap_8 FILLER_80_2722 ();
 sg13g2_decap_8 FILLER_80_2729 ();
 sg13g2_decap_8 FILLER_80_2736 ();
 sg13g2_decap_8 FILLER_80_2743 ();
 sg13g2_decap_8 FILLER_80_2750 ();
 sg13g2_decap_8 FILLER_80_2757 ();
 sg13g2_decap_8 FILLER_80_2764 ();
 sg13g2_decap_8 FILLER_80_2771 ();
 sg13g2_decap_8 FILLER_80_2778 ();
 sg13g2_decap_8 FILLER_80_2785 ();
 sg13g2_decap_8 FILLER_80_2792 ();
 sg13g2_decap_8 FILLER_80_2799 ();
 sg13g2_decap_8 FILLER_80_2806 ();
 sg13g2_decap_8 FILLER_80_2813 ();
 sg13g2_decap_8 FILLER_80_2820 ();
 sg13g2_decap_8 FILLER_80_2827 ();
 sg13g2_decap_8 FILLER_80_2834 ();
 sg13g2_decap_8 FILLER_80_2841 ();
 sg13g2_decap_8 FILLER_80_2848 ();
 sg13g2_decap_8 FILLER_80_2855 ();
 sg13g2_decap_8 FILLER_80_2862 ();
 sg13g2_decap_8 FILLER_80_2869 ();
 sg13g2_decap_8 FILLER_80_2876 ();
 sg13g2_decap_8 FILLER_80_2883 ();
 sg13g2_decap_8 FILLER_80_2890 ();
 sg13g2_decap_8 FILLER_80_2897 ();
 sg13g2_decap_8 FILLER_80_2904 ();
 sg13g2_decap_8 FILLER_80_2911 ();
 sg13g2_decap_8 FILLER_80_2918 ();
 sg13g2_decap_8 FILLER_80_2925 ();
 sg13g2_decap_8 FILLER_80_2932 ();
 sg13g2_decap_8 FILLER_80_2939 ();
 sg13g2_decap_8 FILLER_80_2946 ();
 sg13g2_decap_8 FILLER_80_2953 ();
 sg13g2_decap_8 FILLER_80_2960 ();
 sg13g2_decap_8 FILLER_80_2967 ();
 sg13g2_decap_8 FILLER_80_2974 ();
 sg13g2_decap_8 FILLER_80_2981 ();
 sg13g2_decap_8 FILLER_80_2988 ();
 sg13g2_decap_8 FILLER_80_2995 ();
 sg13g2_decap_8 FILLER_80_3002 ();
 sg13g2_decap_8 FILLER_80_3009 ();
 sg13g2_decap_8 FILLER_80_3016 ();
 sg13g2_decap_8 FILLER_80_3023 ();
 sg13g2_decap_8 FILLER_80_3030 ();
 sg13g2_decap_8 FILLER_80_3037 ();
 sg13g2_decap_8 FILLER_80_3044 ();
 sg13g2_decap_8 FILLER_80_3051 ();
 sg13g2_decap_8 FILLER_80_3058 ();
 sg13g2_decap_8 FILLER_80_3065 ();
 sg13g2_decap_8 FILLER_80_3072 ();
 sg13g2_decap_8 FILLER_80_3079 ();
 sg13g2_decap_8 FILLER_80_3086 ();
 sg13g2_decap_8 FILLER_80_3093 ();
 sg13g2_decap_8 FILLER_80_3100 ();
 sg13g2_decap_8 FILLER_80_3107 ();
 sg13g2_decap_8 FILLER_80_3114 ();
 sg13g2_decap_8 FILLER_80_3121 ();
 sg13g2_decap_8 FILLER_80_3128 ();
 sg13g2_decap_8 FILLER_80_3135 ();
 sg13g2_decap_8 FILLER_80_3142 ();
 sg13g2_decap_8 FILLER_80_3149 ();
 sg13g2_decap_8 FILLER_80_3156 ();
 sg13g2_decap_8 FILLER_80_3163 ();
 sg13g2_decap_8 FILLER_80_3170 ();
 sg13g2_decap_8 FILLER_80_3177 ();
 sg13g2_decap_8 FILLER_80_3184 ();
 sg13g2_decap_8 FILLER_80_3191 ();
 sg13g2_decap_8 FILLER_80_3198 ();
 sg13g2_decap_8 FILLER_80_3205 ();
 sg13g2_decap_8 FILLER_80_3212 ();
 sg13g2_decap_8 FILLER_80_3219 ();
 sg13g2_decap_8 FILLER_80_3226 ();
 sg13g2_decap_8 FILLER_80_3233 ();
 sg13g2_decap_8 FILLER_80_3240 ();
 sg13g2_decap_8 FILLER_80_3247 ();
 sg13g2_decap_8 FILLER_80_3254 ();
 sg13g2_decap_8 FILLER_80_3261 ();
 sg13g2_decap_8 FILLER_80_3268 ();
 sg13g2_decap_8 FILLER_80_3275 ();
 sg13g2_decap_8 FILLER_80_3282 ();
 sg13g2_decap_8 FILLER_80_3289 ();
 sg13g2_decap_8 FILLER_80_3296 ();
 sg13g2_decap_8 FILLER_80_3303 ();
 sg13g2_decap_8 FILLER_80_3310 ();
 sg13g2_decap_8 FILLER_80_3317 ();
 sg13g2_decap_8 FILLER_80_3324 ();
 sg13g2_decap_8 FILLER_80_3331 ();
 sg13g2_decap_8 FILLER_80_3338 ();
 sg13g2_decap_8 FILLER_80_3345 ();
 sg13g2_decap_8 FILLER_80_3352 ();
 sg13g2_decap_8 FILLER_80_3359 ();
 sg13g2_decap_8 FILLER_80_3366 ();
 sg13g2_decap_8 FILLER_80_3373 ();
 sg13g2_decap_8 FILLER_80_3380 ();
 sg13g2_decap_8 FILLER_80_3387 ();
 sg13g2_decap_8 FILLER_80_3394 ();
 sg13g2_decap_8 FILLER_80_3401 ();
 sg13g2_decap_8 FILLER_80_3408 ();
 sg13g2_decap_8 FILLER_80_3415 ();
 sg13g2_decap_8 FILLER_80_3422 ();
 sg13g2_decap_8 FILLER_80_3429 ();
 sg13g2_decap_8 FILLER_80_3436 ();
 sg13g2_decap_8 FILLER_80_3443 ();
 sg13g2_decap_8 FILLER_80_3450 ();
 sg13g2_decap_8 FILLER_80_3457 ();
 sg13g2_decap_8 FILLER_80_3464 ();
 sg13g2_decap_8 FILLER_80_3471 ();
 sg13g2_decap_8 FILLER_80_3478 ();
 sg13g2_decap_8 FILLER_80_3485 ();
 sg13g2_decap_8 FILLER_80_3492 ();
 sg13g2_decap_8 FILLER_80_3499 ();
 sg13g2_decap_8 FILLER_80_3506 ();
 sg13g2_decap_8 FILLER_80_3513 ();
 sg13g2_decap_8 FILLER_80_3520 ();
 sg13g2_decap_8 FILLER_80_3527 ();
 sg13g2_decap_8 FILLER_80_3534 ();
 sg13g2_decap_8 FILLER_80_3541 ();
 sg13g2_decap_8 FILLER_80_3548 ();
 sg13g2_decap_8 FILLER_80_3555 ();
 sg13g2_decap_8 FILLER_80_3562 ();
 sg13g2_decap_8 FILLER_80_3569 ();
 sg13g2_decap_4 FILLER_80_3576 ();
 assign uio_oe[0] = net1061;
 assign uio_oe[1] = net1062;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
