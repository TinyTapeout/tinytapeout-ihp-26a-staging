module tt_um_SotaSoC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire \soc_inst.bus_spi_sclk ;
 wire \soc_inst.core_instr_addr[0] ;
 wire \soc_inst.core_instr_addr[10] ;
 wire \soc_inst.core_instr_addr[11] ;
 wire \soc_inst.core_instr_addr[12] ;
 wire \soc_inst.core_instr_addr[13] ;
 wire \soc_inst.core_instr_addr[14] ;
 wire \soc_inst.core_instr_addr[15] ;
 wire \soc_inst.core_instr_addr[16] ;
 wire \soc_inst.core_instr_addr[17] ;
 wire \soc_inst.core_instr_addr[18] ;
 wire \soc_inst.core_instr_addr[19] ;
 wire \soc_inst.core_instr_addr[1] ;
 wire \soc_inst.core_instr_addr[20] ;
 wire \soc_inst.core_instr_addr[21] ;
 wire \soc_inst.core_instr_addr[22] ;
 wire \soc_inst.core_instr_addr[23] ;
 wire \soc_inst.core_instr_addr[2] ;
 wire \soc_inst.core_instr_addr[3] ;
 wire \soc_inst.core_instr_addr[4] ;
 wire \soc_inst.core_instr_addr[5] ;
 wire \soc_inst.core_instr_addr[6] ;
 wire \soc_inst.core_instr_addr[7] ;
 wire \soc_inst.core_instr_addr[8] ;
 wire \soc_inst.core_instr_addr[9] ;
 wire \soc_inst.core_instr_data[0] ;
 wire \soc_inst.core_instr_data[10] ;
 wire \soc_inst.core_instr_data[11] ;
 wire \soc_inst.core_instr_data[12] ;
 wire \soc_inst.core_instr_data[13] ;
 wire \soc_inst.core_instr_data[14] ;
 wire \soc_inst.core_instr_data[15] ;
 wire \soc_inst.core_instr_data[16] ;
 wire \soc_inst.core_instr_data[17] ;
 wire \soc_inst.core_instr_data[18] ;
 wire \soc_inst.core_instr_data[19] ;
 wire \soc_inst.core_instr_data[1] ;
 wire \soc_inst.core_instr_data[20] ;
 wire \soc_inst.core_instr_data[21] ;
 wire \soc_inst.core_instr_data[22] ;
 wire \soc_inst.core_instr_data[23] ;
 wire \soc_inst.core_instr_data[24] ;
 wire \soc_inst.core_instr_data[25] ;
 wire \soc_inst.core_instr_data[26] ;
 wire \soc_inst.core_instr_data[27] ;
 wire \soc_inst.core_instr_data[28] ;
 wire \soc_inst.core_instr_data[29] ;
 wire \soc_inst.core_instr_data[2] ;
 wire \soc_inst.core_instr_data[30] ;
 wire \soc_inst.core_instr_data[31] ;
 wire \soc_inst.core_instr_data[3] ;
 wire \soc_inst.core_instr_data[4] ;
 wire \soc_inst.core_instr_data[5] ;
 wire \soc_inst.core_instr_data[6] ;
 wire \soc_inst.core_instr_data[7] ;
 wire \soc_inst.core_instr_data[8] ;
 wire \soc_inst.core_instr_data[9] ;
 wire \soc_inst.core_mem_addr[0] ;
 wire \soc_inst.core_mem_addr[10] ;
 wire \soc_inst.core_mem_addr[11] ;
 wire \soc_inst.core_mem_addr[12] ;
 wire \soc_inst.core_mem_addr[13] ;
 wire \soc_inst.core_mem_addr[14] ;
 wire \soc_inst.core_mem_addr[15] ;
 wire \soc_inst.core_mem_addr[16] ;
 wire \soc_inst.core_mem_addr[17] ;
 wire \soc_inst.core_mem_addr[18] ;
 wire \soc_inst.core_mem_addr[19] ;
 wire \soc_inst.core_mem_addr[1] ;
 wire \soc_inst.core_mem_addr[20] ;
 wire \soc_inst.core_mem_addr[21] ;
 wire \soc_inst.core_mem_addr[22] ;
 wire \soc_inst.core_mem_addr[23] ;
 wire \soc_inst.core_mem_addr[24] ;
 wire \soc_inst.core_mem_addr[25] ;
 wire \soc_inst.core_mem_addr[26] ;
 wire \soc_inst.core_mem_addr[27] ;
 wire \soc_inst.core_mem_addr[28] ;
 wire \soc_inst.core_mem_addr[29] ;
 wire \soc_inst.core_mem_addr[2] ;
 wire \soc_inst.core_mem_addr[30] ;
 wire \soc_inst.core_mem_addr[31] ;
 wire \soc_inst.core_mem_addr[3] ;
 wire \soc_inst.core_mem_addr[5] ;
 wire \soc_inst.core_mem_addr[6] ;
 wire \soc_inst.core_mem_addr[7] ;
 wire \soc_inst.core_mem_addr[8] ;
 wire \soc_inst.core_mem_addr[9] ;
 wire \soc_inst.core_mem_flag[0] ;
 wire \soc_inst.core_mem_flag[1] ;
 wire \soc_inst.core_mem_flag[2] ;
 wire \soc_inst.core_mem_rdata[0] ;
 wire \soc_inst.core_mem_rdata[10] ;
 wire \soc_inst.core_mem_rdata[11] ;
 wire \soc_inst.core_mem_rdata[12] ;
 wire \soc_inst.core_mem_rdata[13] ;
 wire \soc_inst.core_mem_rdata[14] ;
 wire \soc_inst.core_mem_rdata[15] ;
 wire \soc_inst.core_mem_rdata[16] ;
 wire \soc_inst.core_mem_rdata[17] ;
 wire \soc_inst.core_mem_rdata[18] ;
 wire \soc_inst.core_mem_rdata[19] ;
 wire \soc_inst.core_mem_rdata[1] ;
 wire \soc_inst.core_mem_rdata[20] ;
 wire \soc_inst.core_mem_rdata[21] ;
 wire \soc_inst.core_mem_rdata[22] ;
 wire \soc_inst.core_mem_rdata[23] ;
 wire \soc_inst.core_mem_rdata[24] ;
 wire \soc_inst.core_mem_rdata[25] ;
 wire \soc_inst.core_mem_rdata[26] ;
 wire \soc_inst.core_mem_rdata[27] ;
 wire \soc_inst.core_mem_rdata[28] ;
 wire \soc_inst.core_mem_rdata[29] ;
 wire \soc_inst.core_mem_rdata[2] ;
 wire \soc_inst.core_mem_rdata[30] ;
 wire \soc_inst.core_mem_rdata[31] ;
 wire \soc_inst.core_mem_rdata[3] ;
 wire \soc_inst.core_mem_rdata[4] ;
 wire \soc_inst.core_mem_rdata[5] ;
 wire \soc_inst.core_mem_rdata[6] ;
 wire \soc_inst.core_mem_rdata[7] ;
 wire \soc_inst.core_mem_rdata[8] ;
 wire \soc_inst.core_mem_rdata[9] ;
 wire \soc_inst.core_mem_re ;
 wire \soc_inst.core_mem_wdata[0] ;
 wire \soc_inst.core_mem_wdata[10] ;
 wire \soc_inst.core_mem_wdata[11] ;
 wire \soc_inst.core_mem_wdata[12] ;
 wire \soc_inst.core_mem_wdata[13] ;
 wire \soc_inst.core_mem_wdata[14] ;
 wire \soc_inst.core_mem_wdata[15] ;
 wire \soc_inst.core_mem_wdata[16] ;
 wire \soc_inst.core_mem_wdata[17] ;
 wire \soc_inst.core_mem_wdata[18] ;
 wire \soc_inst.core_mem_wdata[19] ;
 wire \soc_inst.core_mem_wdata[1] ;
 wire \soc_inst.core_mem_wdata[20] ;
 wire \soc_inst.core_mem_wdata[21] ;
 wire \soc_inst.core_mem_wdata[22] ;
 wire \soc_inst.core_mem_wdata[23] ;
 wire \soc_inst.core_mem_wdata[24] ;
 wire \soc_inst.core_mem_wdata[25] ;
 wire \soc_inst.core_mem_wdata[26] ;
 wire \soc_inst.core_mem_wdata[27] ;
 wire \soc_inst.core_mem_wdata[28] ;
 wire \soc_inst.core_mem_wdata[29] ;
 wire \soc_inst.core_mem_wdata[2] ;
 wire \soc_inst.core_mem_wdata[30] ;
 wire \soc_inst.core_mem_wdata[31] ;
 wire \soc_inst.core_mem_wdata[3] ;
 wire \soc_inst.core_mem_wdata[4] ;
 wire \soc_inst.core_mem_wdata[5] ;
 wire \soc_inst.core_mem_wdata[6] ;
 wire \soc_inst.core_mem_wdata[7] ;
 wire \soc_inst.core_mem_wdata[8] ;
 wire \soc_inst.core_mem_wdata[9] ;
 wire \soc_inst.core_mem_we ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[0] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[1] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[2] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[3] ;
 wire \soc_inst.cpu_core._unused_mem_rd_addr[4] ;
 wire \soc_inst.cpu_core.alu.a[0] ;
 wire \soc_inst.cpu_core.alu.a[10] ;
 wire \soc_inst.cpu_core.alu.a[11] ;
 wire \soc_inst.cpu_core.alu.a[12] ;
 wire \soc_inst.cpu_core.alu.a[13] ;
 wire \soc_inst.cpu_core.alu.a[14] ;
 wire \soc_inst.cpu_core.alu.a[15] ;
 wire \soc_inst.cpu_core.alu.a[16] ;
 wire \soc_inst.cpu_core.alu.a[17] ;
 wire \soc_inst.cpu_core.alu.a[18] ;
 wire \soc_inst.cpu_core.alu.a[19] ;
 wire \soc_inst.cpu_core.alu.a[1] ;
 wire \soc_inst.cpu_core.alu.a[20] ;
 wire \soc_inst.cpu_core.alu.a[21] ;
 wire \soc_inst.cpu_core.alu.a[22] ;
 wire \soc_inst.cpu_core.alu.a[23] ;
 wire \soc_inst.cpu_core.alu.a[24] ;
 wire \soc_inst.cpu_core.alu.a[25] ;
 wire \soc_inst.cpu_core.alu.a[26] ;
 wire \soc_inst.cpu_core.alu.a[27] ;
 wire \soc_inst.cpu_core.alu.a[28] ;
 wire \soc_inst.cpu_core.alu.a[29] ;
 wire \soc_inst.cpu_core.alu.a[2] ;
 wire \soc_inst.cpu_core.alu.a[30] ;
 wire \soc_inst.cpu_core.alu.a[31] ;
 wire \soc_inst.cpu_core.alu.a[3] ;
 wire \soc_inst.cpu_core.alu.a[4] ;
 wire \soc_inst.cpu_core.alu.a[5] ;
 wire \soc_inst.cpu_core.alu.a[6] ;
 wire \soc_inst.cpu_core.alu.a[7] ;
 wire \soc_inst.cpu_core.alu.a[8] ;
 wire \soc_inst.cpu_core.alu.a[9] ;
 wire \soc_inst.cpu_core.alu.b[0] ;
 wire \soc_inst.cpu_core.alu.b[10] ;
 wire \soc_inst.cpu_core.alu.b[11] ;
 wire \soc_inst.cpu_core.alu.b[12] ;
 wire \soc_inst.cpu_core.alu.b[13] ;
 wire \soc_inst.cpu_core.alu.b[14] ;
 wire \soc_inst.cpu_core.alu.b[15] ;
 wire \soc_inst.cpu_core.alu.b[16] ;
 wire \soc_inst.cpu_core.alu.b[17] ;
 wire \soc_inst.cpu_core.alu.b[18] ;
 wire \soc_inst.cpu_core.alu.b[19] ;
 wire \soc_inst.cpu_core.alu.b[1] ;
 wire \soc_inst.cpu_core.alu.b[20] ;
 wire \soc_inst.cpu_core.alu.b[21] ;
 wire \soc_inst.cpu_core.alu.b[22] ;
 wire \soc_inst.cpu_core.alu.b[23] ;
 wire \soc_inst.cpu_core.alu.b[24] ;
 wire \soc_inst.cpu_core.alu.b[25] ;
 wire \soc_inst.cpu_core.alu.b[26] ;
 wire \soc_inst.cpu_core.alu.b[27] ;
 wire \soc_inst.cpu_core.alu.b[28] ;
 wire \soc_inst.cpu_core.alu.b[29] ;
 wire \soc_inst.cpu_core.alu.b[2] ;
 wire \soc_inst.cpu_core.alu.b[30] ;
 wire \soc_inst.cpu_core.alu.b[31] ;
 wire \soc_inst.cpu_core.alu.b[3] ;
 wire \soc_inst.cpu_core.alu.b[4] ;
 wire \soc_inst.cpu_core.alu.b[5] ;
 wire \soc_inst.cpu_core.alu.b[6] ;
 wire \soc_inst.cpu_core.alu.b[7] ;
 wire \soc_inst.cpu_core.alu.b[8] ;
 wire \soc_inst.cpu_core.alu.b[9] ;
 wire \soc_inst.cpu_core.alu.op[0] ;
 wire \soc_inst.cpu_core.alu.op[1] ;
 wire \soc_inst.cpu_core.alu.op[2] ;
 wire \soc_inst.cpu_core.alu.op[3] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[0] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[10] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[11] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[1] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[2] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[3] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[4] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[5] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[6] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[7] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[8] ;
 wire \soc_inst.cpu_core.csr_file.csr_addr[9] ;
 wire \soc_inst.cpu_core.csr_file.external_interrupt ;
 wire \soc_inst.cpu_core.csr_file.mcause[0] ;
 wire \soc_inst.cpu_core.csr_file.mcause[10] ;
 wire \soc_inst.cpu_core.csr_file.mcause[11] ;
 wire \soc_inst.cpu_core.csr_file.mcause[12] ;
 wire \soc_inst.cpu_core.csr_file.mcause[13] ;
 wire \soc_inst.cpu_core.csr_file.mcause[14] ;
 wire \soc_inst.cpu_core.csr_file.mcause[15] ;
 wire \soc_inst.cpu_core.csr_file.mcause[16] ;
 wire \soc_inst.cpu_core.csr_file.mcause[17] ;
 wire \soc_inst.cpu_core.csr_file.mcause[18] ;
 wire \soc_inst.cpu_core.csr_file.mcause[19] ;
 wire \soc_inst.cpu_core.csr_file.mcause[1] ;
 wire \soc_inst.cpu_core.csr_file.mcause[20] ;
 wire \soc_inst.cpu_core.csr_file.mcause[21] ;
 wire \soc_inst.cpu_core.csr_file.mcause[22] ;
 wire \soc_inst.cpu_core.csr_file.mcause[23] ;
 wire \soc_inst.cpu_core.csr_file.mcause[24] ;
 wire \soc_inst.cpu_core.csr_file.mcause[25] ;
 wire \soc_inst.cpu_core.csr_file.mcause[26] ;
 wire \soc_inst.cpu_core.csr_file.mcause[27] ;
 wire \soc_inst.cpu_core.csr_file.mcause[28] ;
 wire \soc_inst.cpu_core.csr_file.mcause[29] ;
 wire \soc_inst.cpu_core.csr_file.mcause[2] ;
 wire \soc_inst.cpu_core.csr_file.mcause[30] ;
 wire \soc_inst.cpu_core.csr_file.mcause[31] ;
 wire \soc_inst.cpu_core.csr_file.mcause[3] ;
 wire \soc_inst.cpu_core.csr_file.mcause[4] ;
 wire \soc_inst.cpu_core.csr_file.mcause[5] ;
 wire \soc_inst.cpu_core.csr_file.mcause[6] ;
 wire \soc_inst.cpu_core.csr_file.mcause[7] ;
 wire \soc_inst.cpu_core.csr_file.mcause[8] ;
 wire \soc_inst.cpu_core.csr_file.mcause[9] ;
 wire \soc_inst.cpu_core.csr_file.mepc[0] ;
 wire \soc_inst.cpu_core.csr_file.mepc[10] ;
 wire \soc_inst.cpu_core.csr_file.mepc[11] ;
 wire \soc_inst.cpu_core.csr_file.mepc[12] ;
 wire \soc_inst.cpu_core.csr_file.mepc[13] ;
 wire \soc_inst.cpu_core.csr_file.mepc[14] ;
 wire \soc_inst.cpu_core.csr_file.mepc[15] ;
 wire \soc_inst.cpu_core.csr_file.mepc[16] ;
 wire \soc_inst.cpu_core.csr_file.mepc[17] ;
 wire \soc_inst.cpu_core.csr_file.mepc[18] ;
 wire \soc_inst.cpu_core.csr_file.mepc[19] ;
 wire \soc_inst.cpu_core.csr_file.mepc[1] ;
 wire \soc_inst.cpu_core.csr_file.mepc[20] ;
 wire \soc_inst.cpu_core.csr_file.mepc[21] ;
 wire \soc_inst.cpu_core.csr_file.mepc[22] ;
 wire \soc_inst.cpu_core.csr_file.mepc[23] ;
 wire \soc_inst.cpu_core.csr_file.mepc[2] ;
 wire \soc_inst.cpu_core.csr_file.mepc[3] ;
 wire \soc_inst.cpu_core.csr_file.mepc[4] ;
 wire \soc_inst.cpu_core.csr_file.mepc[5] ;
 wire \soc_inst.cpu_core.csr_file.mepc[6] ;
 wire \soc_inst.cpu_core.csr_file.mepc[7] ;
 wire \soc_inst.cpu_core.csr_file.mepc[8] ;
 wire \soc_inst.cpu_core.csr_file.mepc[9] ;
 wire \soc_inst.cpu_core.csr_file.mie[11] ;
 wire \soc_inst.cpu_core.csr_file.mie[7] ;
 wire \soc_inst.cpu_core.csr_file.mip_eip ;
 wire \soc_inst.cpu_core.csr_file.mip_tip ;
 wire \soc_inst.cpu_core.csr_file.mret_trigger ;
 wire \soc_inst.cpu_core.csr_file.mscratch[0] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[10] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[11] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[12] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[13] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[14] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[15] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[16] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[17] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[18] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[19] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[1] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[20] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[21] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[22] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[23] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[24] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[25] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[26] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[27] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[28] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[29] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[2] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[30] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[31] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[3] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[4] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[5] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[6] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[7] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[8] ;
 wire \soc_inst.cpu_core.csr_file.mscratch[9] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[0] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[10] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[13] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[14] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[15] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[16] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[17] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[18] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[19] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[1] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[20] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[21] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[22] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[23] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[24] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[25] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[26] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[27] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[28] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[29] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[2] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[30] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[31] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[3] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[4] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[5] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[6] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[7] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[8] ;
 wire \soc_inst.cpu_core.csr_file.mstatus[9] ;
 wire \soc_inst.cpu_core.csr_file.mtime[0] ;
 wire \soc_inst.cpu_core.csr_file.mtime[10] ;
 wire \soc_inst.cpu_core.csr_file.mtime[11] ;
 wire \soc_inst.cpu_core.csr_file.mtime[12] ;
 wire \soc_inst.cpu_core.csr_file.mtime[13] ;
 wire \soc_inst.cpu_core.csr_file.mtime[14] ;
 wire \soc_inst.cpu_core.csr_file.mtime[15] ;
 wire \soc_inst.cpu_core.csr_file.mtime[16] ;
 wire \soc_inst.cpu_core.csr_file.mtime[17] ;
 wire \soc_inst.cpu_core.csr_file.mtime[18] ;
 wire \soc_inst.cpu_core.csr_file.mtime[19] ;
 wire \soc_inst.cpu_core.csr_file.mtime[1] ;
 wire \soc_inst.cpu_core.csr_file.mtime[20] ;
 wire \soc_inst.cpu_core.csr_file.mtime[21] ;
 wire \soc_inst.cpu_core.csr_file.mtime[22] ;
 wire \soc_inst.cpu_core.csr_file.mtime[23] ;
 wire \soc_inst.cpu_core.csr_file.mtime[24] ;
 wire \soc_inst.cpu_core.csr_file.mtime[25] ;
 wire \soc_inst.cpu_core.csr_file.mtime[26] ;
 wire \soc_inst.cpu_core.csr_file.mtime[27] ;
 wire \soc_inst.cpu_core.csr_file.mtime[28] ;
 wire \soc_inst.cpu_core.csr_file.mtime[29] ;
 wire \soc_inst.cpu_core.csr_file.mtime[2] ;
 wire \soc_inst.cpu_core.csr_file.mtime[30] ;
 wire \soc_inst.cpu_core.csr_file.mtime[31] ;
 wire \soc_inst.cpu_core.csr_file.mtime[32] ;
 wire \soc_inst.cpu_core.csr_file.mtime[33] ;
 wire \soc_inst.cpu_core.csr_file.mtime[34] ;
 wire \soc_inst.cpu_core.csr_file.mtime[35] ;
 wire \soc_inst.cpu_core.csr_file.mtime[36] ;
 wire \soc_inst.cpu_core.csr_file.mtime[37] ;
 wire \soc_inst.cpu_core.csr_file.mtime[38] ;
 wire \soc_inst.cpu_core.csr_file.mtime[39] ;
 wire \soc_inst.cpu_core.csr_file.mtime[3] ;
 wire \soc_inst.cpu_core.csr_file.mtime[40] ;
 wire \soc_inst.cpu_core.csr_file.mtime[41] ;
 wire \soc_inst.cpu_core.csr_file.mtime[42] ;
 wire \soc_inst.cpu_core.csr_file.mtime[43] ;
 wire \soc_inst.cpu_core.csr_file.mtime[44] ;
 wire \soc_inst.cpu_core.csr_file.mtime[45] ;
 wire \soc_inst.cpu_core.csr_file.mtime[46] ;
 wire \soc_inst.cpu_core.csr_file.mtime[47] ;
 wire \soc_inst.cpu_core.csr_file.mtime[4] ;
 wire \soc_inst.cpu_core.csr_file.mtime[5] ;
 wire \soc_inst.cpu_core.csr_file.mtime[6] ;
 wire \soc_inst.cpu_core.csr_file.mtime[7] ;
 wire \soc_inst.cpu_core.csr_file.mtime[8] ;
 wire \soc_inst.cpu_core.csr_file.mtime[9] ;
 wire \soc_inst.cpu_core.csr_file.mtval[0] ;
 wire \soc_inst.cpu_core.csr_file.mtval[10] ;
 wire \soc_inst.cpu_core.csr_file.mtval[11] ;
 wire \soc_inst.cpu_core.csr_file.mtval[12] ;
 wire \soc_inst.cpu_core.csr_file.mtval[13] ;
 wire \soc_inst.cpu_core.csr_file.mtval[14] ;
 wire \soc_inst.cpu_core.csr_file.mtval[15] ;
 wire \soc_inst.cpu_core.csr_file.mtval[16] ;
 wire \soc_inst.cpu_core.csr_file.mtval[17] ;
 wire \soc_inst.cpu_core.csr_file.mtval[18] ;
 wire \soc_inst.cpu_core.csr_file.mtval[19] ;
 wire \soc_inst.cpu_core.csr_file.mtval[1] ;
 wire \soc_inst.cpu_core.csr_file.mtval[20] ;
 wire \soc_inst.cpu_core.csr_file.mtval[21] ;
 wire \soc_inst.cpu_core.csr_file.mtval[22] ;
 wire \soc_inst.cpu_core.csr_file.mtval[23] ;
 wire \soc_inst.cpu_core.csr_file.mtval[24] ;
 wire \soc_inst.cpu_core.csr_file.mtval[25] ;
 wire \soc_inst.cpu_core.csr_file.mtval[26] ;
 wire \soc_inst.cpu_core.csr_file.mtval[27] ;
 wire \soc_inst.cpu_core.csr_file.mtval[28] ;
 wire \soc_inst.cpu_core.csr_file.mtval[29] ;
 wire \soc_inst.cpu_core.csr_file.mtval[2] ;
 wire \soc_inst.cpu_core.csr_file.mtval[30] ;
 wire \soc_inst.cpu_core.csr_file.mtval[31] ;
 wire \soc_inst.cpu_core.csr_file.mtval[3] ;
 wire \soc_inst.cpu_core.csr_file.mtval[4] ;
 wire \soc_inst.cpu_core.csr_file.mtval[5] ;
 wire \soc_inst.cpu_core.csr_file.mtval[6] ;
 wire \soc_inst.cpu_core.csr_file.mtval[7] ;
 wire \soc_inst.cpu_core.csr_file.mtval[8] ;
 wire \soc_inst.cpu_core.csr_file.mtval[9] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[0] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[10] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[11] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[12] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[13] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[14] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[15] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[16] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[17] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[18] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[19] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[1] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[20] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[21] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[22] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[23] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[2] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[3] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[4] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[5] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[6] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[7] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[8] ;
 wire \soc_inst.cpu_core.csr_file.mtvec[9] ;
 wire \soc_inst.cpu_core.csr_file.timer_interrupt ;
 wire \soc_inst.cpu_core.error_flag_reg ;
 wire \soc_inst.cpu_core.ex_alu_result[0] ;
 wire \soc_inst.cpu_core.ex_alu_result[10] ;
 wire \soc_inst.cpu_core.ex_alu_result[11] ;
 wire \soc_inst.cpu_core.ex_alu_result[12] ;
 wire \soc_inst.cpu_core.ex_alu_result[13] ;
 wire \soc_inst.cpu_core.ex_alu_result[14] ;
 wire \soc_inst.cpu_core.ex_alu_result[15] ;
 wire \soc_inst.cpu_core.ex_alu_result[16] ;
 wire \soc_inst.cpu_core.ex_alu_result[17] ;
 wire \soc_inst.cpu_core.ex_alu_result[18] ;
 wire \soc_inst.cpu_core.ex_alu_result[19] ;
 wire \soc_inst.cpu_core.ex_alu_result[1] ;
 wire \soc_inst.cpu_core.ex_alu_result[20] ;
 wire \soc_inst.cpu_core.ex_alu_result[21] ;
 wire \soc_inst.cpu_core.ex_alu_result[22] ;
 wire \soc_inst.cpu_core.ex_alu_result[23] ;
 wire \soc_inst.cpu_core.ex_alu_result[24] ;
 wire \soc_inst.cpu_core.ex_alu_result[25] ;
 wire \soc_inst.cpu_core.ex_alu_result[26] ;
 wire \soc_inst.cpu_core.ex_alu_result[27] ;
 wire \soc_inst.cpu_core.ex_alu_result[28] ;
 wire \soc_inst.cpu_core.ex_alu_result[29] ;
 wire \soc_inst.cpu_core.ex_alu_result[2] ;
 wire \soc_inst.cpu_core.ex_alu_result[30] ;
 wire \soc_inst.cpu_core.ex_alu_result[31] ;
 wire \soc_inst.cpu_core.ex_alu_result[3] ;
 wire \soc_inst.cpu_core.ex_alu_result[4] ;
 wire \soc_inst.cpu_core.ex_alu_result[5] ;
 wire \soc_inst.cpu_core.ex_alu_result[6] ;
 wire \soc_inst.cpu_core.ex_alu_result[7] ;
 wire \soc_inst.cpu_core.ex_alu_result[8] ;
 wire \soc_inst.cpu_core.ex_alu_result[9] ;
 wire \soc_inst.cpu_core.ex_branch_target[0] ;
 wire \soc_inst.cpu_core.ex_branch_target[10] ;
 wire \soc_inst.cpu_core.ex_branch_target[11] ;
 wire \soc_inst.cpu_core.ex_branch_target[12] ;
 wire \soc_inst.cpu_core.ex_branch_target[13] ;
 wire \soc_inst.cpu_core.ex_branch_target[14] ;
 wire \soc_inst.cpu_core.ex_branch_target[15] ;
 wire \soc_inst.cpu_core.ex_branch_target[16] ;
 wire \soc_inst.cpu_core.ex_branch_target[17] ;
 wire \soc_inst.cpu_core.ex_branch_target[18] ;
 wire \soc_inst.cpu_core.ex_branch_target[19] ;
 wire \soc_inst.cpu_core.ex_branch_target[1] ;
 wire \soc_inst.cpu_core.ex_branch_target[20] ;
 wire \soc_inst.cpu_core.ex_branch_target[21] ;
 wire \soc_inst.cpu_core.ex_branch_target[22] ;
 wire \soc_inst.cpu_core.ex_branch_target[23] ;
 wire \soc_inst.cpu_core.ex_branch_target[24] ;
 wire \soc_inst.cpu_core.ex_branch_target[25] ;
 wire \soc_inst.cpu_core.ex_branch_target[26] ;
 wire \soc_inst.cpu_core.ex_branch_target[27] ;
 wire \soc_inst.cpu_core.ex_branch_target[28] ;
 wire \soc_inst.cpu_core.ex_branch_target[29] ;
 wire \soc_inst.cpu_core.ex_branch_target[2] ;
 wire \soc_inst.cpu_core.ex_branch_target[30] ;
 wire \soc_inst.cpu_core.ex_branch_target[31] ;
 wire \soc_inst.cpu_core.ex_branch_target[3] ;
 wire \soc_inst.cpu_core.ex_branch_target[4] ;
 wire \soc_inst.cpu_core.ex_branch_target[5] ;
 wire \soc_inst.cpu_core.ex_branch_target[6] ;
 wire \soc_inst.cpu_core.ex_branch_target[7] ;
 wire \soc_inst.cpu_core.ex_branch_target[8] ;
 wire \soc_inst.cpu_core.ex_branch_target[9] ;
 wire \soc_inst.cpu_core.ex_exception_pc[0] ;
 wire \soc_inst.cpu_core.ex_exception_pc[10] ;
 wire \soc_inst.cpu_core.ex_exception_pc[11] ;
 wire \soc_inst.cpu_core.ex_exception_pc[12] ;
 wire \soc_inst.cpu_core.ex_exception_pc[13] ;
 wire \soc_inst.cpu_core.ex_exception_pc[14] ;
 wire \soc_inst.cpu_core.ex_exception_pc[15] ;
 wire \soc_inst.cpu_core.ex_exception_pc[16] ;
 wire \soc_inst.cpu_core.ex_exception_pc[17] ;
 wire \soc_inst.cpu_core.ex_exception_pc[18] ;
 wire \soc_inst.cpu_core.ex_exception_pc[19] ;
 wire \soc_inst.cpu_core.ex_exception_pc[1] ;
 wire \soc_inst.cpu_core.ex_exception_pc[20] ;
 wire \soc_inst.cpu_core.ex_exception_pc[21] ;
 wire \soc_inst.cpu_core.ex_exception_pc[22] ;
 wire \soc_inst.cpu_core.ex_exception_pc[23] ;
 wire \soc_inst.cpu_core.ex_exception_pc[2] ;
 wire \soc_inst.cpu_core.ex_exception_pc[3] ;
 wire \soc_inst.cpu_core.ex_exception_pc[4] ;
 wire \soc_inst.cpu_core.ex_exception_pc[5] ;
 wire \soc_inst.cpu_core.ex_exception_pc[6] ;
 wire \soc_inst.cpu_core.ex_exception_pc[7] ;
 wire \soc_inst.cpu_core.ex_exception_pc[8] ;
 wire \soc_inst.cpu_core.ex_exception_pc[9] ;
 wire \soc_inst.cpu_core.ex_funct3[0] ;
 wire \soc_inst.cpu_core.ex_funct3[1] ;
 wire \soc_inst.cpu_core.ex_funct3[2] ;
 wire \soc_inst.cpu_core.ex_funct7[0] ;
 wire \soc_inst.cpu_core.ex_funct7[1] ;
 wire \soc_inst.cpu_core.ex_funct7[2] ;
 wire \soc_inst.cpu_core.ex_funct7[3] ;
 wire \soc_inst.cpu_core.ex_funct7[4] ;
 wire \soc_inst.cpu_core.ex_funct7[5] ;
 wire \soc_inst.cpu_core.ex_funct7[6] ;
 wire \soc_inst.cpu_core.ex_instr[10] ;
 wire \soc_inst.cpu_core.ex_instr[11] ;
 wire \soc_inst.cpu_core.ex_instr[15] ;
 wire \soc_inst.cpu_core.ex_instr[16] ;
 wire \soc_inst.cpu_core.ex_instr[17] ;
 wire \soc_inst.cpu_core.ex_instr[18] ;
 wire \soc_inst.cpu_core.ex_instr[19] ;
 wire \soc_inst.cpu_core.ex_instr[20] ;
 wire \soc_inst.cpu_core.ex_instr[21] ;
 wire \soc_inst.cpu_core.ex_instr[22] ;
 wire \soc_inst.cpu_core.ex_instr[23] ;
 wire \soc_inst.cpu_core.ex_instr[24] ;
 wire \soc_inst.cpu_core.ex_instr[2] ;
 wire \soc_inst.cpu_core.ex_instr[3] ;
 wire \soc_inst.cpu_core.ex_instr[5] ;
 wire \soc_inst.cpu_core.ex_instr[6] ;
 wire \soc_inst.cpu_core.ex_instr[7] ;
 wire \soc_inst.cpu_core.ex_instr[8] ;
 wire \soc_inst.cpu_core.ex_instr[9] ;
 wire \soc_inst.cpu_core.ex_is_ebreak ;
 wire \soc_inst.cpu_core.ex_is_ecall ;
 wire \soc_inst.cpu_core.ex_mem_re ;
 wire \soc_inst.cpu_core.ex_mem_we ;
 wire \soc_inst.cpu_core.ex_reg_we ;
 wire \soc_inst.cpu_core.ex_rs1_data[0] ;
 wire \soc_inst.cpu_core.ex_rs1_data[10] ;
 wire \soc_inst.cpu_core.ex_rs1_data[11] ;
 wire \soc_inst.cpu_core.ex_rs1_data[12] ;
 wire \soc_inst.cpu_core.ex_rs1_data[13] ;
 wire \soc_inst.cpu_core.ex_rs1_data[14] ;
 wire \soc_inst.cpu_core.ex_rs1_data[15] ;
 wire \soc_inst.cpu_core.ex_rs1_data[16] ;
 wire \soc_inst.cpu_core.ex_rs1_data[17] ;
 wire \soc_inst.cpu_core.ex_rs1_data[18] ;
 wire \soc_inst.cpu_core.ex_rs1_data[19] ;
 wire \soc_inst.cpu_core.ex_rs1_data[1] ;
 wire \soc_inst.cpu_core.ex_rs1_data[20] ;
 wire \soc_inst.cpu_core.ex_rs1_data[21] ;
 wire \soc_inst.cpu_core.ex_rs1_data[22] ;
 wire \soc_inst.cpu_core.ex_rs1_data[23] ;
 wire \soc_inst.cpu_core.ex_rs1_data[24] ;
 wire \soc_inst.cpu_core.ex_rs1_data[25] ;
 wire \soc_inst.cpu_core.ex_rs1_data[26] ;
 wire \soc_inst.cpu_core.ex_rs1_data[27] ;
 wire \soc_inst.cpu_core.ex_rs1_data[28] ;
 wire \soc_inst.cpu_core.ex_rs1_data[29] ;
 wire \soc_inst.cpu_core.ex_rs1_data[2] ;
 wire \soc_inst.cpu_core.ex_rs1_data[30] ;
 wire \soc_inst.cpu_core.ex_rs1_data[31] ;
 wire \soc_inst.cpu_core.ex_rs1_data[3] ;
 wire \soc_inst.cpu_core.ex_rs1_data[4] ;
 wire \soc_inst.cpu_core.ex_rs1_data[5] ;
 wire \soc_inst.cpu_core.ex_rs1_data[6] ;
 wire \soc_inst.cpu_core.ex_rs1_data[7] ;
 wire \soc_inst.cpu_core.ex_rs1_data[8] ;
 wire \soc_inst.cpu_core.ex_rs1_data[9] ;
 wire \soc_inst.cpu_core.ex_rs2_data[0] ;
 wire \soc_inst.cpu_core.ex_rs2_data[10] ;
 wire \soc_inst.cpu_core.ex_rs2_data[11] ;
 wire \soc_inst.cpu_core.ex_rs2_data[12] ;
 wire \soc_inst.cpu_core.ex_rs2_data[13] ;
 wire \soc_inst.cpu_core.ex_rs2_data[14] ;
 wire \soc_inst.cpu_core.ex_rs2_data[15] ;
 wire \soc_inst.cpu_core.ex_rs2_data[16] ;
 wire \soc_inst.cpu_core.ex_rs2_data[17] ;
 wire \soc_inst.cpu_core.ex_rs2_data[18] ;
 wire \soc_inst.cpu_core.ex_rs2_data[19] ;
 wire \soc_inst.cpu_core.ex_rs2_data[1] ;
 wire \soc_inst.cpu_core.ex_rs2_data[20] ;
 wire \soc_inst.cpu_core.ex_rs2_data[21] ;
 wire \soc_inst.cpu_core.ex_rs2_data[22] ;
 wire \soc_inst.cpu_core.ex_rs2_data[23] ;
 wire \soc_inst.cpu_core.ex_rs2_data[24] ;
 wire \soc_inst.cpu_core.ex_rs2_data[25] ;
 wire \soc_inst.cpu_core.ex_rs2_data[26] ;
 wire \soc_inst.cpu_core.ex_rs2_data[27] ;
 wire \soc_inst.cpu_core.ex_rs2_data[28] ;
 wire \soc_inst.cpu_core.ex_rs2_data[29] ;
 wire \soc_inst.cpu_core.ex_rs2_data[2] ;
 wire \soc_inst.cpu_core.ex_rs2_data[30] ;
 wire \soc_inst.cpu_core.ex_rs2_data[31] ;
 wire \soc_inst.cpu_core.ex_rs2_data[3] ;
 wire \soc_inst.cpu_core.ex_rs2_data[4] ;
 wire \soc_inst.cpu_core.ex_rs2_data[5] ;
 wire \soc_inst.cpu_core.ex_rs2_data[6] ;
 wire \soc_inst.cpu_core.ex_rs2_data[7] ;
 wire \soc_inst.cpu_core.ex_rs2_data[8] ;
 wire \soc_inst.cpu_core.ex_rs2_data[9] ;
 wire \soc_inst.cpu_core.i_mem_ready ;
 wire \soc_inst.cpu_core.id_funct3[0] ;
 wire \soc_inst.cpu_core.id_funct3[1] ;
 wire \soc_inst.cpu_core.id_funct3[2] ;
 wire \soc_inst.cpu_core.id_imm12[0] ;
 wire \soc_inst.cpu_core.id_imm12[10] ;
 wire \soc_inst.cpu_core.id_imm12[11] ;
 wire \soc_inst.cpu_core.id_imm12[1] ;
 wire \soc_inst.cpu_core.id_imm12[2] ;
 wire \soc_inst.cpu_core.id_imm12[3] ;
 wire \soc_inst.cpu_core.id_imm12[4] ;
 wire \soc_inst.cpu_core.id_imm12[5] ;
 wire \soc_inst.cpu_core.id_imm12[6] ;
 wire \soc_inst.cpu_core.id_imm12[7] ;
 wire \soc_inst.cpu_core.id_imm12[8] ;
 wire \soc_inst.cpu_core.id_imm12[9] ;
 wire \soc_inst.cpu_core.id_imm[0] ;
 wire \soc_inst.cpu_core.id_imm[10] ;
 wire \soc_inst.cpu_core.id_imm[11] ;
 wire \soc_inst.cpu_core.id_imm[12] ;
 wire \soc_inst.cpu_core.id_imm[13] ;
 wire \soc_inst.cpu_core.id_imm[14] ;
 wire \soc_inst.cpu_core.id_imm[15] ;
 wire \soc_inst.cpu_core.id_imm[16] ;
 wire \soc_inst.cpu_core.id_imm[17] ;
 wire \soc_inst.cpu_core.id_imm[18] ;
 wire \soc_inst.cpu_core.id_imm[19] ;
 wire \soc_inst.cpu_core.id_imm[1] ;
 wire \soc_inst.cpu_core.id_imm[20] ;
 wire \soc_inst.cpu_core.id_imm[21] ;
 wire \soc_inst.cpu_core.id_imm[22] ;
 wire \soc_inst.cpu_core.id_imm[23] ;
 wire \soc_inst.cpu_core.id_imm[24] ;
 wire \soc_inst.cpu_core.id_imm[25] ;
 wire \soc_inst.cpu_core.id_imm[26] ;
 wire \soc_inst.cpu_core.id_imm[27] ;
 wire \soc_inst.cpu_core.id_imm[28] ;
 wire \soc_inst.cpu_core.id_imm[29] ;
 wire \soc_inst.cpu_core.id_imm[2] ;
 wire \soc_inst.cpu_core.id_imm[30] ;
 wire \soc_inst.cpu_core.id_imm[31] ;
 wire \soc_inst.cpu_core.id_imm[3] ;
 wire \soc_inst.cpu_core.id_imm[4] ;
 wire \soc_inst.cpu_core.id_imm[5] ;
 wire \soc_inst.cpu_core.id_imm[6] ;
 wire \soc_inst.cpu_core.id_imm[7] ;
 wire \soc_inst.cpu_core.id_imm[8] ;
 wire \soc_inst.cpu_core.id_imm[9] ;
 wire \soc_inst.cpu_core.id_instr[10] ;
 wire \soc_inst.cpu_core.id_instr[11] ;
 wire \soc_inst.cpu_core.id_instr[15] ;
 wire \soc_inst.cpu_core.id_instr[16] ;
 wire \soc_inst.cpu_core.id_instr[17] ;
 wire \soc_inst.cpu_core.id_instr[18] ;
 wire \soc_inst.cpu_core.id_instr[19] ;
 wire \soc_inst.cpu_core.id_instr[2] ;
 wire \soc_inst.cpu_core.id_instr[3] ;
 wire \soc_inst.cpu_core.id_instr[5] ;
 wire \soc_inst.cpu_core.id_instr[6] ;
 wire \soc_inst.cpu_core.id_instr[7] ;
 wire \soc_inst.cpu_core.id_instr[8] ;
 wire \soc_inst.cpu_core.id_instr[9] ;
 wire \soc_inst.cpu_core.id_int_is_interrupt ;
 wire \soc_inst.cpu_core.id_is_compressed ;
 wire \soc_inst.cpu_core.id_pc[0] ;
 wire \soc_inst.cpu_core.id_pc[10] ;
 wire \soc_inst.cpu_core.id_pc[11] ;
 wire \soc_inst.cpu_core.id_pc[12] ;
 wire \soc_inst.cpu_core.id_pc[13] ;
 wire \soc_inst.cpu_core.id_pc[14] ;
 wire \soc_inst.cpu_core.id_pc[15] ;
 wire \soc_inst.cpu_core.id_pc[16] ;
 wire \soc_inst.cpu_core.id_pc[17] ;
 wire \soc_inst.cpu_core.id_pc[18] ;
 wire \soc_inst.cpu_core.id_pc[19] ;
 wire \soc_inst.cpu_core.id_pc[1] ;
 wire \soc_inst.cpu_core.id_pc[20] ;
 wire \soc_inst.cpu_core.id_pc[21] ;
 wire \soc_inst.cpu_core.id_pc[22] ;
 wire \soc_inst.cpu_core.id_pc[23] ;
 wire \soc_inst.cpu_core.id_pc[2] ;
 wire \soc_inst.cpu_core.id_pc[3] ;
 wire \soc_inst.cpu_core.id_pc[4] ;
 wire \soc_inst.cpu_core.id_pc[5] ;
 wire \soc_inst.cpu_core.id_pc[6] ;
 wire \soc_inst.cpu_core.id_pc[7] ;
 wire \soc_inst.cpu_core.id_pc[8] ;
 wire \soc_inst.cpu_core.id_pc[9] ;
 wire \soc_inst.cpu_core.id_rs1_data[0] ;
 wire \soc_inst.cpu_core.id_rs1_data[10] ;
 wire \soc_inst.cpu_core.id_rs1_data[11] ;
 wire \soc_inst.cpu_core.id_rs1_data[12] ;
 wire \soc_inst.cpu_core.id_rs1_data[13] ;
 wire \soc_inst.cpu_core.id_rs1_data[14] ;
 wire \soc_inst.cpu_core.id_rs1_data[15] ;
 wire \soc_inst.cpu_core.id_rs1_data[16] ;
 wire \soc_inst.cpu_core.id_rs1_data[17] ;
 wire \soc_inst.cpu_core.id_rs1_data[18] ;
 wire \soc_inst.cpu_core.id_rs1_data[19] ;
 wire \soc_inst.cpu_core.id_rs1_data[1] ;
 wire \soc_inst.cpu_core.id_rs1_data[20] ;
 wire \soc_inst.cpu_core.id_rs1_data[21] ;
 wire \soc_inst.cpu_core.id_rs1_data[22] ;
 wire \soc_inst.cpu_core.id_rs1_data[23] ;
 wire \soc_inst.cpu_core.id_rs1_data[24] ;
 wire \soc_inst.cpu_core.id_rs1_data[25] ;
 wire \soc_inst.cpu_core.id_rs1_data[26] ;
 wire \soc_inst.cpu_core.id_rs1_data[27] ;
 wire \soc_inst.cpu_core.id_rs1_data[28] ;
 wire \soc_inst.cpu_core.id_rs1_data[29] ;
 wire \soc_inst.cpu_core.id_rs1_data[2] ;
 wire \soc_inst.cpu_core.id_rs1_data[30] ;
 wire \soc_inst.cpu_core.id_rs1_data[31] ;
 wire \soc_inst.cpu_core.id_rs1_data[3] ;
 wire \soc_inst.cpu_core.id_rs1_data[4] ;
 wire \soc_inst.cpu_core.id_rs1_data[5] ;
 wire \soc_inst.cpu_core.id_rs1_data[6] ;
 wire \soc_inst.cpu_core.id_rs1_data[7] ;
 wire \soc_inst.cpu_core.id_rs1_data[8] ;
 wire \soc_inst.cpu_core.id_rs1_data[9] ;
 wire \soc_inst.cpu_core.id_rs2_data[0] ;
 wire \soc_inst.cpu_core.id_rs2_data[10] ;
 wire \soc_inst.cpu_core.id_rs2_data[11] ;
 wire \soc_inst.cpu_core.id_rs2_data[12] ;
 wire \soc_inst.cpu_core.id_rs2_data[13] ;
 wire \soc_inst.cpu_core.id_rs2_data[14] ;
 wire \soc_inst.cpu_core.id_rs2_data[15] ;
 wire \soc_inst.cpu_core.id_rs2_data[16] ;
 wire \soc_inst.cpu_core.id_rs2_data[17] ;
 wire \soc_inst.cpu_core.id_rs2_data[18] ;
 wire \soc_inst.cpu_core.id_rs2_data[19] ;
 wire \soc_inst.cpu_core.id_rs2_data[1] ;
 wire \soc_inst.cpu_core.id_rs2_data[20] ;
 wire \soc_inst.cpu_core.id_rs2_data[21] ;
 wire \soc_inst.cpu_core.id_rs2_data[22] ;
 wire \soc_inst.cpu_core.id_rs2_data[23] ;
 wire \soc_inst.cpu_core.id_rs2_data[24] ;
 wire \soc_inst.cpu_core.id_rs2_data[25] ;
 wire \soc_inst.cpu_core.id_rs2_data[26] ;
 wire \soc_inst.cpu_core.id_rs2_data[27] ;
 wire \soc_inst.cpu_core.id_rs2_data[28] ;
 wire \soc_inst.cpu_core.id_rs2_data[29] ;
 wire \soc_inst.cpu_core.id_rs2_data[2] ;
 wire \soc_inst.cpu_core.id_rs2_data[30] ;
 wire \soc_inst.cpu_core.id_rs2_data[31] ;
 wire \soc_inst.cpu_core.id_rs2_data[3] ;
 wire \soc_inst.cpu_core.id_rs2_data[4] ;
 wire \soc_inst.cpu_core.id_rs2_data[5] ;
 wire \soc_inst.cpu_core.id_rs2_data[6] ;
 wire \soc_inst.cpu_core.id_rs2_data[7] ;
 wire \soc_inst.cpu_core.id_rs2_data[8] ;
 wire \soc_inst.cpu_core.id_rs2_data[9] ;
 wire \soc_inst.cpu_core.if_funct3[0] ;
 wire \soc_inst.cpu_core.if_funct3[1] ;
 wire \soc_inst.cpu_core.if_funct3[2] ;
 wire \soc_inst.cpu_core.if_funct7[0] ;
 wire \soc_inst.cpu_core.if_funct7[1] ;
 wire \soc_inst.cpu_core.if_funct7[2] ;
 wire \soc_inst.cpu_core.if_funct7[3] ;
 wire \soc_inst.cpu_core.if_funct7[4] ;
 wire \soc_inst.cpu_core.if_funct7[5] ;
 wire \soc_inst.cpu_core.if_funct7[6] ;
 wire \soc_inst.cpu_core.if_imm12[0] ;
 wire \soc_inst.cpu_core.if_imm12[1] ;
 wire \soc_inst.cpu_core.if_imm12[2] ;
 wire \soc_inst.cpu_core.if_imm12[3] ;
 wire \soc_inst.cpu_core.if_imm12[4] ;
 wire \soc_inst.cpu_core.if_instr[10] ;
 wire \soc_inst.cpu_core.if_instr[11] ;
 wire \soc_inst.cpu_core.if_instr[15] ;
 wire \soc_inst.cpu_core.if_instr[16] ;
 wire \soc_inst.cpu_core.if_instr[17] ;
 wire \soc_inst.cpu_core.if_instr[18] ;
 wire \soc_inst.cpu_core.if_instr[19] ;
 wire \soc_inst.cpu_core.if_instr[2] ;
 wire \soc_inst.cpu_core.if_instr[3] ;
 wire \soc_inst.cpu_core.if_instr[5] ;
 wire \soc_inst.cpu_core.if_instr[6] ;
 wire \soc_inst.cpu_core.if_instr[7] ;
 wire \soc_inst.cpu_core.if_instr[8] ;
 wire \soc_inst.cpu_core.if_instr[9] ;
 wire \soc_inst.cpu_core.if_is_compressed ;
 wire \soc_inst.cpu_core.if_pc[0] ;
 wire \soc_inst.cpu_core.if_pc[10] ;
 wire \soc_inst.cpu_core.if_pc[11] ;
 wire \soc_inst.cpu_core.if_pc[12] ;
 wire \soc_inst.cpu_core.if_pc[13] ;
 wire \soc_inst.cpu_core.if_pc[14] ;
 wire \soc_inst.cpu_core.if_pc[15] ;
 wire \soc_inst.cpu_core.if_pc[16] ;
 wire \soc_inst.cpu_core.if_pc[17] ;
 wire \soc_inst.cpu_core.if_pc[18] ;
 wire \soc_inst.cpu_core.if_pc[19] ;
 wire \soc_inst.cpu_core.if_pc[1] ;
 wire \soc_inst.cpu_core.if_pc[20] ;
 wire \soc_inst.cpu_core.if_pc[21] ;
 wire \soc_inst.cpu_core.if_pc[22] ;
 wire \soc_inst.cpu_core.if_pc[23] ;
 wire \soc_inst.cpu_core.if_pc[2] ;
 wire \soc_inst.cpu_core.if_pc[3] ;
 wire \soc_inst.cpu_core.if_pc[4] ;
 wire \soc_inst.cpu_core.if_pc[5] ;
 wire \soc_inst.cpu_core.if_pc[6] ;
 wire \soc_inst.cpu_core.if_pc[7] ;
 wire \soc_inst.cpu_core.if_pc[8] ;
 wire \soc_inst.cpu_core.if_pc[9] ;
 wire \soc_inst.cpu_core.mem_instr[15] ;
 wire \soc_inst.cpu_core.mem_instr[16] ;
 wire \soc_inst.cpu_core.mem_instr[17] ;
 wire \soc_inst.cpu_core.mem_instr[18] ;
 wire \soc_inst.cpu_core.mem_instr[19] ;
 wire \soc_inst.cpu_core.mem_instr[2] ;
 wire \soc_inst.cpu_core.mem_instr[3] ;
 wire \soc_inst.cpu_core.mem_instr[5] ;
 wire \soc_inst.cpu_core.mem_instr[6] ;
 wire \soc_inst.cpu_core.mem_reg_we ;
 wire \soc_inst.cpu_core.mem_rs1_data[0] ;
 wire \soc_inst.cpu_core.mem_rs1_data[10] ;
 wire \soc_inst.cpu_core.mem_rs1_data[11] ;
 wire \soc_inst.cpu_core.mem_rs1_data[12] ;
 wire \soc_inst.cpu_core.mem_rs1_data[13] ;
 wire \soc_inst.cpu_core.mem_rs1_data[14] ;
 wire \soc_inst.cpu_core.mem_rs1_data[15] ;
 wire \soc_inst.cpu_core.mem_rs1_data[16] ;
 wire \soc_inst.cpu_core.mem_rs1_data[17] ;
 wire \soc_inst.cpu_core.mem_rs1_data[18] ;
 wire \soc_inst.cpu_core.mem_rs1_data[19] ;
 wire \soc_inst.cpu_core.mem_rs1_data[1] ;
 wire \soc_inst.cpu_core.mem_rs1_data[20] ;
 wire \soc_inst.cpu_core.mem_rs1_data[21] ;
 wire \soc_inst.cpu_core.mem_rs1_data[22] ;
 wire \soc_inst.cpu_core.mem_rs1_data[23] ;
 wire \soc_inst.cpu_core.mem_rs1_data[24] ;
 wire \soc_inst.cpu_core.mem_rs1_data[25] ;
 wire \soc_inst.cpu_core.mem_rs1_data[26] ;
 wire \soc_inst.cpu_core.mem_rs1_data[27] ;
 wire \soc_inst.cpu_core.mem_rs1_data[28] ;
 wire \soc_inst.cpu_core.mem_rs1_data[29] ;
 wire \soc_inst.cpu_core.mem_rs1_data[2] ;
 wire \soc_inst.cpu_core.mem_rs1_data[30] ;
 wire \soc_inst.cpu_core.mem_rs1_data[31] ;
 wire \soc_inst.cpu_core.mem_rs1_data[3] ;
 wire \soc_inst.cpu_core.mem_rs1_data[4] ;
 wire \soc_inst.cpu_core.mem_rs1_data[5] ;
 wire \soc_inst.cpu_core.mem_rs1_data[6] ;
 wire \soc_inst.cpu_core.mem_rs1_data[7] ;
 wire \soc_inst.cpu_core.mem_rs1_data[8] ;
 wire \soc_inst.cpu_core.mem_rs1_data[9] ;
 wire \soc_inst.cpu_core.mem_stall ;
 wire \soc_inst.cpu_core.register_file.registers[10][0] ;
 wire \soc_inst.cpu_core.register_file.registers[10][10] ;
 wire \soc_inst.cpu_core.register_file.registers[10][11] ;
 wire \soc_inst.cpu_core.register_file.registers[10][12] ;
 wire \soc_inst.cpu_core.register_file.registers[10][13] ;
 wire \soc_inst.cpu_core.register_file.registers[10][14] ;
 wire \soc_inst.cpu_core.register_file.registers[10][15] ;
 wire \soc_inst.cpu_core.register_file.registers[10][16] ;
 wire \soc_inst.cpu_core.register_file.registers[10][17] ;
 wire \soc_inst.cpu_core.register_file.registers[10][18] ;
 wire \soc_inst.cpu_core.register_file.registers[10][19] ;
 wire \soc_inst.cpu_core.register_file.registers[10][1] ;
 wire \soc_inst.cpu_core.register_file.registers[10][20] ;
 wire \soc_inst.cpu_core.register_file.registers[10][21] ;
 wire \soc_inst.cpu_core.register_file.registers[10][22] ;
 wire \soc_inst.cpu_core.register_file.registers[10][23] ;
 wire \soc_inst.cpu_core.register_file.registers[10][24] ;
 wire \soc_inst.cpu_core.register_file.registers[10][25] ;
 wire \soc_inst.cpu_core.register_file.registers[10][26] ;
 wire \soc_inst.cpu_core.register_file.registers[10][27] ;
 wire \soc_inst.cpu_core.register_file.registers[10][28] ;
 wire \soc_inst.cpu_core.register_file.registers[10][29] ;
 wire \soc_inst.cpu_core.register_file.registers[10][2] ;
 wire \soc_inst.cpu_core.register_file.registers[10][30] ;
 wire \soc_inst.cpu_core.register_file.registers[10][31] ;
 wire \soc_inst.cpu_core.register_file.registers[10][3] ;
 wire \soc_inst.cpu_core.register_file.registers[10][4] ;
 wire \soc_inst.cpu_core.register_file.registers[10][5] ;
 wire \soc_inst.cpu_core.register_file.registers[10][6] ;
 wire \soc_inst.cpu_core.register_file.registers[10][7] ;
 wire \soc_inst.cpu_core.register_file.registers[10][8] ;
 wire \soc_inst.cpu_core.register_file.registers[10][9] ;
 wire \soc_inst.cpu_core.register_file.registers[11][0] ;
 wire \soc_inst.cpu_core.register_file.registers[11][10] ;
 wire \soc_inst.cpu_core.register_file.registers[11][11] ;
 wire \soc_inst.cpu_core.register_file.registers[11][12] ;
 wire \soc_inst.cpu_core.register_file.registers[11][13] ;
 wire \soc_inst.cpu_core.register_file.registers[11][14] ;
 wire \soc_inst.cpu_core.register_file.registers[11][15] ;
 wire \soc_inst.cpu_core.register_file.registers[11][16] ;
 wire \soc_inst.cpu_core.register_file.registers[11][17] ;
 wire \soc_inst.cpu_core.register_file.registers[11][18] ;
 wire \soc_inst.cpu_core.register_file.registers[11][19] ;
 wire \soc_inst.cpu_core.register_file.registers[11][1] ;
 wire \soc_inst.cpu_core.register_file.registers[11][20] ;
 wire \soc_inst.cpu_core.register_file.registers[11][21] ;
 wire \soc_inst.cpu_core.register_file.registers[11][22] ;
 wire \soc_inst.cpu_core.register_file.registers[11][23] ;
 wire \soc_inst.cpu_core.register_file.registers[11][24] ;
 wire \soc_inst.cpu_core.register_file.registers[11][25] ;
 wire \soc_inst.cpu_core.register_file.registers[11][26] ;
 wire \soc_inst.cpu_core.register_file.registers[11][27] ;
 wire \soc_inst.cpu_core.register_file.registers[11][28] ;
 wire \soc_inst.cpu_core.register_file.registers[11][29] ;
 wire \soc_inst.cpu_core.register_file.registers[11][2] ;
 wire \soc_inst.cpu_core.register_file.registers[11][30] ;
 wire \soc_inst.cpu_core.register_file.registers[11][31] ;
 wire \soc_inst.cpu_core.register_file.registers[11][3] ;
 wire \soc_inst.cpu_core.register_file.registers[11][4] ;
 wire \soc_inst.cpu_core.register_file.registers[11][5] ;
 wire \soc_inst.cpu_core.register_file.registers[11][6] ;
 wire \soc_inst.cpu_core.register_file.registers[11][7] ;
 wire \soc_inst.cpu_core.register_file.registers[11][8] ;
 wire \soc_inst.cpu_core.register_file.registers[11][9] ;
 wire \soc_inst.cpu_core.register_file.registers[12][0] ;
 wire \soc_inst.cpu_core.register_file.registers[12][10] ;
 wire \soc_inst.cpu_core.register_file.registers[12][11] ;
 wire \soc_inst.cpu_core.register_file.registers[12][12] ;
 wire \soc_inst.cpu_core.register_file.registers[12][13] ;
 wire \soc_inst.cpu_core.register_file.registers[12][14] ;
 wire \soc_inst.cpu_core.register_file.registers[12][15] ;
 wire \soc_inst.cpu_core.register_file.registers[12][16] ;
 wire \soc_inst.cpu_core.register_file.registers[12][17] ;
 wire \soc_inst.cpu_core.register_file.registers[12][18] ;
 wire \soc_inst.cpu_core.register_file.registers[12][19] ;
 wire \soc_inst.cpu_core.register_file.registers[12][1] ;
 wire \soc_inst.cpu_core.register_file.registers[12][20] ;
 wire \soc_inst.cpu_core.register_file.registers[12][21] ;
 wire \soc_inst.cpu_core.register_file.registers[12][22] ;
 wire \soc_inst.cpu_core.register_file.registers[12][23] ;
 wire \soc_inst.cpu_core.register_file.registers[12][24] ;
 wire \soc_inst.cpu_core.register_file.registers[12][25] ;
 wire \soc_inst.cpu_core.register_file.registers[12][26] ;
 wire \soc_inst.cpu_core.register_file.registers[12][27] ;
 wire \soc_inst.cpu_core.register_file.registers[12][28] ;
 wire \soc_inst.cpu_core.register_file.registers[12][29] ;
 wire \soc_inst.cpu_core.register_file.registers[12][2] ;
 wire \soc_inst.cpu_core.register_file.registers[12][30] ;
 wire \soc_inst.cpu_core.register_file.registers[12][31] ;
 wire \soc_inst.cpu_core.register_file.registers[12][3] ;
 wire \soc_inst.cpu_core.register_file.registers[12][4] ;
 wire \soc_inst.cpu_core.register_file.registers[12][5] ;
 wire \soc_inst.cpu_core.register_file.registers[12][6] ;
 wire \soc_inst.cpu_core.register_file.registers[12][7] ;
 wire \soc_inst.cpu_core.register_file.registers[12][8] ;
 wire \soc_inst.cpu_core.register_file.registers[12][9] ;
 wire \soc_inst.cpu_core.register_file.registers[13][0] ;
 wire \soc_inst.cpu_core.register_file.registers[13][10] ;
 wire \soc_inst.cpu_core.register_file.registers[13][11] ;
 wire \soc_inst.cpu_core.register_file.registers[13][12] ;
 wire \soc_inst.cpu_core.register_file.registers[13][13] ;
 wire \soc_inst.cpu_core.register_file.registers[13][14] ;
 wire \soc_inst.cpu_core.register_file.registers[13][15] ;
 wire \soc_inst.cpu_core.register_file.registers[13][16] ;
 wire \soc_inst.cpu_core.register_file.registers[13][17] ;
 wire \soc_inst.cpu_core.register_file.registers[13][18] ;
 wire \soc_inst.cpu_core.register_file.registers[13][19] ;
 wire \soc_inst.cpu_core.register_file.registers[13][1] ;
 wire \soc_inst.cpu_core.register_file.registers[13][20] ;
 wire \soc_inst.cpu_core.register_file.registers[13][21] ;
 wire \soc_inst.cpu_core.register_file.registers[13][22] ;
 wire \soc_inst.cpu_core.register_file.registers[13][23] ;
 wire \soc_inst.cpu_core.register_file.registers[13][24] ;
 wire \soc_inst.cpu_core.register_file.registers[13][25] ;
 wire \soc_inst.cpu_core.register_file.registers[13][26] ;
 wire \soc_inst.cpu_core.register_file.registers[13][27] ;
 wire \soc_inst.cpu_core.register_file.registers[13][28] ;
 wire \soc_inst.cpu_core.register_file.registers[13][29] ;
 wire \soc_inst.cpu_core.register_file.registers[13][2] ;
 wire \soc_inst.cpu_core.register_file.registers[13][30] ;
 wire \soc_inst.cpu_core.register_file.registers[13][31] ;
 wire \soc_inst.cpu_core.register_file.registers[13][3] ;
 wire \soc_inst.cpu_core.register_file.registers[13][4] ;
 wire \soc_inst.cpu_core.register_file.registers[13][5] ;
 wire \soc_inst.cpu_core.register_file.registers[13][6] ;
 wire \soc_inst.cpu_core.register_file.registers[13][7] ;
 wire \soc_inst.cpu_core.register_file.registers[13][8] ;
 wire \soc_inst.cpu_core.register_file.registers[13][9] ;
 wire \soc_inst.cpu_core.register_file.registers[14][0] ;
 wire \soc_inst.cpu_core.register_file.registers[14][10] ;
 wire \soc_inst.cpu_core.register_file.registers[14][11] ;
 wire \soc_inst.cpu_core.register_file.registers[14][12] ;
 wire \soc_inst.cpu_core.register_file.registers[14][13] ;
 wire \soc_inst.cpu_core.register_file.registers[14][14] ;
 wire \soc_inst.cpu_core.register_file.registers[14][15] ;
 wire \soc_inst.cpu_core.register_file.registers[14][16] ;
 wire \soc_inst.cpu_core.register_file.registers[14][17] ;
 wire \soc_inst.cpu_core.register_file.registers[14][18] ;
 wire \soc_inst.cpu_core.register_file.registers[14][19] ;
 wire \soc_inst.cpu_core.register_file.registers[14][1] ;
 wire \soc_inst.cpu_core.register_file.registers[14][20] ;
 wire \soc_inst.cpu_core.register_file.registers[14][21] ;
 wire \soc_inst.cpu_core.register_file.registers[14][22] ;
 wire \soc_inst.cpu_core.register_file.registers[14][23] ;
 wire \soc_inst.cpu_core.register_file.registers[14][24] ;
 wire \soc_inst.cpu_core.register_file.registers[14][25] ;
 wire \soc_inst.cpu_core.register_file.registers[14][26] ;
 wire \soc_inst.cpu_core.register_file.registers[14][27] ;
 wire \soc_inst.cpu_core.register_file.registers[14][28] ;
 wire \soc_inst.cpu_core.register_file.registers[14][29] ;
 wire \soc_inst.cpu_core.register_file.registers[14][2] ;
 wire \soc_inst.cpu_core.register_file.registers[14][30] ;
 wire \soc_inst.cpu_core.register_file.registers[14][31] ;
 wire \soc_inst.cpu_core.register_file.registers[14][3] ;
 wire \soc_inst.cpu_core.register_file.registers[14][4] ;
 wire \soc_inst.cpu_core.register_file.registers[14][5] ;
 wire \soc_inst.cpu_core.register_file.registers[14][6] ;
 wire \soc_inst.cpu_core.register_file.registers[14][7] ;
 wire \soc_inst.cpu_core.register_file.registers[14][8] ;
 wire \soc_inst.cpu_core.register_file.registers[14][9] ;
 wire \soc_inst.cpu_core.register_file.registers[15][0] ;
 wire \soc_inst.cpu_core.register_file.registers[15][10] ;
 wire \soc_inst.cpu_core.register_file.registers[15][11] ;
 wire \soc_inst.cpu_core.register_file.registers[15][12] ;
 wire \soc_inst.cpu_core.register_file.registers[15][13] ;
 wire \soc_inst.cpu_core.register_file.registers[15][14] ;
 wire \soc_inst.cpu_core.register_file.registers[15][15] ;
 wire \soc_inst.cpu_core.register_file.registers[15][16] ;
 wire \soc_inst.cpu_core.register_file.registers[15][17] ;
 wire \soc_inst.cpu_core.register_file.registers[15][18] ;
 wire \soc_inst.cpu_core.register_file.registers[15][19] ;
 wire \soc_inst.cpu_core.register_file.registers[15][1] ;
 wire \soc_inst.cpu_core.register_file.registers[15][20] ;
 wire \soc_inst.cpu_core.register_file.registers[15][21] ;
 wire \soc_inst.cpu_core.register_file.registers[15][22] ;
 wire \soc_inst.cpu_core.register_file.registers[15][23] ;
 wire \soc_inst.cpu_core.register_file.registers[15][24] ;
 wire \soc_inst.cpu_core.register_file.registers[15][25] ;
 wire \soc_inst.cpu_core.register_file.registers[15][26] ;
 wire \soc_inst.cpu_core.register_file.registers[15][27] ;
 wire \soc_inst.cpu_core.register_file.registers[15][28] ;
 wire \soc_inst.cpu_core.register_file.registers[15][29] ;
 wire \soc_inst.cpu_core.register_file.registers[15][2] ;
 wire \soc_inst.cpu_core.register_file.registers[15][30] ;
 wire \soc_inst.cpu_core.register_file.registers[15][31] ;
 wire \soc_inst.cpu_core.register_file.registers[15][3] ;
 wire \soc_inst.cpu_core.register_file.registers[15][4] ;
 wire \soc_inst.cpu_core.register_file.registers[15][5] ;
 wire \soc_inst.cpu_core.register_file.registers[15][6] ;
 wire \soc_inst.cpu_core.register_file.registers[15][7] ;
 wire \soc_inst.cpu_core.register_file.registers[15][8] ;
 wire \soc_inst.cpu_core.register_file.registers[15][9] ;
 wire \soc_inst.cpu_core.register_file.registers[16][0] ;
 wire \soc_inst.cpu_core.register_file.registers[16][10] ;
 wire \soc_inst.cpu_core.register_file.registers[16][11] ;
 wire \soc_inst.cpu_core.register_file.registers[16][12] ;
 wire \soc_inst.cpu_core.register_file.registers[16][13] ;
 wire \soc_inst.cpu_core.register_file.registers[16][14] ;
 wire \soc_inst.cpu_core.register_file.registers[16][15] ;
 wire \soc_inst.cpu_core.register_file.registers[16][16] ;
 wire \soc_inst.cpu_core.register_file.registers[16][17] ;
 wire \soc_inst.cpu_core.register_file.registers[16][18] ;
 wire \soc_inst.cpu_core.register_file.registers[16][19] ;
 wire \soc_inst.cpu_core.register_file.registers[16][1] ;
 wire \soc_inst.cpu_core.register_file.registers[16][20] ;
 wire \soc_inst.cpu_core.register_file.registers[16][21] ;
 wire \soc_inst.cpu_core.register_file.registers[16][22] ;
 wire \soc_inst.cpu_core.register_file.registers[16][23] ;
 wire \soc_inst.cpu_core.register_file.registers[16][24] ;
 wire \soc_inst.cpu_core.register_file.registers[16][25] ;
 wire \soc_inst.cpu_core.register_file.registers[16][26] ;
 wire \soc_inst.cpu_core.register_file.registers[16][27] ;
 wire \soc_inst.cpu_core.register_file.registers[16][28] ;
 wire \soc_inst.cpu_core.register_file.registers[16][29] ;
 wire \soc_inst.cpu_core.register_file.registers[16][2] ;
 wire \soc_inst.cpu_core.register_file.registers[16][30] ;
 wire \soc_inst.cpu_core.register_file.registers[16][31] ;
 wire \soc_inst.cpu_core.register_file.registers[16][3] ;
 wire \soc_inst.cpu_core.register_file.registers[16][4] ;
 wire \soc_inst.cpu_core.register_file.registers[16][5] ;
 wire \soc_inst.cpu_core.register_file.registers[16][6] ;
 wire \soc_inst.cpu_core.register_file.registers[16][7] ;
 wire \soc_inst.cpu_core.register_file.registers[16][8] ;
 wire \soc_inst.cpu_core.register_file.registers[16][9] ;
 wire \soc_inst.cpu_core.register_file.registers[17][0] ;
 wire \soc_inst.cpu_core.register_file.registers[17][10] ;
 wire \soc_inst.cpu_core.register_file.registers[17][11] ;
 wire \soc_inst.cpu_core.register_file.registers[17][12] ;
 wire \soc_inst.cpu_core.register_file.registers[17][13] ;
 wire \soc_inst.cpu_core.register_file.registers[17][14] ;
 wire \soc_inst.cpu_core.register_file.registers[17][15] ;
 wire \soc_inst.cpu_core.register_file.registers[17][16] ;
 wire \soc_inst.cpu_core.register_file.registers[17][17] ;
 wire \soc_inst.cpu_core.register_file.registers[17][18] ;
 wire \soc_inst.cpu_core.register_file.registers[17][19] ;
 wire \soc_inst.cpu_core.register_file.registers[17][1] ;
 wire \soc_inst.cpu_core.register_file.registers[17][20] ;
 wire \soc_inst.cpu_core.register_file.registers[17][21] ;
 wire \soc_inst.cpu_core.register_file.registers[17][22] ;
 wire \soc_inst.cpu_core.register_file.registers[17][23] ;
 wire \soc_inst.cpu_core.register_file.registers[17][24] ;
 wire \soc_inst.cpu_core.register_file.registers[17][25] ;
 wire \soc_inst.cpu_core.register_file.registers[17][26] ;
 wire \soc_inst.cpu_core.register_file.registers[17][27] ;
 wire \soc_inst.cpu_core.register_file.registers[17][28] ;
 wire \soc_inst.cpu_core.register_file.registers[17][29] ;
 wire \soc_inst.cpu_core.register_file.registers[17][2] ;
 wire \soc_inst.cpu_core.register_file.registers[17][30] ;
 wire \soc_inst.cpu_core.register_file.registers[17][31] ;
 wire \soc_inst.cpu_core.register_file.registers[17][3] ;
 wire \soc_inst.cpu_core.register_file.registers[17][4] ;
 wire \soc_inst.cpu_core.register_file.registers[17][5] ;
 wire \soc_inst.cpu_core.register_file.registers[17][6] ;
 wire \soc_inst.cpu_core.register_file.registers[17][7] ;
 wire \soc_inst.cpu_core.register_file.registers[17][8] ;
 wire \soc_inst.cpu_core.register_file.registers[17][9] ;
 wire \soc_inst.cpu_core.register_file.registers[18][0] ;
 wire \soc_inst.cpu_core.register_file.registers[18][10] ;
 wire \soc_inst.cpu_core.register_file.registers[18][11] ;
 wire \soc_inst.cpu_core.register_file.registers[18][12] ;
 wire \soc_inst.cpu_core.register_file.registers[18][13] ;
 wire \soc_inst.cpu_core.register_file.registers[18][14] ;
 wire \soc_inst.cpu_core.register_file.registers[18][15] ;
 wire \soc_inst.cpu_core.register_file.registers[18][16] ;
 wire \soc_inst.cpu_core.register_file.registers[18][17] ;
 wire \soc_inst.cpu_core.register_file.registers[18][18] ;
 wire \soc_inst.cpu_core.register_file.registers[18][19] ;
 wire \soc_inst.cpu_core.register_file.registers[18][1] ;
 wire \soc_inst.cpu_core.register_file.registers[18][20] ;
 wire \soc_inst.cpu_core.register_file.registers[18][21] ;
 wire \soc_inst.cpu_core.register_file.registers[18][22] ;
 wire \soc_inst.cpu_core.register_file.registers[18][23] ;
 wire \soc_inst.cpu_core.register_file.registers[18][24] ;
 wire \soc_inst.cpu_core.register_file.registers[18][25] ;
 wire \soc_inst.cpu_core.register_file.registers[18][26] ;
 wire \soc_inst.cpu_core.register_file.registers[18][27] ;
 wire \soc_inst.cpu_core.register_file.registers[18][28] ;
 wire \soc_inst.cpu_core.register_file.registers[18][29] ;
 wire \soc_inst.cpu_core.register_file.registers[18][2] ;
 wire \soc_inst.cpu_core.register_file.registers[18][30] ;
 wire \soc_inst.cpu_core.register_file.registers[18][31] ;
 wire \soc_inst.cpu_core.register_file.registers[18][3] ;
 wire \soc_inst.cpu_core.register_file.registers[18][4] ;
 wire \soc_inst.cpu_core.register_file.registers[18][5] ;
 wire \soc_inst.cpu_core.register_file.registers[18][6] ;
 wire \soc_inst.cpu_core.register_file.registers[18][7] ;
 wire \soc_inst.cpu_core.register_file.registers[18][8] ;
 wire \soc_inst.cpu_core.register_file.registers[18][9] ;
 wire \soc_inst.cpu_core.register_file.registers[19][0] ;
 wire \soc_inst.cpu_core.register_file.registers[19][10] ;
 wire \soc_inst.cpu_core.register_file.registers[19][11] ;
 wire \soc_inst.cpu_core.register_file.registers[19][12] ;
 wire \soc_inst.cpu_core.register_file.registers[19][13] ;
 wire \soc_inst.cpu_core.register_file.registers[19][14] ;
 wire \soc_inst.cpu_core.register_file.registers[19][15] ;
 wire \soc_inst.cpu_core.register_file.registers[19][16] ;
 wire \soc_inst.cpu_core.register_file.registers[19][17] ;
 wire \soc_inst.cpu_core.register_file.registers[19][18] ;
 wire \soc_inst.cpu_core.register_file.registers[19][19] ;
 wire \soc_inst.cpu_core.register_file.registers[19][1] ;
 wire \soc_inst.cpu_core.register_file.registers[19][20] ;
 wire \soc_inst.cpu_core.register_file.registers[19][21] ;
 wire \soc_inst.cpu_core.register_file.registers[19][22] ;
 wire \soc_inst.cpu_core.register_file.registers[19][23] ;
 wire \soc_inst.cpu_core.register_file.registers[19][24] ;
 wire \soc_inst.cpu_core.register_file.registers[19][25] ;
 wire \soc_inst.cpu_core.register_file.registers[19][26] ;
 wire \soc_inst.cpu_core.register_file.registers[19][27] ;
 wire \soc_inst.cpu_core.register_file.registers[19][28] ;
 wire \soc_inst.cpu_core.register_file.registers[19][29] ;
 wire \soc_inst.cpu_core.register_file.registers[19][2] ;
 wire \soc_inst.cpu_core.register_file.registers[19][30] ;
 wire \soc_inst.cpu_core.register_file.registers[19][31] ;
 wire \soc_inst.cpu_core.register_file.registers[19][3] ;
 wire \soc_inst.cpu_core.register_file.registers[19][4] ;
 wire \soc_inst.cpu_core.register_file.registers[19][5] ;
 wire \soc_inst.cpu_core.register_file.registers[19][6] ;
 wire \soc_inst.cpu_core.register_file.registers[19][7] ;
 wire \soc_inst.cpu_core.register_file.registers[19][8] ;
 wire \soc_inst.cpu_core.register_file.registers[19][9] ;
 wire \soc_inst.cpu_core.register_file.registers[1][0] ;
 wire \soc_inst.cpu_core.register_file.registers[1][10] ;
 wire \soc_inst.cpu_core.register_file.registers[1][11] ;
 wire \soc_inst.cpu_core.register_file.registers[1][12] ;
 wire \soc_inst.cpu_core.register_file.registers[1][13] ;
 wire \soc_inst.cpu_core.register_file.registers[1][14] ;
 wire \soc_inst.cpu_core.register_file.registers[1][15] ;
 wire \soc_inst.cpu_core.register_file.registers[1][16] ;
 wire \soc_inst.cpu_core.register_file.registers[1][17] ;
 wire \soc_inst.cpu_core.register_file.registers[1][18] ;
 wire \soc_inst.cpu_core.register_file.registers[1][19] ;
 wire \soc_inst.cpu_core.register_file.registers[1][1] ;
 wire \soc_inst.cpu_core.register_file.registers[1][20] ;
 wire \soc_inst.cpu_core.register_file.registers[1][21] ;
 wire \soc_inst.cpu_core.register_file.registers[1][22] ;
 wire \soc_inst.cpu_core.register_file.registers[1][23] ;
 wire \soc_inst.cpu_core.register_file.registers[1][24] ;
 wire \soc_inst.cpu_core.register_file.registers[1][25] ;
 wire \soc_inst.cpu_core.register_file.registers[1][26] ;
 wire \soc_inst.cpu_core.register_file.registers[1][27] ;
 wire \soc_inst.cpu_core.register_file.registers[1][28] ;
 wire \soc_inst.cpu_core.register_file.registers[1][29] ;
 wire \soc_inst.cpu_core.register_file.registers[1][2] ;
 wire \soc_inst.cpu_core.register_file.registers[1][30] ;
 wire \soc_inst.cpu_core.register_file.registers[1][31] ;
 wire \soc_inst.cpu_core.register_file.registers[1][3] ;
 wire \soc_inst.cpu_core.register_file.registers[1][4] ;
 wire \soc_inst.cpu_core.register_file.registers[1][5] ;
 wire \soc_inst.cpu_core.register_file.registers[1][6] ;
 wire \soc_inst.cpu_core.register_file.registers[1][7] ;
 wire \soc_inst.cpu_core.register_file.registers[1][8] ;
 wire \soc_inst.cpu_core.register_file.registers[1][9] ;
 wire \soc_inst.cpu_core.register_file.registers[20][0] ;
 wire \soc_inst.cpu_core.register_file.registers[20][10] ;
 wire \soc_inst.cpu_core.register_file.registers[20][11] ;
 wire \soc_inst.cpu_core.register_file.registers[20][12] ;
 wire \soc_inst.cpu_core.register_file.registers[20][13] ;
 wire \soc_inst.cpu_core.register_file.registers[20][14] ;
 wire \soc_inst.cpu_core.register_file.registers[20][15] ;
 wire \soc_inst.cpu_core.register_file.registers[20][16] ;
 wire \soc_inst.cpu_core.register_file.registers[20][17] ;
 wire \soc_inst.cpu_core.register_file.registers[20][18] ;
 wire \soc_inst.cpu_core.register_file.registers[20][19] ;
 wire \soc_inst.cpu_core.register_file.registers[20][1] ;
 wire \soc_inst.cpu_core.register_file.registers[20][20] ;
 wire \soc_inst.cpu_core.register_file.registers[20][21] ;
 wire \soc_inst.cpu_core.register_file.registers[20][22] ;
 wire \soc_inst.cpu_core.register_file.registers[20][23] ;
 wire \soc_inst.cpu_core.register_file.registers[20][24] ;
 wire \soc_inst.cpu_core.register_file.registers[20][25] ;
 wire \soc_inst.cpu_core.register_file.registers[20][26] ;
 wire \soc_inst.cpu_core.register_file.registers[20][27] ;
 wire \soc_inst.cpu_core.register_file.registers[20][28] ;
 wire \soc_inst.cpu_core.register_file.registers[20][29] ;
 wire \soc_inst.cpu_core.register_file.registers[20][2] ;
 wire \soc_inst.cpu_core.register_file.registers[20][30] ;
 wire \soc_inst.cpu_core.register_file.registers[20][31] ;
 wire \soc_inst.cpu_core.register_file.registers[20][3] ;
 wire \soc_inst.cpu_core.register_file.registers[20][4] ;
 wire \soc_inst.cpu_core.register_file.registers[20][5] ;
 wire \soc_inst.cpu_core.register_file.registers[20][6] ;
 wire \soc_inst.cpu_core.register_file.registers[20][7] ;
 wire \soc_inst.cpu_core.register_file.registers[20][8] ;
 wire \soc_inst.cpu_core.register_file.registers[20][9] ;
 wire \soc_inst.cpu_core.register_file.registers[21][0] ;
 wire \soc_inst.cpu_core.register_file.registers[21][10] ;
 wire \soc_inst.cpu_core.register_file.registers[21][11] ;
 wire \soc_inst.cpu_core.register_file.registers[21][12] ;
 wire \soc_inst.cpu_core.register_file.registers[21][13] ;
 wire \soc_inst.cpu_core.register_file.registers[21][14] ;
 wire \soc_inst.cpu_core.register_file.registers[21][15] ;
 wire \soc_inst.cpu_core.register_file.registers[21][16] ;
 wire \soc_inst.cpu_core.register_file.registers[21][17] ;
 wire \soc_inst.cpu_core.register_file.registers[21][18] ;
 wire \soc_inst.cpu_core.register_file.registers[21][19] ;
 wire \soc_inst.cpu_core.register_file.registers[21][1] ;
 wire \soc_inst.cpu_core.register_file.registers[21][20] ;
 wire \soc_inst.cpu_core.register_file.registers[21][21] ;
 wire \soc_inst.cpu_core.register_file.registers[21][22] ;
 wire \soc_inst.cpu_core.register_file.registers[21][23] ;
 wire \soc_inst.cpu_core.register_file.registers[21][24] ;
 wire \soc_inst.cpu_core.register_file.registers[21][25] ;
 wire \soc_inst.cpu_core.register_file.registers[21][26] ;
 wire \soc_inst.cpu_core.register_file.registers[21][27] ;
 wire \soc_inst.cpu_core.register_file.registers[21][28] ;
 wire \soc_inst.cpu_core.register_file.registers[21][29] ;
 wire \soc_inst.cpu_core.register_file.registers[21][2] ;
 wire \soc_inst.cpu_core.register_file.registers[21][30] ;
 wire \soc_inst.cpu_core.register_file.registers[21][31] ;
 wire \soc_inst.cpu_core.register_file.registers[21][3] ;
 wire \soc_inst.cpu_core.register_file.registers[21][4] ;
 wire \soc_inst.cpu_core.register_file.registers[21][5] ;
 wire \soc_inst.cpu_core.register_file.registers[21][6] ;
 wire \soc_inst.cpu_core.register_file.registers[21][7] ;
 wire \soc_inst.cpu_core.register_file.registers[21][8] ;
 wire \soc_inst.cpu_core.register_file.registers[21][9] ;
 wire \soc_inst.cpu_core.register_file.registers[22][0] ;
 wire \soc_inst.cpu_core.register_file.registers[22][10] ;
 wire \soc_inst.cpu_core.register_file.registers[22][11] ;
 wire \soc_inst.cpu_core.register_file.registers[22][12] ;
 wire \soc_inst.cpu_core.register_file.registers[22][13] ;
 wire \soc_inst.cpu_core.register_file.registers[22][14] ;
 wire \soc_inst.cpu_core.register_file.registers[22][15] ;
 wire \soc_inst.cpu_core.register_file.registers[22][16] ;
 wire \soc_inst.cpu_core.register_file.registers[22][17] ;
 wire \soc_inst.cpu_core.register_file.registers[22][18] ;
 wire \soc_inst.cpu_core.register_file.registers[22][19] ;
 wire \soc_inst.cpu_core.register_file.registers[22][1] ;
 wire \soc_inst.cpu_core.register_file.registers[22][20] ;
 wire \soc_inst.cpu_core.register_file.registers[22][21] ;
 wire \soc_inst.cpu_core.register_file.registers[22][22] ;
 wire \soc_inst.cpu_core.register_file.registers[22][23] ;
 wire \soc_inst.cpu_core.register_file.registers[22][24] ;
 wire \soc_inst.cpu_core.register_file.registers[22][25] ;
 wire \soc_inst.cpu_core.register_file.registers[22][26] ;
 wire \soc_inst.cpu_core.register_file.registers[22][27] ;
 wire \soc_inst.cpu_core.register_file.registers[22][28] ;
 wire \soc_inst.cpu_core.register_file.registers[22][29] ;
 wire \soc_inst.cpu_core.register_file.registers[22][2] ;
 wire \soc_inst.cpu_core.register_file.registers[22][30] ;
 wire \soc_inst.cpu_core.register_file.registers[22][31] ;
 wire \soc_inst.cpu_core.register_file.registers[22][3] ;
 wire \soc_inst.cpu_core.register_file.registers[22][4] ;
 wire \soc_inst.cpu_core.register_file.registers[22][5] ;
 wire \soc_inst.cpu_core.register_file.registers[22][6] ;
 wire \soc_inst.cpu_core.register_file.registers[22][7] ;
 wire \soc_inst.cpu_core.register_file.registers[22][8] ;
 wire \soc_inst.cpu_core.register_file.registers[22][9] ;
 wire \soc_inst.cpu_core.register_file.registers[23][0] ;
 wire \soc_inst.cpu_core.register_file.registers[23][10] ;
 wire \soc_inst.cpu_core.register_file.registers[23][11] ;
 wire \soc_inst.cpu_core.register_file.registers[23][12] ;
 wire \soc_inst.cpu_core.register_file.registers[23][13] ;
 wire \soc_inst.cpu_core.register_file.registers[23][14] ;
 wire \soc_inst.cpu_core.register_file.registers[23][15] ;
 wire \soc_inst.cpu_core.register_file.registers[23][16] ;
 wire \soc_inst.cpu_core.register_file.registers[23][17] ;
 wire \soc_inst.cpu_core.register_file.registers[23][18] ;
 wire \soc_inst.cpu_core.register_file.registers[23][19] ;
 wire \soc_inst.cpu_core.register_file.registers[23][1] ;
 wire \soc_inst.cpu_core.register_file.registers[23][20] ;
 wire \soc_inst.cpu_core.register_file.registers[23][21] ;
 wire \soc_inst.cpu_core.register_file.registers[23][22] ;
 wire \soc_inst.cpu_core.register_file.registers[23][23] ;
 wire \soc_inst.cpu_core.register_file.registers[23][24] ;
 wire \soc_inst.cpu_core.register_file.registers[23][25] ;
 wire \soc_inst.cpu_core.register_file.registers[23][26] ;
 wire \soc_inst.cpu_core.register_file.registers[23][27] ;
 wire \soc_inst.cpu_core.register_file.registers[23][28] ;
 wire \soc_inst.cpu_core.register_file.registers[23][29] ;
 wire \soc_inst.cpu_core.register_file.registers[23][2] ;
 wire \soc_inst.cpu_core.register_file.registers[23][30] ;
 wire \soc_inst.cpu_core.register_file.registers[23][31] ;
 wire \soc_inst.cpu_core.register_file.registers[23][3] ;
 wire \soc_inst.cpu_core.register_file.registers[23][4] ;
 wire \soc_inst.cpu_core.register_file.registers[23][5] ;
 wire \soc_inst.cpu_core.register_file.registers[23][6] ;
 wire \soc_inst.cpu_core.register_file.registers[23][7] ;
 wire \soc_inst.cpu_core.register_file.registers[23][8] ;
 wire \soc_inst.cpu_core.register_file.registers[23][9] ;
 wire \soc_inst.cpu_core.register_file.registers[24][0] ;
 wire \soc_inst.cpu_core.register_file.registers[24][10] ;
 wire \soc_inst.cpu_core.register_file.registers[24][11] ;
 wire \soc_inst.cpu_core.register_file.registers[24][12] ;
 wire \soc_inst.cpu_core.register_file.registers[24][13] ;
 wire \soc_inst.cpu_core.register_file.registers[24][14] ;
 wire \soc_inst.cpu_core.register_file.registers[24][15] ;
 wire \soc_inst.cpu_core.register_file.registers[24][16] ;
 wire \soc_inst.cpu_core.register_file.registers[24][17] ;
 wire \soc_inst.cpu_core.register_file.registers[24][18] ;
 wire \soc_inst.cpu_core.register_file.registers[24][19] ;
 wire \soc_inst.cpu_core.register_file.registers[24][1] ;
 wire \soc_inst.cpu_core.register_file.registers[24][20] ;
 wire \soc_inst.cpu_core.register_file.registers[24][21] ;
 wire \soc_inst.cpu_core.register_file.registers[24][22] ;
 wire \soc_inst.cpu_core.register_file.registers[24][23] ;
 wire \soc_inst.cpu_core.register_file.registers[24][24] ;
 wire \soc_inst.cpu_core.register_file.registers[24][25] ;
 wire \soc_inst.cpu_core.register_file.registers[24][26] ;
 wire \soc_inst.cpu_core.register_file.registers[24][27] ;
 wire \soc_inst.cpu_core.register_file.registers[24][28] ;
 wire \soc_inst.cpu_core.register_file.registers[24][29] ;
 wire \soc_inst.cpu_core.register_file.registers[24][2] ;
 wire \soc_inst.cpu_core.register_file.registers[24][30] ;
 wire \soc_inst.cpu_core.register_file.registers[24][31] ;
 wire \soc_inst.cpu_core.register_file.registers[24][3] ;
 wire \soc_inst.cpu_core.register_file.registers[24][4] ;
 wire \soc_inst.cpu_core.register_file.registers[24][5] ;
 wire \soc_inst.cpu_core.register_file.registers[24][6] ;
 wire \soc_inst.cpu_core.register_file.registers[24][7] ;
 wire \soc_inst.cpu_core.register_file.registers[24][8] ;
 wire \soc_inst.cpu_core.register_file.registers[24][9] ;
 wire \soc_inst.cpu_core.register_file.registers[25][0] ;
 wire \soc_inst.cpu_core.register_file.registers[25][10] ;
 wire \soc_inst.cpu_core.register_file.registers[25][11] ;
 wire \soc_inst.cpu_core.register_file.registers[25][12] ;
 wire \soc_inst.cpu_core.register_file.registers[25][13] ;
 wire \soc_inst.cpu_core.register_file.registers[25][14] ;
 wire \soc_inst.cpu_core.register_file.registers[25][15] ;
 wire \soc_inst.cpu_core.register_file.registers[25][16] ;
 wire \soc_inst.cpu_core.register_file.registers[25][17] ;
 wire \soc_inst.cpu_core.register_file.registers[25][18] ;
 wire \soc_inst.cpu_core.register_file.registers[25][19] ;
 wire \soc_inst.cpu_core.register_file.registers[25][1] ;
 wire \soc_inst.cpu_core.register_file.registers[25][20] ;
 wire \soc_inst.cpu_core.register_file.registers[25][21] ;
 wire \soc_inst.cpu_core.register_file.registers[25][22] ;
 wire \soc_inst.cpu_core.register_file.registers[25][23] ;
 wire \soc_inst.cpu_core.register_file.registers[25][24] ;
 wire \soc_inst.cpu_core.register_file.registers[25][25] ;
 wire \soc_inst.cpu_core.register_file.registers[25][26] ;
 wire \soc_inst.cpu_core.register_file.registers[25][27] ;
 wire \soc_inst.cpu_core.register_file.registers[25][28] ;
 wire \soc_inst.cpu_core.register_file.registers[25][29] ;
 wire \soc_inst.cpu_core.register_file.registers[25][2] ;
 wire \soc_inst.cpu_core.register_file.registers[25][30] ;
 wire \soc_inst.cpu_core.register_file.registers[25][31] ;
 wire \soc_inst.cpu_core.register_file.registers[25][3] ;
 wire \soc_inst.cpu_core.register_file.registers[25][4] ;
 wire \soc_inst.cpu_core.register_file.registers[25][5] ;
 wire \soc_inst.cpu_core.register_file.registers[25][6] ;
 wire \soc_inst.cpu_core.register_file.registers[25][7] ;
 wire \soc_inst.cpu_core.register_file.registers[25][8] ;
 wire \soc_inst.cpu_core.register_file.registers[25][9] ;
 wire \soc_inst.cpu_core.register_file.registers[26][0] ;
 wire \soc_inst.cpu_core.register_file.registers[26][10] ;
 wire \soc_inst.cpu_core.register_file.registers[26][11] ;
 wire \soc_inst.cpu_core.register_file.registers[26][12] ;
 wire \soc_inst.cpu_core.register_file.registers[26][13] ;
 wire \soc_inst.cpu_core.register_file.registers[26][14] ;
 wire \soc_inst.cpu_core.register_file.registers[26][15] ;
 wire \soc_inst.cpu_core.register_file.registers[26][16] ;
 wire \soc_inst.cpu_core.register_file.registers[26][17] ;
 wire \soc_inst.cpu_core.register_file.registers[26][18] ;
 wire \soc_inst.cpu_core.register_file.registers[26][19] ;
 wire \soc_inst.cpu_core.register_file.registers[26][1] ;
 wire \soc_inst.cpu_core.register_file.registers[26][20] ;
 wire \soc_inst.cpu_core.register_file.registers[26][21] ;
 wire \soc_inst.cpu_core.register_file.registers[26][22] ;
 wire \soc_inst.cpu_core.register_file.registers[26][23] ;
 wire \soc_inst.cpu_core.register_file.registers[26][24] ;
 wire \soc_inst.cpu_core.register_file.registers[26][25] ;
 wire \soc_inst.cpu_core.register_file.registers[26][26] ;
 wire \soc_inst.cpu_core.register_file.registers[26][27] ;
 wire \soc_inst.cpu_core.register_file.registers[26][28] ;
 wire \soc_inst.cpu_core.register_file.registers[26][29] ;
 wire \soc_inst.cpu_core.register_file.registers[26][2] ;
 wire \soc_inst.cpu_core.register_file.registers[26][30] ;
 wire \soc_inst.cpu_core.register_file.registers[26][31] ;
 wire \soc_inst.cpu_core.register_file.registers[26][3] ;
 wire \soc_inst.cpu_core.register_file.registers[26][4] ;
 wire \soc_inst.cpu_core.register_file.registers[26][5] ;
 wire \soc_inst.cpu_core.register_file.registers[26][6] ;
 wire \soc_inst.cpu_core.register_file.registers[26][7] ;
 wire \soc_inst.cpu_core.register_file.registers[26][8] ;
 wire \soc_inst.cpu_core.register_file.registers[26][9] ;
 wire \soc_inst.cpu_core.register_file.registers[27][0] ;
 wire \soc_inst.cpu_core.register_file.registers[27][10] ;
 wire \soc_inst.cpu_core.register_file.registers[27][11] ;
 wire \soc_inst.cpu_core.register_file.registers[27][12] ;
 wire \soc_inst.cpu_core.register_file.registers[27][13] ;
 wire \soc_inst.cpu_core.register_file.registers[27][14] ;
 wire \soc_inst.cpu_core.register_file.registers[27][15] ;
 wire \soc_inst.cpu_core.register_file.registers[27][16] ;
 wire \soc_inst.cpu_core.register_file.registers[27][17] ;
 wire \soc_inst.cpu_core.register_file.registers[27][18] ;
 wire \soc_inst.cpu_core.register_file.registers[27][19] ;
 wire \soc_inst.cpu_core.register_file.registers[27][1] ;
 wire \soc_inst.cpu_core.register_file.registers[27][20] ;
 wire \soc_inst.cpu_core.register_file.registers[27][21] ;
 wire \soc_inst.cpu_core.register_file.registers[27][22] ;
 wire \soc_inst.cpu_core.register_file.registers[27][23] ;
 wire \soc_inst.cpu_core.register_file.registers[27][24] ;
 wire \soc_inst.cpu_core.register_file.registers[27][25] ;
 wire \soc_inst.cpu_core.register_file.registers[27][26] ;
 wire \soc_inst.cpu_core.register_file.registers[27][27] ;
 wire \soc_inst.cpu_core.register_file.registers[27][28] ;
 wire \soc_inst.cpu_core.register_file.registers[27][29] ;
 wire \soc_inst.cpu_core.register_file.registers[27][2] ;
 wire \soc_inst.cpu_core.register_file.registers[27][30] ;
 wire \soc_inst.cpu_core.register_file.registers[27][31] ;
 wire \soc_inst.cpu_core.register_file.registers[27][3] ;
 wire \soc_inst.cpu_core.register_file.registers[27][4] ;
 wire \soc_inst.cpu_core.register_file.registers[27][5] ;
 wire \soc_inst.cpu_core.register_file.registers[27][6] ;
 wire \soc_inst.cpu_core.register_file.registers[27][7] ;
 wire \soc_inst.cpu_core.register_file.registers[27][8] ;
 wire \soc_inst.cpu_core.register_file.registers[27][9] ;
 wire \soc_inst.cpu_core.register_file.registers[28][0] ;
 wire \soc_inst.cpu_core.register_file.registers[28][10] ;
 wire \soc_inst.cpu_core.register_file.registers[28][11] ;
 wire \soc_inst.cpu_core.register_file.registers[28][12] ;
 wire \soc_inst.cpu_core.register_file.registers[28][13] ;
 wire \soc_inst.cpu_core.register_file.registers[28][14] ;
 wire \soc_inst.cpu_core.register_file.registers[28][15] ;
 wire \soc_inst.cpu_core.register_file.registers[28][16] ;
 wire \soc_inst.cpu_core.register_file.registers[28][17] ;
 wire \soc_inst.cpu_core.register_file.registers[28][18] ;
 wire \soc_inst.cpu_core.register_file.registers[28][19] ;
 wire \soc_inst.cpu_core.register_file.registers[28][1] ;
 wire \soc_inst.cpu_core.register_file.registers[28][20] ;
 wire \soc_inst.cpu_core.register_file.registers[28][21] ;
 wire \soc_inst.cpu_core.register_file.registers[28][22] ;
 wire \soc_inst.cpu_core.register_file.registers[28][23] ;
 wire \soc_inst.cpu_core.register_file.registers[28][24] ;
 wire \soc_inst.cpu_core.register_file.registers[28][25] ;
 wire \soc_inst.cpu_core.register_file.registers[28][26] ;
 wire \soc_inst.cpu_core.register_file.registers[28][27] ;
 wire \soc_inst.cpu_core.register_file.registers[28][28] ;
 wire \soc_inst.cpu_core.register_file.registers[28][29] ;
 wire \soc_inst.cpu_core.register_file.registers[28][2] ;
 wire \soc_inst.cpu_core.register_file.registers[28][30] ;
 wire \soc_inst.cpu_core.register_file.registers[28][31] ;
 wire \soc_inst.cpu_core.register_file.registers[28][3] ;
 wire \soc_inst.cpu_core.register_file.registers[28][4] ;
 wire \soc_inst.cpu_core.register_file.registers[28][5] ;
 wire \soc_inst.cpu_core.register_file.registers[28][6] ;
 wire \soc_inst.cpu_core.register_file.registers[28][7] ;
 wire \soc_inst.cpu_core.register_file.registers[28][8] ;
 wire \soc_inst.cpu_core.register_file.registers[28][9] ;
 wire \soc_inst.cpu_core.register_file.registers[29][0] ;
 wire \soc_inst.cpu_core.register_file.registers[29][10] ;
 wire \soc_inst.cpu_core.register_file.registers[29][11] ;
 wire \soc_inst.cpu_core.register_file.registers[29][12] ;
 wire \soc_inst.cpu_core.register_file.registers[29][13] ;
 wire \soc_inst.cpu_core.register_file.registers[29][14] ;
 wire \soc_inst.cpu_core.register_file.registers[29][15] ;
 wire \soc_inst.cpu_core.register_file.registers[29][16] ;
 wire \soc_inst.cpu_core.register_file.registers[29][17] ;
 wire \soc_inst.cpu_core.register_file.registers[29][18] ;
 wire \soc_inst.cpu_core.register_file.registers[29][19] ;
 wire \soc_inst.cpu_core.register_file.registers[29][1] ;
 wire \soc_inst.cpu_core.register_file.registers[29][20] ;
 wire \soc_inst.cpu_core.register_file.registers[29][21] ;
 wire \soc_inst.cpu_core.register_file.registers[29][22] ;
 wire \soc_inst.cpu_core.register_file.registers[29][23] ;
 wire \soc_inst.cpu_core.register_file.registers[29][24] ;
 wire \soc_inst.cpu_core.register_file.registers[29][25] ;
 wire \soc_inst.cpu_core.register_file.registers[29][26] ;
 wire \soc_inst.cpu_core.register_file.registers[29][27] ;
 wire \soc_inst.cpu_core.register_file.registers[29][28] ;
 wire \soc_inst.cpu_core.register_file.registers[29][29] ;
 wire \soc_inst.cpu_core.register_file.registers[29][2] ;
 wire \soc_inst.cpu_core.register_file.registers[29][30] ;
 wire \soc_inst.cpu_core.register_file.registers[29][31] ;
 wire \soc_inst.cpu_core.register_file.registers[29][3] ;
 wire \soc_inst.cpu_core.register_file.registers[29][4] ;
 wire \soc_inst.cpu_core.register_file.registers[29][5] ;
 wire \soc_inst.cpu_core.register_file.registers[29][6] ;
 wire \soc_inst.cpu_core.register_file.registers[29][7] ;
 wire \soc_inst.cpu_core.register_file.registers[29][8] ;
 wire \soc_inst.cpu_core.register_file.registers[29][9] ;
 wire \soc_inst.cpu_core.register_file.registers[2][0] ;
 wire \soc_inst.cpu_core.register_file.registers[2][10] ;
 wire \soc_inst.cpu_core.register_file.registers[2][11] ;
 wire \soc_inst.cpu_core.register_file.registers[2][12] ;
 wire \soc_inst.cpu_core.register_file.registers[2][13] ;
 wire \soc_inst.cpu_core.register_file.registers[2][14] ;
 wire \soc_inst.cpu_core.register_file.registers[2][15] ;
 wire \soc_inst.cpu_core.register_file.registers[2][16] ;
 wire \soc_inst.cpu_core.register_file.registers[2][17] ;
 wire \soc_inst.cpu_core.register_file.registers[2][18] ;
 wire \soc_inst.cpu_core.register_file.registers[2][19] ;
 wire \soc_inst.cpu_core.register_file.registers[2][1] ;
 wire \soc_inst.cpu_core.register_file.registers[2][20] ;
 wire \soc_inst.cpu_core.register_file.registers[2][21] ;
 wire \soc_inst.cpu_core.register_file.registers[2][22] ;
 wire \soc_inst.cpu_core.register_file.registers[2][23] ;
 wire \soc_inst.cpu_core.register_file.registers[2][24] ;
 wire \soc_inst.cpu_core.register_file.registers[2][25] ;
 wire \soc_inst.cpu_core.register_file.registers[2][26] ;
 wire \soc_inst.cpu_core.register_file.registers[2][27] ;
 wire \soc_inst.cpu_core.register_file.registers[2][28] ;
 wire \soc_inst.cpu_core.register_file.registers[2][29] ;
 wire \soc_inst.cpu_core.register_file.registers[2][2] ;
 wire \soc_inst.cpu_core.register_file.registers[2][30] ;
 wire \soc_inst.cpu_core.register_file.registers[2][31] ;
 wire \soc_inst.cpu_core.register_file.registers[2][3] ;
 wire \soc_inst.cpu_core.register_file.registers[2][4] ;
 wire \soc_inst.cpu_core.register_file.registers[2][5] ;
 wire \soc_inst.cpu_core.register_file.registers[2][6] ;
 wire \soc_inst.cpu_core.register_file.registers[2][7] ;
 wire \soc_inst.cpu_core.register_file.registers[2][8] ;
 wire \soc_inst.cpu_core.register_file.registers[2][9] ;
 wire \soc_inst.cpu_core.register_file.registers[30][0] ;
 wire \soc_inst.cpu_core.register_file.registers[30][10] ;
 wire \soc_inst.cpu_core.register_file.registers[30][11] ;
 wire \soc_inst.cpu_core.register_file.registers[30][12] ;
 wire \soc_inst.cpu_core.register_file.registers[30][13] ;
 wire \soc_inst.cpu_core.register_file.registers[30][14] ;
 wire \soc_inst.cpu_core.register_file.registers[30][15] ;
 wire \soc_inst.cpu_core.register_file.registers[30][16] ;
 wire \soc_inst.cpu_core.register_file.registers[30][17] ;
 wire \soc_inst.cpu_core.register_file.registers[30][18] ;
 wire \soc_inst.cpu_core.register_file.registers[30][19] ;
 wire \soc_inst.cpu_core.register_file.registers[30][1] ;
 wire \soc_inst.cpu_core.register_file.registers[30][20] ;
 wire \soc_inst.cpu_core.register_file.registers[30][21] ;
 wire \soc_inst.cpu_core.register_file.registers[30][22] ;
 wire \soc_inst.cpu_core.register_file.registers[30][23] ;
 wire \soc_inst.cpu_core.register_file.registers[30][24] ;
 wire \soc_inst.cpu_core.register_file.registers[30][25] ;
 wire \soc_inst.cpu_core.register_file.registers[30][26] ;
 wire \soc_inst.cpu_core.register_file.registers[30][27] ;
 wire \soc_inst.cpu_core.register_file.registers[30][28] ;
 wire \soc_inst.cpu_core.register_file.registers[30][29] ;
 wire \soc_inst.cpu_core.register_file.registers[30][2] ;
 wire \soc_inst.cpu_core.register_file.registers[30][30] ;
 wire \soc_inst.cpu_core.register_file.registers[30][31] ;
 wire \soc_inst.cpu_core.register_file.registers[30][3] ;
 wire \soc_inst.cpu_core.register_file.registers[30][4] ;
 wire \soc_inst.cpu_core.register_file.registers[30][5] ;
 wire \soc_inst.cpu_core.register_file.registers[30][6] ;
 wire \soc_inst.cpu_core.register_file.registers[30][7] ;
 wire \soc_inst.cpu_core.register_file.registers[30][8] ;
 wire \soc_inst.cpu_core.register_file.registers[30][9] ;
 wire \soc_inst.cpu_core.register_file.registers[31][0] ;
 wire \soc_inst.cpu_core.register_file.registers[31][10] ;
 wire \soc_inst.cpu_core.register_file.registers[31][11] ;
 wire \soc_inst.cpu_core.register_file.registers[31][12] ;
 wire \soc_inst.cpu_core.register_file.registers[31][13] ;
 wire \soc_inst.cpu_core.register_file.registers[31][14] ;
 wire \soc_inst.cpu_core.register_file.registers[31][15] ;
 wire \soc_inst.cpu_core.register_file.registers[31][16] ;
 wire \soc_inst.cpu_core.register_file.registers[31][17] ;
 wire \soc_inst.cpu_core.register_file.registers[31][18] ;
 wire \soc_inst.cpu_core.register_file.registers[31][19] ;
 wire \soc_inst.cpu_core.register_file.registers[31][1] ;
 wire \soc_inst.cpu_core.register_file.registers[31][20] ;
 wire \soc_inst.cpu_core.register_file.registers[31][21] ;
 wire \soc_inst.cpu_core.register_file.registers[31][22] ;
 wire \soc_inst.cpu_core.register_file.registers[31][23] ;
 wire \soc_inst.cpu_core.register_file.registers[31][24] ;
 wire \soc_inst.cpu_core.register_file.registers[31][25] ;
 wire \soc_inst.cpu_core.register_file.registers[31][26] ;
 wire \soc_inst.cpu_core.register_file.registers[31][27] ;
 wire \soc_inst.cpu_core.register_file.registers[31][28] ;
 wire \soc_inst.cpu_core.register_file.registers[31][29] ;
 wire \soc_inst.cpu_core.register_file.registers[31][2] ;
 wire \soc_inst.cpu_core.register_file.registers[31][30] ;
 wire \soc_inst.cpu_core.register_file.registers[31][31] ;
 wire \soc_inst.cpu_core.register_file.registers[31][3] ;
 wire \soc_inst.cpu_core.register_file.registers[31][4] ;
 wire \soc_inst.cpu_core.register_file.registers[31][5] ;
 wire \soc_inst.cpu_core.register_file.registers[31][6] ;
 wire \soc_inst.cpu_core.register_file.registers[31][7] ;
 wire \soc_inst.cpu_core.register_file.registers[31][8] ;
 wire \soc_inst.cpu_core.register_file.registers[31][9] ;
 wire \soc_inst.cpu_core.register_file.registers[3][0] ;
 wire \soc_inst.cpu_core.register_file.registers[3][10] ;
 wire \soc_inst.cpu_core.register_file.registers[3][11] ;
 wire \soc_inst.cpu_core.register_file.registers[3][12] ;
 wire \soc_inst.cpu_core.register_file.registers[3][13] ;
 wire \soc_inst.cpu_core.register_file.registers[3][14] ;
 wire \soc_inst.cpu_core.register_file.registers[3][15] ;
 wire \soc_inst.cpu_core.register_file.registers[3][16] ;
 wire \soc_inst.cpu_core.register_file.registers[3][17] ;
 wire \soc_inst.cpu_core.register_file.registers[3][18] ;
 wire \soc_inst.cpu_core.register_file.registers[3][19] ;
 wire \soc_inst.cpu_core.register_file.registers[3][1] ;
 wire \soc_inst.cpu_core.register_file.registers[3][20] ;
 wire \soc_inst.cpu_core.register_file.registers[3][21] ;
 wire \soc_inst.cpu_core.register_file.registers[3][22] ;
 wire \soc_inst.cpu_core.register_file.registers[3][23] ;
 wire \soc_inst.cpu_core.register_file.registers[3][24] ;
 wire \soc_inst.cpu_core.register_file.registers[3][25] ;
 wire \soc_inst.cpu_core.register_file.registers[3][26] ;
 wire \soc_inst.cpu_core.register_file.registers[3][27] ;
 wire \soc_inst.cpu_core.register_file.registers[3][28] ;
 wire \soc_inst.cpu_core.register_file.registers[3][29] ;
 wire \soc_inst.cpu_core.register_file.registers[3][2] ;
 wire \soc_inst.cpu_core.register_file.registers[3][30] ;
 wire \soc_inst.cpu_core.register_file.registers[3][31] ;
 wire \soc_inst.cpu_core.register_file.registers[3][3] ;
 wire \soc_inst.cpu_core.register_file.registers[3][4] ;
 wire \soc_inst.cpu_core.register_file.registers[3][5] ;
 wire \soc_inst.cpu_core.register_file.registers[3][6] ;
 wire \soc_inst.cpu_core.register_file.registers[3][7] ;
 wire \soc_inst.cpu_core.register_file.registers[3][8] ;
 wire \soc_inst.cpu_core.register_file.registers[3][9] ;
 wire \soc_inst.cpu_core.register_file.registers[4][0] ;
 wire \soc_inst.cpu_core.register_file.registers[4][10] ;
 wire \soc_inst.cpu_core.register_file.registers[4][11] ;
 wire \soc_inst.cpu_core.register_file.registers[4][12] ;
 wire \soc_inst.cpu_core.register_file.registers[4][13] ;
 wire \soc_inst.cpu_core.register_file.registers[4][14] ;
 wire \soc_inst.cpu_core.register_file.registers[4][15] ;
 wire \soc_inst.cpu_core.register_file.registers[4][16] ;
 wire \soc_inst.cpu_core.register_file.registers[4][17] ;
 wire \soc_inst.cpu_core.register_file.registers[4][18] ;
 wire \soc_inst.cpu_core.register_file.registers[4][19] ;
 wire \soc_inst.cpu_core.register_file.registers[4][1] ;
 wire \soc_inst.cpu_core.register_file.registers[4][20] ;
 wire \soc_inst.cpu_core.register_file.registers[4][21] ;
 wire \soc_inst.cpu_core.register_file.registers[4][22] ;
 wire \soc_inst.cpu_core.register_file.registers[4][23] ;
 wire \soc_inst.cpu_core.register_file.registers[4][24] ;
 wire \soc_inst.cpu_core.register_file.registers[4][25] ;
 wire \soc_inst.cpu_core.register_file.registers[4][26] ;
 wire \soc_inst.cpu_core.register_file.registers[4][27] ;
 wire \soc_inst.cpu_core.register_file.registers[4][28] ;
 wire \soc_inst.cpu_core.register_file.registers[4][29] ;
 wire \soc_inst.cpu_core.register_file.registers[4][2] ;
 wire \soc_inst.cpu_core.register_file.registers[4][30] ;
 wire \soc_inst.cpu_core.register_file.registers[4][31] ;
 wire \soc_inst.cpu_core.register_file.registers[4][3] ;
 wire \soc_inst.cpu_core.register_file.registers[4][4] ;
 wire \soc_inst.cpu_core.register_file.registers[4][5] ;
 wire \soc_inst.cpu_core.register_file.registers[4][6] ;
 wire \soc_inst.cpu_core.register_file.registers[4][7] ;
 wire \soc_inst.cpu_core.register_file.registers[4][8] ;
 wire \soc_inst.cpu_core.register_file.registers[4][9] ;
 wire \soc_inst.cpu_core.register_file.registers[5][0] ;
 wire \soc_inst.cpu_core.register_file.registers[5][10] ;
 wire \soc_inst.cpu_core.register_file.registers[5][11] ;
 wire \soc_inst.cpu_core.register_file.registers[5][12] ;
 wire \soc_inst.cpu_core.register_file.registers[5][13] ;
 wire \soc_inst.cpu_core.register_file.registers[5][14] ;
 wire \soc_inst.cpu_core.register_file.registers[5][15] ;
 wire \soc_inst.cpu_core.register_file.registers[5][16] ;
 wire \soc_inst.cpu_core.register_file.registers[5][17] ;
 wire \soc_inst.cpu_core.register_file.registers[5][18] ;
 wire \soc_inst.cpu_core.register_file.registers[5][19] ;
 wire \soc_inst.cpu_core.register_file.registers[5][1] ;
 wire \soc_inst.cpu_core.register_file.registers[5][20] ;
 wire \soc_inst.cpu_core.register_file.registers[5][21] ;
 wire \soc_inst.cpu_core.register_file.registers[5][22] ;
 wire \soc_inst.cpu_core.register_file.registers[5][23] ;
 wire \soc_inst.cpu_core.register_file.registers[5][24] ;
 wire \soc_inst.cpu_core.register_file.registers[5][25] ;
 wire \soc_inst.cpu_core.register_file.registers[5][26] ;
 wire \soc_inst.cpu_core.register_file.registers[5][27] ;
 wire \soc_inst.cpu_core.register_file.registers[5][28] ;
 wire \soc_inst.cpu_core.register_file.registers[5][29] ;
 wire \soc_inst.cpu_core.register_file.registers[5][2] ;
 wire \soc_inst.cpu_core.register_file.registers[5][30] ;
 wire \soc_inst.cpu_core.register_file.registers[5][31] ;
 wire \soc_inst.cpu_core.register_file.registers[5][3] ;
 wire \soc_inst.cpu_core.register_file.registers[5][4] ;
 wire \soc_inst.cpu_core.register_file.registers[5][5] ;
 wire \soc_inst.cpu_core.register_file.registers[5][6] ;
 wire \soc_inst.cpu_core.register_file.registers[5][7] ;
 wire \soc_inst.cpu_core.register_file.registers[5][8] ;
 wire \soc_inst.cpu_core.register_file.registers[5][9] ;
 wire \soc_inst.cpu_core.register_file.registers[6][0] ;
 wire \soc_inst.cpu_core.register_file.registers[6][10] ;
 wire \soc_inst.cpu_core.register_file.registers[6][11] ;
 wire \soc_inst.cpu_core.register_file.registers[6][12] ;
 wire \soc_inst.cpu_core.register_file.registers[6][13] ;
 wire \soc_inst.cpu_core.register_file.registers[6][14] ;
 wire \soc_inst.cpu_core.register_file.registers[6][15] ;
 wire \soc_inst.cpu_core.register_file.registers[6][16] ;
 wire \soc_inst.cpu_core.register_file.registers[6][17] ;
 wire \soc_inst.cpu_core.register_file.registers[6][18] ;
 wire \soc_inst.cpu_core.register_file.registers[6][19] ;
 wire \soc_inst.cpu_core.register_file.registers[6][1] ;
 wire \soc_inst.cpu_core.register_file.registers[6][20] ;
 wire \soc_inst.cpu_core.register_file.registers[6][21] ;
 wire \soc_inst.cpu_core.register_file.registers[6][22] ;
 wire \soc_inst.cpu_core.register_file.registers[6][23] ;
 wire \soc_inst.cpu_core.register_file.registers[6][24] ;
 wire \soc_inst.cpu_core.register_file.registers[6][25] ;
 wire \soc_inst.cpu_core.register_file.registers[6][26] ;
 wire \soc_inst.cpu_core.register_file.registers[6][27] ;
 wire \soc_inst.cpu_core.register_file.registers[6][28] ;
 wire \soc_inst.cpu_core.register_file.registers[6][29] ;
 wire \soc_inst.cpu_core.register_file.registers[6][2] ;
 wire \soc_inst.cpu_core.register_file.registers[6][30] ;
 wire \soc_inst.cpu_core.register_file.registers[6][31] ;
 wire \soc_inst.cpu_core.register_file.registers[6][3] ;
 wire \soc_inst.cpu_core.register_file.registers[6][4] ;
 wire \soc_inst.cpu_core.register_file.registers[6][5] ;
 wire \soc_inst.cpu_core.register_file.registers[6][6] ;
 wire \soc_inst.cpu_core.register_file.registers[6][7] ;
 wire \soc_inst.cpu_core.register_file.registers[6][8] ;
 wire \soc_inst.cpu_core.register_file.registers[6][9] ;
 wire \soc_inst.cpu_core.register_file.registers[7][0] ;
 wire \soc_inst.cpu_core.register_file.registers[7][10] ;
 wire \soc_inst.cpu_core.register_file.registers[7][11] ;
 wire \soc_inst.cpu_core.register_file.registers[7][12] ;
 wire \soc_inst.cpu_core.register_file.registers[7][13] ;
 wire \soc_inst.cpu_core.register_file.registers[7][14] ;
 wire \soc_inst.cpu_core.register_file.registers[7][15] ;
 wire \soc_inst.cpu_core.register_file.registers[7][16] ;
 wire \soc_inst.cpu_core.register_file.registers[7][17] ;
 wire \soc_inst.cpu_core.register_file.registers[7][18] ;
 wire \soc_inst.cpu_core.register_file.registers[7][19] ;
 wire \soc_inst.cpu_core.register_file.registers[7][1] ;
 wire \soc_inst.cpu_core.register_file.registers[7][20] ;
 wire \soc_inst.cpu_core.register_file.registers[7][21] ;
 wire \soc_inst.cpu_core.register_file.registers[7][22] ;
 wire \soc_inst.cpu_core.register_file.registers[7][23] ;
 wire \soc_inst.cpu_core.register_file.registers[7][24] ;
 wire \soc_inst.cpu_core.register_file.registers[7][25] ;
 wire \soc_inst.cpu_core.register_file.registers[7][26] ;
 wire \soc_inst.cpu_core.register_file.registers[7][27] ;
 wire \soc_inst.cpu_core.register_file.registers[7][28] ;
 wire \soc_inst.cpu_core.register_file.registers[7][29] ;
 wire \soc_inst.cpu_core.register_file.registers[7][2] ;
 wire \soc_inst.cpu_core.register_file.registers[7][30] ;
 wire \soc_inst.cpu_core.register_file.registers[7][31] ;
 wire \soc_inst.cpu_core.register_file.registers[7][3] ;
 wire \soc_inst.cpu_core.register_file.registers[7][4] ;
 wire \soc_inst.cpu_core.register_file.registers[7][5] ;
 wire \soc_inst.cpu_core.register_file.registers[7][6] ;
 wire \soc_inst.cpu_core.register_file.registers[7][7] ;
 wire \soc_inst.cpu_core.register_file.registers[7][8] ;
 wire \soc_inst.cpu_core.register_file.registers[7][9] ;
 wire \soc_inst.cpu_core.register_file.registers[8][0] ;
 wire \soc_inst.cpu_core.register_file.registers[8][10] ;
 wire \soc_inst.cpu_core.register_file.registers[8][11] ;
 wire \soc_inst.cpu_core.register_file.registers[8][12] ;
 wire \soc_inst.cpu_core.register_file.registers[8][13] ;
 wire \soc_inst.cpu_core.register_file.registers[8][14] ;
 wire \soc_inst.cpu_core.register_file.registers[8][15] ;
 wire \soc_inst.cpu_core.register_file.registers[8][16] ;
 wire \soc_inst.cpu_core.register_file.registers[8][17] ;
 wire \soc_inst.cpu_core.register_file.registers[8][18] ;
 wire \soc_inst.cpu_core.register_file.registers[8][19] ;
 wire \soc_inst.cpu_core.register_file.registers[8][1] ;
 wire \soc_inst.cpu_core.register_file.registers[8][20] ;
 wire \soc_inst.cpu_core.register_file.registers[8][21] ;
 wire \soc_inst.cpu_core.register_file.registers[8][22] ;
 wire \soc_inst.cpu_core.register_file.registers[8][23] ;
 wire \soc_inst.cpu_core.register_file.registers[8][24] ;
 wire \soc_inst.cpu_core.register_file.registers[8][25] ;
 wire \soc_inst.cpu_core.register_file.registers[8][26] ;
 wire \soc_inst.cpu_core.register_file.registers[8][27] ;
 wire \soc_inst.cpu_core.register_file.registers[8][28] ;
 wire \soc_inst.cpu_core.register_file.registers[8][29] ;
 wire \soc_inst.cpu_core.register_file.registers[8][2] ;
 wire \soc_inst.cpu_core.register_file.registers[8][30] ;
 wire \soc_inst.cpu_core.register_file.registers[8][31] ;
 wire \soc_inst.cpu_core.register_file.registers[8][3] ;
 wire \soc_inst.cpu_core.register_file.registers[8][4] ;
 wire \soc_inst.cpu_core.register_file.registers[8][5] ;
 wire \soc_inst.cpu_core.register_file.registers[8][6] ;
 wire \soc_inst.cpu_core.register_file.registers[8][7] ;
 wire \soc_inst.cpu_core.register_file.registers[8][8] ;
 wire \soc_inst.cpu_core.register_file.registers[8][9] ;
 wire \soc_inst.cpu_core.register_file.registers[9][0] ;
 wire \soc_inst.cpu_core.register_file.registers[9][10] ;
 wire \soc_inst.cpu_core.register_file.registers[9][11] ;
 wire \soc_inst.cpu_core.register_file.registers[9][12] ;
 wire \soc_inst.cpu_core.register_file.registers[9][13] ;
 wire \soc_inst.cpu_core.register_file.registers[9][14] ;
 wire \soc_inst.cpu_core.register_file.registers[9][15] ;
 wire \soc_inst.cpu_core.register_file.registers[9][16] ;
 wire \soc_inst.cpu_core.register_file.registers[9][17] ;
 wire \soc_inst.cpu_core.register_file.registers[9][18] ;
 wire \soc_inst.cpu_core.register_file.registers[9][19] ;
 wire \soc_inst.cpu_core.register_file.registers[9][1] ;
 wire \soc_inst.cpu_core.register_file.registers[9][20] ;
 wire \soc_inst.cpu_core.register_file.registers[9][21] ;
 wire \soc_inst.cpu_core.register_file.registers[9][22] ;
 wire \soc_inst.cpu_core.register_file.registers[9][23] ;
 wire \soc_inst.cpu_core.register_file.registers[9][24] ;
 wire \soc_inst.cpu_core.register_file.registers[9][25] ;
 wire \soc_inst.cpu_core.register_file.registers[9][26] ;
 wire \soc_inst.cpu_core.register_file.registers[9][27] ;
 wire \soc_inst.cpu_core.register_file.registers[9][28] ;
 wire \soc_inst.cpu_core.register_file.registers[9][29] ;
 wire \soc_inst.cpu_core.register_file.registers[9][2] ;
 wire \soc_inst.cpu_core.register_file.registers[9][30] ;
 wire \soc_inst.cpu_core.register_file.registers[9][31] ;
 wire \soc_inst.cpu_core.register_file.registers[9][3] ;
 wire \soc_inst.cpu_core.register_file.registers[9][4] ;
 wire \soc_inst.cpu_core.register_file.registers[9][5] ;
 wire \soc_inst.cpu_core.register_file.registers[9][6] ;
 wire \soc_inst.cpu_core.register_file.registers[9][7] ;
 wire \soc_inst.cpu_core.register_file.registers[9][8] ;
 wire \soc_inst.cpu_core.register_file.registers[9][9] ;
 wire \soc_inst.flash_cs_n ;
 wire \soc_inst.gpio_inst.gpio_out[0] ;
 wire \soc_inst.gpio_inst.gpio_out[1] ;
 wire \soc_inst.gpio_inst.gpio_out[2] ;
 wire \soc_inst.gpio_inst.gpio_out[3] ;
 wire \soc_inst.gpio_inst.gpio_out[4] ;
 wire \soc_inst.gpio_inst.gpio_out[5] ;
 wire \soc_inst.gpio_inst.gpio_sync1[0] ;
 wire \soc_inst.gpio_inst.gpio_sync1[1] ;
 wire \soc_inst.gpio_inst.gpio_sync1[2] ;
 wire \soc_inst.gpio_inst.gpio_sync1[3] ;
 wire \soc_inst.gpio_inst.gpio_sync1[4] ;
 wire \soc_inst.gpio_inst.gpio_sync1[5] ;
 wire \soc_inst.gpio_inst.gpio_sync1[6] ;
 wire \soc_inst.gpio_inst.gpio_sync2[0] ;
 wire \soc_inst.gpio_inst.gpio_sync2[1] ;
 wire \soc_inst.gpio_inst.gpio_sync2[2] ;
 wire \soc_inst.gpio_inst.gpio_sync2[3] ;
 wire \soc_inst.gpio_inst.gpio_sync2[4] ;
 wire \soc_inst.gpio_inst.gpio_sync2[5] ;
 wire \soc_inst.gpio_inst.gpio_sync2[6] ;
 wire \soc_inst.gpio_inst.int_en_reg[0] ;
 wire \soc_inst.gpio_inst.int_en_reg[1] ;
 wire \soc_inst.gpio_inst.int_en_reg[2] ;
 wire \soc_inst.gpio_inst.int_en_reg[3] ;
 wire \soc_inst.gpio_inst.int_en_reg[4] ;
 wire \soc_inst.gpio_inst.int_en_reg[5] ;
 wire \soc_inst.gpio_inst.int_en_reg[6] ;
 wire \soc_inst.gpio_inst.int_pend_reg[0] ;
 wire \soc_inst.gpio_inst.int_pend_reg[1] ;
 wire \soc_inst.gpio_inst.int_pend_reg[2] ;
 wire \soc_inst.gpio_inst.int_pend_reg[3] ;
 wire \soc_inst.gpio_inst.int_pend_reg[4] ;
 wire \soc_inst.gpio_inst.int_pend_reg[5] ;
 wire \soc_inst.gpio_inst.int_pend_reg[6] ;
 wire \soc_inst.i2c_ena ;
 wire \soc_inst.i2c_inst.ack_enable ;
 wire \soc_inst.i2c_inst.ack_received ;
 wire \soc_inst.i2c_inst.arb_lost ;
 wire \soc_inst.i2c_inst.bit_cnt[0] ;
 wire \soc_inst.i2c_inst.bit_cnt[1] ;
 wire \soc_inst.i2c_inst.bit_cnt[2] ;
 wire \soc_inst.i2c_inst.bit_cnt[3] ;
 wire \soc_inst.i2c_inst.clk_cnt[0] ;
 wire \soc_inst.i2c_inst.clk_cnt[1] ;
 wire \soc_inst.i2c_inst.clk_cnt[2] ;
 wire \soc_inst.i2c_inst.clk_cnt[3] ;
 wire \soc_inst.i2c_inst.clk_cnt[4] ;
 wire \soc_inst.i2c_inst.clk_cnt[5] ;
 wire \soc_inst.i2c_inst.clk_cnt[6] ;
 wire \soc_inst.i2c_inst.clk_cnt[7] ;
 wire \soc_inst.i2c_inst.ctrl_reg[2] ;
 wire \soc_inst.i2c_inst.ctrl_reg[4] ;
 wire \soc_inst.i2c_inst.data_reg[0] ;
 wire \soc_inst.i2c_inst.data_reg[1] ;
 wire \soc_inst.i2c_inst.data_reg[2] ;
 wire \soc_inst.i2c_inst.data_reg[3] ;
 wire \soc_inst.i2c_inst.data_reg[4] ;
 wire \soc_inst.i2c_inst.data_reg[5] ;
 wire \soc_inst.i2c_inst.data_reg[6] ;
 wire \soc_inst.i2c_inst.data_reg[7] ;
 wire \soc_inst.i2c_inst.prescale_reg[5] ;
 wire \soc_inst.i2c_inst.prescale_reg[6] ;
 wire \soc_inst.i2c_inst.restart_pending ;
 wire \soc_inst.i2c_inst.shift_reg[0] ;
 wire \soc_inst.i2c_inst.shift_reg[1] ;
 wire \soc_inst.i2c_inst.shift_reg[2] ;
 wire \soc_inst.i2c_inst.shift_reg[3] ;
 wire \soc_inst.i2c_inst.shift_reg[4] ;
 wire \soc_inst.i2c_inst.shift_reg[5] ;
 wire \soc_inst.i2c_inst.shift_reg[6] ;
 wire \soc_inst.i2c_inst.shift_reg[7] ;
 wire \soc_inst.i2c_inst.start_pending ;
 wire \soc_inst.i2c_inst.state[0] ;
 wire \soc_inst.i2c_inst.state[1] ;
 wire \soc_inst.i2c_inst.state[2] ;
 wire \soc_inst.i2c_inst.state[3] ;
 wire \soc_inst.i2c_inst.status_reg[0] ;
 wire \soc_inst.i2c_inst.status_reg[1] ;
 wire \soc_inst.i2c_inst.status_reg[2] ;
 wire \soc_inst.i2c_inst.status_reg[3] ;
 wire \soc_inst.i2c_inst.stop_pending ;
 wire \soc_inst.i2c_inst.transfer_done ;
 wire \soc_inst.mem_ctrl.access_state[1] ;
 wire \soc_inst.mem_ctrl.access_state[2] ;
 wire \soc_inst.mem_ctrl.access_state[3] ;
 wire \soc_inst.mem_ctrl.access_state[4] ;
 wire \soc_inst.mem_ctrl.instr_ready_reg ;
 wire \soc_inst.mem_ctrl.next_instr_addr[0] ;
 wire \soc_inst.mem_ctrl.next_instr_data[0] ;
 wire \soc_inst.mem_ctrl.next_instr_data[10] ;
 wire \soc_inst.mem_ctrl.next_instr_data[11] ;
 wire \soc_inst.mem_ctrl.next_instr_data[12] ;
 wire \soc_inst.mem_ctrl.next_instr_data[13] ;
 wire \soc_inst.mem_ctrl.next_instr_data[14] ;
 wire \soc_inst.mem_ctrl.next_instr_data[15] ;
 wire \soc_inst.mem_ctrl.next_instr_data[16] ;
 wire \soc_inst.mem_ctrl.next_instr_data[17] ;
 wire \soc_inst.mem_ctrl.next_instr_data[18] ;
 wire \soc_inst.mem_ctrl.next_instr_data[19] ;
 wire \soc_inst.mem_ctrl.next_instr_data[1] ;
 wire \soc_inst.mem_ctrl.next_instr_data[20] ;
 wire \soc_inst.mem_ctrl.next_instr_data[21] ;
 wire \soc_inst.mem_ctrl.next_instr_data[22] ;
 wire \soc_inst.mem_ctrl.next_instr_data[23] ;
 wire \soc_inst.mem_ctrl.next_instr_data[24] ;
 wire \soc_inst.mem_ctrl.next_instr_data[25] ;
 wire \soc_inst.mem_ctrl.next_instr_data[26] ;
 wire \soc_inst.mem_ctrl.next_instr_data[27] ;
 wire \soc_inst.mem_ctrl.next_instr_data[28] ;
 wire \soc_inst.mem_ctrl.next_instr_data[29] ;
 wire \soc_inst.mem_ctrl.next_instr_data[2] ;
 wire \soc_inst.mem_ctrl.next_instr_data[30] ;
 wire \soc_inst.mem_ctrl.next_instr_data[31] ;
 wire \soc_inst.mem_ctrl.next_instr_data[3] ;
 wire \soc_inst.mem_ctrl.next_instr_data[4] ;
 wire \soc_inst.mem_ctrl.next_instr_data[5] ;
 wire \soc_inst.mem_ctrl.next_instr_data[6] ;
 wire \soc_inst.mem_ctrl.next_instr_data[7] ;
 wire \soc_inst.mem_ctrl.next_instr_data[8] ;
 wire \soc_inst.mem_ctrl.next_instr_data[9] ;
 wire \soc_inst.mem_ctrl.next_instr_ready_reg ;
 wire \soc_inst.mem_ctrl.ram_cs_n ;
 wire \soc_inst.mem_ctrl.spi_addr[10] ;
 wire \soc_inst.mem_ctrl.spi_addr[11] ;
 wire \soc_inst.mem_ctrl.spi_addr[12] ;
 wire \soc_inst.mem_ctrl.spi_addr[13] ;
 wire \soc_inst.mem_ctrl.spi_addr[14] ;
 wire \soc_inst.mem_ctrl.spi_addr[15] ;
 wire \soc_inst.mem_ctrl.spi_addr[16] ;
 wire \soc_inst.mem_ctrl.spi_addr[17] ;
 wire \soc_inst.mem_ctrl.spi_addr[18] ;
 wire \soc_inst.mem_ctrl.spi_addr[19] ;
 wire \soc_inst.mem_ctrl.spi_addr[1] ;
 wire \soc_inst.mem_ctrl.spi_addr[20] ;
 wire \soc_inst.mem_ctrl.spi_addr[21] ;
 wire \soc_inst.mem_ctrl.spi_addr[22] ;
 wire \soc_inst.mem_ctrl.spi_addr[23] ;
 wire \soc_inst.mem_ctrl.spi_addr[2] ;
 wire \soc_inst.mem_ctrl.spi_addr[3] ;
 wire \soc_inst.mem_ctrl.spi_addr[4] ;
 wire \soc_inst.mem_ctrl.spi_addr[5] ;
 wire \soc_inst.mem_ctrl.spi_addr[6] ;
 wire \soc_inst.mem_ctrl.spi_addr[7] ;
 wire \soc_inst.mem_ctrl.spi_addr[8] ;
 wire \soc_inst.mem_ctrl.spi_addr[9] ;
 wire \soc_inst.mem_ctrl.spi_data_in[0] ;
 wire \soc_inst.mem_ctrl.spi_data_in[10] ;
 wire \soc_inst.mem_ctrl.spi_data_in[11] ;
 wire \soc_inst.mem_ctrl.spi_data_in[12] ;
 wire \soc_inst.mem_ctrl.spi_data_in[13] ;
 wire \soc_inst.mem_ctrl.spi_data_in[14] ;
 wire \soc_inst.mem_ctrl.spi_data_in[15] ;
 wire \soc_inst.mem_ctrl.spi_data_in[16] ;
 wire \soc_inst.mem_ctrl.spi_data_in[17] ;
 wire \soc_inst.mem_ctrl.spi_data_in[18] ;
 wire \soc_inst.mem_ctrl.spi_data_in[19] ;
 wire \soc_inst.mem_ctrl.spi_data_in[1] ;
 wire \soc_inst.mem_ctrl.spi_data_in[20] ;
 wire \soc_inst.mem_ctrl.spi_data_in[21] ;
 wire \soc_inst.mem_ctrl.spi_data_in[22] ;
 wire \soc_inst.mem_ctrl.spi_data_in[23] ;
 wire \soc_inst.mem_ctrl.spi_data_in[24] ;
 wire \soc_inst.mem_ctrl.spi_data_in[25] ;
 wire \soc_inst.mem_ctrl.spi_data_in[26] ;
 wire \soc_inst.mem_ctrl.spi_data_in[27] ;
 wire \soc_inst.mem_ctrl.spi_data_in[28] ;
 wire \soc_inst.mem_ctrl.spi_data_in[29] ;
 wire \soc_inst.mem_ctrl.spi_data_in[2] ;
 wire \soc_inst.mem_ctrl.spi_data_in[30] ;
 wire \soc_inst.mem_ctrl.spi_data_in[31] ;
 wire \soc_inst.mem_ctrl.spi_data_in[3] ;
 wire \soc_inst.mem_ctrl.spi_data_in[4] ;
 wire \soc_inst.mem_ctrl.spi_data_in[5] ;
 wire \soc_inst.mem_ctrl.spi_data_in[6] ;
 wire \soc_inst.mem_ctrl.spi_data_in[7] ;
 wire \soc_inst.mem_ctrl.spi_data_in[8] ;
 wire \soc_inst.mem_ctrl.spi_data_in[9] ;
 wire \soc_inst.mem_ctrl.spi_data_len[3] ;
 wire \soc_inst.mem_ctrl.spi_data_len[4] ;
 wire \soc_inst.mem_ctrl.spi_data_len[5] ;
 wire \soc_inst.mem_ctrl.spi_data_out[0] ;
 wire \soc_inst.mem_ctrl.spi_data_out[10] ;
 wire \soc_inst.mem_ctrl.spi_data_out[11] ;
 wire \soc_inst.mem_ctrl.spi_data_out[12] ;
 wire \soc_inst.mem_ctrl.spi_data_out[13] ;
 wire \soc_inst.mem_ctrl.spi_data_out[14] ;
 wire \soc_inst.mem_ctrl.spi_data_out[15] ;
 wire \soc_inst.mem_ctrl.spi_data_out[16] ;
 wire \soc_inst.mem_ctrl.spi_data_out[17] ;
 wire \soc_inst.mem_ctrl.spi_data_out[18] ;
 wire \soc_inst.mem_ctrl.spi_data_out[19] ;
 wire \soc_inst.mem_ctrl.spi_data_out[1] ;
 wire \soc_inst.mem_ctrl.spi_data_out[20] ;
 wire \soc_inst.mem_ctrl.spi_data_out[21] ;
 wire \soc_inst.mem_ctrl.spi_data_out[22] ;
 wire \soc_inst.mem_ctrl.spi_data_out[23] ;
 wire \soc_inst.mem_ctrl.spi_data_out[24] ;
 wire \soc_inst.mem_ctrl.spi_data_out[25] ;
 wire \soc_inst.mem_ctrl.spi_data_out[26] ;
 wire \soc_inst.mem_ctrl.spi_data_out[27] ;
 wire \soc_inst.mem_ctrl.spi_data_out[28] ;
 wire \soc_inst.mem_ctrl.spi_data_out[29] ;
 wire \soc_inst.mem_ctrl.spi_data_out[2] ;
 wire \soc_inst.mem_ctrl.spi_data_out[30] ;
 wire \soc_inst.mem_ctrl.spi_data_out[31] ;
 wire \soc_inst.mem_ctrl.spi_data_out[3] ;
 wire \soc_inst.mem_ctrl.spi_data_out[4] ;
 wire \soc_inst.mem_ctrl.spi_data_out[5] ;
 wire \soc_inst.mem_ctrl.spi_data_out[6] ;
 wire \soc_inst.mem_ctrl.spi_data_out[7] ;
 wire \soc_inst.mem_ctrl.spi_data_out[8] ;
 wire \soc_inst.mem_ctrl.spi_data_out[9] ;
 wire \soc_inst.mem_ctrl.spi_done ;
 wire \soc_inst.mem_ctrl.spi_is_instr ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.boot_mode_latched ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.initialized ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.is_write_op ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.sample_trigger ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d1 ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d2 ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d3 ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.start ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.stop ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.write_enable ;
 wire \soc_inst.mem_ctrl.spi_mem_inst.write_mosi ;
 wire \soc_inst.mem_ctrl.spi_read_enable ;
 wire \soc_inst.pwm_inst.channel_counter[0][0] ;
 wire \soc_inst.pwm_inst.channel_counter[0][10] ;
 wire \soc_inst.pwm_inst.channel_counter[0][11] ;
 wire \soc_inst.pwm_inst.channel_counter[0][12] ;
 wire \soc_inst.pwm_inst.channel_counter[0][13] ;
 wire \soc_inst.pwm_inst.channel_counter[0][14] ;
 wire \soc_inst.pwm_inst.channel_counter[0][15] ;
 wire \soc_inst.pwm_inst.channel_counter[0][1] ;
 wire \soc_inst.pwm_inst.channel_counter[0][2] ;
 wire \soc_inst.pwm_inst.channel_counter[0][3] ;
 wire \soc_inst.pwm_inst.channel_counter[0][4] ;
 wire \soc_inst.pwm_inst.channel_counter[0][5] ;
 wire \soc_inst.pwm_inst.channel_counter[0][6] ;
 wire \soc_inst.pwm_inst.channel_counter[0][7] ;
 wire \soc_inst.pwm_inst.channel_counter[0][8] ;
 wire \soc_inst.pwm_inst.channel_counter[0][9] ;
 wire \soc_inst.pwm_inst.channel_duty[0][0] ;
 wire \soc_inst.pwm_inst.channel_duty[0][10] ;
 wire \soc_inst.pwm_inst.channel_duty[0][11] ;
 wire \soc_inst.pwm_inst.channel_duty[0][12] ;
 wire \soc_inst.pwm_inst.channel_duty[0][13] ;
 wire \soc_inst.pwm_inst.channel_duty[0][14] ;
 wire \soc_inst.pwm_inst.channel_duty[0][15] ;
 wire \soc_inst.pwm_inst.channel_duty[0][1] ;
 wire \soc_inst.pwm_inst.channel_duty[0][2] ;
 wire \soc_inst.pwm_inst.channel_duty[0][3] ;
 wire \soc_inst.pwm_inst.channel_duty[0][4] ;
 wire \soc_inst.pwm_inst.channel_duty[0][5] ;
 wire \soc_inst.pwm_inst.channel_duty[0][6] ;
 wire \soc_inst.pwm_inst.channel_duty[0][7] ;
 wire \soc_inst.pwm_inst.channel_duty[0][8] ;
 wire \soc_inst.pwm_inst.channel_duty[0][9] ;
 wire \soc_inst.spi_ena ;
 wire \soc_inst.spi_inst.bit_counter[0] ;
 wire \soc_inst.spi_inst.bit_counter[1] ;
 wire \soc_inst.spi_inst.bit_counter[2] ;
 wire \soc_inst.spi_inst.bit_counter[3] ;
 wire \soc_inst.spi_inst.bit_counter[4] ;
 wire \soc_inst.spi_inst.bit_counter[5] ;
 wire \soc_inst.spi_inst.busy ;
 wire \soc_inst.spi_inst.clk_counter[0] ;
 wire \soc_inst.spi_inst.clk_counter[1] ;
 wire \soc_inst.spi_inst.clk_counter[2] ;
 wire \soc_inst.spi_inst.clk_counter[3] ;
 wire \soc_inst.spi_inst.clk_counter[4] ;
 wire \soc_inst.spi_inst.clk_counter[5] ;
 wire \soc_inst.spi_inst.clk_counter[6] ;
 wire \soc_inst.spi_inst.clk_counter[7] ;
 wire \soc_inst.spi_inst.clock_divider[5] ;
 wire \soc_inst.spi_inst.clock_divider[6] ;
 wire \soc_inst.spi_inst.clock_divider[7] ;
 wire \soc_inst.spi_inst.cpha ;
 wire \soc_inst.spi_inst.cpol ;
 wire \soc_inst.spi_inst.done ;
 wire \soc_inst.spi_inst.len_sel[0] ;
 wire \soc_inst.spi_inst.len_sel[1] ;
 wire \soc_inst.spi_inst.next_state[0] ;
 wire \soc_inst.spi_inst.next_state[1] ;
 wire \soc_inst.spi_inst.rx_shift_reg[0] ;
 wire \soc_inst.spi_inst.rx_shift_reg[10] ;
 wire \soc_inst.spi_inst.rx_shift_reg[11] ;
 wire \soc_inst.spi_inst.rx_shift_reg[12] ;
 wire \soc_inst.spi_inst.rx_shift_reg[13] ;
 wire \soc_inst.spi_inst.rx_shift_reg[14] ;
 wire \soc_inst.spi_inst.rx_shift_reg[15] ;
 wire \soc_inst.spi_inst.rx_shift_reg[16] ;
 wire \soc_inst.spi_inst.rx_shift_reg[17] ;
 wire \soc_inst.spi_inst.rx_shift_reg[18] ;
 wire \soc_inst.spi_inst.rx_shift_reg[19] ;
 wire \soc_inst.spi_inst.rx_shift_reg[1] ;
 wire \soc_inst.spi_inst.rx_shift_reg[20] ;
 wire \soc_inst.spi_inst.rx_shift_reg[21] ;
 wire \soc_inst.spi_inst.rx_shift_reg[22] ;
 wire \soc_inst.spi_inst.rx_shift_reg[23] ;
 wire \soc_inst.spi_inst.rx_shift_reg[24] ;
 wire \soc_inst.spi_inst.rx_shift_reg[25] ;
 wire \soc_inst.spi_inst.rx_shift_reg[26] ;
 wire \soc_inst.spi_inst.rx_shift_reg[27] ;
 wire \soc_inst.spi_inst.rx_shift_reg[28] ;
 wire \soc_inst.spi_inst.rx_shift_reg[29] ;
 wire \soc_inst.spi_inst.rx_shift_reg[2] ;
 wire \soc_inst.spi_inst.rx_shift_reg[30] ;
 wire \soc_inst.spi_inst.rx_shift_reg[31] ;
 wire \soc_inst.spi_inst.rx_shift_reg[3] ;
 wire \soc_inst.spi_inst.rx_shift_reg[4] ;
 wire \soc_inst.spi_inst.rx_shift_reg[5] ;
 wire \soc_inst.spi_inst.rx_shift_reg[6] ;
 wire \soc_inst.spi_inst.rx_shift_reg[7] ;
 wire \soc_inst.spi_inst.rx_shift_reg[8] ;
 wire \soc_inst.spi_inst.rx_shift_reg[9] ;
 wire \soc_inst.spi_inst.spi_clk_en ;
 wire \soc_inst.spi_inst.spi_mosi ;
 wire \soc_inst.spi_inst.spi_sclk ;
 wire \soc_inst.spi_inst.start_pending ;
 wire \soc_inst.spi_inst.state[0] ;
 wire \soc_inst.spi_inst.state[1] ;
 wire \soc_inst.spi_inst.tx_shift_reg[0] ;
 wire \soc_inst.spi_inst.tx_shift_reg[10] ;
 wire \soc_inst.spi_inst.tx_shift_reg[11] ;
 wire \soc_inst.spi_inst.tx_shift_reg[12] ;
 wire \soc_inst.spi_inst.tx_shift_reg[13] ;
 wire \soc_inst.spi_inst.tx_shift_reg[14] ;
 wire \soc_inst.spi_inst.tx_shift_reg[15] ;
 wire \soc_inst.spi_inst.tx_shift_reg[16] ;
 wire \soc_inst.spi_inst.tx_shift_reg[17] ;
 wire \soc_inst.spi_inst.tx_shift_reg[18] ;
 wire \soc_inst.spi_inst.tx_shift_reg[19] ;
 wire \soc_inst.spi_inst.tx_shift_reg[1] ;
 wire \soc_inst.spi_inst.tx_shift_reg[20] ;
 wire \soc_inst.spi_inst.tx_shift_reg[21] ;
 wire \soc_inst.spi_inst.tx_shift_reg[22] ;
 wire \soc_inst.spi_inst.tx_shift_reg[23] ;
 wire \soc_inst.spi_inst.tx_shift_reg[24] ;
 wire \soc_inst.spi_inst.tx_shift_reg[25] ;
 wire \soc_inst.spi_inst.tx_shift_reg[26] ;
 wire \soc_inst.spi_inst.tx_shift_reg[27] ;
 wire \soc_inst.spi_inst.tx_shift_reg[28] ;
 wire \soc_inst.spi_inst.tx_shift_reg[29] ;
 wire \soc_inst.spi_inst.tx_shift_reg[2] ;
 wire \soc_inst.spi_inst.tx_shift_reg[30] ;
 wire \soc_inst.spi_inst.tx_shift_reg[31] ;
 wire \soc_inst.spi_inst.tx_shift_reg[3] ;
 wire \soc_inst.spi_inst.tx_shift_reg[4] ;
 wire \soc_inst.spi_inst.tx_shift_reg[5] ;
 wire \soc_inst.spi_inst.tx_shift_reg[6] ;
 wire \soc_inst.spi_inst.tx_shift_reg[7] ;
 wire \soc_inst.spi_inst.tx_shift_reg[8] ;
 wire \soc_inst.spi_inst.tx_shift_reg[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ;
 wire \soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ;
 wire net78;
 wire net79;
 wire clknet_leaf_0_clk;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire [0:0] _11835_;
 wire [0:0] _11836_;
 wire [0:0] _11837_;
 wire [0:0] \soc_inst.gpio_bidir_oe ;
 wire [0:0] \soc_inst.gpio_bidir_out ;
 wire [0:0] \soc_inst.pwm_ena ;
 wire [0:0] \soc_inst.pwm_inst.channel_idx ;
 wire [0:0] \soc_inst.uart_tx ;

 sg13g2_inv_1 _11838_ (.Y(_07763_),
    .A(net1838));
 sg13g2_inv_1 _11839_ (.Y(_07764_),
    .A(net738));
 sg13g2_inv_1 _11840_ (.Y(_07765_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ));
 sg13g2_inv_1 _11841_ (.Y(_07766_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ));
 sg13g2_inv_1 _11842_ (.Y(_07767_),
    .A(net303));
 sg13g2_inv_1 _11843_ (.Y(_07768_),
    .A(net1888));
 sg13g2_inv_1 _11844_ (.Y(_07769_),
    .A(net2489));
 sg13g2_inv_1 _11845_ (.Y(_07770_),
    .A(net1417));
 sg13g2_inv_1 _11846_ (.Y(_07771_),
    .A(net746));
 sg13g2_inv_2 _11847_ (.Y(_07772_),
    .A(net670));
 sg13g2_inv_1 _11848_ (.Y(_07773_),
    .A(net1018));
 sg13g2_inv_1 _11849_ (.Y(_07774_),
    .A(net921));
 sg13g2_inv_1 _11850_ (.Y(_07775_),
    .A(net665));
 sg13g2_inv_1 _11851_ (.Y(_07776_),
    .A(net529));
 sg13g2_inv_1 _11852_ (.Y(_07777_),
    .A(net6178));
 sg13g2_inv_2 _11853_ (.Y(_07778_),
    .A(_00318_));
 sg13g2_inv_1 _11854_ (.Y(_07779_),
    .A(_00317_));
 sg13g2_inv_1 _11855_ (.Y(_07780_),
    .A(_00316_));
 sg13g2_inv_1 _11856_ (.Y(_07781_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ));
 sg13g2_inv_1 _11857_ (.Y(_07782_),
    .A(net2406));
 sg13g2_inv_1 _11858_ (.Y(_07783_),
    .A(_00290_));
 sg13g2_inv_8 _11859_ (.Y(_07784_),
    .A(net6468));
 sg13g2_inv_8 _11860_ (.Y(_07785_),
    .A(net6471));
 sg13g2_inv_1 _11861_ (.Y(_07786_),
    .A(_00274_));
 sg13g2_inv_1 _11862_ (.Y(_07787_),
    .A(_00271_));
 sg13g2_inv_1 _11863_ (.Y(_07788_),
    .A(_00267_));
 sg13g2_inv_1 _11864_ (.Y(_07789_),
    .A(net2771));
 sg13g2_inv_1 _11865_ (.Y(_07790_),
    .A(net2792));
 sg13g2_inv_2 _11866_ (.Y(_07791_),
    .A(net2418));
 sg13g2_inv_1 _11867_ (.Y(_07792_),
    .A(_00257_));
 sg13g2_inv_1 _11868_ (.Y(_07793_),
    .A(_00238_));
 sg13g2_inv_1 _11869_ (.Y(_07794_),
    .A(_00235_));
 sg13g2_inv_1 _11870_ (.Y(_07795_),
    .A(_00225_));
 sg13g2_inv_1 _11871_ (.Y(_07796_),
    .A(_00224_));
 sg13g2_inv_1 _11872_ (.Y(_07797_),
    .A(_00223_));
 sg13g2_inv_1 _11873_ (.Y(_07798_),
    .A(net2237));
 sg13g2_inv_1 _11874_ (.Y(_00173_),
    .A(net770));
 sg13g2_inv_1 _11875_ (.Y(_07799_),
    .A(net2919));
 sg13g2_inv_1 _11876_ (.Y(_07800_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ));
 sg13g2_inv_2 _11877_ (.Y(_07801_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ));
 sg13g2_inv_1 _11878_ (.Y(_07802_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ));
 sg13g2_inv_2 _11879_ (.Y(_07803_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ));
 sg13g2_inv_1 _11880_ (.Y(_07804_),
    .A(\soc_inst.spi_inst.state[1] ));
 sg13g2_inv_1 _11881_ (.Y(_07805_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[2] ));
 sg13g2_inv_1 _11882_ (.Y(_07806_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[4] ));
 sg13g2_inv_1 _11883_ (.Y(_07807_),
    .A(net2564));
 sg13g2_inv_1 _11884_ (.Y(_07808_),
    .A(net6303));
 sg13g2_inv_2 _11885_ (.Y(_07809_),
    .A(net6294));
 sg13g2_inv_4 _11886_ (.A(net3318),
    .Y(_07810_));
 sg13g2_inv_1 _11887_ (.Y(_07811_),
    .A(net6212));
 sg13g2_inv_2 _11888_ (.Y(_07812_),
    .A(net1538));
 sg13g2_inv_8 _11889_ (.Y(_07813_),
    .A(net3388));
 sg13g2_inv_1 _11890_ (.Y(_07814_),
    .A(net2365));
 sg13g2_inv_4 _11891_ (.A(net3263),
    .Y(_07815_));
 sg13g2_inv_2 _11892_ (.Y(_07816_),
    .A(net6505));
 sg13g2_inv_1 _11893_ (.Y(_07817_),
    .A(net2949));
 sg13g2_inv_1 _11894_ (.Y(_07818_),
    .A(net2927));
 sg13g2_inv_1 _11895_ (.Y(_07819_),
    .A(net2904));
 sg13g2_inv_4 _11896_ (.A(net2685),
    .Y(_07820_));
 sg13g2_inv_1 _11897_ (.Y(_07821_),
    .A(net3031));
 sg13g2_inv_2 _11898_ (.Y(_07822_),
    .A(net3076));
 sg13g2_inv_1 _11899_ (.Y(_07823_),
    .A(net2831));
 sg13g2_inv_4 _11900_ (.A(net2492),
    .Y(_07824_));
 sg13g2_inv_1 _11901_ (.Y(_07825_),
    .A(net2967));
 sg13g2_inv_1 _11902_ (.Y(_07826_),
    .A(net2738));
 sg13g2_inv_1 _11903_ (.Y(_07827_),
    .A(net3310));
 sg13g2_inv_2 _11904_ (.Y(_07828_),
    .A(net2703));
 sg13g2_inv_1 _11905_ (.Y(_07829_),
    .A(net3125));
 sg13g2_inv_2 _11906_ (.Y(_07830_),
    .A(net2713));
 sg13g2_inv_1 _11907_ (.Y(_07831_),
    .A(net3166));
 sg13g2_inv_2 _11908_ (.Y(_07832_),
    .A(net2807));
 sg13g2_inv_1 _11909_ (.Y(_07833_),
    .A(net2968));
 sg13g2_inv_2 _11910_ (.Y(_07834_),
    .A(net2493));
 sg13g2_inv_1 _11911_ (.Y(_07835_),
    .A(net3321));
 sg13g2_inv_2 _11912_ (.Y(_07836_),
    .A(net3044));
 sg13g2_inv_1 _11913_ (.Y(_07837_),
    .A(net2954));
 sg13g2_inv_2 _11914_ (.Y(_07838_),
    .A(net3010));
 sg13g2_inv_1 _11915_ (.Y(_07839_),
    .A(net3140));
 sg13g2_inv_2 _11916_ (.Y(_07840_),
    .A(\soc_inst.core_instr_addr[11] ));
 sg13g2_inv_2 _11917_ (.Y(_07841_),
    .A(net2820));
 sg13g2_inv_2 _11918_ (.Y(_07842_),
    .A(net3247));
 sg13g2_inv_1 _11919_ (.Y(_07843_),
    .A(net3082));
 sg13g2_inv_1 _11920_ (.Y(_07844_),
    .A(net3311));
 sg13g2_inv_1 _11921_ (.Y(_07845_),
    .A(net2865));
 sg13g2_inv_1 _11922_ (.Y(_07846_),
    .A(net3299));
 sg13g2_inv_1 _11923_ (.Y(_07847_),
    .A(net2657));
 sg13g2_inv_1 _11924_ (.Y(_07848_),
    .A(net2704));
 sg13g2_inv_1 _11925_ (.Y(_07849_),
    .A(net3177));
 sg13g2_inv_2 _11926_ (.Y(_07850_),
    .A(net3138));
 sg13g2_inv_1 _11927_ (.Y(_07851_),
    .A(net3265));
 sg13g2_inv_1 _11928_ (.Y(_07852_),
    .A(net3092));
 sg13g2_inv_1 _11929_ (.Y(_07853_),
    .A(net3181));
 sg13g2_inv_2 _11930_ (.Y(_07854_),
    .A(net2925));
 sg13g2_inv_1 _11931_ (.Y(_07855_),
    .A(net3054));
 sg13g2_inv_1 _11932_ (.Y(_07856_),
    .A(net3133));
 sg13g2_inv_1 _11933_ (.Y(_07857_),
    .A(net3096));
 sg13g2_inv_2 _11934_ (.Y(_07858_),
    .A(net3129));
 sg13g2_inv_1 _11935_ (.Y(_07859_),
    .A(net3004));
 sg13g2_inv_4 _11936_ (.A(net2693),
    .Y(_07860_));
 sg13g2_inv_1 _11937_ (.Y(_07861_),
    .A(net3078));
 sg13g2_inv_4 _11938_ (.A(net3315),
    .Y(_07862_));
 sg13g2_inv_1 _11939_ (.Y(_07863_),
    .A(net2797));
 sg13g2_inv_2 _11940_ (.Y(_07864_),
    .A(net3173));
 sg13g2_inv_1 _11941_ (.Y(_07865_),
    .A(net6194));
 sg13g2_inv_2 _11942_ (.Y(_07866_),
    .A(net6181));
 sg13g2_inv_1 _11943_ (.Y(_07867_),
    .A(net6179));
 sg13g2_inv_1 _11944_ (.Y(_07868_),
    .A(net6473));
 sg13g2_inv_2 _11945_ (.Y(_07869_),
    .A(net1756));
 sg13g2_inv_1 _11946_ (.Y(_07870_),
    .A(net3205));
 sg13g2_inv_4 _11947_ (.A(net6480),
    .Y(_07871_));
 sg13g2_inv_1 _11948_ (.Y(_07872_),
    .A(net6399));
 sg13g2_inv_1 _11949_ (.Y(_07873_),
    .A(net6488));
 sg13g2_inv_2 _11950_ (.Y(_07874_),
    .A(net6482));
 sg13g2_inv_4 _11951_ (.A(net6490),
    .Y(_07875_));
 sg13g2_inv_1 _11952_ (.Y(_07876_),
    .A(net2659));
 sg13g2_inv_1 _11953_ (.Y(_07877_),
    .A(net1077));
 sg13g2_inv_2 _11954_ (.Y(_07878_),
    .A(net6486));
 sg13g2_inv_2 _11955_ (.Y(_07879_),
    .A(net6485));
 sg13g2_inv_1 _11956_ (.Y(_07880_),
    .A(net3334));
 sg13g2_inv_1 _11957_ (.Y(_07881_),
    .A(net6484));
 sg13g2_inv_2 _11958_ (.Y(_07882_),
    .A(net3366));
 sg13g2_inv_1 _11959_ (.Y(_07883_),
    .A(net1812));
 sg13g2_inv_4 _11960_ (.A(net6552),
    .Y(_07884_));
 sg13g2_inv_1 _11961_ (.Y(_07885_),
    .A(net3207));
 sg13g2_inv_1 _11962_ (.Y(_07886_),
    .A(net3297));
 sg13g2_inv_8 _11963_ (.Y(_07887_),
    .A(net6211));
 sg13g2_inv_8 _11964_ (.Y(_07888_),
    .A(net6208));
 sg13g2_inv_1 _11965_ (.Y(_07889_),
    .A(net2908));
 sg13g2_inv_1 _11966_ (.Y(_07890_),
    .A(net3038));
 sg13g2_inv_1 _11967_ (.Y(_07891_),
    .A(net3104));
 sg13g2_inv_1 _11968_ (.Y(_07892_),
    .A(net2958));
 sg13g2_inv_1 _11969_ (.Y(_07893_),
    .A(net6540));
 sg13g2_inv_1 _11970_ (.Y(_07894_),
    .A(\soc_inst.i2c_inst.start_pending ));
 sg13g2_inv_1 _11971_ (.Y(_07895_),
    .A(net13));
 sg13g2_inv_1 _11972_ (.Y(_07896_),
    .A(net2803));
 sg13g2_inv_1 _11973_ (.Y(_07897_),
    .A(\soc_inst.spi_inst.spi_clk_en ));
 sg13g2_inv_2 _11974_ (.Y(_07898_),
    .A(net2653));
 sg13g2_inv_1 _11975_ (.Y(_07899_),
    .A(net3175));
 sg13g2_inv_1 _11976_ (.Y(_07900_),
    .A(net1842));
 sg13g2_inv_2 _11977_ (.Y(_07901_),
    .A(net400));
 sg13g2_inv_1 _11978_ (.Y(_07902_),
    .A(net3255));
 sg13g2_inv_1 _11979_ (.Y(_07903_),
    .A(net3380));
 sg13g2_inv_1 _11980_ (.Y(_07904_),
    .A(net2464));
 sg13g2_inv_2 _11981_ (.Y(_07905_),
    .A(net3120));
 sg13g2_inv_1 _11982_ (.Y(_07906_),
    .A(\soc_inst.cpu_core.csr_file.mtime[34] ));
 sg13g2_inv_1 _11983_ (.Y(_07907_),
    .A(net358));
 sg13g2_inv_1 _11984_ (.Y(_07908_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ));
 sg13g2_inv_1 _11985_ (.Y(_07909_),
    .A(net2093));
 sg13g2_inv_1 _11986_ (.Y(_07910_),
    .A(net2809));
 sg13g2_inv_1 _11987_ (.Y(_07911_),
    .A(net2324));
 sg13g2_inv_1 _11988_ (.Y(_07912_),
    .A(net1316));
 sg13g2_inv_1 _11989_ (.Y(_07913_),
    .A(net2046));
 sg13g2_inv_1 _11990_ (.Y(_07914_),
    .A(net1748));
 sg13g2_inv_1 _11991_ (.Y(_07915_),
    .A(net1946));
 sg13g2_inv_1 _11992_ (.Y(_07916_),
    .A(net2271));
 sg13g2_inv_1 _11993_ (.Y(_07917_),
    .A(net2258));
 sg13g2_inv_1 _11994_ (.Y(_07918_),
    .A(net2834));
 sg13g2_inv_1 _11995_ (.Y(_07919_),
    .A(net2767));
 sg13g2_inv_1 _11996_ (.Y(_07920_),
    .A(net2342));
 sg13g2_inv_1 _11997_ (.Y(_07921_),
    .A(net2763));
 sg13g2_inv_1 _11998_ (.Y(_07922_),
    .A(net2590));
 sg13g2_inv_1 _11999_ (.Y(_07923_),
    .A(net2483));
 sg13g2_inv_1 _12000_ (.Y(_07924_),
    .A(net2411));
 sg13g2_inv_1 _12001_ (.Y(_07925_),
    .A(net2400));
 sg13g2_inv_1 _12002_ (.Y(_07926_),
    .A(net2349));
 sg13g2_inv_1 _12003_ (.Y(_07927_),
    .A(net2679));
 sg13g2_inv_1 _12004_ (.Y(_07928_),
    .A(net2765));
 sg13g2_inv_1 _12005_ (.Y(_07929_),
    .A(net2558));
 sg13g2_inv_1 _12006_ (.Y(_07930_),
    .A(net2078));
 sg13g2_inv_1 _12007_ (.Y(_07931_),
    .A(net2382));
 sg13g2_inv_1 _12008_ (.Y(_07932_),
    .A(net2947));
 sg13g2_inv_2 _12009_ (.Y(_07933_),
    .A(net1177));
 sg13g2_inv_1 _12010_ (.Y(_07934_),
    .A(\soc_inst.spi_inst.rx_shift_reg[10] ));
 sg13g2_inv_1 _12011_ (.Y(_07935_),
    .A(\soc_inst.spi_inst.rx_shift_reg[11] ));
 sg13g2_inv_1 _12012_ (.Y(_07936_),
    .A(\soc_inst.spi_inst.rx_shift_reg[13] ));
 sg13g2_inv_1 _12013_ (.Y(_07937_),
    .A(\soc_inst.spi_inst.rx_shift_reg[14] ));
 sg13g2_inv_1 _12014_ (.Y(_07938_),
    .A(\soc_inst.spi_inst.rx_shift_reg[15] ));
 sg13g2_inv_1 _12015_ (.Y(_07939_),
    .A(\soc_inst.spi_inst.rx_shift_reg[24] ));
 sg13g2_inv_1 _12016_ (.Y(_07940_),
    .A(\soc_inst.spi_inst.rx_shift_reg[28] ));
 sg13g2_inv_1 _12017_ (.Y(_07941_),
    .A(\soc_inst.pwm_inst.channel_counter[0][15] ));
 sg13g2_inv_1 _12018_ (.Y(_07942_),
    .A(\soc_inst.pwm_inst.channel_counter[0][12] ));
 sg13g2_inv_1 _12019_ (.Y(_07943_),
    .A(\soc_inst.pwm_inst.channel_counter[0][10] ));
 sg13g2_inv_1 _12020_ (.Y(_07944_),
    .A(\soc_inst.pwm_inst.channel_counter[0][9] ));
 sg13g2_inv_1 _12021_ (.Y(_07945_),
    .A(\soc_inst.pwm_inst.channel_counter[0][8] ));
 sg13g2_inv_1 _12022_ (.Y(_07946_),
    .A(\soc_inst.pwm_inst.channel_counter[0][5] ));
 sg13g2_inv_1 _12023_ (.Y(_07947_),
    .A(\soc_inst.pwm_inst.channel_counter[0][4] ));
 sg13g2_inv_1 _12024_ (.Y(_07948_),
    .A(\soc_inst.pwm_inst.channel_counter[0][3] ));
 sg13g2_inv_2 _12025_ (.Y(_07949_),
    .A(net1105));
 sg13g2_inv_1 _12026_ (.Y(_07950_),
    .A(\soc_inst.mem_ctrl.spi_data_out[0] ));
 sg13g2_inv_1 _12027_ (.Y(_07951_),
    .A(\soc_inst.mem_ctrl.spi_data_out[1] ));
 sg13g2_inv_1 _12028_ (.Y(_07952_),
    .A(\soc_inst.mem_ctrl.spi_data_out[2] ));
 sg13g2_inv_1 _12029_ (.Y(_07953_),
    .A(\soc_inst.mem_ctrl.spi_data_out[5] ));
 sg13g2_inv_1 _12030_ (.Y(_07954_),
    .A(\soc_inst.pwm_inst.channel_duty[0][1] ));
 sg13g2_inv_1 _12031_ (.Y(_07955_),
    .A(net2348));
 sg13g2_inv_1 _12032_ (.Y(_07956_),
    .A(net1560));
 sg13g2_inv_1 _12033_ (.Y(_07957_),
    .A(net2249));
 sg13g2_inv_1 _12034_ (.Y(_07958_),
    .A(net1215));
 sg13g2_inv_1 _12035_ (.Y(_07959_),
    .A(net1730));
 sg13g2_inv_2 _12036_ (.Y(_07960_),
    .A(net1386));
 sg13g2_inv_1 _12037_ (.Y(_07961_),
    .A(net782));
 sg13g2_inv_1 _12038_ (.Y(_07962_),
    .A(\soc_inst.pwm_inst.channel_duty[0][6] ));
 sg13g2_inv_1 _12039_ (.Y(_07963_),
    .A(\soc_inst.pwm_inst.channel_duty[0][7] ));
 sg13g2_inv_1 _12040_ (.Y(_07964_),
    .A(net2601));
 sg13g2_inv_1 _12041_ (.Y(_07965_),
    .A(net2431));
 sg13g2_inv_1 _12042_ (.Y(_07966_),
    .A(net2405));
 sg13g2_inv_1 _12043_ (.Y(_07967_),
    .A(net689));
 sg13g2_inv_1 _12044_ (.Y(_07968_),
    .A(net762));
 sg13g2_inv_1 _12045_ (.Y(_07969_),
    .A(net1114));
 sg13g2_inv_1 _12046_ (.Y(_07970_),
    .A(net468));
 sg13g2_inv_1 _12047_ (.Y(_07971_),
    .A(net615));
 sg13g2_inv_1 _12048_ (.Y(_07972_),
    .A(net822));
 sg13g2_inv_1 _12049_ (.Y(_07973_),
    .A(net774));
 sg13g2_inv_1 _12050_ (.Y(_07974_),
    .A(net945));
 sg13g2_inv_1 _12051_ (.Y(_07975_),
    .A(net558));
 sg13g2_inv_1 _12052_ (.Y(_07976_),
    .A(net1226));
 sg13g2_inv_1 _12053_ (.Y(_07977_),
    .A(net1009));
 sg13g2_inv_1 _12054_ (.Y(_07978_),
    .A(net655));
 sg13g2_inv_1 _12055_ (.Y(_07979_),
    .A(net1065));
 sg13g2_inv_1 _12056_ (.Y(_07980_),
    .A(net1132));
 sg13g2_inv_1 _12057_ (.Y(_07981_),
    .A(net642));
 sg13g2_inv_1 _12058_ (.Y(_07982_),
    .A(net795));
 sg13g2_inv_1 _12059_ (.Y(_07983_),
    .A(net883));
 sg13g2_inv_1 _12060_ (.Y(_07984_),
    .A(net551));
 sg13g2_inv_1 _12061_ (.Y(_07985_),
    .A(net901));
 sg13g2_inv_1 _12062_ (.Y(_07986_),
    .A(net736));
 sg13g2_inv_1 _12063_ (.Y(_07987_),
    .A(net764));
 sg13g2_inv_1 _12064_ (.Y(_07988_),
    .A(net661));
 sg13g2_inv_1 _12065_ (.Y(_07989_),
    .A(net497));
 sg13g2_inv_1 _12066_ (.Y(_07990_),
    .A(net680));
 sg13g2_inv_1 _12067_ (.Y(_07991_),
    .A(net906));
 sg13g2_inv_1 _12068_ (.Y(_07992_),
    .A(net1031));
 sg13g2_inv_1 _12069_ (.Y(_07993_),
    .A(net556));
 sg13g2_inv_1 _12070_ (.Y(_07994_),
    .A(net976));
 sg13g2_inv_1 _12071_ (.Y(_07995_),
    .A(net486));
 sg13g2_inv_1 _12072_ (.Y(_07996_),
    .A(net724));
 sg13g2_inv_1 _12073_ (.Y(_07997_),
    .A(net903));
 sg13g2_inv_1 _12074_ (.Y(_07998_),
    .A(net663));
 sg13g2_inv_1 _12075_ (.Y(_07999_),
    .A(net3195));
 sg13g2_inv_1 _12076_ (.Y(_08000_),
    .A(net1985));
 sg13g2_inv_1 _12077_ (.Y(_08001_),
    .A(net2150));
 sg13g2_inv_1 _12078_ (.Y(_08002_),
    .A(net1967));
 sg13g2_inv_1 _12079_ (.Y(_08003_),
    .A(net3213));
 sg13g2_inv_1 _12080_ (.Y(_08004_),
    .A(net1420));
 sg13g2_inv_1 _12081_ (.Y(_08005_),
    .A(net2706));
 sg13g2_inv_1 _12082_ (.Y(_08006_),
    .A(net1261));
 sg13g2_inv_1 _12083_ (.Y(_08007_),
    .A(net1292));
 sg13g2_inv_1 _12084_ (.Y(_08008_),
    .A(net1216));
 sg13g2_inv_1 _12085_ (.Y(_08009_),
    .A(net2077));
 sg13g2_inv_1 _12086_ (.Y(_08010_),
    .A(net693));
 sg13g2_inv_1 _12087_ (.Y(_08011_),
    .A(net2346));
 sg13g2_inv_1 _12088_ (.Y(_08012_),
    .A(net708));
 sg13g2_inv_1 _12089_ (.Y(_08013_),
    .A(net2510));
 sg13g2_inv_1 _12090_ (.Y(_08014_),
    .A(net516));
 sg13g2_inv_1 _12091_ (.Y(_08015_),
    .A(net2449));
 sg13g2_inv_1 _12092_ (.Y(_08016_),
    .A(net2114));
 sg13g2_inv_1 _12093_ (.Y(_08017_),
    .A(net1966));
 sg13g2_inv_1 _12094_ (.Y(_08018_),
    .A(net2534));
 sg13g2_inv_1 _12095_ (.Y(_08019_),
    .A(net2796));
 sg13g2_inv_1 _12096_ (.Y(_08020_),
    .A(net1576));
 sg13g2_inv_1 _12097_ (.Y(_08021_),
    .A(net2586));
 sg13g2_inv_1 _12098_ (.Y(_08022_),
    .A(net842));
 sg13g2_inv_1 _12099_ (.Y(_08023_),
    .A(net2133));
 sg13g2_inv_1 _12100_ (.Y(_08024_),
    .A(net1181));
 sg13g2_inv_1 _12101_ (.Y(_08025_),
    .A(net2460));
 sg13g2_inv_2 _12102_ (.Y(_08026_),
    .A(net3358));
 sg13g2_inv_2 _12103_ (.Y(_08027_),
    .A(net6520));
 sg13g2_inv_2 _12104_ (.Y(_08028_),
    .A(net6515));
 sg13g2_inv_2 _12105_ (.Y(_08029_),
    .A(net2977));
 sg13g2_inv_2 _12106_ (.Y(_08030_),
    .A(\soc_inst.cpu_core.id_rs1_data[1] ));
 sg13g2_inv_2 _12107_ (.Y(_08031_),
    .A(net2858));
 sg13g2_inv_8 _12108_ (.Y(_08032_),
    .A(net2895));
 sg13g2_inv_4 _12109_ (.A(net2846),
    .Y(_08033_));
 sg13g2_inv_8 _12110_ (.Y(_08034_),
    .A(net2990));
 sg13g2_inv_4 _12111_ (.A(net2532),
    .Y(_08035_));
 sg13g2_inv_8 _12112_ (.Y(_08036_),
    .A(net3039));
 sg13g2_inv_2 _12113_ (.Y(_08037_),
    .A(net3081));
 sg13g2_inv_8 _12114_ (.Y(_08038_),
    .A(net2937));
 sg13g2_inv_4 _12115_ (.A(net2597),
    .Y(_08039_));
 sg13g2_inv_8 _12116_ (.Y(_08040_),
    .A(net2855));
 sg13g2_inv_2 _12117_ (.Y(_08041_),
    .A(net3214));
 sg13g2_inv_4 _12118_ (.A(net2869),
    .Y(_08042_));
 sg13g2_inv_4 _12119_ (.A(net3072),
    .Y(_08043_));
 sg13g2_inv_8 _12120_ (.Y(_08044_),
    .A(net2871));
 sg13g2_inv_4 _12121_ (.A(net2953),
    .Y(_08045_));
 sg13g2_inv_8 _12122_ (.Y(_08046_),
    .A(net2881));
 sg13g2_inv_4 _12123_ (.A(net3020),
    .Y(_08047_));
 sg13g2_inv_4 _12124_ (.A(net2650),
    .Y(_08048_));
 sg13g2_inv_2 _12125_ (.Y(_08049_),
    .A(net3089));
 sg13g2_inv_2 _12126_ (.Y(_08050_),
    .A(net3000));
 sg13g2_inv_4 _12127_ (.A(net2669),
    .Y(_08051_));
 sg13g2_inv_4 _12128_ (.A(net2987),
    .Y(_08052_));
 sg13g2_inv_8 _12129_ (.Y(_08053_),
    .A(net2880));
 sg13g2_inv_2 _12130_ (.Y(_08054_),
    .A(net3170));
 sg13g2_inv_4 _12131_ (.A(net2567),
    .Y(_08055_));
 sg13g2_inv_8 _12132_ (.Y(_08056_),
    .A(net2358));
 sg13g2_inv_2 _12133_ (.Y(_08057_),
    .A(net2711));
 sg13g2_inv_4 _12134_ (.A(net2728),
    .Y(_08058_));
 sg13g2_inv_2 _12135_ (.Y(_08059_),
    .A(\soc_inst.cpu_core.id_rs1_data[29] ));
 sg13g2_inv_2 _12136_ (.Y(_08060_),
    .A(net3123));
 sg13g2_inv_4 _12137_ (.A(net2971),
    .Y(_08061_));
 sg13g2_inv_4 _12138_ (.A(\soc_inst.cpu_core.id_rs2_data[27] ),
    .Y(_08062_));
 sg13g2_inv_1 _12139_ (.Y(_08063_),
    .A(net3250));
 sg13g2_inv_8 _12140_ (.Y(_08064_),
    .A(\soc_inst.cpu_core.id_rs2_data[26] ));
 sg13g2_inv_4 _12141_ (.A(net2912),
    .Y(_08065_));
 sg13g2_inv_1 _12142_ (.Y(_08066_),
    .A(net2852));
 sg13g2_inv_8 _12143_ (.Y(_08067_),
    .A(\soc_inst.cpu_core.id_rs2_data[24] ));
 sg13g2_inv_2 _12144_ (.Y(_08068_),
    .A(net3007));
 sg13g2_inv_4 _12145_ (.A(\soc_inst.cpu_core.id_rs2_data[23] ),
    .Y(_08069_));
 sg13g2_inv_2 _12146_ (.Y(_08070_),
    .A(net2804));
 sg13g2_inv_4 _12147_ (.A(\soc_inst.cpu_core.id_rs2_data[22] ),
    .Y(_08071_));
 sg13g2_inv_8 _12148_ (.Y(_08072_),
    .A(\soc_inst.cpu_core.id_rs2_data[21] ));
 sg13g2_inv_2 _12149_ (.Y(_08073_),
    .A(net2939));
 sg13g2_inv_2 _12150_ (.Y(_08074_),
    .A(net3219));
 sg13g2_inv_8 _12151_ (.Y(_08075_),
    .A(net2802));
 sg13g2_inv_4 _12152_ (.A(net2901),
    .Y(_08076_));
 sg13g2_inv_4 _12153_ (.A(net2956),
    .Y(_08077_));
 sg13g2_inv_2 _12154_ (.Y(_08078_),
    .A(net3059));
 sg13g2_inv_4 _12155_ (.A(net2748),
    .Y(_08079_));
 sg13g2_inv_1 _12156_ (.Y(_08080_),
    .A(net3135));
 sg13g2_inv_8 _12157_ (.Y(_08081_),
    .A(net2750));
 sg13g2_inv_2 _12158_ (.Y(_08082_),
    .A(\soc_inst.cpu_core.id_pc[0] ));
 sg13g2_inv_2 _12159_ (.Y(_08083_),
    .A(\soc_inst.cpu_core.id_pc[1] ));
 sg13g2_inv_1 _12160_ (.Y(_08084_),
    .A(\soc_inst.cpu_core.id_pc[2] ));
 sg13g2_inv_2 _12161_ (.Y(_08085_),
    .A(\soc_inst.cpu_core.id_pc[3] ));
 sg13g2_inv_1 _12162_ (.Y(_08086_),
    .A(net2816));
 sg13g2_inv_2 _12163_ (.Y(_08087_),
    .A(\soc_inst.cpu_core.id_pc[4] ));
 sg13g2_inv_2 _12164_ (.Y(_08088_),
    .A(net2648));
 sg13g2_inv_4 _12165_ (.A(\soc_inst.cpu_core.id_pc[5] ),
    .Y(_08089_));
 sg13g2_inv_1 _12166_ (.Y(_08090_),
    .A(net3086));
 sg13g2_inv_2 _12167_ (.Y(_08091_),
    .A(\soc_inst.cpu_core.id_pc[6] ));
 sg13g2_inv_1 _12168_ (.Y(_08092_),
    .A(net2794));
 sg13g2_inv_2 _12169_ (.Y(_08093_),
    .A(\soc_inst.cpu_core.id_pc[7] ));
 sg13g2_inv_1 _12170_ (.Y(_08094_),
    .A(net2707));
 sg13g2_inv_2 _12171_ (.Y(_08095_),
    .A(\soc_inst.cpu_core.id_pc[8] ));
 sg13g2_inv_1 _12172_ (.Y(_08096_),
    .A(net2426));
 sg13g2_inv_4 _12173_ (.A(\soc_inst.cpu_core.id_pc[9] ),
    .Y(_08097_));
 sg13g2_inv_1 _12174_ (.Y(_08098_),
    .A(net3080));
 sg13g2_inv_2 _12175_ (.Y(_08099_),
    .A(\soc_inst.cpu_core.id_pc[10] ));
 sg13g2_inv_1 _12176_ (.Y(_08100_),
    .A(net2478));
 sg13g2_inv_4 _12177_ (.A(\soc_inst.cpu_core.id_pc[11] ),
    .Y(_08101_));
 sg13g2_inv_1 _12178_ (.Y(_08102_),
    .A(\soc_inst.cpu_core.id_imm[11] ));
 sg13g2_inv_2 _12179_ (.Y(_08103_),
    .A(\soc_inst.cpu_core.id_pc[12] ));
 sg13g2_inv_1 _12180_ (.Y(_08104_),
    .A(\soc_inst.cpu_core.id_imm[12] ));
 sg13g2_inv_1 _12181_ (.Y(_08105_),
    .A(\soc_inst.cpu_core.id_pc[13] ));
 sg13g2_inv_2 _12182_ (.Y(_08106_),
    .A(\soc_inst.cpu_core.id_pc[14] ));
 sg13g2_inv_4 _12183_ (.A(\soc_inst.cpu_core.id_pc[15] ),
    .Y(_08107_));
 sg13g2_inv_2 _12184_ (.Y(_08108_),
    .A(\soc_inst.cpu_core.id_pc[16] ));
 sg13g2_inv_2 _12185_ (.Y(_08109_),
    .A(\soc_inst.cpu_core.id_pc[17] ));
 sg13g2_inv_2 _12186_ (.Y(_08110_),
    .A(\soc_inst.cpu_core.id_pc[18] ));
 sg13g2_inv_1 _12187_ (.Y(_08111_),
    .A(\soc_inst.cpu_core.id_pc[19] ));
 sg13g2_inv_2 _12188_ (.Y(_08112_),
    .A(\soc_inst.cpu_core.id_pc[20] ));
 sg13g2_inv_4 _12189_ (.A(\soc_inst.cpu_core.id_pc[21] ),
    .Y(_08113_));
 sg13g2_inv_1 _12190_ (.Y(_08114_),
    .A(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_inv_2 _12191_ (.Y(_08115_),
    .A(net3410));
 sg13g2_inv_4 _12192_ (.A(net2628),
    .Y(_08116_));
 sg13g2_inv_1 _12193_ (.Y(_08117_),
    .A(\soc_inst.cpu_core.id_imm[27] ));
 sg13g2_inv_1 _12194_ (.Y(_08118_),
    .A(net2876));
 sg13g2_inv_1 _12195_ (.Y(_08119_),
    .A(net2910));
 sg13g2_inv_1 _12196_ (.Y(_08120_),
    .A(net2446));
 sg13g2_inv_1 _12197_ (.Y(_08121_),
    .A(net2818));
 sg13g2_inv_1 _12198_ (.Y(_08122_),
    .A(net2859));
 sg13g2_inv_1 _12199_ (.Y(_08123_),
    .A(net3034));
 sg13g2_inv_1 _12200_ (.Y(_08124_),
    .A(net2476));
 sg13g2_inv_1 _12201_ (.Y(_08125_),
    .A(net2441));
 sg13g2_inv_2 _12202_ (.Y(_08126_),
    .A(net2719));
 sg13g2_inv_1 _12203_ (.Y(_08127_),
    .A(net2754));
 sg13g2_inv_2 _12204_ (.Y(_08128_),
    .A(net2830));
 sg13g2_inv_1 _12205_ (.Y(_08129_),
    .A(net2238));
 sg13g2_inv_2 _12206_ (.Y(_08130_),
    .A(net1251));
 sg13g2_inv_2 _12207_ (.Y(_08131_),
    .A(net6430));
 sg13g2_inv_1 _12208_ (.Y(_08132_),
    .A(net6436));
 sg13g2_inv_1 _12209_ (.Y(_08133_),
    .A(net6452));
 sg13g2_inv_1 _12210_ (.Y(_08134_),
    .A(net2924));
 sg13g2_inv_2 _12211_ (.Y(_08135_),
    .A(net6441));
 sg13g2_inv_1 _12212_ (.Y(_08136_),
    .A(net1672));
 sg13g2_inv_1 _12213_ (.Y(_08137_),
    .A(net2368));
 sg13g2_inv_1 _12214_ (.Y(_08138_),
    .A(net2356));
 sg13g2_inv_1 _12215_ (.Y(_08139_),
    .A(net1923));
 sg13g2_inv_1 _12216_ (.Y(_08140_),
    .A(net2219));
 sg13g2_inv_1 _12217_ (.Y(_08141_),
    .A(net1268));
 sg13g2_inv_1 _12218_ (.Y(_08142_),
    .A(net1384));
 sg13g2_inv_1 _12219_ (.Y(_08143_),
    .A(net1697));
 sg13g2_inv_1 _12220_ (.Y(_08144_),
    .A(net1881));
 sg13g2_inv_1 _12221_ (.Y(_08145_),
    .A(net2102));
 sg13g2_inv_1 _12222_ (.Y(_08146_),
    .A(net1401));
 sg13g2_inv_1 _12223_ (.Y(_08147_),
    .A(net2292));
 sg13g2_inv_1 _12224_ (.Y(_08148_),
    .A(net1453));
 sg13g2_inv_1 _12225_ (.Y(_08149_),
    .A(net1867));
 sg13g2_inv_1 _12226_ (.Y(_08150_),
    .A(net1382));
 sg13g2_inv_1 _12227_ (.Y(_08151_),
    .A(net1822));
 sg13g2_inv_1 _12228_ (.Y(_08152_),
    .A(net2231));
 sg13g2_inv_1 _12229_ (.Y(_08153_),
    .A(net1778));
 sg13g2_inv_1 _12230_ (.Y(_08154_),
    .A(net2643));
 sg13g2_inv_1 _12231_ (.Y(_08155_),
    .A(net1764));
 sg13g2_inv_1 _12232_ (.Y(_08156_),
    .A(net1562));
 sg13g2_inv_1 _12233_ (.Y(_08157_),
    .A(net1801));
 sg13g2_inv_1 _12234_ (.Y(_08158_),
    .A(net1853));
 sg13g2_inv_1 _12235_ (.Y(_08159_),
    .A(net1668));
 sg13g2_inv_1 _12236_ (.Y(_08160_),
    .A(net3266));
 sg13g2_inv_1 _12237_ (.Y(_08161_),
    .A(net3279));
 sg13g2_inv_1 _12238_ (.Y(_08162_),
    .A(net3110));
 sg13g2_inv_1 _12239_ (.Y(_08163_),
    .A(net2938));
 sg13g2_inv_1 _12240_ (.Y(_08164_),
    .A(net2900));
 sg13g2_inv_1 _12241_ (.Y(_08165_),
    .A(net2656));
 sg13g2_inv_4 _12242_ (.A(net3215),
    .Y(_08166_));
 sg13g2_inv_4 _12243_ (.A(net3160),
    .Y(_08167_));
 sg13g2_inv_4 _12244_ (.A(net3208),
    .Y(_08168_));
 sg13g2_inv_1 _12245_ (.Y(_08169_),
    .A(net3210));
 sg13g2_inv_1 _12246_ (.Y(_08170_),
    .A(net2800));
 sg13g2_inv_1 _12247_ (.Y(_08171_),
    .A(net3287));
 sg13g2_inv_1 _12248_ (.Y(_08172_),
    .A(net3289));
 sg13g2_inv_4 _12249_ (.A(\soc_inst.cpu_core.ex_instr[15] ),
    .Y(_08173_));
 sg13g2_inv_1 _12250_ (.Y(_08174_),
    .A(net3212));
 sg13g2_inv_2 _12251_ (.Y(_08175_),
    .A(net1158));
 sg13g2_inv_2 _12252_ (.Y(_08176_),
    .A(net603));
 sg13g2_inv_1 _12253_ (.Y(_08177_),
    .A(net1281));
 sg13g2_inv_2 _12254_ (.Y(_08178_),
    .A(net2523));
 sg13g2_inv_2 _12255_ (.Y(_08179_),
    .A(net917));
 sg13g2_inv_1 _12256_ (.Y(_08180_),
    .A(net2681));
 sg13g2_inv_1 _12257_ (.Y(_08181_),
    .A(net2617));
 sg13g2_inv_1 _12258_ (.Y(_08182_),
    .A(net2469));
 sg13g2_inv_1 _12259_ (.Y(_08183_),
    .A(net2414));
 sg13g2_inv_4 _12260_ (.A(\soc_inst.cpu_core.ex_alu_result[31] ),
    .Y(_08184_));
 sg13g2_inv_1 _12261_ (.Y(_08185_),
    .A(net1904));
 sg13g2_inv_1 _12262_ (.Y(_08186_),
    .A(\soc_inst.spi_inst.spi_mosi ));
 sg13g2_inv_1 _12263_ (.Y(_08187_),
    .A(net2975));
 sg13g2_inv_1 _12264_ (.Y(_08188_),
    .A(\soc_inst.cpu_core.alu.a[30] ));
 sg13g2_inv_1 _12265_ (.Y(_08189_),
    .A(net3171));
 sg13g2_inv_1 _12266_ (.Y(_08190_),
    .A(net2605));
 sg13g2_inv_1 _12267_ (.Y(_08191_),
    .A(net2072));
 sg13g2_inv_1 _12268_ (.Y(_08192_),
    .A(net2678));
 sg13g2_inv_1 _12269_ (.Y(_08193_),
    .A(net2557));
 sg13g2_inv_1 _12270_ (.Y(_08194_),
    .A(net3003));
 sg13g2_inv_2 _12271_ (.Y(_08195_),
    .A(net6279));
 sg13g2_inv_1 _12272_ (.Y(_08196_),
    .A(net6281));
 sg13g2_inv_1 _12273_ (.Y(_08197_),
    .A(\soc_inst.cpu_core.alu.b[15] ));
 sg13g2_inv_1 _12274_ (.Y(_08198_),
    .A(net6283));
 sg13g2_inv_1 _12275_ (.Y(_08199_),
    .A(\soc_inst.cpu_core.alu.b[13] ));
 sg13g2_inv_1 _12276_ (.Y(_08200_),
    .A(\soc_inst.cpu_core.alu.a[13] ));
 sg13g2_inv_2 _12277_ (.Y(_08201_),
    .A(net3290));
 sg13g2_inv_1 _12278_ (.Y(_08202_),
    .A(net2828));
 sg13g2_inv_1 _12279_ (.Y(_08203_),
    .A(\soc_inst.cpu_core.alu.a[10] ));
 sg13g2_inv_2 _12280_ (.Y(_08204_),
    .A(\soc_inst.cpu_core.alu.a[9] ));
 sg13g2_inv_2 _12281_ (.Y(_08205_),
    .A(net2923));
 sg13g2_inv_2 _12282_ (.Y(_08206_),
    .A(net6222));
 sg13g2_inv_2 _12283_ (.Y(_08207_),
    .A(net6231));
 sg13g2_inv_1 _12284_ (.Y(_08208_),
    .A(net6238));
 sg13g2_inv_1 _12285_ (.Y(_08209_),
    .A(\soc_inst.cpu_core.alu.a[2] ));
 sg13g2_inv_1 _12286_ (.Y(_08210_),
    .A(net6244));
 sg13g2_inv_1 _12287_ (.Y(_08211_),
    .A(net6254));
 sg13g2_inv_1 _12288_ (.Y(_08212_),
    .A(net605));
 sg13g2_inv_1 _12289_ (.Y(_08213_),
    .A(net352));
 sg13g2_inv_1 _12290_ (.Y(_08214_),
    .A(net376));
 sg13g2_inv_1 _12291_ (.Y(_08215_),
    .A(net309));
 sg13g2_inv_1 _12292_ (.Y(_08216_),
    .A(net379));
 sg13g2_inv_1 _12293_ (.Y(_08217_),
    .A(net701));
 sg13g2_inv_1 _12294_ (.Y(_08218_),
    .A(net431));
 sg13g2_inv_1 _12295_ (.Y(_08219_),
    .A(net898));
 sg13g2_inv_1 _12296_ (.Y(_08220_),
    .A(net342));
 sg13g2_inv_1 _12297_ (.Y(_08221_),
    .A(net2991));
 sg13g2_inv_1 _12298_ (.Y(_08222_),
    .A(net2862));
 sg13g2_nand2_1 _12299_ (.Y(_08223_),
    .A(net6179),
    .B(\soc_inst.mem_ctrl.spi_done ));
 sg13g2_nor4_2 _12300_ (.A(\soc_inst.core_mem_addr[25] ),
    .B(\soc_inst.core_mem_addr[24] ),
    .C(\soc_inst.core_mem_addr[27] ),
    .Y(_08224_),
    .D(\soc_inst.core_mem_addr[26] ));
 sg13g2_nor3_1 _12301_ (.A(\soc_inst.core_mem_addr[29] ),
    .B(\soc_inst.core_mem_addr[28] ),
    .C(\soc_inst.core_mem_addr[31] ),
    .Y(_08225_));
 sg13g2_nand3_1 _12302_ (.B(_08224_),
    .C(_08225_),
    .A(\soc_inst.core_mem_addr[30] ),
    .Y(_08226_));
 sg13g2_nor3_1 _12303_ (.A(\soc_inst.core_mem_addr[8] ),
    .B(\soc_inst.core_mem_addr[9] ),
    .C(\soc_inst.core_mem_addr[10] ),
    .Y(_08227_));
 sg13g2_nand3_1 _12304_ (.B(_07814_),
    .C(_08227_),
    .A(_07812_),
    .Y(_08228_));
 sg13g2_nor4_2 _12305_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(_07815_),
    .C(_08226_),
    .Y(_08229_),
    .D(_08228_));
 sg13g2_nor3_2 _12306_ (.A(net3263),
    .B(_08226_),
    .C(_08228_),
    .Y(_08230_));
 sg13g2_inv_1 _12307_ (.Y(_08231_),
    .A(_08230_));
 sg13g2_or2_1 _12308_ (.X(_08232_),
    .B(_08230_),
    .A(_08229_));
 sg13g2_nor4_1 _12309_ (.A(\soc_inst.core_mem_addr[21] ),
    .B(\soc_inst.core_mem_addr[20] ),
    .C(\soc_inst.core_mem_addr[23] ),
    .D(\soc_inst.core_mem_addr[22] ),
    .Y(_08233_));
 sg13g2_nor4_1 _12310_ (.A(\soc_inst.core_mem_addr[17] ),
    .B(\soc_inst.core_mem_addr[16] ),
    .C(\soc_inst.core_mem_addr[19] ),
    .D(\soc_inst.core_mem_addr[18] ),
    .Y(_08234_));
 sg13g2_and2_1 _12311_ (.A(_08233_),
    .B(_08234_),
    .X(_08235_));
 sg13g2_or2_1 _12312_ (.X(_08236_),
    .B(net6205),
    .A(net6212));
 sg13g2_nor2_1 _12313_ (.A(\soc_inst.core_mem_addr[14] ),
    .B(_08226_),
    .Y(_08237_));
 sg13g2_nor3_1 _12314_ (.A(\soc_inst.core_mem_addr[14] ),
    .B(_08226_),
    .C(_08228_),
    .Y(_08238_));
 sg13g2_o21ai_1 _12315_ (.B1(_08235_),
    .Y(_08239_),
    .A1(_08229_),
    .A2(_08238_));
 sg13g2_nor2b_2 _12316_ (.A(_08239_),
    .B_N(_08236_),
    .Y(_08240_));
 sg13g2_nand3_1 _12317_ (.B(_08235_),
    .C(_08236_),
    .A(_08232_),
    .Y(_08241_));
 sg13g2_o21ai_1 _12318_ (.B1(net5188),
    .Y(_08242_),
    .A1(net6504),
    .A2(_08223_));
 sg13g2_nand2_1 _12319_ (.Y(_08243_),
    .A(net1222),
    .B(net5197));
 sg13g2_nor2_2 _12320_ (.A(\soc_inst.core_mem_re ),
    .B(net1438),
    .Y(_08244_));
 sg13g2_nor2_2 _12321_ (.A(net6205),
    .B(net6507),
    .Y(_08245_));
 sg13g2_nand2_2 _12322_ (.Y(_08246_),
    .A(_08244_),
    .B(_08245_));
 sg13g2_a21oi_2 _12323_ (.B1(_07816_),
    .Y(_08247_),
    .A2(_08245_),
    .A1(_08244_));
 sg13g2_nand2_2 _12324_ (.Y(_08248_),
    .A(net6504),
    .B(_08246_));
 sg13g2_nor2_2 _12325_ (.A(net5194),
    .B(_08247_),
    .Y(_08249_));
 sg13g2_nand2_2 _12326_ (.Y(_08250_),
    .A(net5190),
    .B(_08248_));
 sg13g2_xor2_1 _12327_ (.B(\soc_inst.core_instr_addr[21] ),
    .A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .X(_08251_));
 sg13g2_xor2_1 _12328_ (.B(\soc_inst.core_instr_addr[10] ),
    .A(\soc_inst.mem_ctrl.spi_addr[10] ),
    .X(_08252_));
 sg13g2_xor2_1 _12329_ (.B(\soc_inst.core_instr_addr[5] ),
    .A(\soc_inst.mem_ctrl.spi_addr[5] ),
    .X(_08253_));
 sg13g2_xor2_1 _12330_ (.B(\soc_inst.core_instr_addr[4] ),
    .A(\soc_inst.mem_ctrl.spi_addr[4] ),
    .X(_08254_));
 sg13g2_xor2_1 _12331_ (.B(\soc_inst.core_instr_addr[12] ),
    .A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .X(_08255_));
 sg13g2_xor2_1 _12332_ (.B(\soc_inst.core_instr_addr[7] ),
    .A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .X(_08256_));
 sg13g2_xor2_1 _12333_ (.B(\soc_inst.core_instr_addr[3] ),
    .A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .X(_08257_));
 sg13g2_inv_1 _12334_ (.Y(_08258_),
    .A(_08257_));
 sg13g2_xor2_1 _12335_ (.B(\soc_inst.core_instr_addr[15] ),
    .A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .X(_08259_));
 sg13g2_xor2_1 _12336_ (.B(\soc_inst.core_instr_addr[13] ),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .X(_08260_));
 sg13g2_xor2_1 _12337_ (.B(\soc_inst.core_instr_addr[1] ),
    .A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(_08261_));
 sg13g2_xnor2_1 _12338_ (.Y(_08262_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .B(\soc_inst.core_instr_addr[2] ));
 sg13g2_xor2_1 _12339_ (.B(\soc_inst.core_instr_addr[23] ),
    .A(\soc_inst.mem_ctrl.spi_addr[23] ),
    .X(_08263_));
 sg13g2_a21oi_1 _12340_ (.A1(_07861_),
    .A2(\soc_inst.core_instr_addr[22] ),
    .Y(_08264_),
    .B1(_08263_));
 sg13g2_nand2_1 _12341_ (.Y(_08265_),
    .A(\soc_inst.mem_ctrl.spi_addr[22] ),
    .B(_07862_));
 sg13g2_xnor2_1 _12342_ (.Y(_08266_),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .B(\soc_inst.core_instr_addr[9] ));
 sg13g2_xnor2_1 _12343_ (.Y(_08267_),
    .A(\soc_inst.mem_ctrl.spi_addr[8] ),
    .B(\soc_inst.core_instr_addr[8] ));
 sg13g2_xnor2_1 _12344_ (.Y(_08268_),
    .A(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .B(\soc_inst.core_instr_addr[0] ));
 sg13g2_xnor2_1 _12345_ (.Y(_08269_),
    .A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .B(\soc_inst.core_instr_addr[19] ));
 sg13g2_xor2_1 _12346_ (.B(\soc_inst.core_instr_addr[18] ),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .X(_08270_));
 sg13g2_inv_2 _12347_ (.Y(_08271_),
    .A(_08270_));
 sg13g2_xor2_1 _12348_ (.B(\soc_inst.core_instr_addr[17] ),
    .A(\soc_inst.mem_ctrl.spi_addr[17] ),
    .X(_08272_));
 sg13g2_xor2_1 _12349_ (.B(\soc_inst.core_instr_addr[11] ),
    .A(\soc_inst.mem_ctrl.spi_addr[11] ),
    .X(_08273_));
 sg13g2_xor2_1 _12350_ (.B(\soc_inst.core_instr_addr[20] ),
    .A(\soc_inst.mem_ctrl.spi_addr[20] ),
    .X(_08274_));
 sg13g2_xor2_1 _12351_ (.B(\soc_inst.core_instr_addr[16] ),
    .A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .X(_08275_));
 sg13g2_xor2_1 _12352_ (.B(\soc_inst.core_instr_addr[14] ),
    .A(\soc_inst.mem_ctrl.spi_addr[14] ),
    .X(_08276_));
 sg13g2_xnor2_1 _12353_ (.Y(_08277_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(\soc_inst.core_instr_addr[6] ));
 sg13g2_nor2b_1 _12354_ (.A(_08253_),
    .B_N(_08277_),
    .Y(_08278_));
 sg13g2_nor2_1 _12355_ (.A(_08252_),
    .B(_08256_),
    .Y(_08279_));
 sg13g2_nand2_1 _12356_ (.Y(_08280_),
    .A(_08269_),
    .B(_08279_));
 sg13g2_nor4_1 _12357_ (.A(_08257_),
    .B(_08259_),
    .C(_08261_),
    .D(_08276_),
    .Y(_08281_));
 sg13g2_nor3_1 _12358_ (.A(_08251_),
    .B(_08272_),
    .C(_08274_),
    .Y(_08282_));
 sg13g2_nand3_1 _12359_ (.B(_08281_),
    .C(_08282_),
    .A(_08262_),
    .Y(_08283_));
 sg13g2_or2_1 _12360_ (.X(_08284_),
    .B(_08283_),
    .A(_08280_));
 sg13g2_nand4_1 _12361_ (.B(_08265_),
    .C(_08267_),
    .A(_08264_),
    .Y(_08285_),
    .D(_08278_));
 sg13g2_nor4_1 _12362_ (.A(_08254_),
    .B(_08255_),
    .C(_08273_),
    .D(_08275_),
    .Y(_08286_));
 sg13g2_nor2b_1 _12363_ (.A(_08260_),
    .B_N(_08266_),
    .Y(_08287_));
 sg13g2_nand4_1 _12364_ (.B(_08271_),
    .C(_08286_),
    .A(_08268_),
    .Y(_08288_),
    .D(_08287_));
 sg13g2_nor3_2 _12365_ (.A(_08284_),
    .B(_08285_),
    .C(_08288_),
    .Y(_08289_));
 sg13g2_nand2_2 _12366_ (.Y(_08290_),
    .A(net3148),
    .B(_08289_));
 sg13g2_nor2_1 _12367_ (.A(net1222),
    .B(_08246_),
    .Y(_08291_));
 sg13g2_nor2_1 _12368_ (.A(_08246_),
    .B(_08290_),
    .Y(_08292_));
 sg13g2_nor3_2 _12369_ (.A(net1222),
    .B(_08246_),
    .C(_08290_),
    .Y(_08293_));
 sg13g2_a221oi_1 _12370_ (.B2(net2751),
    .C1(_08293_),
    .B1(_08249_),
    .A1(_08242_),
    .Y(_00320_),
    .A2(_08243_));
 sg13g2_nor2_1 _12371_ (.A(net1568),
    .B(_00251_),
    .Y(_08294_));
 sg13g2_nor3_1 _12372_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(net6543),
    .C(net1569),
    .Y(_00319_));
 sg13g2_a22oi_1 _12373_ (.Y(_08295_),
    .B1(net703),
    .B2(net2505),
    .A2(net2783),
    .A1(net978));
 sg13g2_nand2_1 _12374_ (.Y(_08296_),
    .A(net290),
    .B(net2466));
 sg13g2_a22oi_1 _12375_ (.Y(_08297_),
    .B1(net3339),
    .B2(net2536),
    .A2(net2782),
    .A1(\soc_inst.gpio_inst.int_pend_reg[3] ));
 sg13g2_a22oi_1 _12376_ (.Y(_08298_),
    .B1(net407),
    .B2(net2499),
    .A2(net2898),
    .A1(net428));
 sg13g2_nand4_1 _12377_ (.B(_08296_),
    .C(net3340),
    .A(_08295_),
    .Y(_00088_),
    .D(_08298_));
 sg13g2_a21o_2 _12378_ (.A2(net6533),
    .A1(net6532),
    .B1(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(_08299_));
 sg13g2_nand3_1 _12379_ (.B(\soc_inst.mem_ctrl.spi_addr[3] ),
    .C(_08299_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .Y(_08300_));
 sg13g2_nand4_1 _12380_ (.B(\soc_inst.mem_ctrl.spi_addr[3] ),
    .C(\soc_inst.mem_ctrl.spi_addr[4] ),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .Y(_08301_),
    .D(_08299_));
 sg13g2_nor2_2 _12381_ (.A(_07827_),
    .B(_08301_),
    .Y(_08302_));
 sg13g2_nand2_1 _12382_ (.Y(_08303_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(_08302_));
 sg13g2_nand3_1 _12383_ (.B(\soc_inst.mem_ctrl.spi_addr[7] ),
    .C(_08302_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .Y(_08304_));
 sg13g2_and4_1 _12384_ (.A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(\soc_inst.mem_ctrl.spi_addr[7] ),
    .C(\soc_inst.mem_ctrl.spi_addr[8] ),
    .D(_08302_),
    .X(_08305_));
 sg13g2_nand2_1 _12385_ (.Y(_08306_),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .B(_08305_));
 sg13g2_nand3_1 _12386_ (.B(\soc_inst.mem_ctrl.spi_addr[10] ),
    .C(_08305_),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .Y(_08307_));
 sg13g2_and4_1 _12387_ (.A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .B(\soc_inst.mem_ctrl.spi_addr[10] ),
    .C(\soc_inst.mem_ctrl.spi_addr[11] ),
    .D(_08305_),
    .X(_08308_));
 sg13g2_and2_1 _12388_ (.A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .B(_08308_),
    .X(_08309_));
 sg13g2_nand2_1 _12389_ (.Y(_08310_),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .B(_08309_));
 sg13g2_nand3_1 _12390_ (.B(\soc_inst.mem_ctrl.spi_addr[14] ),
    .C(_08309_),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .Y(_08311_));
 sg13g2_nand4_1 _12391_ (.B(\soc_inst.mem_ctrl.spi_addr[14] ),
    .C(\soc_inst.mem_ctrl.spi_addr[15] ),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .Y(_08312_),
    .D(_08309_));
 sg13g2_or2_1 _12392_ (.X(_08313_),
    .B(_08312_),
    .A(_07849_));
 sg13g2_nor2_2 _12393_ (.A(_07851_),
    .B(_08313_),
    .Y(_08314_));
 sg13g2_nand3_1 _12394_ (.B(\soc_inst.mem_ctrl.spi_addr[19] ),
    .C(_08314_),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .Y(_08315_));
 sg13g2_and4_1 _12395_ (.A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .B(\soc_inst.mem_ctrl.spi_addr[19] ),
    .C(\soc_inst.mem_ctrl.spi_addr[20] ),
    .D(_08314_),
    .X(_08316_));
 sg13g2_nand2_1 _12396_ (.Y(_08317_),
    .A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .B(_08316_));
 sg13g2_o21ai_1 _12397_ (.B1(_08265_),
    .Y(_08318_),
    .A1(_08263_),
    .A2(_08317_));
 sg13g2_or2_1 _12398_ (.X(_08319_),
    .B(_08318_),
    .A(_08264_));
 sg13g2_o21ai_1 _12399_ (.B1(_08318_),
    .Y(_08320_),
    .A1(_08264_),
    .A2(_08317_));
 sg13g2_xnor2_1 _12400_ (.Y(_08321_),
    .A(_08251_),
    .B(_08316_));
 sg13g2_xnor2_1 _12401_ (.Y(_08322_),
    .A(_08274_),
    .B(_08315_));
 sg13g2_and3_1 _12402_ (.X(_08323_),
    .A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .B(_08269_),
    .C(_08314_));
 sg13g2_a21oi_1 _12403_ (.A1(\soc_inst.mem_ctrl.spi_addr[18] ),
    .A2(_08314_),
    .Y(_08324_),
    .B1(_08269_));
 sg13g2_or2_1 _12404_ (.X(_08325_),
    .B(_08324_),
    .A(_08323_));
 sg13g2_xnor2_1 _12405_ (.Y(_08326_),
    .A(_08271_),
    .B(_08314_));
 sg13g2_or2_1 _12406_ (.X(_08327_),
    .B(_08313_),
    .A(_08272_));
 sg13g2_nand2_1 _12407_ (.Y(_08328_),
    .A(_08272_),
    .B(_08313_));
 sg13g2_and2_1 _12408_ (.A(_08327_),
    .B(_08328_),
    .X(_08329_));
 sg13g2_xor2_1 _12409_ (.B(_08312_),
    .A(_08275_),
    .X(_08330_));
 sg13g2_xor2_1 _12410_ (.B(_08311_),
    .A(_08259_),
    .X(_08331_));
 sg13g2_and2_1 _12411_ (.A(_08276_),
    .B(_08310_),
    .X(_08332_));
 sg13g2_nand2_1 _12412_ (.Y(_08333_),
    .A(_08276_),
    .B(_08310_));
 sg13g2_o21ai_1 _12413_ (.B1(_08260_),
    .Y(_08334_),
    .A1(_07843_),
    .A2(_08276_));
 sg13g2_mux2_1 _12414_ (.A0(_08260_),
    .A1(_08334_),
    .S(_08309_),
    .X(_08335_));
 sg13g2_xor2_1 _12415_ (.B(_08308_),
    .A(_08255_),
    .X(_08336_));
 sg13g2_xor2_1 _12416_ (.B(_08305_),
    .A(_08266_),
    .X(_08337_));
 sg13g2_o21ai_1 _12417_ (.B1(_08252_),
    .Y(_08338_),
    .A1(\soc_inst.core_instr_addr[10] ),
    .A2(_08273_));
 sg13g2_nand3_1 _12418_ (.B(_08305_),
    .C(_08338_),
    .A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .Y(_08339_));
 sg13g2_nand2_1 _12419_ (.Y(_08340_),
    .A(_08252_),
    .B(_08306_));
 sg13g2_nand3_1 _12420_ (.B(_08339_),
    .C(_08340_),
    .A(_08337_),
    .Y(_08341_));
 sg13g2_and2_1 _12421_ (.A(_08273_),
    .B(_08307_),
    .X(_08342_));
 sg13g2_and3_1 _12422_ (.X(_08343_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .B(_08258_),
    .C(_08299_));
 sg13g2_a21oi_1 _12423_ (.A1(\soc_inst.mem_ctrl.spi_addr[2] ),
    .A2(_08299_),
    .Y(_08344_),
    .B1(_08258_));
 sg13g2_nand3_1 _12424_ (.B(net6533),
    .C(_08261_),
    .A(net6532),
    .Y(_08345_));
 sg13g2_nand2_1 _12425_ (.Y(_08346_),
    .A(_08268_),
    .B(_08345_));
 sg13g2_nor3_1 _12426_ (.A(_08343_),
    .B(_08344_),
    .C(_08346_),
    .Y(_08347_));
 sg13g2_o21ai_1 _12427_ (.B1(_08347_),
    .Y(_08348_),
    .A1(_08253_),
    .A2(_08301_));
 sg13g2_a221oi_1 _12428_ (.B2(_08256_),
    .C1(_08348_),
    .B1(_08303_),
    .A1(_08253_),
    .Y(_08349_),
    .A2(_08301_));
 sg13g2_o21ai_1 _12429_ (.B1(_08349_),
    .Y(_08350_),
    .A1(_08256_),
    .A2(_08303_));
 sg13g2_nand2b_1 _12430_ (.Y(_08351_),
    .B(_08267_),
    .A_N(_08304_));
 sg13g2_nand2b_1 _12431_ (.Y(_08352_),
    .B(_08304_),
    .A_N(_08267_));
 sg13g2_and2_1 _12432_ (.A(_08277_),
    .B(_08302_),
    .X(_08353_));
 sg13g2_a21o_1 _12433_ (.A2(net6533),
    .A1(net6532),
    .B1(_08261_),
    .X(_08354_));
 sg13g2_o21ai_1 _12434_ (.B1(_08354_),
    .Y(_08355_),
    .A1(_08262_),
    .A2(_08299_));
 sg13g2_a21oi_1 _12435_ (.A1(_08262_),
    .A2(_08299_),
    .Y(_08356_),
    .B1(_08355_));
 sg13g2_o21ai_1 _12436_ (.B1(_08356_),
    .Y(_08357_),
    .A1(_08254_),
    .A2(_08300_));
 sg13g2_a21oi_1 _12437_ (.A1(_08254_),
    .A2(_08300_),
    .Y(_08358_),
    .B1(_08357_));
 sg13g2_o21ai_1 _12438_ (.B1(_08358_),
    .Y(_08359_),
    .A1(_08277_),
    .A2(_08302_));
 sg13g2_nor2_1 _12439_ (.A(_08353_),
    .B(_08359_),
    .Y(_08360_));
 sg13g2_nand3_1 _12440_ (.B(_08352_),
    .C(_08360_),
    .A(_08351_),
    .Y(_08361_));
 sg13g2_or4_1 _12441_ (.A(_08341_),
    .B(_08342_),
    .C(_08350_),
    .D(_08361_),
    .X(_08362_));
 sg13g2_nor4_1 _12442_ (.A(_08332_),
    .B(_08335_),
    .C(_08336_),
    .D(_08362_),
    .Y(_08363_));
 sg13g2_nand4_1 _12443_ (.B(_08330_),
    .C(_08331_),
    .A(_08329_),
    .Y(_08364_),
    .D(_08363_));
 sg13g2_nor4_1 _12444_ (.A(_08322_),
    .B(_08325_),
    .C(_08326_),
    .D(_08364_),
    .Y(_08365_));
 sg13g2_and4_1 _12445_ (.A(_08319_),
    .B(_08320_),
    .C(_08321_),
    .D(_08365_),
    .X(_08366_));
 sg13g2_xnor2_1 _12446_ (.Y(_08367_),
    .A(_08262_),
    .B(_08299_));
 sg13g2_xor2_1 _12447_ (.B(_08303_),
    .A(_08256_),
    .X(_08368_));
 sg13g2_xnor2_1 _12448_ (.Y(_08369_),
    .A(_08254_),
    .B(_08300_));
 sg13g2_nand3_1 _12449_ (.B(_08345_),
    .C(_08354_),
    .A(_08268_),
    .Y(_08370_));
 sg13g2_nor4_1 _12450_ (.A(_08343_),
    .B(_08344_),
    .C(_08369_),
    .D(_08370_),
    .Y(_08371_));
 sg13g2_o21ai_1 _12451_ (.B1(_08371_),
    .Y(_08372_),
    .A1(_08277_),
    .A2(_08302_));
 sg13g2_xnor2_1 _12452_ (.Y(_08373_),
    .A(_08253_),
    .B(_08301_));
 sg13g2_nor4_1 _12453_ (.A(_08353_),
    .B(_08367_),
    .C(_08372_),
    .D(_08373_),
    .Y(_08374_));
 sg13g2_nand4_1 _12454_ (.B(_08352_),
    .C(_08368_),
    .A(_08351_),
    .Y(_08375_),
    .D(_08374_));
 sg13g2_nor4_1 _12455_ (.A(_08336_),
    .B(_08341_),
    .C(_08342_),
    .D(_08375_),
    .Y(_08376_));
 sg13g2_nor2b_1 _12456_ (.A(_08335_),
    .B_N(_08376_),
    .Y(_08377_));
 sg13g2_and4_1 _12457_ (.A(_08327_),
    .B(_08331_),
    .C(_08333_),
    .D(_08377_),
    .X(_08378_));
 sg13g2_nand3_1 _12458_ (.B(_08330_),
    .C(_08378_),
    .A(_08328_),
    .Y(_08379_));
 sg13g2_a21oi_1 _12459_ (.A1(_08274_),
    .A2(_08315_),
    .Y(_08380_),
    .B1(_08379_));
 sg13g2_o21ai_1 _12460_ (.B1(_08380_),
    .Y(_08381_),
    .A1(_08274_),
    .A2(_08315_));
 sg13g2_nor4_1 _12461_ (.A(_08323_),
    .B(_08324_),
    .C(_08326_),
    .D(_08381_),
    .Y(_08382_));
 sg13g2_nand4_1 _12462_ (.B(_08320_),
    .C(_08321_),
    .A(_08319_),
    .Y(_08383_),
    .D(_08382_));
 sg13g2_nor2_2 _12463_ (.A(_08289_),
    .B(_08366_),
    .Y(_08384_));
 sg13g2_nand2_2 _12464_ (.Y(_08385_),
    .A(net6194),
    .B(_08384_));
 sg13g2_nor3_1 _12465_ (.A(_07866_),
    .B(_08289_),
    .C(_08366_),
    .Y(_08386_));
 sg13g2_nand2b_1 _12466_ (.Y(_08387_),
    .B(_08249_),
    .A_N(_08386_));
 sg13g2_o21ai_1 _12467_ (.B1(_08387_),
    .Y(_08388_),
    .A1(net2751),
    .A2(net5190));
 sg13g2_o21ai_1 _12468_ (.B1(_08388_),
    .Y(_00009_),
    .A1(_08250_),
    .A2(_08385_));
 sg13g2_a21oi_1 _12469_ (.A1(_08244_),
    .A2(_08245_),
    .Y(_08389_),
    .B1(net1222));
 sg13g2_inv_1 _12470_ (.Y(_08390_),
    .A(_08389_));
 sg13g2_nand2b_1 _12471_ (.Y(_08391_),
    .B(net6179),
    .A_N(net3281));
 sg13g2_nor2_1 _12472_ (.A(_08247_),
    .B(_08391_),
    .Y(_08392_));
 sg13g2_a221oi_1 _12473_ (.B2(_08291_),
    .C1(_08392_),
    .B1(_08290_),
    .A1(net6179),
    .Y(_08393_),
    .A2(net5194));
 sg13g2_o21ai_1 _12474_ (.B1(_08393_),
    .Y(_00008_),
    .A1(_08250_),
    .A2(_08390_));
 sg13g2_nand2b_1 _12475_ (.Y(_08394_),
    .B(net6193),
    .A_N(\soc_inst.mem_ctrl.spi_done ));
 sg13g2_nand2_1 _12476_ (.Y(_08395_),
    .A(net6181),
    .B(_08366_));
 sg13g2_nand3_1 _12477_ (.B(net1812),
    .C(_08366_),
    .A(net6181),
    .Y(_08396_));
 sg13g2_o21ai_1 _12478_ (.B1(_08396_),
    .Y(_08397_),
    .A1(_08384_),
    .A2(_08394_));
 sg13g2_nand3_1 _12479_ (.B(net6179),
    .C(net3281),
    .A(net6504),
    .Y(_08398_));
 sg13g2_nor2_1 _12480_ (.A(_08246_),
    .B(_08398_),
    .Y(_08399_));
 sg13g2_a221oi_1 _12481_ (.B2(_08397_),
    .C1(_08399_),
    .B1(_08249_),
    .A1(net6193),
    .Y(_08400_),
    .A2(net5195));
 sg13g2_inv_1 _12482_ (.Y(_00006_),
    .A(_08400_));
 sg13g2_nor2_1 _12483_ (.A(net6539),
    .B(net6535),
    .Y(_08401_));
 sg13g2_nor3_1 _12484_ (.A(net6539),
    .B(net6537),
    .C(net6535),
    .Y(_08402_));
 sg13g2_nor2_2 _12485_ (.A(net6540),
    .B(net6537),
    .Y(_08403_));
 sg13g2_nor3_1 _12486_ (.A(net3217),
    .B(net3384),
    .C(net3240),
    .Y(_08404_));
 sg13g2_nor2b_2 _12487_ (.A(net6536),
    .B_N(_08404_),
    .Y(_08405_));
 sg13g2_inv_2 _12488_ (.Y(\soc_inst.i2c_ena ),
    .A(_08405_));
 sg13g2_nor2_1 _12489_ (.A(net1812),
    .B(_08395_),
    .Y(_08406_));
 sg13g2_nor2_1 _12490_ (.A(_07865_),
    .B(_08384_),
    .Y(_08407_));
 sg13g2_a21oi_1 _12491_ (.A1(net3281),
    .A2(_08407_),
    .Y(_08408_),
    .B1(_08406_));
 sg13g2_and2_1 _12492_ (.A(_08248_),
    .B(_08289_),
    .X(_08409_));
 sg13g2_o21ai_1 _12493_ (.B1(net6181),
    .Y(_08410_),
    .A1(net5194),
    .A2(_08409_));
 sg13g2_o21ai_1 _12494_ (.B1(_08410_),
    .Y(_00007_),
    .A1(_08250_),
    .A2(_08408_));
 sg13g2_nor2_1 _12495_ (.A(net6202),
    .B(net6201),
    .Y(_08411_));
 sg13g2_nor2_2 _12496_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .B(net6484),
    .Y(_08412_));
 sg13g2_nor3_2 _12497_ (.A(net6202),
    .B(net6201),
    .C(net6486),
    .Y(_08413_));
 sg13g2_nand3_1 _12498_ (.B(_08412_),
    .C(_08413_),
    .A(net6485),
    .Y(_08414_));
 sg13g2_a21oi_1 _12499_ (.A1(net6501),
    .A2(_08414_),
    .Y(_08415_),
    .B1(net2882));
 sg13g2_nor2b_2 _12500_ (.A(\soc_inst.core_mem_addr[30] ),
    .B_N(_08225_),
    .Y(_08416_));
 sg13g2_a21oi_2 _12501_ (.B1(\soc_inst.mem_ctrl.spi_is_instr ),
    .Y(_08417_),
    .A2(_08416_),
    .A1(_08224_));
 sg13g2_a21o_2 _12502_ (.A2(_08416_),
    .A1(_08224_),
    .B1(net6504),
    .X(_08418_));
 sg13g2_and2_1 _12503_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .B(net1309),
    .X(_08419_));
 sg13g2_nor2_2 _12504_ (.A(net6543),
    .B(net3009),
    .Y(_08420_));
 sg13g2_nand2_1 _12505_ (.Y(_08421_),
    .A(_08419_),
    .B(_08420_));
 sg13g2_or3_1 _12506_ (.A(net436),
    .B(_08417_),
    .C(_08421_),
    .X(_08422_));
 sg13g2_o21ai_1 _12507_ (.B1(_08422_),
    .Y(_00013_),
    .A1(net6542),
    .A2(_08415_));
 sg13g2_nand2b_2 _12508_ (.Y(_08423_),
    .B(net850),
    .A_N(net2811));
 sg13g2_xor2_1 _12509_ (.B(net2811),
    .A(net850),
    .X(_00127_));
 sg13g2_nand2_1 _12510_ (.Y(_08424_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(_00315_));
 sg13g2_and2_1 _12511_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B(_00317_),
    .X(_08425_));
 sg13g2_nand2_1 _12512_ (.Y(_08426_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B(_00317_));
 sg13g2_nand2b_1 _12513_ (.Y(_08427_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .A_N(net6175));
 sg13g2_nand4_1 _12514_ (.B(_08424_),
    .C(_08426_),
    .A(_07765_),
    .Y(_08428_),
    .D(_08427_));
 sg13g2_xnor2_1 _12515_ (.Y(_08429_),
    .A(net1742),
    .B(_00318_));
 sg13g2_xnor2_1 _12516_ (.Y(_08430_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .B(_00316_));
 sg13g2_nand2b_1 _12517_ (.Y(_08431_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ));
 sg13g2_nor2_1 _12518_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(_00315_),
    .Y(_08432_));
 sg13g2_a21oi_1 _12519_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .A2(_07802_),
    .Y(_08433_),
    .B1(_08432_));
 sg13g2_nor2_1 _12520_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .B(_07803_),
    .Y(_08434_));
 sg13g2_nor2b_1 _12521_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .Y(_08435_));
 sg13g2_nand2_1 _12522_ (.Y(_08436_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .B(_07803_));
 sg13g2_nor2b_1 _12523_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .B_N(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .Y(_08437_));
 sg13g2_nor2_1 _12524_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .B(_07802_),
    .Y(_08438_));
 sg13g2_nor4_1 _12525_ (.A(_08434_),
    .B(_08435_),
    .C(_08437_),
    .D(_08438_),
    .Y(_08439_));
 sg13g2_nor2b_1 _12526_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .B_N(net6175),
    .Y(_08440_));
 sg13g2_nor2_1 _12527_ (.A(_07766_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .Y(_08441_));
 sg13g2_nor2_1 _12528_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B(_00317_),
    .Y(_08442_));
 sg13g2_nor2_1 _12529_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .B(_07801_),
    .Y(_08443_));
 sg13g2_nor4_1 _12530_ (.A(_08440_),
    .B(_08441_),
    .C(_08442_),
    .D(_08443_),
    .Y(_08444_));
 sg13g2_nand4_1 _12531_ (.B(_08433_),
    .C(_08439_),
    .A(_08431_),
    .Y(_08445_),
    .D(_08444_));
 sg13g2_nor4_1 _12532_ (.A(_08428_),
    .B(_08429_),
    .C(_08430_),
    .D(_08445_),
    .Y(_08446_));
 sg13g2_xnor2_1 _12533_ (.Y(_08447_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ));
 sg13g2_or2_1 _12534_ (.X(_08448_),
    .B(_00317_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ));
 sg13g2_nand2_1 _12535_ (.Y(_08449_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .B(_00317_));
 sg13g2_nand3_1 _12536_ (.B(_08448_),
    .C(_08449_),
    .A(_08447_),
    .Y(_08450_));
 sg13g2_xnor2_1 _12537_ (.Y(_08451_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .B(_00315_));
 sg13g2_xnor2_1 _12538_ (.Y(_08452_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ));
 sg13g2_nand2b_1 _12539_ (.Y(_08453_),
    .B(_08452_),
    .A_N(_08451_));
 sg13g2_nor2_1 _12540_ (.A(_08450_),
    .B(_08453_),
    .Y(_08454_));
 sg13g2_nand2_1 _12541_ (.Y(_08455_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .B(_00318_));
 sg13g2_nand2b_1 _12542_ (.Y(_08456_),
    .B(net6175),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ));
 sg13g2_nand2b_1 _12543_ (.Y(_08457_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ));
 sg13g2_nand2b_1 _12544_ (.Y(_08458_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .A_N(net6175));
 sg13g2_nand4_1 _12545_ (.B(_08456_),
    .C(_08457_),
    .A(_08455_),
    .Y(_08459_),
    .D(_08458_));
 sg13g2_xor2_1 _12546_ (.B(_00316_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .X(_08460_));
 sg13g2_nand2_1 _12547_ (.Y(_08461_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .B(_07802_));
 sg13g2_nand2_1 _12548_ (.Y(_08462_),
    .A(_07765_),
    .B(_07778_));
 sg13g2_nand3_1 _12549_ (.B(_08461_),
    .C(_08462_),
    .A(_08460_),
    .Y(_08463_));
 sg13g2_nand2b_1 _12550_ (.Y(_08464_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ));
 sg13g2_o21ai_1 _12551_ (.B1(_08464_),
    .Y(_08465_),
    .A1(_07766_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ));
 sg13g2_nand2_1 _12552_ (.Y(_08466_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(_07801_));
 sg13g2_o21ai_1 _12553_ (.B1(_08466_),
    .Y(_08467_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .A2(_07800_));
 sg13g2_nor4_1 _12554_ (.A(_08459_),
    .B(_08463_),
    .C(_08465_),
    .D(_08467_),
    .Y(_08468_));
 sg13g2_a22oi_1 _12555_ (.Y(_08469_),
    .B1(_08454_),
    .B2(_08468_),
    .A2(_08446_),
    .A1(net6178));
 sg13g2_xnor2_1 _12556_ (.Y(_08470_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ));
 sg13g2_and2_1 _12557_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .B(_00316_),
    .X(_08471_));
 sg13g2_nand4_1 _12558_ (.B(_08427_),
    .C(_08431_),
    .A(_08424_),
    .Y(_08472_),
    .D(_08436_));
 sg13g2_nor4_1 _12559_ (.A(_08432_),
    .B(_08437_),
    .C(_08471_),
    .D(_08472_),
    .Y(_08473_));
 sg13g2_nor4_1 _12560_ (.A(_08434_),
    .B(_08440_),
    .C(_08441_),
    .D(_08443_),
    .Y(_08474_));
 sg13g2_o21ai_1 _12561_ (.B1(_07765_),
    .Y(_08475_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .A2(_00316_));
 sg13g2_nor4_1 _12562_ (.A(_08425_),
    .B(_08429_),
    .C(_08442_),
    .D(_08475_),
    .Y(_08476_));
 sg13g2_and4_1 _12563_ (.A(_08470_),
    .B(_08473_),
    .C(_08474_),
    .D(_08476_),
    .X(_08477_));
 sg13g2_xnor2_1 _12564_ (.Y(_08478_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ));
 sg13g2_nand2_1 _12565_ (.Y(_08479_),
    .A(_08461_),
    .B(_08464_));
 sg13g2_xnor2_1 _12566_ (.Y(_08480_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ));
 sg13g2_nand4_1 _12567_ (.B(_08452_),
    .C(_08455_),
    .A(_08448_),
    .Y(_08481_),
    .D(_08480_));
 sg13g2_xnor2_1 _12568_ (.Y(_08482_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .B(net6175));
 sg13g2_nand4_1 _12569_ (.B(_08449_),
    .C(_08462_),
    .A(_08447_),
    .Y(_08483_),
    .D(_08482_));
 sg13g2_nor4_1 _12570_ (.A(_08451_),
    .B(_08479_),
    .C(_08481_),
    .D(_08483_),
    .Y(_08484_));
 sg13g2_and3_1 _12571_ (.X(_08485_),
    .A(_08460_),
    .B(_08478_),
    .C(_08484_));
 sg13g2_a21oi_2 _12572_ (.B1(_08485_),
    .Y(_08486_),
    .A2(_08477_),
    .A1(net6178));
 sg13g2_nand2_2 _12573_ (.Y(_08487_),
    .A(net6553),
    .B(_08486_));
 sg13g2_inv_1 _12574_ (.Y(_08488_),
    .A(net5049));
 sg13g2_nor4_1 _12575_ (.A(_07768_),
    .B(net824),
    .C(net2420),
    .D(net2089),
    .Y(_08489_));
 sg13g2_nand2_1 _12576_ (.Y(_08490_),
    .A(net6553),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ));
 sg13g2_nand3_1 _12577_ (.B(net2009),
    .C(_08489_),
    .A(net6553),
    .Y(_08491_));
 sg13g2_o21ai_1 _12578_ (.B1(_08491_),
    .Y(_00022_),
    .A1(_07777_),
    .A2(net5049));
 sg13g2_nor2b_1 _12579_ (.A(net1838),
    .B_N(net2106),
    .Y(_08492_));
 sg13g2_a22oi_1 _12580_ (.Y(_08493_),
    .B1(_08492_),
    .B2(net6553),
    .A2(_08488_),
    .A1(net1842));
 sg13g2_inv_1 _12581_ (.Y(_00021_),
    .A(_08493_));
 sg13g2_nand3b_1 _12582_ (.B(net1842),
    .C(net6553),
    .Y(_08494_),
    .A_N(_08486_));
 sg13g2_o21ai_1 _12583_ (.B1(_08494_),
    .Y(_00020_),
    .A1(_08489_),
    .A2(_08490_));
 sg13g2_a22oi_1 _12584_ (.Y(_08495_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .B2(_00275_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .A1(_00276_));
 sg13g2_a22oi_1 _12585_ (.Y(_08496_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .B2(_00278_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .A1(_00279_));
 sg13g2_nor2_1 _12586_ (.A(_00279_),
    .B(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .Y(_08497_));
 sg13g2_nor2_1 _12587_ (.A(_00280_),
    .B(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .Y(_08498_));
 sg13g2_nor2_1 _12588_ (.A(_08497_),
    .B(_08498_),
    .Y(_08499_));
 sg13g2_or2_1 _12589_ (.X(_08500_),
    .B(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .A(_00276_));
 sg13g2_nor2_1 _12590_ (.A(_00277_),
    .B(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .Y(_08501_));
 sg13g2_nand2_1 _12591_ (.Y(_08502_),
    .A(_00277_),
    .B(\soc_inst.cpu_core.csr_file.mtime[42] ));
 sg13g2_nor2_1 _12592_ (.A(_00278_),
    .B(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .Y(_08503_));
 sg13g2_nor2_1 _12593_ (.A(_08501_),
    .B(_08503_),
    .Y(_08504_));
 sg13g2_nand3_1 _12594_ (.B(_08502_),
    .C(_08504_),
    .A(_08500_),
    .Y(_08505_));
 sg13g2_nor2_1 _12595_ (.A(_00282_),
    .B(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .Y(_08506_));
 sg13g2_a21oi_1 _12596_ (.A1(_00281_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .Y(_08507_),
    .B1(_08506_));
 sg13g2_o21ai_1 _12597_ (.B1(_08507_),
    .Y(_08508_),
    .A1(_00281_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[46] ));
 sg13g2_nand2_1 _12598_ (.Y(_08509_),
    .A(_00280_),
    .B(\soc_inst.cpu_core.csr_file.mtime[45] ));
 sg13g2_a22oi_1 _12599_ (.Y(_08510_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .B2(_00280_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .A1(_00282_));
 sg13g2_o21ai_1 _12600_ (.B1(_08510_),
    .Y(_08511_),
    .A1(_00275_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[40] ));
 sg13g2_nor3_1 _12601_ (.A(_08505_),
    .B(_08508_),
    .C(_08511_),
    .Y(_08512_));
 sg13g2_nand4_1 _12602_ (.B(_08496_),
    .C(_08499_),
    .A(_08495_),
    .Y(_08513_),
    .D(_08512_));
 sg13g2_nor2_1 _12603_ (.A(_00273_),
    .B(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .Y(_08514_));
 sg13g2_a21oi_1 _12604_ (.A1(_07786_),
    .A2(_07905_),
    .Y(_08515_),
    .B1(_08514_));
 sg13g2_a22oi_1 _12605_ (.Y(_08516_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .B2(_00272_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .A1(_00273_));
 sg13g2_or2_1 _12606_ (.X(_08517_),
    .B(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .A(_00272_));
 sg13g2_o21ai_1 _12607_ (.B1(_08517_),
    .Y(_08518_),
    .A1(_00271_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[36] ));
 sg13g2_nand2_1 _12608_ (.Y(_08519_),
    .A(_00269_),
    .B(\soc_inst.cpu_core.csr_file.mtime[34] ));
 sg13g2_nor2_1 _12609_ (.A(_00270_),
    .B(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .Y(_08520_));
 sg13g2_a21oi_1 _12610_ (.A1(_00269_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .Y(_08521_),
    .B1(_08520_));
 sg13g2_o21ai_1 _12611_ (.B1(_08521_),
    .Y(_08522_),
    .A1(_00269_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[34] ));
 sg13g2_nor2_1 _12612_ (.A(_00268_),
    .B(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .Y(_08523_));
 sg13g2_a22oi_1 _12613_ (.Y(_08524_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .B2(_00267_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .A1(_00268_));
 sg13g2_nor3_1 _12614_ (.A(_08522_),
    .B(_08523_),
    .C(_08524_),
    .Y(_08525_));
 sg13g2_a22oi_1 _12615_ (.Y(_08526_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .B2(_00270_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .A1(_00271_));
 sg13g2_o21ai_1 _12616_ (.B1(_08526_),
    .Y(_08527_),
    .A1(_08519_),
    .A2(_08520_));
 sg13g2_nor2_1 _12617_ (.A(_08525_),
    .B(_08527_),
    .Y(_08528_));
 sg13g2_o21ai_1 _12618_ (.B1(_08516_),
    .Y(_08529_),
    .A1(_08518_),
    .A2(_08528_));
 sg13g2_a22oi_1 _12619_ (.Y(_08530_),
    .B1(_08515_),
    .B2(_08529_),
    .A2(net3398),
    .A1(net1641));
 sg13g2_a22oi_1 _12620_ (.Y(_08531_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .B2(_00281_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .A1(_00282_));
 sg13g2_nor2_1 _12621_ (.A(_08506_),
    .B(_08531_),
    .Y(_08532_));
 sg13g2_nor2_1 _12622_ (.A(_08495_),
    .B(_08505_),
    .Y(_08533_));
 sg13g2_o21ai_1 _12623_ (.B1(_08496_),
    .Y(_08534_),
    .A1(_08502_),
    .A2(_08503_));
 sg13g2_o21ai_1 _12624_ (.B1(_08499_),
    .Y(_08535_),
    .A1(_08533_),
    .A2(_08534_));
 sg13g2_a21oi_1 _12625_ (.A1(_08509_),
    .A2(_08535_),
    .Y(_08536_),
    .B1(_08508_));
 sg13g2_nor2_1 _12626_ (.A(_08532_),
    .B(_08536_),
    .Y(_08537_));
 sg13g2_o21ai_1 _12627_ (.B1(_08537_),
    .Y(_08538_),
    .A1(_08513_),
    .A2(_08530_));
 sg13g2_a22oi_1 _12628_ (.Y(_08539_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .B2(_00297_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .A1(_00298_));
 sg13g2_a22oi_1 _12629_ (.Y(_08540_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .B2(_00295_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .A1(_00296_));
 sg13g2_nor2_1 _12630_ (.A(_00298_),
    .B(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .Y(_08541_));
 sg13g2_or2_1 _12631_ (.X(_08542_),
    .B(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .A(_00297_));
 sg13g2_o21ai_1 _12632_ (.B1(_08542_),
    .Y(_08543_),
    .A1(_00296_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[13] ));
 sg13g2_o21ai_1 _12633_ (.B1(_08539_),
    .Y(_08544_),
    .A1(_08540_),
    .A2(_08543_));
 sg13g2_nand2b_1 _12634_ (.Y(_08545_),
    .B(_08544_),
    .A_N(_08541_));
 sg13g2_nand2_1 _12635_ (.Y(_08546_),
    .A(_00289_),
    .B(\soc_inst.cpu_core.csr_file.mtime[6] ));
 sg13g2_or2_1 _12636_ (.X(_08547_),
    .B(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .A(_00287_));
 sg13g2_nor2_1 _12637_ (.A(_00284_),
    .B(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .Y(_08548_));
 sg13g2_nor2_1 _12638_ (.A(_00283_),
    .B(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .Y(_08549_));
 sg13g2_a22oi_1 _12639_ (.Y(_08550_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .B2(_00285_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .A1(_00284_));
 sg13g2_o21ai_1 _12640_ (.B1(_08550_),
    .Y(_08551_),
    .A1(_08548_),
    .A2(_08549_));
 sg13g2_or2_1 _12641_ (.X(_08552_),
    .B(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .A(_00285_));
 sg13g2_a22oi_1 _12642_ (.Y(_08553_),
    .B1(_08551_),
    .B2(_08552_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .A1(_00286_));
 sg13g2_o21ai_1 _12643_ (.B1(_08547_),
    .Y(_08554_),
    .A1(_00286_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[3] ));
 sg13g2_a22oi_1 _12644_ (.Y(_08555_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .B2(_00287_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .A1(_00288_));
 sg13g2_o21ai_1 _12645_ (.B1(_08555_),
    .Y(_08556_),
    .A1(_08553_),
    .A2(_08554_));
 sg13g2_o21ai_1 _12646_ (.B1(_08556_),
    .Y(_08557_),
    .A1(_00288_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[5] ));
 sg13g2_nor2_1 _12647_ (.A(_00289_),
    .B(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .Y(_08558_));
 sg13g2_a21oi_1 _12648_ (.A1(_08546_),
    .A2(_08557_),
    .Y(_08559_),
    .B1(_08558_));
 sg13g2_o21ai_1 _12649_ (.B1(_08559_),
    .Y(_08560_),
    .A1(_00290_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[7] ));
 sg13g2_o21ai_1 _12650_ (.B1(_08560_),
    .Y(_08561_),
    .A1(_07783_),
    .A2(_07901_));
 sg13g2_o21ai_1 _12651_ (.B1(_08561_),
    .Y(_08562_),
    .A1(_00291_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[8] ));
 sg13g2_a22oi_1 _12652_ (.Y(_08563_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .B2(_00291_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .A1(_00292_));
 sg13g2_or2_1 _12653_ (.X(_08564_),
    .B(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .A(_00293_));
 sg13g2_o21ai_1 _12654_ (.B1(_08564_),
    .Y(_08565_),
    .A1(_00292_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[9] ));
 sg13g2_a21oi_1 _12655_ (.A1(_08562_),
    .A2(_08563_),
    .Y(_08566_),
    .B1(_08565_));
 sg13g2_a221oi_1 _12656_ (.B2(_00293_),
    .C1(_08566_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .A1(_00294_),
    .Y(_08567_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[11] ));
 sg13g2_nor2_1 _12657_ (.A(_00294_),
    .B(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .Y(_08568_));
 sg13g2_nor2_1 _12658_ (.A(_00295_),
    .B(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .Y(_08569_));
 sg13g2_nor4_1 _12659_ (.A(_08541_),
    .B(_08543_),
    .C(_08568_),
    .D(_08569_),
    .Y(_08570_));
 sg13g2_nand3_1 _12660_ (.B(_08540_),
    .C(_08570_),
    .A(_08539_),
    .Y(_08571_));
 sg13g2_o21ai_1 _12661_ (.B1(_08545_),
    .Y(_08572_),
    .A1(_08567_),
    .A2(_08571_));
 sg13g2_or2_1 _12662_ (.X(_08573_),
    .B(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A(_00303_));
 sg13g2_o21ai_1 _12663_ (.B1(_08573_),
    .Y(_08574_),
    .A1(_00304_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[21] ));
 sg13g2_a22oi_1 _12664_ (.Y(_08575_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .B2(_00300_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .A1(_00301_));
 sg13g2_nand2b_1 _12665_ (.Y(_08576_),
    .B(_08575_),
    .A_N(_08574_));
 sg13g2_or2_1 _12666_ (.X(_08577_),
    .B(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .A(_00306_));
 sg13g2_o21ai_1 _12667_ (.B1(_08577_),
    .Y(_08578_),
    .A1(_00305_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[22] ));
 sg13g2_or2_1 _12668_ (.X(_08579_),
    .B(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .A(_00302_));
 sg13g2_o21ai_1 _12669_ (.B1(_08579_),
    .Y(_08580_),
    .A1(_00301_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[18] ));
 sg13g2_nor2_1 _12670_ (.A(_00300_),
    .B(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .Y(_08581_));
 sg13g2_a21oi_1 _12671_ (.A1(_00306_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .Y(_08582_),
    .B1(_08581_));
 sg13g2_or2_1 _12672_ (.X(_08583_),
    .B(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .A(_00299_));
 sg13g2_nand2_1 _12673_ (.Y(_08584_),
    .A(_00299_),
    .B(\soc_inst.cpu_core.csr_file.mtime[16] ));
 sg13g2_a22oi_1 _12674_ (.Y(_08585_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .B2(_00302_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .A1(_00303_));
 sg13g2_a22oi_1 _12675_ (.Y(_08586_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .B2(_00304_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .A1(_00305_));
 sg13g2_and2_1 _12676_ (.A(_08585_),
    .B(_08586_),
    .X(_08587_));
 sg13g2_nand4_1 _12677_ (.B(_08583_),
    .C(_08584_),
    .A(_08582_),
    .Y(_08588_),
    .D(_08587_));
 sg13g2_nor4_1 _12678_ (.A(_08576_),
    .B(_08578_),
    .C(_08580_),
    .D(_08588_),
    .Y(_08589_));
 sg13g2_o21ai_1 _12679_ (.B1(_08575_),
    .Y(_08590_),
    .A1(_08581_),
    .A2(_08584_));
 sg13g2_nand2b_1 _12680_ (.Y(_08591_),
    .B(_08590_),
    .A_N(_08580_));
 sg13g2_a221oi_1 _12681_ (.B2(_08591_),
    .C1(_08578_),
    .B1(_08587_),
    .A1(_08574_),
    .Y(_08592_),
    .A2(_08586_));
 sg13g2_a221oi_1 _12682_ (.B2(_08589_),
    .C1(_08592_),
    .B1(_08572_),
    .A1(_00306_),
    .Y(_08593_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[23] ));
 sg13g2_or2_1 _12683_ (.X(_08594_),
    .B(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .A(_00311_));
 sg13g2_o21ai_1 _12684_ (.B1(_08594_),
    .Y(_08595_),
    .A1(_00312_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[29] ));
 sg13g2_a22oi_1 _12685_ (.Y(_08596_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .B2(_00307_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .A1(_00308_));
 sg13g2_a22oi_1 _12686_ (.Y(_08597_),
    .B1(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .B2(_00310_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .A1(_00311_));
 sg13g2_nand2_1 _12687_ (.Y(_08598_),
    .A(_08596_),
    .B(_08597_));
 sg13g2_nand2_1 _12688_ (.Y(_08599_),
    .A(_00313_),
    .B(\soc_inst.cpu_core.csr_file.mtime[30] ));
 sg13g2_nor2_1 _12689_ (.A(_00314_),
    .B(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .Y(_08600_));
 sg13g2_xnor2_1 _12690_ (.Y(_08601_),
    .A(_00313_),
    .B(\soc_inst.cpu_core.csr_file.mtime[30] ));
 sg13g2_nor2_1 _12691_ (.A(_08600_),
    .B(_08601_),
    .Y(_08602_));
 sg13g2_nand2_1 _12692_ (.Y(_08603_),
    .A(_00312_),
    .B(\soc_inst.cpu_core.csr_file.mtime[29] ));
 sg13g2_o21ai_1 _12693_ (.B1(_08603_),
    .Y(_08604_),
    .A1(_00307_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[24] ));
 sg13g2_a21oi_1 _12694_ (.A1(_00314_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .Y(_08605_),
    .B1(_08604_));
 sg13g2_nor2_1 _12695_ (.A(_00308_),
    .B(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .Y(_08606_));
 sg13g2_or2_1 _12696_ (.X(_08607_),
    .B(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .A(_00309_));
 sg13g2_nor2_1 _12697_ (.A(_00310_),
    .B(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .Y(_08608_));
 sg13g2_nand2_1 _12698_ (.Y(_08609_),
    .A(_00309_),
    .B(\soc_inst.cpu_core.csr_file.mtime[26] ));
 sg13g2_nor2_1 _12699_ (.A(_08606_),
    .B(_08608_),
    .Y(_08610_));
 sg13g2_nand3_1 _12700_ (.B(_08609_),
    .C(_08610_),
    .A(_08607_),
    .Y(_08611_));
 sg13g2_nor3_1 _12701_ (.A(_08595_),
    .B(_08598_),
    .C(_08611_),
    .Y(_08612_));
 sg13g2_nand3_1 _12702_ (.B(_08605_),
    .C(_08612_),
    .A(_08602_),
    .Y(_08613_));
 sg13g2_nor2_1 _12703_ (.A(_08608_),
    .B(_08609_),
    .Y(_08614_));
 sg13g2_o21ai_1 _12704_ (.B1(_08597_),
    .Y(_08615_),
    .A1(_08596_),
    .A2(_08611_));
 sg13g2_nor2_1 _12705_ (.A(_08614_),
    .B(_08615_),
    .Y(_08616_));
 sg13g2_o21ai_1 _12706_ (.B1(_08603_),
    .Y(_08617_),
    .A1(_08595_),
    .A2(_08616_));
 sg13g2_nor2_1 _12707_ (.A(_08599_),
    .B(_08600_),
    .Y(_08618_));
 sg13g2_a221oi_1 _12708_ (.B2(_08617_),
    .C1(_08618_),
    .B1(_08602_),
    .A1(_00314_),
    .Y(_08619_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[31] ));
 sg13g2_o21ai_1 _12709_ (.B1(_08619_),
    .Y(_08620_),
    .A1(_08593_),
    .A2(_08613_));
 sg13g2_nand3b_1 _12710_ (.B(_08524_),
    .C(_08526_),
    .Y(_08621_),
    .A_N(_08518_));
 sg13g2_a21oi_1 _12711_ (.A1(_00274_),
    .A2(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .Y(_08622_),
    .B1(_08523_));
 sg13g2_or2_1 _12712_ (.X(_08623_),
    .B(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .A(_00267_));
 sg13g2_nand4_1 _12713_ (.B(_08516_),
    .C(_08622_),
    .A(_08515_),
    .Y(_08624_),
    .D(_08623_));
 sg13g2_nor4_1 _12714_ (.A(_08513_),
    .B(_08522_),
    .C(_08621_),
    .D(_08624_),
    .Y(_08625_));
 sg13g2_a21o_2 _12715_ (.A2(_08625_),
    .A1(_08620_),
    .B1(_08538_),
    .X(_00023_));
 sg13g2_a21oi_1 _12716_ (.A1(net1838),
    .A2(net2106),
    .Y(_08626_),
    .B1(_07884_));
 sg13g2_o21ai_1 _12717_ (.B1(_08626_),
    .Y(_00019_),
    .A1(_07777_),
    .A2(_08486_));
 sg13g2_nand2_1 _12718_ (.Y(_08627_),
    .A(net3344),
    .B(_08414_));
 sg13g2_a21oi_1 _12719_ (.A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .A2(_08414_),
    .Y(_08628_),
    .B1(net1375));
 sg13g2_nand4_1 _12720_ (.B(_08417_),
    .C(_08419_),
    .A(net227),
    .Y(_08629_),
    .D(_08420_));
 sg13g2_o21ai_1 _12721_ (.B1(_08629_),
    .Y(_00011_),
    .A1(net6542),
    .A2(net1376));
 sg13g2_nor2_1 _12722_ (.A(_07878_),
    .B(net6485),
    .Y(_08630_));
 sg13g2_nand3_1 _12723_ (.B(_08412_),
    .C(_08630_),
    .A(net6201),
    .Y(_08631_));
 sg13g2_o21ai_1 _12724_ (.B1(net6488),
    .Y(_08632_),
    .A1(net6202),
    .A2(_08631_));
 sg13g2_nand4_1 _12725_ (.B(_07880_),
    .C(net6484),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .Y(_08633_),
    .D(_08413_));
 sg13g2_nor2_2 _12726_ (.A(_07882_),
    .B(_08633_),
    .Y(_08634_));
 sg13g2_nand2b_1 _12727_ (.Y(_08635_),
    .B(net3367),
    .A_N(net6507));
 sg13g2_a21oi_1 _12728_ (.A1(_08632_),
    .A2(_08635_),
    .Y(_00010_),
    .B1(net6542));
 sg13g2_nand4_1 _12729_ (.B(net6201),
    .C(_08412_),
    .A(net6202),
    .Y(_08636_),
    .D(_08630_));
 sg13g2_a21oi_1 _12730_ (.A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .A2(_08636_),
    .Y(_08637_),
    .B1(net1134));
 sg13g2_nand2b_1 _12731_ (.Y(_08638_),
    .B(net2273),
    .A_N(net6541));
 sg13g2_nor2_1 _12732_ (.A(net6541),
    .B(net1135),
    .Y(_00018_));
 sg13g2_nand2b_1 _12733_ (.Y(_08639_),
    .B(net311),
    .A_N(net6541));
 sg13g2_nand4_1 _12734_ (.B(net354),
    .C(net388),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .Y(_08640_),
    .D(net144));
 sg13g2_nand4_1 _12735_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .C(net363),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .Y(_08641_),
    .D(net358));
 sg13g2_nand4_1 _12736_ (.B(net1638),
    .C(net338),
    .A(net253),
    .Y(_08642_),
    .D(net562));
 sg13g2_nor3_1 _12737_ (.A(_08640_),
    .B(_08641_),
    .C(_08642_),
    .Y(_08643_));
 sg13g2_nand3b_1 _12738_ (.B(_08420_),
    .C(net1568),
    .Y(_08644_),
    .A_N(net1309));
 sg13g2_o21ai_1 _12739_ (.B1(_08644_),
    .Y(_00017_),
    .A1(_08639_),
    .A2(net1639));
 sg13g2_nand2_1 _12740_ (.Y(_08645_),
    .A(net6203),
    .B(_08412_));
 sg13g2_nor2_1 _12741_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .B(_08645_),
    .Y(_08646_));
 sg13g2_nand3_1 _12742_ (.B(net6485),
    .C(_08646_),
    .A(_07878_),
    .Y(_08647_));
 sg13g2_nand2_1 _12743_ (.Y(_08648_),
    .A(net1027),
    .B(_08647_));
 sg13g2_a21oi_1 _12744_ (.A1(_07876_),
    .A2(_08648_),
    .Y(_00016_),
    .B1(net6541));
 sg13g2_xnor2_1 _12745_ (.Y(_08649_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .B(net2851));
 sg13g2_xnor2_1 _12746_ (.Y(_08650_),
    .A(net6485),
    .B(net2779));
 sg13g2_xnor2_1 _12747_ (.Y(_08651_),
    .A(net6484),
    .B(\soc_inst.mem_ctrl.spi_data_len[4] ));
 sg13g2_nand4_1 _12748_ (.B(_08649_),
    .C(_08650_),
    .A(_08413_),
    .Y(_08652_),
    .D(_08651_));
 sg13g2_nor2_1 _12749_ (.A(net6543),
    .B(net6505),
    .Y(_08653_));
 sg13g2_nand3_1 _12750_ (.B(_08652_),
    .C(_08653_),
    .A(net6494),
    .Y(_08654_));
 sg13g2_nor3_1 _12751_ (.A(_07873_),
    .B(net6203),
    .C(_08631_),
    .Y(_08655_));
 sg13g2_a221oi_1 _12752_ (.B2(net3190),
    .C1(_08655_),
    .B1(_08634_),
    .A1(net6505),
    .Y(_08656_),
    .A2(net6489));
 sg13g2_o21ai_1 _12753_ (.B1(_08654_),
    .Y(_00015_),
    .A1(net6543),
    .A2(net3191));
 sg13g2_nor2_2 _12754_ (.A(_07878_),
    .B(_07879_),
    .Y(_08657_));
 sg13g2_nand2_1 _12755_ (.Y(_08658_),
    .A(_08646_),
    .B(_08657_));
 sg13g2_nand3b_1 _12756_ (.B(net1077),
    .C(_08658_),
    .Y(_08659_),
    .A_N(net6541));
 sg13g2_o21ai_1 _12757_ (.B1(_08659_),
    .Y(_00014_),
    .A1(_08636_),
    .A2(_08638_));
 sg13g2_nand2_2 _12758_ (.Y(_08660_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .B(_08633_));
 sg13g2_nor2_1 _12759_ (.A(net6501),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .Y(_08661_));
 sg13g2_o21ai_1 _12760_ (.B1(_08660_),
    .Y(_08662_),
    .A1(_08414_),
    .A2(_08661_));
 sg13g2_inv_1 _12761_ (.Y(_08663_),
    .A(_08662_));
 sg13g2_nand4_1 _12762_ (.B(net5568),
    .C(_08419_),
    .A(net436),
    .Y(_08664_),
    .D(_08420_));
 sg13g2_o21ai_1 _12763_ (.B1(net437),
    .Y(_00012_),
    .A1(net6542),
    .A2(_08663_));
 sg13g2_nor2_1 _12764_ (.A(_07875_),
    .B(net6506),
    .Y(_08665_));
 sg13g2_nand2b_2 _12765_ (.Y(_08666_),
    .B(net6490),
    .A_N(net6506));
 sg13g2_nor2_1 _12766_ (.A(net95),
    .B(net98),
    .Y(_00109_));
 sg13g2_nor4_2 _12767_ (.A(net2908),
    .B(net3038),
    .C(net3104),
    .Y(_08667_),
    .D(net2958));
 sg13g2_nor2_2 _12768_ (.A(\soc_inst.core_mem_addr[1] ),
    .B(\soc_inst.core_mem_addr[0] ),
    .Y(_08668_));
 sg13g2_and2_1 _12769_ (.A(net6211),
    .B(_08668_),
    .X(_08669_));
 sg13g2_nand2_1 _12770_ (.Y(_08670_),
    .A(net6211),
    .B(_08668_));
 sg13g2_nand2_1 _12771_ (.Y(_08671_),
    .A(net6206),
    .B(_08668_));
 sg13g2_nand2_2 _12772_ (.Y(_08672_),
    .A(net6206),
    .B(net6067));
 sg13g2_and3_2 _12773_ (.X(_08673_),
    .A(net6209),
    .B(_08667_),
    .C(net6068));
 sg13g2_inv_1 _12774_ (.Y(_08674_),
    .A(net5566));
 sg13g2_and2_1 _12775_ (.A(\soc_inst.core_mem_addr[12] ),
    .B(_08235_),
    .X(_08675_));
 sg13g2_nand2_2 _12776_ (.Y(_08676_),
    .A(\soc_inst.core_mem_addr[12] ),
    .B(_08235_));
 sg13g2_nand3_1 _12777_ (.B(_08229_),
    .C(_08675_),
    .A(net6204),
    .Y(_08677_));
 sg13g2_nor3_1 _12778_ (.A(\soc_inst.spi_inst.busy ),
    .B(_08674_),
    .C(_08677_),
    .Y(_08678_));
 sg13g2_nor2b_1 _12779_ (.A(net5183),
    .B_N(net187),
    .Y(_08679_));
 sg13g2_a21oi_1 _12780_ (.A1(net268),
    .A2(net5181),
    .Y(_08680_),
    .B1(_08679_));
 sg13g2_xnor2_1 _12781_ (.Y(_08681_),
    .A(\soc_inst.spi_inst.clk_counter[6] ),
    .B(\soc_inst.spi_inst.clock_divider[6] ));
 sg13g2_xnor2_1 _12782_ (.Y(_08682_),
    .A(\soc_inst.spi_inst.clk_counter[5] ),
    .B(\soc_inst.spi_inst.clock_divider[5] ));
 sg13g2_nand2_1 _12783_ (.Y(_08683_),
    .A(_08681_),
    .B(_08682_));
 sg13g2_xor2_1 _12784_ (.B(\soc_inst.spi_inst.clk_counter[3] ),
    .A(_00224_),
    .X(_08684_));
 sg13g2_inv_1 _12785_ (.Y(_08685_),
    .A(_08684_));
 sg13g2_nor2b_1 _12786_ (.A(\soc_inst.spi_inst.clock_divider[7] ),
    .B_N(\soc_inst.spi_inst.clk_counter[7] ),
    .Y(_08686_));
 sg13g2_xor2_1 _12787_ (.B(\soc_inst.spi_inst.clock_divider[7] ),
    .A(\soc_inst.spi_inst.clk_counter[7] ),
    .X(_08687_));
 sg13g2_xor2_1 _12788_ (.B(\soc_inst.spi_inst.clk_counter[0] ),
    .A(_00221_),
    .X(_08688_));
 sg13g2_xor2_1 _12789_ (.B(\soc_inst.spi_inst.clk_counter[1] ),
    .A(_00222_),
    .X(_08689_));
 sg13g2_xor2_1 _12790_ (.B(\soc_inst.spi_inst.clk_counter[2] ),
    .A(_00223_),
    .X(_08690_));
 sg13g2_xor2_1 _12791_ (.B(\soc_inst.spi_inst.clk_counter[4] ),
    .A(_00225_),
    .X(_08691_));
 sg13g2_nand4_1 _12792_ (.B(_08689_),
    .C(_08690_),
    .A(_08688_),
    .Y(_08692_),
    .D(_08691_));
 sg13g2_nor4_1 _12793_ (.A(_08683_),
    .B(_08685_),
    .C(_08687_),
    .D(_08692_),
    .Y(_08693_));
 sg13g2_nand2_1 _12794_ (.Y(_08694_),
    .A(\soc_inst.spi_inst.spi_clk_en ),
    .B(_08693_));
 sg13g2_nor2_1 _12795_ (.A(_07898_),
    .B(_08694_),
    .Y(_08695_));
 sg13g2_nor2_1 _12796_ (.A(net2653),
    .B(_08694_),
    .Y(_08696_));
 sg13g2_mux2_1 _12797_ (.A0(_08696_),
    .A1(_08695_),
    .S(\soc_inst.spi_inst.cpol ),
    .X(_08697_));
 sg13g2_nor2_1 _12798_ (.A(\soc_inst.spi_inst.cpha ),
    .B(_08697_),
    .Y(_08698_));
 sg13g2_nor3_1 _12799_ (.A(\soc_inst.spi_inst.cpol ),
    .B(_07898_),
    .C(_08694_),
    .Y(_08699_));
 sg13g2_a21oi_1 _12800_ (.A1(\soc_inst.spi_inst.cpol ),
    .A2(_08696_),
    .Y(_08700_),
    .B1(_08699_));
 sg13g2_and2_1 _12801_ (.A(\soc_inst.spi_inst.cpha ),
    .B(_08700_),
    .X(_08701_));
 sg13g2_nor3_1 _12802_ (.A(net6110),
    .B(_08698_),
    .C(_08701_),
    .Y(_08702_));
 sg13g2_nor3_2 _12803_ (.A(_08423_),
    .B(_08698_),
    .C(_08701_),
    .Y(_08703_));
 sg13g2_nor2_1 _12804_ (.A(_08680_),
    .B(net5013),
    .Y(_00138_));
 sg13g2_nand2b_1 _12805_ (.Y(_08704_),
    .B(net5183),
    .A_N(\soc_inst.core_mem_wdata[25] ));
 sg13g2_o21ai_1 _12806_ (.B1(_08704_),
    .Y(_08705_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[1] ),
    .A2(net5181));
 sg13g2_nand2_1 _12807_ (.Y(_08706_),
    .A(net187),
    .B(net5013));
 sg13g2_o21ai_1 _12808_ (.B1(_08706_),
    .Y(_00149_),
    .A1(net5014),
    .A2(_08705_));
 sg13g2_nand2b_1 _12809_ (.Y(_08707_),
    .B(net5183),
    .A_N(\soc_inst.core_mem_wdata[26] ));
 sg13g2_o21ai_1 _12810_ (.B1(_08707_),
    .Y(_08708_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[2] ),
    .A2(net5181));
 sg13g2_nand2_1 _12811_ (.Y(_08709_),
    .A(net189),
    .B(net5013));
 sg13g2_o21ai_1 _12812_ (.B1(_08709_),
    .Y(_00160_),
    .A1(net5013),
    .A2(_08708_));
 sg13g2_mux2_1 _12813_ (.A0(net286),
    .A1(net712),
    .S(net5183),
    .X(_08710_));
 sg13g2_mux2_1 _12814_ (.A0(_08710_),
    .A1(net1445),
    .S(net5013),
    .X(_00163_));
 sg13g2_nand2b_1 _12815_ (.Y(_08711_),
    .B(net5182),
    .A_N(\soc_inst.core_mem_wdata[28] ));
 sg13g2_o21ai_1 _12816_ (.B1(_08711_),
    .Y(_08712_),
    .A1(net155),
    .A2(net5182));
 sg13g2_nand2_1 _12817_ (.Y(_08713_),
    .A(net286),
    .B(net5012));
 sg13g2_o21ai_1 _12818_ (.B1(_08713_),
    .Y(_00164_),
    .A1(net5012),
    .A2(_08712_));
 sg13g2_nand2b_1 _12819_ (.Y(_08714_),
    .B(net5182),
    .A_N(\soc_inst.core_mem_wdata[29] ));
 sg13g2_o21ai_1 _12820_ (.B1(_08714_),
    .Y(_08715_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[5] ),
    .A2(net5182));
 sg13g2_nand2_1 _12821_ (.Y(_08716_),
    .A(net155),
    .B(net5012));
 sg13g2_o21ai_1 _12822_ (.B1(_08716_),
    .Y(_00165_),
    .A1(net5012),
    .A2(_08715_));
 sg13g2_mux2_1 _12823_ (.A0(net330),
    .A1(net734),
    .S(net5181),
    .X(_08717_));
 sg13g2_mux2_1 _12824_ (.A0(_08717_),
    .A1(net1526),
    .S(net5012),
    .X(_00166_));
 sg13g2_nand2b_1 _12825_ (.Y(_08718_),
    .B(net5183),
    .A_N(\soc_inst.core_mem_wdata[31] ));
 sg13g2_o21ai_1 _12826_ (.B1(_08718_),
    .Y(_08719_),
    .A1(net174),
    .A2(net5181));
 sg13g2_nand2_1 _12827_ (.Y(_08720_),
    .A(net330),
    .B(net5012));
 sg13g2_o21ai_1 _12828_ (.B1(_08720_),
    .Y(_00167_),
    .A1(net5013),
    .A2(_08719_));
 sg13g2_nand2b_1 _12829_ (.Y(_08721_),
    .B(net5181),
    .A_N(\soc_inst.core_mem_wdata[16] ));
 sg13g2_o21ai_1 _12830_ (.B1(_08721_),
    .Y(_08722_),
    .A1(net163),
    .A2(net5181));
 sg13g2_nand2_1 _12831_ (.Y(_08723_),
    .A(net174),
    .B(net5012));
 sg13g2_o21ai_1 _12832_ (.B1(_08723_),
    .Y(_00168_),
    .A1(net5013),
    .A2(_08722_));
 sg13g2_nand2b_1 _12833_ (.Y(_08724_),
    .B(net5181),
    .A_N(net160));
 sg13g2_o21ai_1 _12834_ (.B1(_08724_),
    .Y(_08725_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .A2(net5182));
 sg13g2_nand2_1 _12835_ (.Y(_08726_),
    .A(net163),
    .B(net5012));
 sg13g2_o21ai_1 _12836_ (.B1(_08726_),
    .Y(_00169_),
    .A1(net5014),
    .A2(_08725_));
 sg13g2_nand2b_1 _12837_ (.Y(_08727_),
    .B(net5182),
    .A_N(\soc_inst.core_mem_wdata[18] ));
 sg13g2_o21ai_1 _12838_ (.B1(_08727_),
    .Y(_08728_),
    .A1(net413),
    .A2(net5184));
 sg13g2_nand2_1 _12839_ (.Y(_08729_),
    .A(net596),
    .B(net5014));
 sg13g2_o21ai_1 _12840_ (.B1(_08729_),
    .Y(_00139_),
    .A1(net5015),
    .A2(_08728_));
 sg13g2_nand2b_1 _12841_ (.Y(_08730_),
    .B(net5182),
    .A_N(net295));
 sg13g2_o21ai_1 _12842_ (.B1(_08730_),
    .Y(_08731_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[11] ),
    .A2(net5184));
 sg13g2_nand2_1 _12843_ (.Y(_08732_),
    .A(net413),
    .B(net5015));
 sg13g2_o21ai_1 _12844_ (.B1(_08732_),
    .Y(_00140_),
    .A1(net5015),
    .A2(_08731_));
 sg13g2_mux2_1 _12845_ (.A0(net158),
    .A1(net548),
    .S(net5184),
    .X(_08733_));
 sg13g2_mux2_1 _12846_ (.A0(_08733_),
    .A1(net1428),
    .S(net5015),
    .X(_00141_));
 sg13g2_nand2b_1 _12847_ (.Y(_08734_),
    .B(net5182),
    .A_N(\soc_inst.core_mem_wdata[21] ));
 sg13g2_o21ai_1 _12848_ (.B1(_08734_),
    .Y(_08735_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[13] ),
    .A2(net5184));
 sg13g2_nand2_1 _12849_ (.Y(_08736_),
    .A(net158),
    .B(net5015));
 sg13g2_o21ai_1 _12850_ (.B1(_08736_),
    .Y(_00142_),
    .A1(net5015),
    .A2(_08735_));
 sg13g2_mux2_1 _12851_ (.A0(net204),
    .A1(net1311),
    .S(net5184),
    .X(_08737_));
 sg13g2_mux2_1 _12852_ (.A0(_08737_),
    .A1(net2246),
    .S(net5015),
    .X(_00143_));
 sg13g2_nand2b_1 _12853_ (.Y(_08738_),
    .B(net5180),
    .A_N(\soc_inst.core_mem_wdata[23] ));
 sg13g2_o21ai_1 _12854_ (.B1(_08738_),
    .Y(_08739_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[15] ),
    .A2(net5180));
 sg13g2_nand2_1 _12855_ (.Y(_08740_),
    .A(net204),
    .B(net5010));
 sg13g2_o21ai_1 _12856_ (.B1(_08740_),
    .Y(_00144_),
    .A1(net5010),
    .A2(_08739_));
 sg13g2_mux2_1 _12857_ (.A0(net323),
    .A1(net6454),
    .S(net5179),
    .X(_08741_));
 sg13g2_mux2_1 _12858_ (.A0(_08741_),
    .A1(net1769),
    .S(net5009),
    .X(_00145_));
 sg13g2_nand2b_1 _12859_ (.Y(_08742_),
    .B(net5179),
    .A_N(net6453));
 sg13g2_o21ai_1 _12860_ (.B1(_08742_),
    .Y(_08743_),
    .A1(net307),
    .A2(net5179));
 sg13g2_nand2_1 _12861_ (.Y(_08744_),
    .A(net323),
    .B(net5009));
 sg13g2_o21ai_1 _12862_ (.B1(_08744_),
    .Y(_00146_),
    .A1(net5009),
    .A2(_08743_));
 sg13g2_nand2b_1 _12863_ (.Y(_08745_),
    .B(net5179),
    .A_N(\soc_inst.core_mem_wdata[10] ));
 sg13g2_o21ai_1 _12864_ (.B1(_08745_),
    .Y(_08746_),
    .A1(net200),
    .A2(net5179));
 sg13g2_nand2_1 _12865_ (.Y(_08747_),
    .A(net307),
    .B(net5009));
 sg13g2_o21ai_1 _12866_ (.B1(_08747_),
    .Y(_00147_),
    .A1(net5009),
    .A2(_08746_));
 sg13g2_nand2b_1 _12867_ (.Y(_08748_),
    .B(net5179),
    .A_N(\soc_inst.core_mem_wdata[11] ));
 sg13g2_o21ai_1 _12868_ (.B1(_08748_),
    .Y(_08749_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[19] ),
    .A2(net5179));
 sg13g2_nand2_1 _12869_ (.Y(_08750_),
    .A(net200),
    .B(net5009));
 sg13g2_o21ai_1 _12870_ (.B1(_08750_),
    .Y(_00148_),
    .A1(net5009),
    .A2(_08749_));
 sg13g2_mux2_1 _12871_ (.A0(\soc_inst.spi_inst.tx_shift_reg[20] ),
    .A1(\soc_inst.core_mem_wdata[12] ),
    .S(net5179),
    .X(_08751_));
 sg13g2_mux2_1 _12872_ (.A0(_08751_),
    .A1(net1493),
    .S(net5009),
    .X(_00150_));
 sg13g2_mux2_1 _12873_ (.A0(net1335),
    .A1(net1321),
    .S(net5180),
    .X(_08752_));
 sg13g2_mux2_1 _12874_ (.A0(_08752_),
    .A1(net1950),
    .S(net5010),
    .X(_00151_));
 sg13g2_mux2_1 _12875_ (.A0(net1103),
    .A1(\soc_inst.core_mem_wdata[14] ),
    .S(net5180),
    .X(_08753_));
 sg13g2_mux2_1 _12876_ (.A0(_08753_),
    .A1(net1335),
    .S(net5011),
    .X(_00152_));
 sg13g2_mux2_1 _12877_ (.A0(net249),
    .A1(\soc_inst.core_mem_wdata[15] ),
    .S(net5180),
    .X(_08754_));
 sg13g2_mux2_1 _12878_ (.A0(_08754_),
    .A1(net1103),
    .S(net5010),
    .X(_00153_));
 sg13g2_nand2_1 _12879_ (.Y(_08755_),
    .A(_07785_),
    .B(net5180));
 sg13g2_o21ai_1 _12880_ (.B1(_08755_),
    .Y(_08756_),
    .A1(net210),
    .A2(net5180));
 sg13g2_nand2_1 _12881_ (.Y(_08757_),
    .A(net249),
    .B(net5010));
 sg13g2_o21ai_1 _12882_ (.B1(_08757_),
    .Y(_00154_),
    .A1(net5010),
    .A2(_08756_));
 sg13g2_nand2_1 _12883_ (.Y(_08758_),
    .A(_07784_),
    .B(net5185));
 sg13g2_o21ai_1 _12884_ (.B1(_08758_),
    .Y(_08759_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .A2(net5185));
 sg13g2_nand2_1 _12885_ (.Y(_08760_),
    .A(net210),
    .B(net5010));
 sg13g2_o21ai_1 _12886_ (.B1(_08760_),
    .Y(_00155_),
    .A1(net5011),
    .A2(_08759_));
 sg13g2_nand2b_1 _12887_ (.Y(_08761_),
    .B(net5186),
    .A_N(net6466));
 sg13g2_o21ai_1 _12888_ (.B1(_08761_),
    .Y(_08762_),
    .A1(net1341),
    .A2(net5186));
 sg13g2_nand2_2 _12889_ (.Y(_08763_),
    .A(net2008),
    .B(net5011));
 sg13g2_o21ai_1 _12890_ (.B1(_08763_),
    .Y(_00156_),
    .A1(net5023),
    .A2(_08762_));
 sg13g2_mux2_1 _12891_ (.A0(net229),
    .A1(net6464),
    .S(net5186),
    .X(_08764_));
 sg13g2_mux2_1 _12892_ (.A0(_08764_),
    .A1(net1341),
    .S(net5023),
    .X(_00157_));
 sg13g2_nand2b_1 _12893_ (.Y(_08765_),
    .B(net5186),
    .A_N(net6462));
 sg13g2_o21ai_1 _12894_ (.B1(_08765_),
    .Y(_08766_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[28] ),
    .A2(net5187));
 sg13g2_nand2_1 _12895_ (.Y(_08767_),
    .A(net229),
    .B(net5016));
 sg13g2_o21ai_1 _12896_ (.B1(_08767_),
    .Y(_00158_),
    .A1(net5017),
    .A2(_08766_));
 sg13g2_mux2_1 _12897_ (.A0(net262),
    .A1(net6460),
    .S(net5187),
    .X(_08768_));
 sg13g2_mux2_1 _12898_ (.A0(_08768_),
    .A1(net1737),
    .S(net5016),
    .X(_00159_));
 sg13g2_nand2b_1 _12899_ (.Y(_08769_),
    .B(net5186),
    .A_N(net6458));
 sg13g2_o21ai_1 _12900_ (.B1(_08769_),
    .Y(_08770_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .A2(net5186));
 sg13g2_nand2_1 _12901_ (.Y(_08771_),
    .A(net262),
    .B(net5016));
 sg13g2_o21ai_1 _12902_ (.B1(_08771_),
    .Y(_00161_),
    .A1(net5017),
    .A2(_08770_));
 sg13g2_nand2b_1 _12903_ (.Y(_08772_),
    .B(net5186),
    .A_N(net6455));
 sg13g2_o21ai_1 _12904_ (.B1(_08772_),
    .Y(_08773_),
    .A1(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .A2(net5186));
 sg13g2_nand2_1 _12905_ (.Y(_08774_),
    .A(net365),
    .B(net5017));
 sg13g2_o21ai_1 _12906_ (.B1(_08774_),
    .Y(_00162_),
    .A1(net5017),
    .A2(_08773_));
 sg13g2_nand2b_2 _12907_ (.Y(_08775_),
    .B(\soc_inst.spi_inst.spi_clk_en ),
    .A_N(_08693_));
 sg13g2_inv_1 _12908_ (.Y(_08776_),
    .A(_08775_));
 sg13g2_nor2_1 _12909_ (.A(net167),
    .B(_08775_),
    .Y(_00128_));
 sg13g2_o21ai_1 _12910_ (.B1(_08776_),
    .Y(_08777_),
    .A1(net167),
    .A2(net577));
 sg13g2_a21oi_1 _12911_ (.A1(net167),
    .A2(net577),
    .Y(_00129_),
    .B1(_08777_));
 sg13g2_and3_1 _12912_ (.X(_08778_),
    .A(net167),
    .B(net577),
    .C(net760));
 sg13g2_a21oi_1 _12913_ (.A1(net167),
    .A2(net577),
    .Y(_08779_),
    .B1(net760));
 sg13g2_nor3_1 _12914_ (.A(_08775_),
    .B(_08778_),
    .C(_08779_),
    .Y(_00130_));
 sg13g2_and2_1 _12915_ (.A(net1901),
    .B(_08778_),
    .X(_08780_));
 sg13g2_nor2_1 _12916_ (.A(net1901),
    .B(_08778_),
    .Y(_08781_));
 sg13g2_nor3_1 _12917_ (.A(_08775_),
    .B(_08780_),
    .C(_08781_),
    .Y(_00131_));
 sg13g2_and2_1 _12918_ (.A(net2777),
    .B(_08780_),
    .X(_08782_));
 sg13g2_nor2_1 _12919_ (.A(net2777),
    .B(_08780_),
    .Y(_08783_));
 sg13g2_nor3_1 _12920_ (.A(_08775_),
    .B(_08782_),
    .C(_08783_),
    .Y(_00132_));
 sg13g2_nor2_1 _12921_ (.A(net2206),
    .B(_08782_),
    .Y(_08784_));
 sg13g2_and2_1 _12922_ (.A(net2206),
    .B(_08782_),
    .X(_08785_));
 sg13g2_nor3_1 _12923_ (.A(_08775_),
    .B(net2207),
    .C(_08785_),
    .Y(_00133_));
 sg13g2_nor2_1 _12924_ (.A(net2620),
    .B(_08785_),
    .Y(_08786_));
 sg13g2_and2_1 _12925_ (.A(net2620),
    .B(_08785_),
    .X(_08787_));
 sg13g2_nor3_1 _12926_ (.A(_08775_),
    .B(net2621),
    .C(_08787_),
    .Y(_00134_));
 sg13g2_o21ai_1 _12927_ (.B1(_08776_),
    .Y(_08788_),
    .A1(net462),
    .A2(_08787_));
 sg13g2_a21oi_1 _12928_ (.A1(net462),
    .A2(_08787_),
    .Y(_00135_),
    .B1(_08788_));
 sg13g2_a21oi_1 _12929_ (.A1(\soc_inst.spi_inst.cpol ),
    .A2(_07897_),
    .Y(_08789_),
    .B1(_08696_));
 sg13g2_o21ai_1 _12930_ (.B1(_08789_),
    .Y(_00136_),
    .A1(_07898_),
    .A2(_08775_));
 sg13g2_nor3_2 _12931_ (.A(\soc_inst.core_mem_addr[1] ),
    .B(\soc_inst.core_mem_addr[0] ),
    .C(net6210),
    .Y(_08790_));
 sg13g2_and2_1 _12932_ (.A(_07887_),
    .B(net6108),
    .X(_08791_));
 sg13g2_nand2_2 _12933_ (.Y(_08792_),
    .A(_07887_),
    .B(net6109));
 sg13g2_nor2b_2 _12934_ (.A(\soc_inst.core_mem_addr[12] ),
    .B_N(_08235_),
    .Y(_08793_));
 sg13g2_nand3_1 _12935_ (.B(_08229_),
    .C(_08793_),
    .A(net6204),
    .Y(_08794_));
 sg13g2_nor2_2 _12936_ (.A(_08792_),
    .B(_08794_),
    .Y(_08795_));
 sg13g2_a21oi_1 _12937_ (.A1(net6468),
    .A2(_08795_),
    .Y(_08796_),
    .B1(net1565));
 sg13g2_nand2b_1 _12938_ (.Y(_08797_),
    .B(net6539),
    .A_N(net6535));
 sg13g2_nor2_2 _12939_ (.A(net6537),
    .B(_08797_),
    .Y(_08798_));
 sg13g2_nand2_1 _12940_ (.Y(_08799_),
    .A(net6534),
    .B(_08798_));
 sg13g2_xnor2_1 _12941_ (.Y(_08800_),
    .A(_00229_),
    .B(\soc_inst.i2c_inst.clk_cnt[3] ));
 sg13g2_xor2_1 _12942_ (.B(\soc_inst.i2c_inst.clk_cnt[5] ),
    .A(\soc_inst.i2c_inst.prescale_reg[5] ),
    .X(_08801_));
 sg13g2_nor2_1 _12943_ (.A(_08800_),
    .B(_08801_),
    .Y(_08802_));
 sg13g2_xor2_1 _12944_ (.B(\soc_inst.i2c_inst.clk_cnt[0] ),
    .A(_00226_),
    .X(_08803_));
 sg13g2_xnor2_1 _12945_ (.Y(_08804_),
    .A(_00228_),
    .B(\soc_inst.i2c_inst.clk_cnt[2] ));
 sg13g2_inv_1 _12946_ (.Y(_08805_),
    .A(_08804_));
 sg13g2_xnor2_1 _12947_ (.Y(_08806_),
    .A(_00230_),
    .B(\soc_inst.i2c_inst.clk_cnt[4] ));
 sg13g2_inv_1 _12948_ (.Y(_08807_),
    .A(_08806_));
 sg13g2_xor2_1 _12949_ (.B(\soc_inst.i2c_inst.clk_cnt[6] ),
    .A(\soc_inst.i2c_inst.prescale_reg[6] ),
    .X(_08808_));
 sg13g2_xnor2_1 _12950_ (.Y(_08809_),
    .A(_00231_),
    .B(\soc_inst.i2c_inst.clk_cnt[7] ));
 sg13g2_xnor2_1 _12951_ (.Y(_08810_),
    .A(_00227_),
    .B(\soc_inst.i2c_inst.clk_cnt[1] ));
 sg13g2_nor4_1 _12952_ (.A(_08806_),
    .B(_08808_),
    .C(_08809_),
    .D(_08810_),
    .Y(_08811_));
 sg13g2_nand4_1 _12953_ (.B(_08803_),
    .C(_08805_),
    .A(_08802_),
    .Y(_08812_),
    .D(_08811_));
 sg13g2_nor4_1 _12954_ (.A(_08804_),
    .B(_08808_),
    .C(_08809_),
    .D(_08810_),
    .Y(_08813_));
 sg13g2_nand4_1 _12955_ (.B(_08803_),
    .C(_08807_),
    .A(_08802_),
    .Y(_08814_),
    .D(_08813_));
 sg13g2_nor2_1 _12956_ (.A(_08799_),
    .B(net5565),
    .Y(_08815_));
 sg13g2_nor2_1 _12957_ (.A(_08800_),
    .B(_08809_),
    .Y(_08816_));
 sg13g2_nor4_1 _12958_ (.A(_08801_),
    .B(_08804_),
    .C(_08808_),
    .D(_08810_),
    .Y(_08817_));
 sg13g2_nand4_1 _12959_ (.B(_08807_),
    .C(_08816_),
    .A(_08803_),
    .Y(_08818_),
    .D(_08817_));
 sg13g2_nor2_1 _12960_ (.A(net1566),
    .B(_08815_),
    .Y(_00105_));
 sg13g2_nor2_2 _12961_ (.A(net6211),
    .B(_08671_),
    .Y(_08819_));
 sg13g2_nand3_1 _12962_ (.B(net6210),
    .C(_08668_),
    .A(_07887_),
    .Y(_08820_));
 sg13g2_nor2_1 _12963_ (.A(_08794_),
    .B(net6051),
    .Y(_08821_));
 sg13g2_nand2b_2 _12964_ (.Y(_08822_),
    .B(net5563),
    .A_N(_08794_));
 sg13g2_nand2_1 _12965_ (.Y(_08823_),
    .A(net82),
    .B(net5175));
 sg13g2_a21oi_1 _12966_ (.A1(net6470),
    .A2(_08795_),
    .Y(_08824_),
    .B1(_08823_));
 sg13g2_nor2b_2 _12967_ (.A(net6534),
    .B_N(net6538),
    .Y(_08825_));
 sg13g2_nand2b_1 _12968_ (.Y(_08826_),
    .B(net6537),
    .A_N(net6534));
 sg13g2_nor2b_2 _12969_ (.A(net6534),
    .B_N(net6535),
    .Y(_08827_));
 sg13g2_nand2b_2 _12970_ (.Y(_08828_),
    .B(net6535),
    .A_N(\soc_inst.i2c_inst.state[3] ));
 sg13g2_nand2_2 _12971_ (.Y(_08829_),
    .A(net6537),
    .B(_08827_));
 sg13g2_inv_1 _12972_ (.Y(_08830_),
    .A(_08829_));
 sg13g2_nor2_2 _12973_ (.A(net6539),
    .B(_08829_),
    .Y(_08831_));
 sg13g2_nor2b_1 _12974_ (.A(_08812_),
    .B_N(_08831_),
    .Y(_08832_));
 sg13g2_or2_1 _12975_ (.X(_00106_),
    .B(net5367),
    .A(_08824_));
 sg13g2_nor2_1 _12976_ (.A(\soc_inst.i2c_inst.data_reg[0] ),
    .B(net5178),
    .Y(_08833_));
 sg13g2_nor2_1 _12977_ (.A(net6470),
    .B(_08822_),
    .Y(_08834_));
 sg13g2_nor3_1 _12978_ (.A(net5368),
    .B(_08833_),
    .C(_08834_),
    .Y(_08835_));
 sg13g2_a21o_1 _12979_ (.A2(net5368),
    .A1(net2250),
    .B1(_08835_),
    .X(_00097_));
 sg13g2_nor2_1 _12980_ (.A(\soc_inst.i2c_inst.data_reg[1] ),
    .B(net5177),
    .Y(_08836_));
 sg13g2_nor2_1 _12981_ (.A(net6468),
    .B(net5175),
    .Y(_08837_));
 sg13g2_nor3_1 _12982_ (.A(net5367),
    .B(_08836_),
    .C(_08837_),
    .Y(_08838_));
 sg13g2_a21o_1 _12983_ (.A2(net5367),
    .A1(net1718),
    .B1(_08838_),
    .X(_00098_));
 sg13g2_nor2_1 _12984_ (.A(\soc_inst.i2c_inst.data_reg[2] ),
    .B(net5176),
    .Y(_08839_));
 sg13g2_nor2_1 _12985_ (.A(net6465),
    .B(net5175),
    .Y(_08840_));
 sg13g2_nor3_1 _12986_ (.A(net5366),
    .B(_08839_),
    .C(_08840_),
    .Y(_08841_));
 sg13g2_a21o_1 _12987_ (.A2(net5366),
    .A1(net1836),
    .B1(_08841_),
    .X(_00099_));
 sg13g2_nor2_1 _12988_ (.A(\soc_inst.i2c_inst.data_reg[3] ),
    .B(net5176),
    .Y(_08842_));
 sg13g2_nor2_1 _12989_ (.A(net6463),
    .B(net5175),
    .Y(_08843_));
 sg13g2_nor3_1 _12990_ (.A(net5366),
    .B(_08842_),
    .C(_08843_),
    .Y(_08844_));
 sg13g2_a21o_1 _12991_ (.A2(net5366),
    .A1(net2017),
    .B1(_08844_),
    .X(_00100_));
 sg13g2_nor2_1 _12992_ (.A(\soc_inst.i2c_inst.data_reg[4] ),
    .B(net5176),
    .Y(_08845_));
 sg13g2_nor2_1 _12993_ (.A(net6461),
    .B(net5175),
    .Y(_08846_));
 sg13g2_nor3_1 _12994_ (.A(net5366),
    .B(_08845_),
    .C(_08846_),
    .Y(_08847_));
 sg13g2_a21o_1 _12995_ (.A2(net5366),
    .A1(net2086),
    .B1(_08847_),
    .X(_00101_));
 sg13g2_nor2_1 _12996_ (.A(\soc_inst.i2c_inst.data_reg[5] ),
    .B(net5176),
    .Y(_08848_));
 sg13g2_nor2_1 _12997_ (.A(net6459),
    .B(net5175),
    .Y(_08849_));
 sg13g2_nor3_1 _12998_ (.A(net5366),
    .B(_08848_),
    .C(_08849_),
    .Y(_08850_));
 sg13g2_a21o_1 _12999_ (.A2(net5366),
    .A1(net2199),
    .B1(_08850_),
    .X(_00102_));
 sg13g2_nor2_1 _13000_ (.A(\soc_inst.i2c_inst.data_reg[6] ),
    .B(net5177),
    .Y(_08851_));
 sg13g2_nor2_1 _13001_ (.A(net6457),
    .B(net5175),
    .Y(_08852_));
 sg13g2_nor3_1 _13002_ (.A(net5367),
    .B(_08851_),
    .C(_08852_),
    .Y(_08853_));
 sg13g2_a21o_1 _13003_ (.A2(net5367),
    .A1(net1912),
    .B1(_08853_),
    .X(_00103_));
 sg13g2_nor2_1 _13004_ (.A(\soc_inst.i2c_inst.data_reg[7] ),
    .B(net5178),
    .Y(_08854_));
 sg13g2_nor2_1 _13005_ (.A(net6455),
    .B(net5175),
    .Y(_08855_));
 sg13g2_nor3_1 _13006_ (.A(net5368),
    .B(_08854_),
    .C(_08855_),
    .Y(_08856_));
 sg13g2_a21o_1 _13007_ (.A2(net5368),
    .A1(net2049),
    .B1(_08856_),
    .X(_00104_));
 sg13g2_nand2_1 _13008_ (.Y(_08857_),
    .A(\soc_inst.i2c_ena ),
    .B(_08812_));
 sg13g2_nor2_1 _13009_ (.A(net216),
    .B(net5365),
    .Y(_00089_));
 sg13g2_xnor2_1 _13010_ (.Y(_08858_),
    .A(net216),
    .B(net2594));
 sg13g2_nor2_1 _13011_ (.A(net5365),
    .B(_08858_),
    .Y(_00090_));
 sg13g2_and3_1 _13012_ (.X(_08859_),
    .A(net216),
    .B(net3407),
    .C(net1230));
 sg13g2_a21oi_1 _13013_ (.A1(net216),
    .A2(\soc_inst.i2c_inst.clk_cnt[1] ),
    .Y(_08860_),
    .B1(net1230));
 sg13g2_nor3_1 _13014_ (.A(net5365),
    .B(_08859_),
    .C(net1231),
    .Y(_00091_));
 sg13g2_and2_1 _13015_ (.A(net2073),
    .B(_08859_),
    .X(_08861_));
 sg13g2_nor2_1 _13016_ (.A(net2073),
    .B(_08859_),
    .Y(_08862_));
 sg13g2_nor3_1 _13017_ (.A(net5365),
    .B(_08861_),
    .C(net2074),
    .Y(_00092_));
 sg13g2_and2_1 _13018_ (.A(net2244),
    .B(_08861_),
    .X(_08863_));
 sg13g2_nor2_1 _13019_ (.A(net2244),
    .B(_08861_),
    .Y(_08864_));
 sg13g2_nor3_1 _13020_ (.A(net5365),
    .B(_08863_),
    .C(_08864_),
    .Y(_00093_));
 sg13g2_and2_1 _13021_ (.A(net2569),
    .B(_08863_),
    .X(_08865_));
 sg13g2_nor2_1 _13022_ (.A(net2569),
    .B(_08863_),
    .Y(_08866_));
 sg13g2_nor3_1 _13023_ (.A(net5365),
    .B(_08865_),
    .C(_08866_),
    .Y(_00094_));
 sg13g2_nor2_1 _13024_ (.A(net2529),
    .B(_08865_),
    .Y(_08867_));
 sg13g2_and2_1 _13025_ (.A(net2529),
    .B(_08865_),
    .X(_08868_));
 sg13g2_nor3_1 _13026_ (.A(net5365),
    .B(net2530),
    .C(_08868_),
    .Y(_00095_));
 sg13g2_xnor2_1 _13027_ (.Y(_08869_),
    .A(net2560),
    .B(_08868_));
 sg13g2_nor2_1 _13028_ (.A(net5365),
    .B(net2561),
    .Y(_00096_));
 sg13g2_nand2_1 _13029_ (.Y(_08870_),
    .A(_00237_),
    .B(\soc_inst.pwm_inst.channel_counter[0][3] ));
 sg13g2_nor2_1 _13030_ (.A(_00235_),
    .B(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .Y(_08871_));
 sg13g2_nor2_1 _13031_ (.A(_00234_),
    .B(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .Y(_08872_));
 sg13g2_a22oi_1 _13032_ (.Y(_08873_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .B2(_00235_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .A1(_00236_));
 sg13g2_o21ai_1 _13033_ (.B1(_08873_),
    .Y(_08874_),
    .A1(_08871_),
    .A2(_08872_));
 sg13g2_o21ai_1 _13034_ (.B1(_08874_),
    .Y(_08875_),
    .A1(_00236_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][2] ));
 sg13g2_a22oi_1 _13035_ (.Y(_08876_),
    .B1(_08870_),
    .B2(_08875_),
    .A2(_07947_),
    .A1(_07793_));
 sg13g2_o21ai_1 _13036_ (.B1(_08876_),
    .Y(_08877_),
    .A1(_00237_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][3] ));
 sg13g2_a22oi_1 _13037_ (.Y(_08878_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .B2(_00238_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .A1(_00239_));
 sg13g2_or2_1 _13038_ (.X(_08879_),
    .B(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .A(_00240_));
 sg13g2_o21ai_1 _13039_ (.B1(_08879_),
    .Y(_08880_),
    .A1(_00239_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][5] ));
 sg13g2_a21oi_1 _13040_ (.A1(_08877_),
    .A2(_08878_),
    .Y(_08881_),
    .B1(_08880_));
 sg13g2_a221oi_1 _13041_ (.B2(_00240_),
    .C1(_08881_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .A1(_00241_),
    .Y(_08882_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][7] ));
 sg13g2_nor2_1 _13042_ (.A(_00241_),
    .B(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .Y(_08883_));
 sg13g2_nor2_1 _13043_ (.A(_00243_),
    .B(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .Y(_08884_));
 sg13g2_nor2_1 _13044_ (.A(_00242_),
    .B(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .Y(_08885_));
 sg13g2_nor4_1 _13045_ (.A(_08882_),
    .B(_08883_),
    .C(_08884_),
    .D(_08885_),
    .Y(_08886_));
 sg13g2_a221oi_1 _13046_ (.B2(_00242_),
    .C1(_08886_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .A1(_00243_),
    .Y(_08887_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][9] ));
 sg13g2_nand3_1 _13047_ (.B(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .C(_08884_),
    .A(_00242_),
    .Y(_08888_));
 sg13g2_o21ai_1 _13048_ (.B1(_08888_),
    .Y(_08889_),
    .A1(_00244_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][10] ));
 sg13g2_a22oi_1 _13049_ (.Y(_08890_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .B2(_00244_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .A1(_00245_));
 sg13g2_o21ai_1 _13050_ (.B1(_08890_),
    .Y(_08891_),
    .A1(_08887_),
    .A2(_08889_));
 sg13g2_nor2_1 _13051_ (.A(net2055),
    .B(net1071),
    .Y(_08892_));
 sg13g2_or2_1 _13052_ (.X(_08893_),
    .B(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .A(_00245_));
 sg13g2_o21ai_1 _13053_ (.B1(_08893_),
    .Y(_08894_),
    .A1(_00246_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][12] ));
 sg13g2_a22oi_1 _13054_ (.Y(_08895_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .B2(_00246_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .A1(_00247_));
 sg13g2_a22oi_1 _13055_ (.Y(_08896_),
    .B1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .B2(_00248_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .A1(_00249_));
 sg13g2_nor2_1 _13056_ (.A(_00248_),
    .B(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .Y(_08897_));
 sg13g2_nor2_1 _13057_ (.A(_00247_),
    .B(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .Y(_08898_));
 sg13g2_nand2b_1 _13058_ (.Y(_08899_),
    .B(_08896_),
    .A_N(_08897_));
 sg13g2_nor4_1 _13059_ (.A(_08892_),
    .B(_08894_),
    .C(_08898_),
    .D(_08899_),
    .Y(_08900_));
 sg13g2_and3_1 _13060_ (.X(_08901_),
    .A(_08891_),
    .B(_08895_),
    .C(_08900_));
 sg13g2_or3_1 _13061_ (.A(_08895_),
    .B(_08897_),
    .C(_08898_),
    .X(_08902_));
 sg13g2_a21oi_1 _13062_ (.A1(_08896_),
    .A2(_08902_),
    .Y(_08903_),
    .B1(_08892_));
 sg13g2_nor2_1 _13063_ (.A(net6206),
    .B(net6064),
    .Y(_08904_));
 sg13g2_nand2_1 _13064_ (.Y(_08905_),
    .A(net6211),
    .B(net6109));
 sg13g2_and2_1 _13065_ (.A(_08667_),
    .B(net5559),
    .X(_08906_));
 sg13g2_nand2_2 _13066_ (.Y(_08907_),
    .A(_08667_),
    .B(net5559));
 sg13g2_and4_1 _13067_ (.A(net6204),
    .B(\soc_inst.core_mem_addr[13] ),
    .C(_08230_),
    .D(_08675_),
    .X(_08908_));
 sg13g2_and2_1 _13068_ (.A(net5364),
    .B(_08908_),
    .X(_08909_));
 sg13g2_or4_1 _13069_ (.A(_07949_),
    .B(_08901_),
    .C(_08903_),
    .D(net5170),
    .X(_08910_));
 sg13g2_nor2_1 _13070_ (.A(net264),
    .B(net4740),
    .Y(_00111_));
 sg13g2_xnor2_1 _13071_ (.Y(_08911_),
    .A(net3025),
    .B(net264));
 sg13g2_nor2_1 _13072_ (.A(net4740),
    .B(_08911_),
    .Y(_00118_));
 sg13g2_and3_1 _13073_ (.X(_08912_),
    .A(net2638),
    .B(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .C(net264));
 sg13g2_a21oi_1 _13074_ (.A1(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .A2(net264),
    .Y(_08913_),
    .B1(net2638));
 sg13g2_nor3_1 _13075_ (.A(net4740),
    .B(_08912_),
    .C(net2639),
    .Y(_00119_));
 sg13g2_nor2_1 _13076_ (.A(net2872),
    .B(_08912_),
    .Y(_08914_));
 sg13g2_and2_1 _13077_ (.A(net2872),
    .B(_08912_),
    .X(_08915_));
 sg13g2_nor3_1 _13078_ (.A(net4740),
    .B(net2873),
    .C(_08915_),
    .Y(_00120_));
 sg13g2_and2_1 _13079_ (.A(net2525),
    .B(_08915_),
    .X(_08916_));
 sg13g2_nor2_1 _13080_ (.A(net2525),
    .B(_08915_),
    .Y(_08917_));
 sg13g2_nor3_1 _13081_ (.A(net4740),
    .B(_08916_),
    .C(net2526),
    .Y(_00121_));
 sg13g2_nor2_1 _13082_ (.A(net2691),
    .B(_08916_),
    .Y(_08918_));
 sg13g2_and2_1 _13083_ (.A(net2691),
    .B(_08916_),
    .X(_08919_));
 sg13g2_nor3_1 _13084_ (.A(_08910_),
    .B(net2692),
    .C(_08919_),
    .Y(_00122_));
 sg13g2_and2_1 _13085_ (.A(net3013),
    .B(_08919_),
    .X(_08920_));
 sg13g2_nor2_1 _13086_ (.A(net3013),
    .B(_08919_),
    .Y(_08921_));
 sg13g2_nor3_1 _13087_ (.A(net4740),
    .B(_08920_),
    .C(_08921_),
    .Y(_00123_));
 sg13g2_and2_1 _13088_ (.A(net2929),
    .B(_08920_),
    .X(_08922_));
 sg13g2_nor2_1 _13089_ (.A(net2929),
    .B(_08920_),
    .Y(_08923_));
 sg13g2_nor3_1 _13090_ (.A(net4739),
    .B(_08922_),
    .C(net2930),
    .Y(_00124_));
 sg13g2_nor2_1 _13091_ (.A(net2940),
    .B(_08922_),
    .Y(_08924_));
 sg13g2_and2_1 _13092_ (.A(net2940),
    .B(_08922_),
    .X(_08925_));
 sg13g2_nor3_1 _13093_ (.A(net4739),
    .B(net2941),
    .C(_08925_),
    .Y(_00125_));
 sg13g2_xnor2_1 _13094_ (.Y(_08926_),
    .A(net3143),
    .B(_08925_));
 sg13g2_nor2_1 _13095_ (.A(net4740),
    .B(_08926_),
    .Y(_00126_));
 sg13g2_a21oi_1 _13096_ (.A1(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .A2(_08925_),
    .Y(_08927_),
    .B1(net2471));
 sg13g2_and3_1 _13097_ (.X(_08928_),
    .A(net2471),
    .B(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .C(_08925_));
 sg13g2_nor3_1 _13098_ (.A(net4739),
    .B(net2472),
    .C(_08928_),
    .Y(_00112_));
 sg13g2_and2_1 _13099_ (.A(net2787),
    .B(_08928_),
    .X(_08929_));
 sg13g2_nor2_1 _13100_ (.A(net2787),
    .B(_08928_),
    .Y(_08930_));
 sg13g2_nor3_1 _13101_ (.A(net4739),
    .B(_08929_),
    .C(net2788),
    .Y(_00113_));
 sg13g2_and2_1 _13102_ (.A(net3022),
    .B(_08929_),
    .X(_08931_));
 sg13g2_nor2_1 _13103_ (.A(net3022),
    .B(_08929_),
    .Y(_08932_));
 sg13g2_nor3_1 _13104_ (.A(net4739),
    .B(_08931_),
    .C(_08932_),
    .Y(_00114_));
 sg13g2_and2_1 _13105_ (.A(net2994),
    .B(_08931_),
    .X(_08933_));
 sg13g2_nor2_1 _13106_ (.A(net2994),
    .B(_08931_),
    .Y(_08934_));
 sg13g2_nor3_1 _13107_ (.A(net4739),
    .B(_08933_),
    .C(net2995),
    .Y(_00115_));
 sg13g2_xnor2_1 _13108_ (.Y(_08935_),
    .A(net3188),
    .B(_08933_));
 sg13g2_nor2_1 _13109_ (.A(net4739),
    .B(_08935_),
    .Y(_00116_));
 sg13g2_a21oi_1 _13110_ (.A1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .A2(_08933_),
    .Y(_08936_),
    .B1(net1071));
 sg13g2_nor2_1 _13111_ (.A(net4739),
    .B(net1072),
    .Y(_00117_));
 sg13g2_nand3b_1 _13112_ (.B(_08418_),
    .C(_00250_),
    .Y(\soc_inst.flash_cs_n ),
    .A_N(net6542));
 sg13g2_nand3_1 _13113_ (.B(\soc_inst.core_mem_addr[24] ),
    .C(_08653_),
    .A(_00250_),
    .Y(_08937_));
 sg13g2_nor4_1 _13114_ (.A(\soc_inst.core_mem_addr[25] ),
    .B(\soc_inst.core_mem_addr[27] ),
    .C(\soc_inst.core_mem_addr[26] ),
    .D(_08937_),
    .Y(_08938_));
 sg13g2_nand2_1 _13115_ (.Y(\soc_inst.mem_ctrl.ram_cs_n ),
    .A(_08416_),
    .B(_08938_));
 sg13g2_nor2_1 _13116_ (.A(_08247_),
    .B(_08386_),
    .Y(_08939_));
 sg13g2_a21oi_1 _13117_ (.A1(_08385_),
    .A2(_08939_),
    .Y(_00108_),
    .B1(net5195));
 sg13g2_nor3_1 _13118_ (.A(net1222),
    .B(_08250_),
    .C(_08292_),
    .Y(_00107_));
 sg13g2_nor2_1 _13119_ (.A(_00262_),
    .B(_00261_),
    .Y(_08940_));
 sg13g2_nand2b_1 _13120_ (.Y(_08941_),
    .B(_08940_),
    .A_N(\soc_inst.cpu_core.ex_instr[3] ));
 sg13g2_nor2_1 _13121_ (.A(\soc_inst.cpu_core.ex_instr[2] ),
    .B(_08941_),
    .Y(_08942_));
 sg13g2_nor2_1 _13122_ (.A(_07791_),
    .B(\soc_inst.cpu_core.ex_instr[6] ),
    .Y(_08943_));
 sg13g2_nand2_2 _13123_ (.Y(_08944_),
    .A(_08942_),
    .B(_08943_));
 sg13g2_nand3b_1 _13124_ (.B(\soc_inst.cpu_core.ex_alu_result[0] ),
    .C(\soc_inst.cpu_core.ex_funct3[0] ),
    .Y(_08945_),
    .A_N(\soc_inst.cpu_core.ex_funct3[1] ));
 sg13g2_nor2b_1 _13125_ (.A(\soc_inst.cpu_core.ex_funct3[0] ),
    .B_N(\soc_inst.cpu_core.ex_funct3[1] ),
    .Y(_08946_));
 sg13g2_o21ai_1 _13126_ (.B1(_08946_),
    .Y(_08947_),
    .A1(\soc_inst.cpu_core.ex_alu_result[1] ),
    .A2(\soc_inst.cpu_core.ex_alu_result[0] ));
 sg13g2_a21o_1 _13127_ (.A2(_08947_),
    .A1(_08945_),
    .B1(\soc_inst.cpu_core.ex_funct3[2] ),
    .X(_08948_));
 sg13g2_o21ai_1 _13128_ (.B1(_08948_),
    .Y(_08949_),
    .A1(net6213),
    .A2(_08945_));
 sg13g2_nor2b_2 _13129_ (.A(_08944_),
    .B_N(_08949_),
    .Y(_08950_));
 sg13g2_nand2b_1 _13130_ (.Y(_08951_),
    .B(_08949_),
    .A_N(_08944_));
 sg13g2_nand2_1 _13131_ (.Y(_08952_),
    .A(\soc_inst.cpu_core.ex_instr[2] ),
    .B(_08940_));
 sg13g2_nand2_1 _13132_ (.Y(_08953_),
    .A(_08941_),
    .B(_08952_));
 sg13g2_and4_1 _13133_ (.A(_00263_),
    .B(net6213),
    .C(\soc_inst.cpu_core.ex_instr[6] ),
    .D(_08953_),
    .X(_08954_));
 sg13g2_nand4_1 _13134_ (.B(net6213),
    .C(\soc_inst.cpu_core.ex_instr[6] ),
    .A(_00263_),
    .Y(_08955_),
    .D(_08953_));
 sg13g2_nor2b_1 _13135_ (.A(net6213),
    .B_N(\soc_inst.cpu_core.ex_instr[3] ),
    .Y(_08956_));
 sg13g2_nand4_1 _13136_ (.B(_08940_),
    .C(_08943_),
    .A(\soc_inst.cpu_core.ex_instr[2] ),
    .Y(_08957_),
    .D(_08956_));
 sg13g2_nand3_1 _13137_ (.B(net5354),
    .C(_08957_),
    .A(_08944_),
    .Y(_08958_));
 sg13g2_nand2_1 _13138_ (.Y(_08959_),
    .A(net6213),
    .B(_08942_));
 sg13g2_nand2_1 _13139_ (.Y(_08960_),
    .A(\soc_inst.cpu_core.ex_instr[6] ),
    .B(_08959_));
 sg13g2_nor2_1 _13140_ (.A(_00263_),
    .B(_08941_),
    .Y(_08961_));
 sg13g2_a21oi_1 _13141_ (.A1(_08960_),
    .A2(_08961_),
    .Y(_08962_),
    .B1(_08958_));
 sg13g2_a21o_1 _13142_ (.A2(_08961_),
    .A1(_08960_),
    .B1(_08958_),
    .X(_08963_));
 sg13g2_and2_1 _13143_ (.A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .B(net5360),
    .X(_08964_));
 sg13g2_nand2_1 _13144_ (.Y(_08965_),
    .A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .B(net5360));
 sg13g2_nand3_1 _13145_ (.B(net5071),
    .C(net5158),
    .A(net5167),
    .Y(_08966_));
 sg13g2_nor3_1 _13146_ (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .B(\soc_inst.cpu_core.ex_is_ebreak ),
    .C(net5047),
    .Y(_08967_));
 sg13g2_or3_1 _13147_ (.A(net2455),
    .B(net2562),
    .C(net5047),
    .X(_08968_));
 sg13g2_and3_2 _13148_ (.X(_00025_),
    .A(net6145),
    .B(net2128),
    .C(net5007));
 sg13g2_nor3_2 _13149_ (.A(net6370),
    .B(_08130_),
    .C(net4999),
    .Y(_00024_));
 sg13g2_nor2_1 _13150_ (.A(net6158),
    .B(net421),
    .Y(_08969_));
 sg13g2_or3_1 _13151_ (.A(_00025_),
    .B(_00024_),
    .C(_08969_),
    .X(_00026_));
 sg13g2_nor2_1 _13152_ (.A(net6480),
    .B(net4999),
    .Y(_08970_));
 sg13g2_nand2_2 _13153_ (.Y(_08971_),
    .A(_07871_),
    .B(net5002));
 sg13g2_nand2_1 _13154_ (.Y(_08972_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[9] ));
 sg13g2_nor2_1 _13155_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .Y(_08973_));
 sg13g2_nand2b_2 _13156_ (.Y(_08974_),
    .B(_08973_),
    .A_N(_08972_));
 sg13g2_nor2_1 _13157_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .Y(_08975_));
 sg13g2_or4_1 _13158_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .C(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .D(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .X(_08976_));
 sg13g2_nor2_2 _13159_ (.A(_08974_),
    .B(_08976_),
    .Y(_08977_));
 sg13g2_inv_1 _13160_ (.Y(_08978_),
    .A(_08977_));
 sg13g2_nor2_2 _13161_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .Y(_08979_));
 sg13g2_nor2_2 _13162_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .Y(_08980_));
 sg13g2_and2_1 _13163_ (.A(_08979_),
    .B(_08980_),
    .X(_08981_));
 sg13g2_nand2_2 _13164_ (.Y(_08982_),
    .A(_08979_),
    .B(_08980_));
 sg13g2_nor2_2 _13165_ (.A(net6298),
    .B(net6304),
    .Y(_08983_));
 sg13g2_or2_1 _13166_ (.X(_08984_),
    .B(net6304),
    .A(net6298));
 sg13g2_nor4_2 _13167_ (.A(_00259_),
    .B(_00258_),
    .C(\soc_inst.cpu_core.mem_instr[3] ),
    .Y(_08985_),
    .D(\soc_inst.cpu_core.mem_instr[2] ));
 sg13g2_nor2b_1 _13168_ (.A(_00260_),
    .B_N(\soc_inst.cpu_core.mem_instr[5] ),
    .Y(_08986_));
 sg13g2_nor2_2 _13169_ (.A(net6298),
    .B(net6289),
    .Y(_08987_));
 sg13g2_nor2_2 _13170_ (.A(net6289),
    .B(net6106),
    .Y(_08988_));
 sg13g2_nand2_1 _13171_ (.Y(_08989_),
    .A(net6168),
    .B(net6107));
 sg13g2_and4_1 _13172_ (.A(\soc_inst.cpu_core.mem_instr[6] ),
    .B(_08985_),
    .C(_08986_),
    .D(net6046),
    .X(_08990_));
 sg13g2_nand4_1 _13173_ (.B(_08985_),
    .C(_08986_),
    .A(\soc_inst.cpu_core.mem_instr[6] ),
    .Y(_08991_),
    .D(_08989_));
 sg13g2_nand2_1 _13174_ (.Y(_08992_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .B(_08979_));
 sg13g2_or2_1 _13175_ (.X(_08993_),
    .B(_08992_),
    .A(_08976_));
 sg13g2_nor2b_1 _13176_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .B_N(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .Y(_08994_));
 sg13g2_nand3_1 _13177_ (.B(_08981_),
    .C(_08994_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .Y(_08995_));
 sg13g2_a21oi_1 _13178_ (.A1(_08993_),
    .A2(_08995_),
    .Y(_08996_),
    .B1(_08972_));
 sg13g2_nand2_1 _13179_ (.Y(_08997_),
    .A(_08975_),
    .B(_08994_));
 sg13g2_nor4_1 _13180_ (.A(_07807_),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .C(_08982_),
    .D(_08997_),
    .Y(_08998_));
 sg13g2_nor2_1 _13181_ (.A(_08996_),
    .B(_08998_),
    .Y(_08999_));
 sg13g2_nor2b_1 _13182_ (.A(_08999_),
    .B_N(_08973_),
    .Y(_09000_));
 sg13g2_nand3b_1 _13183_ (.B(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .C(_08980_),
    .Y(_09001_),
    .A_N(\soc_inst.cpu_core.csr_file.csr_addr[3] ));
 sg13g2_nand3b_1 _13184_ (.B(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .C(_08975_),
    .Y(_09002_),
    .A_N(\soc_inst.cpu_core.csr_file.csr_addr[7] ));
 sg13g2_or2_1 _13185_ (.X(_09003_),
    .B(_09002_),
    .A(_08974_));
 sg13g2_nand2_1 _13186_ (.Y(_09004_),
    .A(_08980_),
    .B(_09003_));
 sg13g2_nand2_1 _13187_ (.Y(_09005_),
    .A(_08979_),
    .B(_09004_));
 sg13g2_nor4_1 _13188_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B(_07806_),
    .C(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .D(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .Y(_09006_));
 sg13g2_nand3_1 _13189_ (.B(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .C(_09006_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .Y(_09007_));
 sg13g2_or2_1 _13190_ (.X(_09008_),
    .B(_09007_),
    .A(_08972_));
 sg13g2_a22oi_1 _13191_ (.Y(_09009_),
    .B1(_09008_),
    .B2(_09003_),
    .A2(_09005_),
    .A1(_09001_));
 sg13g2_nor4_1 _13192_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .C(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .D(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .Y(_09010_));
 sg13g2_nand2_1 _13193_ (.Y(_09011_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[0] ));
 sg13g2_nand4_1 _13194_ (.B(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .C(_09010_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .Y(_09012_),
    .D(_09011_));
 sg13g2_nor2_1 _13195_ (.A(_08997_),
    .B(_09012_),
    .Y(_09013_));
 sg13g2_nor2_2 _13196_ (.A(_08976_),
    .B(_09012_),
    .Y(_09014_));
 sg13g2_nand2b_1 _13197_ (.Y(_09015_),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .A_N(\soc_inst.cpu_core.csr_file.csr_addr[1] ));
 sg13g2_nor3_1 _13198_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B(_07805_),
    .C(_09015_),
    .Y(_09016_));
 sg13g2_and2_1 _13199_ (.A(_08977_),
    .B(_09016_),
    .X(_09017_));
 sg13g2_inv_1 _13200_ (.Y(_09018_),
    .A(net5350));
 sg13g2_nor3_1 _13201_ (.A(net5544),
    .B(net5540),
    .C(net5350),
    .Y(_09019_));
 sg13g2_nor3_1 _13202_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .C(_09015_),
    .Y(_09020_));
 sg13g2_nand2_2 _13203_ (.Y(_09021_),
    .A(_08977_),
    .B(_09020_));
 sg13g2_nor2_2 _13204_ (.A(_08978_),
    .B(_08982_),
    .Y(_09022_));
 sg13g2_nand2_2 _13205_ (.Y(_09023_),
    .A(_08977_),
    .B(_08981_));
 sg13g2_nor2_1 _13206_ (.A(_08976_),
    .B(_09001_),
    .Y(_09024_));
 sg13g2_nor3_1 _13207_ (.A(_08974_),
    .B(_08976_),
    .C(_09001_),
    .Y(_09025_));
 sg13g2_nand2b_1 _13208_ (.Y(_09026_),
    .B(_09024_),
    .A_N(_08974_));
 sg13g2_nand4_1 _13209_ (.B(_09021_),
    .C(_09023_),
    .A(_09019_),
    .Y(_09027_),
    .D(_09026_));
 sg13g2_nor3_1 _13210_ (.A(_09000_),
    .B(_09009_),
    .C(_09027_),
    .Y(_09028_));
 sg13g2_nor2_2 _13211_ (.A(net5546),
    .B(_09028_),
    .Y(_09029_));
 sg13g2_nor3_1 _13212_ (.A(net6107),
    .B(net5546),
    .C(_09028_),
    .Y(_09030_));
 sg13g2_nor4_1 _13213_ (.A(_07807_),
    .B(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .C(_08982_),
    .D(_08997_),
    .Y(_09031_));
 sg13g2_o21ai_1 _13214_ (.B1(_08973_),
    .Y(_09032_),
    .A1(_08996_),
    .A2(_09031_));
 sg13g2_o21ai_1 _13215_ (.B1(_09021_),
    .Y(_09033_),
    .A1(_08978_),
    .A2(_09001_));
 sg13g2_nor2_1 _13216_ (.A(net5350),
    .B(_09033_),
    .Y(_09034_));
 sg13g2_nor4_1 _13217_ (.A(_09009_),
    .B(net5544),
    .C(net5540),
    .D(net5153),
    .Y(_09035_));
 sg13g2_nand3_1 _13218_ (.B(_09034_),
    .C(_09035_),
    .A(_09032_),
    .Y(_09036_));
 sg13g2_and3_2 _13219_ (.X(_09037_),
    .A(net6106),
    .B(net5551),
    .C(_09036_));
 sg13g2_and2_1 _13220_ (.A(net5156),
    .B(_09037_),
    .X(_09038_));
 sg13g2_nor3_1 _13221_ (.A(net5544),
    .B(net5539),
    .C(net5153),
    .Y(_09039_));
 sg13g2_nand4_1 _13222_ (.B(_09021_),
    .C(_09026_),
    .A(_09018_),
    .Y(_09040_),
    .D(_09039_));
 sg13g2_nor3_1 _13223_ (.A(_09000_),
    .B(_09009_),
    .C(_09040_),
    .Y(_09041_));
 sg13g2_nor2_2 _13224_ (.A(net5546),
    .B(_09041_),
    .Y(_09042_));
 sg13g2_nor3_2 _13225_ (.A(net6107),
    .B(net5546),
    .C(_09041_),
    .Y(_09043_));
 sg13g2_nand2_2 _13226_ (.Y(_09044_),
    .A(_08984_),
    .B(_09042_));
 sg13g2_o21ai_1 _13227_ (.B1(net4945),
    .Y(_09045_),
    .A1(_09023_),
    .A2(_09044_));
 sg13g2_inv_1 _13228_ (.Y(_09046_),
    .A(_09045_));
 sg13g2_nand2b_1 _13229_ (.Y(_09047_),
    .B(net6472),
    .A_N(net2626));
 sg13g2_o21ai_1 _13230_ (.B1(_09047_),
    .Y(_09048_),
    .A1(net6477),
    .A2(net3270));
 sg13g2_and2_1 _13231_ (.A(net6303),
    .B(net6304),
    .X(_09049_));
 sg13g2_or2_1 _13232_ (.X(_09050_),
    .B(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .A(net6293));
 sg13g2_o21ai_1 _13233_ (.B1(_09050_),
    .Y(_09051_),
    .A1(net6169),
    .A2(\soc_inst.cpu_core.mem_instr[18] ));
 sg13g2_inv_1 _13234_ (.Y(_09052_),
    .A(_09051_));
 sg13g2_nor2_1 _13235_ (.A(net6105),
    .B(_09051_),
    .Y(_09053_));
 sg13g2_and3_1 _13236_ (.X(_09054_),
    .A(net6301),
    .B(net3270),
    .C(_09051_));
 sg13g2_a21oi_1 _13237_ (.A1(net6301),
    .A2(_09051_),
    .Y(_09055_),
    .B1(_09053_));
 sg13g2_o21ai_1 _13238_ (.B1(net4792),
    .Y(_09056_),
    .A1(_09053_),
    .A2(_09054_));
 sg13g2_o21ai_1 _13239_ (.B1(_09056_),
    .Y(_00082_),
    .A1(_09045_),
    .A2(_09048_));
 sg13g2_and3_1 _13240_ (.X(_00063_),
    .A(net6159),
    .B(net515),
    .C(net4736));
 sg13g2_and3_1 _13241_ (.X(_00064_),
    .A(net6160),
    .B(net373),
    .C(net4737));
 sg13g2_and3_1 _13242_ (.X(_00065_),
    .A(net6160),
    .B(net391),
    .C(net4737));
 sg13g2_and3_1 _13243_ (.X(_00066_),
    .A(net6160),
    .B(net334),
    .C(net4737));
 sg13g2_and3_1 _13244_ (.X(_00067_),
    .A(net6162),
    .B(net124),
    .C(net4737));
 sg13g2_and3_1 _13245_ (.X(_00068_),
    .A(net6165),
    .B(net125),
    .C(net4737));
 sg13g2_and3_1 _13246_ (.X(_00069_),
    .A(net6159),
    .B(net118),
    .C(net4736));
 sg13g2_and3_1 _13247_ (.X(_00070_),
    .A(net6159),
    .B(net221),
    .C(net4736));
 sg13g2_and3_1 _13248_ (.X(_00071_),
    .A(net6160),
    .B(net349),
    .C(net4737));
 sg13g2_and3_1 _13249_ (.X(_00072_),
    .A(net6160),
    .B(net340),
    .C(net4737));
 sg13g2_and3_1 _13250_ (.X(_00073_),
    .A(net6160),
    .B(net265),
    .C(net4737));
 sg13g2_and3_1 _13251_ (.X(_00074_),
    .A(net6159),
    .B(net322),
    .C(net4736));
 sg13g2_and3_1 _13252_ (.X(_00075_),
    .A(net6161),
    .B(net146),
    .C(net4738));
 sg13g2_and3_1 _13253_ (.X(_00076_),
    .A(net6159),
    .B(net259),
    .C(net4736));
 sg13g2_and3_1 _13254_ (.X(_00077_),
    .A(net6161),
    .B(net143),
    .C(net4738));
 sg13g2_and3_1 _13255_ (.X(_00078_),
    .A(net6159),
    .B(net179),
    .C(net4736));
 sg13g2_and3_1 _13256_ (.X(_00079_),
    .A(net6159),
    .B(net151),
    .C(net4736));
 sg13g2_and3_1 _13257_ (.X(_00080_),
    .A(net6159),
    .B(net371),
    .C(net4736));
 sg13g2_and3_1 _13258_ (.X(_00081_),
    .A(net6161),
    .B(net180),
    .C(net4738));
 sg13g2_nor2b_1 _13259_ (.A(_09003_),
    .B_N(_09020_),
    .Y(_09057_));
 sg13g2_inv_4 _13260_ (.A(net5345),
    .Y(_09058_));
 sg13g2_nor2_2 _13261_ (.A(_09044_),
    .B(_09058_),
    .Y(_09059_));
 sg13g2_nand2_1 _13262_ (.Y(_09060_),
    .A(net4936),
    .B(net5345));
 sg13g2_nand2_2 _13263_ (.Y(_09061_),
    .A(net4948),
    .B(net4789));
 sg13g2_a21oi_1 _13264_ (.A1(net6480),
    .A2(_08082_),
    .Y(_09062_),
    .B1(net4999));
 sg13g2_a21oi_1 _13265_ (.A1(net1672),
    .A2(net4999),
    .Y(_09063_),
    .B1(_09062_));
 sg13g2_nand2b_2 _13266_ (.Y(_09064_),
    .B(net6303),
    .A_N(net6305));
 sg13g2_nor2b_1 _13267_ (.A(net6296),
    .B_N(net6304),
    .Y(_09065_));
 sg13g2_nand2_2 _13268_ (.Y(_09066_),
    .A(net6172),
    .B(net6304));
 sg13g2_and2_1 _13269_ (.A(_09064_),
    .B(_09066_),
    .X(_09067_));
 sg13g2_nand2_2 _13270_ (.Y(_09068_),
    .A(_09064_),
    .B(_09066_));
 sg13g2_or2_1 _13271_ (.X(_09069_),
    .B(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .A(net6293));
 sg13g2_o21ai_1 _13272_ (.B1(_09069_),
    .Y(_09070_),
    .A1(net6168),
    .A2(\soc_inst.cpu_core.mem_instr[15] ));
 sg13g2_inv_1 _13273_ (.Y(_09071_),
    .A(_09070_));
 sg13g2_nand2_1 _13274_ (.Y(_09072_),
    .A(net5348),
    .B(_09070_));
 sg13g2_a21oi_2 _13275_ (.B1(net6172),
    .Y(_09073_),
    .A2(_09071_),
    .A1(net6304));
 sg13g2_a22oi_1 _13276_ (.Y(_09074_),
    .B1(_09073_),
    .B2(net3021),
    .A2(_09072_),
    .A1(net5533));
 sg13g2_nand2_1 _13277_ (.Y(_09075_),
    .A(_09029_),
    .B(net5533));
 sg13g2_o21ai_1 _13278_ (.B1(net4789),
    .Y(_09076_),
    .A1(_09044_),
    .A2(net6105));
 sg13g2_a22oi_1 _13279_ (.Y(_09077_),
    .B1(_09074_),
    .B2(_09076_),
    .A2(_09063_),
    .A1(net4789));
 sg13g2_o21ai_1 _13280_ (.B1(_09077_),
    .Y(_09078_),
    .A1(net3021),
    .A2(_09061_));
 sg13g2_inv_1 _13281_ (.Y(_00058_),
    .A(_09078_));
 sg13g2_o21ai_1 _13282_ (.B1(net5007),
    .Y(_09079_),
    .A1(_07871_),
    .A2(\soc_inst.cpu_core.id_pc[1] ));
 sg13g2_o21ai_1 _13283_ (.B1(_09079_),
    .Y(_09080_),
    .A1(_08137_),
    .A2(net5007));
 sg13g2_or2_1 _13284_ (.X(_09081_),
    .B(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .A(net6293));
 sg13g2_o21ai_1 _13285_ (.B1(_09081_),
    .Y(_09082_),
    .A1(net6168),
    .A2(\soc_inst.cpu_core.mem_instr[16] ));
 sg13g2_inv_1 _13286_ (.Y(_09083_),
    .A(_09082_));
 sg13g2_nand2_1 _13287_ (.Y(_09084_),
    .A(net5347),
    .B(_09082_));
 sg13g2_a21oi_2 _13288_ (.B1(net6172),
    .Y(_09085_),
    .A2(_09083_),
    .A1(net6305));
 sg13g2_a22oi_1 _13289_ (.Y(_09086_),
    .B1(_09085_),
    .B2(net3149),
    .A2(_09084_),
    .A1(net5533));
 sg13g2_o21ai_1 _13290_ (.B1(_09080_),
    .Y(_09087_),
    .A1(net3149),
    .A2(net4940));
 sg13g2_a22oi_1 _13291_ (.Y(_00059_),
    .B1(_09087_),
    .B2(net4789),
    .A2(_09086_),
    .A1(_09076_));
 sg13g2_nor3_1 _13292_ (.A(_07871_),
    .B(\soc_inst.cpu_core.id_pc[2] ),
    .C(net4999),
    .Y(_09088_));
 sg13g2_a21oi_1 _13293_ (.A1(_08138_),
    .A2(net5000),
    .Y(_09089_),
    .B1(_09088_));
 sg13g2_or2_1 _13294_ (.X(_09090_),
    .B(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .A(net6293));
 sg13g2_o21ai_1 _13295_ (.B1(_09090_),
    .Y(_09091_),
    .A1(net6169),
    .A2(\soc_inst.cpu_core.mem_instr[17] ));
 sg13g2_inv_1 _13296_ (.Y(_09092_),
    .A(_09091_));
 sg13g2_a21oi_2 _13297_ (.B1(net6172),
    .Y(_09093_),
    .A2(_09092_),
    .A1(net6305));
 sg13g2_nand2_1 _13298_ (.Y(_09094_),
    .A(net5347),
    .B(_09091_));
 sg13g2_a22oi_1 _13299_ (.Y(_09095_),
    .B1(_09094_),
    .B2(net5535),
    .A2(_09093_),
    .A1(net3246));
 sg13g2_o21ai_1 _13300_ (.B1(_09089_),
    .Y(_09096_),
    .A1(net3246),
    .A2(net4940));
 sg13g2_and2_1 _13301_ (.A(net4789),
    .B(_09096_),
    .X(_09097_));
 sg13g2_a21oi_1 _13302_ (.A1(_09076_),
    .A2(_09095_),
    .Y(_00060_),
    .B1(_09097_));
 sg13g2_nor3_1 _13303_ (.A(_07871_),
    .B(\soc_inst.cpu_core.id_pc[3] ),
    .C(net5000),
    .Y(_09098_));
 sg13g2_a21oi_1 _13304_ (.A1(_08139_),
    .A2(net4999),
    .Y(_09099_),
    .B1(_09098_));
 sg13g2_a21oi_1 _13305_ (.A1(net6305),
    .A2(_09052_),
    .Y(_09100_),
    .B1(net6172));
 sg13g2_nand2_1 _13306_ (.Y(_09101_),
    .A(_09051_),
    .B(net5347));
 sg13g2_a22oi_1 _13307_ (.Y(_09102_),
    .B1(_09101_),
    .B2(net5534),
    .A2(_09100_),
    .A1(net3245));
 sg13g2_o21ai_1 _13308_ (.B1(_09099_),
    .Y(_09103_),
    .A1(net3245),
    .A2(net4941));
 sg13g2_and2_1 _13309_ (.A(net4789),
    .B(_09103_),
    .X(_09104_));
 sg13g2_a21oi_1 _13310_ (.A1(_09076_),
    .A2(_09102_),
    .Y(_00061_),
    .B1(_09104_));
 sg13g2_o21ai_1 _13311_ (.B1(net5007),
    .Y(_09105_),
    .A1(_07871_),
    .A2(\soc_inst.cpu_core.id_pc[4] ));
 sg13g2_o21ai_1 _13312_ (.B1(_09105_),
    .Y(_09106_),
    .A1(_08140_),
    .A2(net5008));
 sg13g2_or2_1 _13313_ (.X(_09107_),
    .B(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .A(net6293));
 sg13g2_o21ai_1 _13314_ (.B1(_09107_),
    .Y(_09108_),
    .A1(net6169),
    .A2(\soc_inst.cpu_core.mem_instr[19] ));
 sg13g2_inv_1 _13315_ (.Y(_09109_),
    .A(_09108_));
 sg13g2_nand2_1 _13316_ (.Y(_09110_),
    .A(net5348),
    .B(_09108_));
 sg13g2_a21oi_2 _13317_ (.B1(net6172),
    .Y(_09111_),
    .A2(_09109_),
    .A1(net6304));
 sg13g2_a22oi_1 _13318_ (.Y(_09112_),
    .B1(_09111_),
    .B2(net2959),
    .A2(_09110_),
    .A1(net5533));
 sg13g2_o21ai_1 _13319_ (.B1(_09106_),
    .Y(_09113_),
    .A1(net2959),
    .A2(net4940));
 sg13g2_a22oi_1 _13320_ (.Y(_00062_),
    .B1(_09113_),
    .B2(net4790),
    .A2(_09112_),
    .A1(_09076_));
 sg13g2_a21oi_1 _13321_ (.A1(_07999_),
    .A2(net4949),
    .Y(_09114_),
    .B1(net5048));
 sg13g2_nor2_1 _13322_ (.A(_08992_),
    .B(_09003_),
    .Y(_09115_));
 sg13g2_nor3_1 _13323_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(_08992_),
    .C(_09003_),
    .Y(_09116_));
 sg13g2_nand2b_2 _13324_ (.Y(_09117_),
    .B(_09115_),
    .A_N(\soc_inst.cpu_core.csr_file.csr_addr[0] ));
 sg13g2_nand2_1 _13325_ (.Y(_09118_),
    .A(_09030_),
    .B(net5340));
 sg13g2_nor2_1 _13326_ (.A(_09044_),
    .B(_09117_),
    .Y(_09119_));
 sg13g2_nor2_1 _13327_ (.A(_09114_),
    .B(_09119_),
    .Y(_09120_));
 sg13g2_nand2_1 _13328_ (.Y(_09121_),
    .A(_09070_),
    .B(net5342));
 sg13g2_a22oi_1 _13329_ (.Y(_09122_),
    .B1(_09121_),
    .B2(net5535),
    .A2(_09073_),
    .A1(net3195));
 sg13g2_nand2_2 _13330_ (.Y(_09123_),
    .A(_09075_),
    .B(net4934));
 sg13g2_a21oi_1 _13331_ (.A1(_09122_),
    .A2(_09123_),
    .Y(_00027_),
    .B1(_09120_));
 sg13g2_and2_1 _13332_ (.A(_08945_),
    .B(_08948_),
    .X(_09124_));
 sg13g2_nor3_1 _13333_ (.A(net6213),
    .B(_08944_),
    .C(_09124_),
    .Y(_09125_));
 sg13g2_nor3_1 _13334_ (.A(net5163),
    .B(net4950),
    .C(_09125_),
    .Y(_09126_));
 sg13g2_a221oi_1 _13335_ (.B2(net5341),
    .C1(_09126_),
    .B1(_09037_),
    .A1(net3128),
    .Y(_09127_),
    .A2(net4945));
 sg13g2_nand2_1 _13336_ (.Y(_09128_),
    .A(_09082_),
    .B(net5342));
 sg13g2_a22oi_1 _13337_ (.Y(_09129_),
    .B1(_09128_),
    .B2(net5535),
    .A2(_09085_),
    .A1(net3128));
 sg13g2_a21oi_1 _13338_ (.A1(_09123_),
    .A2(_09129_),
    .Y(_00038_),
    .B1(_09127_));
 sg13g2_and2_1 _13339_ (.A(\soc_inst.cpu_core.csr_file.mie[7] ),
    .B(\soc_inst.cpu_core.csr_file.mip_tip ),
    .X(_09130_));
 sg13g2_o21ai_1 _13340_ (.B1(net5001),
    .Y(_09131_),
    .A1(_07871_),
    .A2(_09130_));
 sg13g2_a22oi_1 _13341_ (.Y(_09132_),
    .B1(_09131_),
    .B2(net5166),
    .A2(net4948),
    .A1(_08003_));
 sg13g2_nor2_1 _13342_ (.A(_09119_),
    .B(_09132_),
    .Y(_09133_));
 sg13g2_nand2_1 _13343_ (.Y(_09134_),
    .A(_09091_),
    .B(net5342));
 sg13g2_a22oi_1 _13344_ (.Y(_09135_),
    .B1(_09134_),
    .B2(net5535),
    .A2(_09093_),
    .A1(net3213));
 sg13g2_a21oi_1 _13345_ (.A1(_09123_),
    .A2(_09135_),
    .Y(_00049_),
    .B1(_09133_));
 sg13g2_nor2b_1 _13346_ (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .B_N(\soc_inst.cpu_core.ex_is_ebreak ),
    .Y(_09136_));
 sg13g2_nor2_2 _13347_ (.A(net5046),
    .B(net6099),
    .Y(_09137_));
 sg13g2_a221oi_1 _13348_ (.B2(_09137_),
    .C1(_09119_),
    .B1(_09131_),
    .A1(net3116),
    .Y(_09138_),
    .A2(net4948));
 sg13g2_nand2_1 _13349_ (.Y(_09139_),
    .A(_09051_),
    .B(net5343));
 sg13g2_a22oi_1 _13350_ (.Y(_09140_),
    .B1(_09139_),
    .B2(net5535),
    .A2(_09100_),
    .A1(net3116));
 sg13g2_a21oi_1 _13351_ (.A1(_09123_),
    .A2(_09140_),
    .Y(_00051_),
    .B1(_09138_));
 sg13g2_and3_1 _13352_ (.X(_00052_),
    .A(net99),
    .B(net4945),
    .C(net4933));
 sg13g2_and3_1 _13353_ (.X(_00053_),
    .A(net116),
    .B(net4945),
    .C(net4933));
 sg13g2_and3_1 _13354_ (.X(_00054_),
    .A(net130),
    .B(net4952),
    .C(net4935));
 sg13g2_and3_1 _13355_ (.X(_00055_),
    .A(net114),
    .B(net4951),
    .C(net4935));
 sg13g2_and3_1 _13356_ (.X(_00056_),
    .A(net120),
    .B(net4953),
    .C(net4933));
 sg13g2_and3_1 _13357_ (.X(_00057_),
    .A(net122),
    .B(net4952),
    .C(net4934));
 sg13g2_and3_1 _13358_ (.X(_00028_),
    .A(net147),
    .B(net4947),
    .C(net4934));
 sg13g2_and3_1 _13359_ (.X(_00029_),
    .A(net107),
    .B(net4951),
    .C(net4935));
 sg13g2_and3_1 _13360_ (.X(_00030_),
    .A(net109),
    .B(net4947),
    .C(net4934));
 sg13g2_and3_1 _13361_ (.X(_00031_),
    .A(net152),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13362_ (.X(_00032_),
    .A(net121),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13363_ (.X(_00033_),
    .A(net106),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13364_ (.X(_00034_),
    .A(net105),
    .B(net4946),
    .C(net4934));
 sg13g2_and3_1 _13365_ (.X(_00035_),
    .A(net108),
    .B(net4944),
    .C(net4932));
 sg13g2_and3_1 _13366_ (.X(_00036_),
    .A(net101),
    .B(net4947),
    .C(net4934));
 sg13g2_and3_1 _13367_ (.X(_00037_),
    .A(net157),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13368_ (.X(_00039_),
    .A(net186),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13369_ (.X(_00040_),
    .A(net110),
    .B(net4947),
    .C(net4934));
 sg13g2_and3_1 _13370_ (.X(_00041_),
    .A(net123),
    .B(net4944),
    .C(net4932));
 sg13g2_and3_1 _13371_ (.X(_00042_),
    .A(net117),
    .B(net4945),
    .C(net4932));
 sg13g2_and3_1 _13372_ (.X(_00043_),
    .A(net119),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13373_ (.X(_00044_),
    .A(net103),
    .B(net4944),
    .C(net4931));
 sg13g2_and3_1 _13374_ (.X(_00045_),
    .A(net102),
    .B(net4943),
    .C(net4931));
 sg13g2_and3_1 _13375_ (.X(_00046_),
    .A(net100),
    .B(net4944),
    .C(net4932));
 sg13g2_and3_1 _13376_ (.X(_00047_),
    .A(net115),
    .B(net4944),
    .C(net4932));
 sg13g2_and3_1 _13377_ (.X(_00048_),
    .A(net104),
    .B(net4943),
    .C(net4932));
 sg13g2_and3_1 _13378_ (.X(_00050_),
    .A(net129),
    .B(net4944),
    .C(net4932));
 sg13g2_and2_1 _13379_ (.A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(_09115_),
    .X(_09141_));
 sg13g2_nand2_1 _13380_ (.Y(_09142_),
    .A(_09030_),
    .B(net5146));
 sg13g2_and2_1 _13381_ (.A(net4936),
    .B(net5145),
    .X(_09143_));
 sg13g2_nand2_2 _13382_ (.Y(_09144_),
    .A(net4936),
    .B(net5145));
 sg13g2_nor3_1 _13383_ (.A(net3091),
    .B(net4941),
    .C(_09143_),
    .Y(_09145_));
 sg13g2_nand3_1 _13384_ (.B(net5166),
    .C(net6100),
    .A(\soc_inst.cpu_core.ex_exception_pc[0] ),
    .Y(_09146_));
 sg13g2_a21oi_1 _13385_ (.A1(\soc_inst.cpu_core.ex_alu_result[0] ),
    .A2(net5169),
    .Y(_09147_),
    .B1(net5076));
 sg13g2_a21oi_1 _13386_ (.A1(_09146_),
    .A2(_09147_),
    .Y(_09148_),
    .B1(_00261_));
 sg13g2_nor3_1 _13387_ (.A(net5163),
    .B(net4949),
    .C(_09148_),
    .Y(_09149_));
 sg13g2_nand2_1 _13388_ (.Y(_09150_),
    .A(_09070_),
    .B(net5148));
 sg13g2_a22oi_1 _13389_ (.Y(_09151_),
    .B1(_09150_),
    .B2(net5533),
    .A2(_09073_),
    .A1(net3091));
 sg13g2_nand2_2 _13390_ (.Y(_09152_),
    .A(_09075_),
    .B(net4929));
 sg13g2_a22oi_1 _13391_ (.Y(_09153_),
    .B1(_09151_),
    .B2(_09152_),
    .A2(_09149_),
    .A1(net4929));
 sg13g2_nor2b_1 _13392_ (.A(_09145_),
    .B_N(_09153_),
    .Y(_00083_));
 sg13g2_a21oi_1 _13393_ (.A1(net2368),
    .A2(net6100),
    .Y(_09154_),
    .B1(net5048));
 sg13g2_nor2_1 _13394_ (.A(net3401),
    .B(net5166),
    .Y(_09155_));
 sg13g2_nor2_1 _13395_ (.A(net3012),
    .B(net5158),
    .Y(_09156_));
 sg13g2_nor4_1 _13396_ (.A(net2888),
    .B(_09154_),
    .C(_09155_),
    .D(_09156_),
    .Y(_09157_));
 sg13g2_a21oi_1 _13397_ (.A1(net3172),
    .A2(net4949),
    .Y(_09158_),
    .B1(_09157_));
 sg13g2_nand2_1 _13398_ (.Y(_09159_),
    .A(_09082_),
    .B(net5148));
 sg13g2_a22oi_1 _13399_ (.Y(_09160_),
    .B1(_09159_),
    .B2(net5534),
    .A2(_09085_),
    .A1(net3172));
 sg13g2_a22oi_1 _13400_ (.Y(_00084_),
    .B1(_09160_),
    .B2(_09152_),
    .A2(_09158_),
    .A1(net4785));
 sg13g2_nand2_1 _13401_ (.Y(_09161_),
    .A(\soc_inst.cpu_core.ex_alu_result[2] ),
    .B(_08950_));
 sg13g2_nand3_1 _13402_ (.B(net5167),
    .C(net6100),
    .A(\soc_inst.cpu_core.ex_exception_pc[2] ),
    .Y(_09162_));
 sg13g2_nand3_1 _13403_ (.B(_09161_),
    .C(_09162_),
    .A(net5071),
    .Y(_09163_));
 sg13g2_o21ai_1 _13404_ (.B1(_09163_),
    .Y(_09164_),
    .A1(\soc_inst.cpu_core.ex_instr[2] ),
    .A2(net5071));
 sg13g2_nor2_1 _13405_ (.A(net5163),
    .B(_09164_),
    .Y(_09165_));
 sg13g2_a221oi_1 _13406_ (.B2(net3260),
    .C1(_09165_),
    .B1(net4949),
    .A1(net1784),
    .Y(_09166_),
    .A2(net5163));
 sg13g2_nand2_1 _13407_ (.Y(_09167_),
    .A(_09091_),
    .B(net5148));
 sg13g2_a22oi_1 _13408_ (.Y(_09168_),
    .B1(_09167_),
    .B2(net5535),
    .A2(_09093_),
    .A1(net3260));
 sg13g2_a22oi_1 _13409_ (.Y(_00085_),
    .B1(_09168_),
    .B2(_09152_),
    .A2(_09166_),
    .A1(net4785));
 sg13g2_a21oi_1 _13410_ (.A1(net1923),
    .A2(net6100),
    .Y(_09169_),
    .B1(net5047));
 sg13g2_nor2_1 _13411_ (.A(\soc_inst.cpu_core.ex_instr[3] ),
    .B(net5071),
    .Y(_09170_));
 sg13g2_nor2_1 _13412_ (.A(net2914),
    .B(net5158),
    .Y(_09171_));
 sg13g2_nor2_1 _13413_ (.A(\soc_inst.cpu_core.ex_alu_result[3] ),
    .B(net5166),
    .Y(_09172_));
 sg13g2_nor4_1 _13414_ (.A(_09169_),
    .B(_09170_),
    .C(_09171_),
    .D(_09172_),
    .Y(_09173_));
 sg13g2_a21oi_1 _13415_ (.A1(net3101),
    .A2(net4949),
    .Y(_09174_),
    .B1(_09173_));
 sg13g2_nand2_1 _13416_ (.Y(_09175_),
    .A(_09051_),
    .B(net5148));
 sg13g2_a22oi_1 _13417_ (.Y(_09176_),
    .B1(_09175_),
    .B2(net5534),
    .A2(_09100_),
    .A1(net3101));
 sg13g2_a22oi_1 _13418_ (.Y(_00086_),
    .B1(_09176_),
    .B2(_09152_),
    .A2(_09174_),
    .A1(net4785));
 sg13g2_a21oi_1 _13419_ (.A1(net2219),
    .A2(net6100),
    .Y(_09177_),
    .B1(net5047));
 sg13g2_nor2_1 _13420_ (.A(_07791_),
    .B(_08958_),
    .Y(_09178_));
 sg13g2_nor2_1 _13421_ (.A(\soc_inst.cpu_core.ex_alu_result[4] ),
    .B(net5167),
    .Y(_09179_));
 sg13g2_nor2_1 _13422_ (.A(net2876),
    .B(_08965_),
    .Y(_09180_));
 sg13g2_nor4_2 _13423_ (.A(_09177_),
    .B(_09178_),
    .C(_09179_),
    .Y(_09181_),
    .D(_09180_));
 sg13g2_a21oi_1 _13424_ (.A1(net3026),
    .A2(net4945),
    .Y(_09182_),
    .B1(_09181_));
 sg13g2_nand2_1 _13425_ (.Y(_09183_),
    .A(_09108_),
    .B(net5149));
 sg13g2_a22oi_1 _13426_ (.Y(_09184_),
    .B1(_09183_),
    .B2(net5533),
    .A2(_09111_),
    .A1(net3026));
 sg13g2_a22oi_1 _13427_ (.Y(_00087_),
    .B1(_09184_),
    .B2(_09152_),
    .A2(net3027),
    .A1(net4785));
 sg13g2_mux2_1 _13428_ (.A0(_00232_),
    .A1(\soc_inst.gpio_bidir_oe [0]),
    .S(_08405_),
    .X(uio_oe[7]));
 sg13g2_and2_1 _13429_ (.A(\soc_inst.gpio_bidir_out [0]),
    .B(_08405_),
    .X(uio_out[7]));
 sg13g2_nand2b_1 _13430_ (.Y(_09185_),
    .B(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][11] ));
 sg13g2_nand2b_1 _13431_ (.Y(_09186_),
    .B(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][10] ));
 sg13g2_nor2b_1 _13432_ (.A(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .B_N(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .Y(_09187_));
 sg13g2_a21oi_1 _13433_ (.A1(_09185_),
    .A2(_09186_),
    .Y(_09188_),
    .B1(_09187_));
 sg13g2_nand2b_1 _13434_ (.Y(_09189_),
    .B(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .A_N(\soc_inst.pwm_inst.channel_counter[0][6] ));
 sg13g2_nor2_1 _13435_ (.A(_07946_),
    .B(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .Y(_09190_));
 sg13g2_nor2_1 _13436_ (.A(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .B(_07954_),
    .Y(_09191_));
 sg13g2_nor2b_1 _13437_ (.A(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .B_N(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .Y(_09192_));
 sg13g2_a22oi_1 _13438_ (.Y(_09193_),
    .B1(_07955_),
    .B2(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .A2(_07954_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][1] ));
 sg13g2_o21ai_1 _13439_ (.B1(_09193_),
    .Y(_09194_),
    .A1(_09191_),
    .A2(_09192_));
 sg13g2_o21ai_1 _13440_ (.B1(_09194_),
    .Y(_09195_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .A2(_07955_));
 sg13g2_a21oi_1 _13441_ (.A1(_07948_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .Y(_09196_),
    .B1(_09195_));
 sg13g2_a221oi_1 _13442_ (.B2(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .C1(_09196_),
    .B1(_07959_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .Y(_09197_),
    .A2(_07957_));
 sg13g2_a221oi_1 _13443_ (.B2(_07946_),
    .C1(_09197_),
    .B1(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .A1(_07947_),
    .Y(_09198_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][4] ));
 sg13g2_o21ai_1 _13444_ (.B1(_09189_),
    .Y(_09199_),
    .A1(_09190_),
    .A2(_09198_));
 sg13g2_a22oi_1 _13445_ (.Y(_09200_),
    .B1(_07963_),
    .B2(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .A2(_07962_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][6] ));
 sg13g2_nor2_1 _13446_ (.A(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .B(_07963_),
    .Y(_09201_));
 sg13g2_a221oi_1 _13447_ (.B2(_09200_),
    .C1(_09201_),
    .B1(_09199_),
    .A1(_07945_),
    .Y(_09202_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][8] ));
 sg13g2_nand2b_1 _13448_ (.Y(_09203_),
    .B(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .A_N(\soc_inst.pwm_inst.channel_duty[0][9] ));
 sg13g2_o21ai_1 _13449_ (.B1(_09203_),
    .Y(_09204_),
    .A1(_07945_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][8] ));
 sg13g2_or2_1 _13450_ (.X(_09205_),
    .B(_09204_),
    .A(_09202_));
 sg13g2_a221oi_1 _13451_ (.B2(_07943_),
    .C1(_09187_),
    .B1(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .A1(_07944_),
    .Y(_09206_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][9] ));
 sg13g2_nand4_1 _13452_ (.B(_09186_),
    .C(_09205_),
    .A(_09185_),
    .Y(_09207_),
    .D(_09206_));
 sg13g2_nand2b_1 _13453_ (.Y(_09208_),
    .B(_09207_),
    .A_N(_09188_));
 sg13g2_nand2_1 _13454_ (.Y(_09209_),
    .A(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .B(_07966_));
 sg13g2_o21ai_1 _13455_ (.B1(_09209_),
    .Y(_09210_),
    .A1(_07941_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][15] ));
 sg13g2_nand2_1 _13456_ (.Y(_09211_),
    .A(_07941_),
    .B(\soc_inst.pwm_inst.channel_duty[0][15] ));
 sg13g2_o21ai_1 _13457_ (.B1(_09211_),
    .Y(_09212_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .A2(_07966_));
 sg13g2_nor2_1 _13458_ (.A(_09210_),
    .B(_09212_),
    .Y(_09213_));
 sg13g2_a22oi_1 _13459_ (.Y(_09214_),
    .B1(_07965_),
    .B2(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .A2(_07964_),
    .A1(\soc_inst.pwm_inst.channel_counter[0][12] ));
 sg13g2_nor2_1 _13460_ (.A(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .B(_07965_),
    .Y(_09215_));
 sg13g2_a21oi_1 _13461_ (.A1(_07942_),
    .A2(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .Y(_09216_),
    .B1(_09215_));
 sg13g2_nand4_1 _13462_ (.B(_09213_),
    .C(_09214_),
    .A(_09208_),
    .Y(_09217_),
    .D(_09216_));
 sg13g2_nor2_1 _13463_ (.A(_09214_),
    .B(_09215_),
    .Y(_09218_));
 sg13g2_a22oi_1 _13464_ (.Y(_09219_),
    .B1(_09213_),
    .B2(_09218_),
    .A2(_09211_),
    .A1(_09210_));
 sg13g2_nand3_1 _13465_ (.B(_09217_),
    .C(_09219_),
    .A(\soc_inst.pwm_ena [0]),
    .Y(_09220_));
 sg13g2_o21ai_1 _13466_ (.B1(_09220_),
    .Y(uo_out[6]),
    .A1(\soc_inst.pwm_ena [0]),
    .A2(_07960_));
 sg13g2_nor2_1 _13467_ (.A(\soc_inst.spi_ena ),
    .B(\soc_inst.gpio_inst.gpio_out[3] ),
    .Y(_09221_));
 sg13g2_a21oi_2 _13468_ (.B1(_09221_),
    .Y(uo_out[5]),
    .A2(_08186_),
    .A1(\soc_inst.spi_ena ));
 sg13g2_nor2_1 _13469_ (.A(\soc_inst.spi_ena ),
    .B(\soc_inst.gpio_inst.gpio_out[2] ),
    .Y(_09222_));
 sg13g2_a21oi_2 _13470_ (.B1(_09222_),
    .Y(uo_out[4]),
    .A2(\soc_inst.spi_ena ),
    .A1(_07898_));
 sg13g2_nand2_1 _13471_ (.Y(_09223_),
    .A(\soc_inst.gpio_inst.gpio_out[0] ),
    .B(_08405_));
 sg13g2_o21ai_1 _13472_ (.B1(_09223_),
    .Y(uo_out[2]),
    .A1(_00233_),
    .A2(_08405_));
 sg13g2_a21oi_1 _13473_ (.A1(net6461),
    .A2(_08795_),
    .Y(_09224_),
    .B1(net594));
 sg13g2_nand2_1 _13474_ (.Y(_09225_),
    .A(net6536),
    .B(_08403_));
 sg13g2_and3_2 _13475_ (.X(_09226_),
    .A(net6534),
    .B(net6535),
    .C(_08403_));
 sg13g2_nand3_1 _13476_ (.B(net6535),
    .C(_08403_),
    .A(net6534),
    .Y(_09227_));
 sg13g2_nand2b_2 _13477_ (.Y(_09228_),
    .B(net6534),
    .A_N(net6535));
 sg13g2_a21oi_1 _13478_ (.A1(_08798_),
    .A2(_09228_),
    .Y(_09229_),
    .B1(_09226_));
 sg13g2_nor2_1 _13479_ (.A(net820),
    .B(_09227_),
    .Y(_09230_));
 sg13g2_nand2_1 _13480_ (.Y(_09231_),
    .A(_07894_),
    .B(_09226_));
 sg13g2_nor3_1 _13481_ (.A(net5565),
    .B(_09229_),
    .C(_09230_),
    .Y(_09232_));
 sg13g2_o21ai_1 _13482_ (.B1(_09232_),
    .Y(_09233_),
    .A1(net594),
    .A2(_09227_));
 sg13g2_nor2b_1 _13483_ (.A(_09224_),
    .B_N(_09233_),
    .Y(_11835_[0]));
 sg13g2_nand2_1 _13484_ (.Y(_09234_),
    .A(_07804_),
    .B(net183));
 sg13g2_and2_1 _13485_ (.A(_00222_),
    .B(_00221_),
    .X(_09235_));
 sg13g2_and2_1 _13486_ (.A(_00223_),
    .B(_09235_),
    .X(_09236_));
 sg13g2_nand2_1 _13487_ (.Y(_09237_),
    .A(_00224_),
    .B(_09236_));
 sg13g2_nand3_1 _13488_ (.B(_00224_),
    .C(_09236_),
    .A(_00225_),
    .Y(_09238_));
 sg13g2_nor2_1 _13489_ (.A(net2996),
    .B(_09238_),
    .Y(_09239_));
 sg13g2_nor2_1 _13490_ (.A(_00221_),
    .B(_08689_),
    .Y(_09240_));
 sg13g2_a21oi_1 _13491_ (.A1(_08690_),
    .A2(_09235_),
    .Y(_09241_),
    .B1(_09240_));
 sg13g2_xor2_1 _13492_ (.B(net6545),
    .A(\soc_inst.spi_inst.bit_counter[5] ),
    .X(_09242_));
 sg13g2_nor2b_2 _13493_ (.A(net6545),
    .B_N(\soc_inst.spi_inst.len_sel[0] ),
    .Y(_09243_));
 sg13g2_nand2b_2 _13494_ (.Y(_09244_),
    .B(\soc_inst.spi_inst.len_sel[0] ),
    .A_N(net6545));
 sg13g2_o21ai_1 _13495_ (.B1(\soc_inst.spi_inst.bit_counter[4] ),
    .Y(_09245_),
    .A1(\soc_inst.spi_inst.bit_counter[3] ),
    .A2(_09244_));
 sg13g2_nor4_1 _13496_ (.A(\soc_inst.spi_inst.bit_counter[0] ),
    .B(\soc_inst.spi_inst.bit_counter[1] ),
    .C(net3356),
    .D(_08688_),
    .Y(_09246_));
 sg13g2_nor3_1 _13497_ (.A(\soc_inst.spi_inst.bit_counter[3] ),
    .B(\soc_inst.spi_inst.bit_counter[4] ),
    .C(net6545),
    .Y(_09247_));
 sg13g2_or2_1 _13498_ (.X(_09248_),
    .B(\soc_inst.spi_inst.len_sel[0] ),
    .A(net6545));
 sg13g2_a21oi_1 _13499_ (.A1(\soc_inst.spi_inst.bit_counter[3] ),
    .A2(_09248_),
    .Y(_09249_),
    .B1(_09247_));
 sg13g2_nor3_1 _13500_ (.A(\soc_inst.spi_inst.clock_divider[5] ),
    .B(\soc_inst.spi_inst.clock_divider[6] ),
    .C(_09238_),
    .Y(_09250_));
 sg13g2_nor2b_1 _13501_ (.A(_08687_),
    .B_N(_09250_),
    .Y(_09251_));
 sg13g2_nor3_1 _13502_ (.A(\soc_inst.spi_inst.clk_counter[7] ),
    .B(_07896_),
    .C(_09250_),
    .Y(_09252_));
 sg13g2_nor2_1 _13503_ (.A(_08684_),
    .B(_09236_),
    .Y(_09253_));
 sg13g2_or2_1 _13504_ (.X(_09254_),
    .B(_09235_),
    .A(_08690_));
 sg13g2_a22oi_1 _13505_ (.Y(_09255_),
    .B1(_09236_),
    .B2(_08684_),
    .A2(_08689_),
    .A1(_00221_));
 sg13g2_nor4_1 _13506_ (.A(net6110),
    .B(_08686_),
    .C(_09242_),
    .D(_09253_),
    .Y(_09256_));
 sg13g2_xnor2_1 _13507_ (.Y(_09257_),
    .A(_08682_),
    .B(_09238_));
 sg13g2_xor2_1 _13508_ (.B(_09239_),
    .A(_08681_),
    .X(_09258_));
 sg13g2_nand4_1 _13509_ (.B(_09249_),
    .C(_09255_),
    .A(net3357),
    .Y(_09259_),
    .D(_09256_));
 sg13g2_xnor2_1 _13510_ (.Y(_09260_),
    .A(_08691_),
    .B(_09237_));
 sg13g2_nand4_1 _13511_ (.B(_09245_),
    .C(_09254_),
    .A(_09241_),
    .Y(_09261_),
    .D(_09260_));
 sg13g2_nor4_1 _13512_ (.A(_09251_),
    .B(_09252_),
    .C(_09259_),
    .D(_09261_),
    .Y(_09262_));
 sg13g2_nand3_1 _13513_ (.B(_09258_),
    .C(_09262_),
    .A(_09257_),
    .Y(_09263_));
 sg13g2_o21ai_1 _13514_ (.B1(_09263_),
    .Y(\soc_inst.spi_inst.next_state[0] ),
    .A1(\soc_inst.spi_inst.state[0] ),
    .A2(net184));
 sg13g2_and2_1 _13515_ (.A(_00127_),
    .B(_09263_),
    .X(_11837_[0]));
 sg13g2_a21oi_1 _13516_ (.A1(net6470),
    .A2(_08795_),
    .Y(_09264_),
    .B1(net820));
 sg13g2_nor2_1 _13517_ (.A(_09232_),
    .B(net821),
    .Y(_11836_[0]));
 sg13g2_nor2_2 _13518_ (.A(net6537),
    .B(_08828_),
    .Y(_09265_));
 sg13g2_and2_1 _13519_ (.A(_08403_),
    .B(_08827_),
    .X(_09266_));
 sg13g2_a22oi_1 _13520_ (.Y(_09267_),
    .B1(net5565),
    .B2(_09266_),
    .A2(_08405_),
    .A1(_07894_));
 sg13g2_nand2_1 _13521_ (.Y(_09268_),
    .A(net5565),
    .B(_09226_));
 sg13g2_nand2_1 _13522_ (.Y(_09269_),
    .A(_08403_),
    .B(_09228_));
 sg13g2_nor4_1 _13523_ (.A(\soc_inst.i2c_inst.clk_cnt[4] ),
    .B(\soc_inst.i2c_inst.clk_cnt[5] ),
    .C(\soc_inst.i2c_inst.clk_cnt[6] ),
    .D(\soc_inst.i2c_inst.clk_cnt[7] ),
    .Y(_09270_));
 sg13g2_nor4_1 _13524_ (.A(\soc_inst.i2c_inst.clk_cnt[0] ),
    .B(\soc_inst.i2c_inst.clk_cnt[1] ),
    .C(\soc_inst.i2c_inst.clk_cnt[2] ),
    .D(\soc_inst.i2c_inst.clk_cnt[3] ),
    .Y(_09271_));
 sg13g2_and2_1 _13525_ (.A(_09270_),
    .B(_09271_),
    .X(_09272_));
 sg13g2_nand2b_2 _13526_ (.Y(_09273_),
    .B(_08825_),
    .A_N(_08797_));
 sg13g2_inv_1 _13527_ (.Y(_09274_),
    .A(_09273_));
 sg13g2_nand3_1 _13528_ (.B(_09272_),
    .C(_09274_),
    .A(net6546),
    .Y(_09275_));
 sg13g2_inv_1 _13529_ (.Y(_09276_),
    .A(_09275_));
 sg13g2_a22oi_1 _13530_ (.Y(_09277_),
    .B1(_09269_),
    .B2(_09275_),
    .A2(_09266_),
    .A1(net6546));
 sg13g2_nand4_1 _13531_ (.B(_09267_),
    .C(_09268_),
    .A(_09231_),
    .Y(_09278_),
    .D(_09277_));
 sg13g2_o21ai_1 _13532_ (.B1(_09278_),
    .Y(_09279_),
    .A1(net2250),
    .A2(net5178));
 sg13g2_nand2_1 _13533_ (.Y(_09280_),
    .A(\soc_inst.i2c_ena ),
    .B(_09227_));
 sg13g2_and3_2 _13534_ (.X(_09281_),
    .A(net820),
    .B(_08857_),
    .C(_09280_));
 sg13g2_a22oi_1 _13535_ (.Y(_09282_),
    .B1(_09281_),
    .B2(net2985),
    .A2(_09276_),
    .A1(net13));
 sg13g2_o21ai_1 _13536_ (.B1(_09282_),
    .Y(_02599_),
    .A1(_08834_),
    .A2(_09279_));
 sg13g2_o21ai_1 _13537_ (.B1(_09278_),
    .Y(_09283_),
    .A1(net1718),
    .A2(net5177));
 sg13g2_nand2b_1 _13538_ (.Y(_09284_),
    .B(_09266_),
    .A_N(net6546));
 sg13g2_o21ai_1 _13539_ (.B1(_09275_),
    .Y(_09285_),
    .A1(_08818_),
    .A2(_09284_));
 sg13g2_a22oi_1 _13540_ (.Y(_09286_),
    .B1(_09285_),
    .B2(net2250),
    .A2(_09281_),
    .A1(net2864));
 sg13g2_o21ai_1 _13541_ (.B1(_09286_),
    .Y(_02600_),
    .A1(_08837_),
    .A2(_09283_));
 sg13g2_o21ai_1 _13542_ (.B1(_09278_),
    .Y(_09287_),
    .A1(net1836),
    .A2(net5176));
 sg13g2_a22oi_1 _13543_ (.Y(_09288_),
    .B1(_09285_),
    .B2(net1718),
    .A2(_09281_),
    .A1(net2355));
 sg13g2_o21ai_1 _13544_ (.B1(_09288_),
    .Y(_02601_),
    .A1(_08840_),
    .A2(_09287_));
 sg13g2_o21ai_1 _13545_ (.B1(_09278_),
    .Y(_09289_),
    .A1(net2017),
    .A2(net5176));
 sg13g2_a22oi_1 _13546_ (.Y(_09290_),
    .B1(_09285_),
    .B2(net1836),
    .A2(_09281_),
    .A1(net2375));
 sg13g2_o21ai_1 _13547_ (.B1(_09290_),
    .Y(_02602_),
    .A1(_08843_),
    .A2(_09289_));
 sg13g2_nor2_1 _13548_ (.A(net2086),
    .B(net5176),
    .Y(_09291_));
 sg13g2_nand2b_1 _13549_ (.Y(_09292_),
    .B(_09278_),
    .A_N(_08846_));
 sg13g2_a22oi_1 _13550_ (.Y(_09293_),
    .B1(_09285_),
    .B2(net2017),
    .A2(_09281_),
    .A1(net2584));
 sg13g2_o21ai_1 _13551_ (.B1(_09293_),
    .Y(_02603_),
    .A1(_09291_),
    .A2(_09292_));
 sg13g2_o21ai_1 _13552_ (.B1(_09278_),
    .Y(_09294_),
    .A1(net2199),
    .A2(net5176));
 sg13g2_a22oi_1 _13553_ (.Y(_09295_),
    .B1(_09285_),
    .B2(net2086),
    .A2(_09281_),
    .A1(net2490));
 sg13g2_o21ai_1 _13554_ (.B1(_09295_),
    .Y(_02604_),
    .A1(_08849_),
    .A2(_09294_));
 sg13g2_o21ai_1 _13555_ (.B1(_09278_),
    .Y(_09296_),
    .A1(net1912),
    .A2(net5177));
 sg13g2_a22oi_1 _13556_ (.Y(_09297_),
    .B1(_09285_),
    .B2(net2199),
    .A2(_09281_),
    .A1(net2984));
 sg13g2_o21ai_1 _13557_ (.B1(_09297_),
    .Y(_02605_),
    .A1(_08852_),
    .A2(_09296_));
 sg13g2_o21ai_1 _13558_ (.B1(_09278_),
    .Y(_09298_),
    .A1(net2049),
    .A2(net5178));
 sg13g2_a22oi_1 _13559_ (.Y(_09299_),
    .B1(_09285_),
    .B2(net1912),
    .A2(_09281_),
    .A1(net2378));
 sg13g2_o21ai_1 _13560_ (.B1(_09299_),
    .Y(_02606_),
    .A1(_08855_),
    .A2(_09298_));
 sg13g2_nand4_1 _13561_ (.B(_07813_),
    .C(_08230_),
    .A(net6204),
    .Y(_09300_),
    .D(_08793_));
 sg13g2_nor2_2 _13562_ (.A(_08674_),
    .B(_09300_),
    .Y(_09301_));
 sg13g2_nor3_1 _13563_ (.A(net1842),
    .B(net2009),
    .C(_08492_),
    .Y(_09302_));
 sg13g2_nand3b_1 _13564_ (.B(_09302_),
    .C(net6178),
    .Y(_09303_),
    .A_N(_08469_));
 sg13g2_nor4_1 _13565_ (.A(net1018),
    .B(net921),
    .C(net665),
    .D(net529),
    .Y(_09304_));
 sg13g2_nor3_1 _13566_ (.A(net2489),
    .B(net1417),
    .C(net746),
    .Y(_09305_));
 sg13g2_nand3_1 _13567_ (.B(_09304_),
    .C(_09305_),
    .A(_07772_),
    .Y(_09306_));
 sg13g2_nand2_1 _13568_ (.Y(_09307_),
    .A(_08230_),
    .B(_08793_));
 sg13g2_nor2_2 _13569_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(_09307_),
    .Y(_09308_));
 sg13g2_nor3_1 _13570_ (.A(_09301_),
    .B(_09303_),
    .C(_09306_),
    .Y(_09309_));
 sg13g2_a21o_1 _13571_ (.A2(_09301_),
    .A1(net6465),
    .B1(_09309_),
    .X(_00170_));
 sg13g2_nor2_1 _13572_ (.A(net2623),
    .B(_09301_),
    .Y(_09310_));
 sg13g2_a22oi_1 _13573_ (.Y(_00171_),
    .B1(_09303_),
    .B2(_09310_),
    .A2(_09301_),
    .A1(_07785_));
 sg13g2_nand3_1 _13574_ (.B(\soc_inst.spi_ena ),
    .C(net5362),
    .A(\soc_inst.core_mem_wdata[0] ),
    .Y(_09311_));
 sg13g2_nor3_2 _13575_ (.A(net721),
    .B(_08677_),
    .C(_09311_),
    .Y(_00137_));
 sg13g2_inv_1 _13576_ (.Y(_09312_),
    .A(net722));
 sg13g2_nor2b_1 _13577_ (.A(_08639_),
    .B_N(net1639),
    .Y(_00000_));
 sg13g2_nor2b_1 _13578_ (.A(net95),
    .B_N(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .Y(_00110_));
 sg13g2_xor2_1 _13579_ (.B(net1353),
    .A(net770),
    .X(_00184_));
 sg13g2_nand3_1 _13580_ (.B(net1353),
    .C(net3379),
    .A(net770),
    .Y(_09313_));
 sg13g2_a21o_1 _13581_ (.A2(net1353),
    .A1(net770),
    .B1(net3379),
    .X(_09314_));
 sg13g2_and2_1 _13582_ (.A(_09313_),
    .B(_09314_),
    .X(_00195_));
 sg13g2_and4_1 _13583_ (.A(net770),
    .B(net1353),
    .C(net1179),
    .D(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .X(_09315_));
 sg13g2_xnor2_1 _13584_ (.Y(_00206_),
    .A(net1179),
    .B(_09313_));
 sg13g2_xnor2_1 _13585_ (.Y(_00215_),
    .A(_07902_),
    .B(_09315_));
 sg13g2_nand3_1 _13586_ (.B(net3255),
    .C(_09315_),
    .A(net3335),
    .Y(_09316_));
 sg13g2_a21o_1 _13587_ (.A2(_09315_),
    .A1(net3255),
    .B1(net3335),
    .X(_09317_));
 sg13g2_and2_1 _13588_ (.A(_09316_),
    .B(_09317_),
    .X(_00216_));
 sg13g2_nand4_1 _13589_ (.B(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .C(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .A(net1090),
    .Y(_09318_),
    .D(_09315_));
 sg13g2_xnor2_1 _13590_ (.Y(_00217_),
    .A(net1090),
    .B(_09316_));
 sg13g2_nor2_2 _13591_ (.A(_07901_),
    .B(_09318_),
    .Y(_09319_));
 sg13g2_xnor2_1 _13592_ (.Y(_00218_),
    .A(net400),
    .B(_09318_));
 sg13g2_xor2_1 _13593_ (.B(_09319_),
    .A(net3164),
    .X(_00219_));
 sg13g2_nand3_1 _13594_ (.B(net3164),
    .C(_09319_),
    .A(net3317),
    .Y(_09320_));
 sg13g2_a21o_1 _13595_ (.A2(_09319_),
    .A1(net3164),
    .B1(net3317),
    .X(_09321_));
 sg13g2_and2_1 _13596_ (.A(_09320_),
    .B(_09321_),
    .X(_00220_));
 sg13g2_and4_1 _13597_ (.A(net988),
    .B(net3406),
    .C(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .D(_09319_),
    .X(_09322_));
 sg13g2_xnor2_1 _13598_ (.Y(_00174_),
    .A(net988),
    .B(_09320_));
 sg13g2_xor2_1 _13599_ (.B(_09322_),
    .A(net1081),
    .X(_00175_));
 sg13g2_and3_2 _13600_ (.X(_09323_),
    .A(net1166),
    .B(net1081),
    .C(_09322_));
 sg13g2_a21oi_1 _13601_ (.A1(net1081),
    .A2(_09322_),
    .Y(_09324_),
    .B1(net1166));
 sg13g2_nor2_1 _13602_ (.A(_09323_),
    .B(net1167),
    .Y(_00176_));
 sg13g2_and2_1 _13603_ (.A(net1323),
    .B(_09323_),
    .X(_09325_));
 sg13g2_xor2_1 _13604_ (.B(_09323_),
    .A(net1323),
    .X(_00177_));
 sg13g2_xor2_1 _13605_ (.B(_09325_),
    .A(net1245),
    .X(_00178_));
 sg13g2_nand4_1 _13606_ (.B(net1245),
    .C(net1323),
    .A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .Y(_09326_),
    .D(_09323_));
 sg13g2_a21o_1 _13607_ (.A2(_09325_),
    .A1(net1245),
    .B1(net3333),
    .X(_09327_));
 sg13g2_and2_1 _13608_ (.A(_09326_),
    .B(_09327_),
    .X(_00179_));
 sg13g2_xnor2_1 _13609_ (.Y(_00180_),
    .A(net2464),
    .B(_09326_));
 sg13g2_nor3_2 _13610_ (.A(_07903_),
    .B(_07904_),
    .C(_09326_),
    .Y(_09328_));
 sg13g2_o21ai_1 _13611_ (.B1(_07903_),
    .Y(_09329_),
    .A1(_07904_),
    .A2(_09326_));
 sg13g2_nor2b_1 _13612_ (.A(_09328_),
    .B_N(_09329_),
    .Y(_00181_));
 sg13g2_xor2_1 _13613_ (.B(_09328_),
    .A(net2717),
    .X(_00182_));
 sg13g2_a21oi_1 _13614_ (.A1(net2717),
    .A2(_09328_),
    .Y(_09330_),
    .B1(net2789));
 sg13g2_nand3_1 _13615_ (.B(net2717),
    .C(_09328_),
    .A(net2789),
    .Y(_09331_));
 sg13g2_nand4_1 _13616_ (.B(net2717),
    .C(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .A(net2789),
    .Y(_09332_),
    .D(net2464));
 sg13g2_nor2_2 _13617_ (.A(_09326_),
    .B(_09332_),
    .Y(_09333_));
 sg13g2_nor2_1 _13618_ (.A(net2790),
    .B(_09333_),
    .Y(_00183_));
 sg13g2_xor2_1 _13619_ (.B(_09333_),
    .A(net2388),
    .X(_00185_));
 sg13g2_a21oi_1 _13620_ (.A1(net2388),
    .A2(_09333_),
    .Y(_09334_),
    .B1(net2934));
 sg13g2_nand2_1 _13621_ (.Y(_09335_),
    .A(net2934),
    .B(net2388));
 sg13g2_nor2_1 _13622_ (.A(_09331_),
    .B(_09335_),
    .Y(_09336_));
 sg13g2_nand3_1 _13623_ (.B(net2388),
    .C(_09333_),
    .A(net2934),
    .Y(_09337_));
 sg13g2_nor2_1 _13624_ (.A(net2935),
    .B(_09336_),
    .Y(_00186_));
 sg13g2_xnor2_1 _13625_ (.Y(_00187_),
    .A(net2769),
    .B(_09337_));
 sg13g2_a21oi_1 _13626_ (.A1(net2769),
    .A2(_09336_),
    .Y(_09338_),
    .B1(net2980));
 sg13g2_nand2_1 _13627_ (.Y(_09339_),
    .A(net2980),
    .B(net2769));
 sg13g2_nor2_1 _13628_ (.A(_09337_),
    .B(_09339_),
    .Y(_09340_));
 sg13g2_or4_1 _13629_ (.A(_09326_),
    .B(_09332_),
    .C(_09335_),
    .D(_09339_),
    .X(_09341_));
 sg13g2_nor2_1 _13630_ (.A(_09338_),
    .B(_09340_),
    .Y(_00188_));
 sg13g2_xnor2_1 _13631_ (.Y(_00189_),
    .A(net2570),
    .B(_09341_));
 sg13g2_a21oi_1 _13632_ (.A1(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .A2(_09340_),
    .Y(_09342_),
    .B1(net2516));
 sg13g2_nand2_1 _13633_ (.Y(_09343_),
    .A(net2516),
    .B(\soc_inst.cpu_core.csr_file.mtime[24] ));
 sg13g2_nor2_2 _13634_ (.A(_09341_),
    .B(_09343_),
    .Y(_09344_));
 sg13g2_nor2_1 _13635_ (.A(net2517),
    .B(_09344_),
    .Y(_00190_));
 sg13g2_nand2_1 _13636_ (.Y(_09345_),
    .A(net2075),
    .B(_09344_));
 sg13g2_xor2_1 _13637_ (.B(_09344_),
    .A(net2075),
    .X(_00191_));
 sg13g2_xnor2_1 _13638_ (.Y(_00192_),
    .A(net2318),
    .B(_09345_));
 sg13g2_nand3_1 _13639_ (.B(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .C(_09344_),
    .A(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .Y(_09346_));
 sg13g2_and4_1 _13640_ (.A(net1980),
    .B(net2318),
    .C(net2075),
    .D(_09344_),
    .X(_09347_));
 sg13g2_xnor2_1 _13641_ (.Y(_00193_),
    .A(net1980),
    .B(_09346_));
 sg13g2_xor2_1 _13642_ (.B(_09347_),
    .A(net2632),
    .X(_00194_));
 sg13g2_nand3_1 _13643_ (.B(net2632),
    .C(_09347_),
    .A(net3371),
    .Y(_09348_));
 sg13g2_a21o_1 _13644_ (.A2(_09347_),
    .A1(net2632),
    .B1(net3371),
    .X(_09349_));
 sg13g2_and2_1 _13645_ (.A(_09348_),
    .B(_09349_),
    .X(_00196_));
 sg13g2_and4_1 _13646_ (.A(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .B(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .C(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .D(_09347_),
    .X(_09350_));
 sg13g2_xnor2_1 _13647_ (.Y(_00197_),
    .A(net2891),
    .B(_09348_));
 sg13g2_xor2_1 _13648_ (.B(_09350_),
    .A(net2135),
    .X(_00198_));
 sg13g2_nand3_1 _13649_ (.B(net2135),
    .C(_09350_),
    .A(net3229),
    .Y(_09351_));
 sg13g2_a21o_1 _13650_ (.A2(_09350_),
    .A1(net2135),
    .B1(net3229),
    .X(_09352_));
 sg13g2_and2_1 _13651_ (.A(_09351_),
    .B(_09352_),
    .X(_00199_));
 sg13g2_and4_1 _13652_ (.A(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .B(net3229),
    .C(net2135),
    .D(_09350_),
    .X(_09353_));
 sg13g2_a21oi_1 _13653_ (.A1(_07906_),
    .A2(_09351_),
    .Y(_00200_),
    .B1(_09353_));
 sg13g2_and2_1 _13654_ (.A(net1199),
    .B(_09353_),
    .X(_09354_));
 sg13g2_xor2_1 _13655_ (.B(_09353_),
    .A(net1199),
    .X(_00201_));
 sg13g2_xor2_1 _13656_ (.B(_09354_),
    .A(net1482),
    .X(_00202_));
 sg13g2_and3_2 _13657_ (.X(_09355_),
    .A(net2058),
    .B(net1482),
    .C(_09354_));
 sg13g2_a21oi_1 _13658_ (.A1(net1482),
    .A2(_09354_),
    .Y(_09356_),
    .B1(net2058));
 sg13g2_nor2_1 _13659_ (.A(_09355_),
    .B(_09356_),
    .Y(_00203_));
 sg13g2_and2_1 _13660_ (.A(net1331),
    .B(_09355_),
    .X(_09357_));
 sg13g2_xor2_1 _13661_ (.B(_09355_),
    .A(net1331),
    .X(_00204_));
 sg13g2_xnor2_1 _13662_ (.Y(_00205_),
    .A(_07905_),
    .B(_09357_));
 sg13g2_nand3_1 _13663_ (.B(net3120),
    .C(_09357_),
    .A(net3377),
    .Y(_09358_));
 sg13g2_a21o_1 _13664_ (.A2(_09357_),
    .A1(net3120),
    .B1(net3377),
    .X(_09359_));
 sg13g2_and2_1 _13665_ (.A(_09358_),
    .B(_09359_),
    .X(_00207_));
 sg13g2_and4_1 _13666_ (.A(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .B(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .C(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .D(_09357_),
    .X(_09360_));
 sg13g2_xnor2_1 _13667_ (.Y(_00208_),
    .A(net1372),
    .B(_09358_));
 sg13g2_nand2_1 _13668_ (.Y(_09361_),
    .A(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .B(_09360_));
 sg13g2_xor2_1 _13669_ (.B(_09360_),
    .A(net1169),
    .X(_00209_));
 sg13g2_xnor2_1 _13670_ (.Y(_00210_),
    .A(net941),
    .B(_09361_));
 sg13g2_and3_1 _13671_ (.X(_09362_),
    .A(net941),
    .B(net1169),
    .C(_09360_));
 sg13g2_and2_1 _13672_ (.A(net627),
    .B(_09362_),
    .X(_09363_));
 sg13g2_xor2_1 _13673_ (.B(_09362_),
    .A(net627),
    .X(_00211_));
 sg13g2_xor2_1 _13674_ (.B(_09363_),
    .A(net1857),
    .X(_00212_));
 sg13g2_a21oi_1 _13675_ (.A1(net1857),
    .A2(_09363_),
    .Y(_09364_),
    .B1(net2011));
 sg13g2_nand3_1 _13676_ (.B(net1857),
    .C(_09363_),
    .A(net2011),
    .Y(_09365_));
 sg13g2_nor2b_1 _13677_ (.A(_09364_),
    .B_N(_09365_),
    .Y(_00213_));
 sg13g2_xnor2_1 _13678_ (.Y(_00214_),
    .A(net1140),
    .B(_09365_));
 sg13g2_nor2b_1 _13679_ (.A(net6543),
    .B_N(net405),
    .Y(_00001_));
 sg13g2_nand4_1 _13680_ (.B(_07878_),
    .C(net6485),
    .A(net1027),
    .Y(_09366_),
    .D(_08646_));
 sg13g2_nor2_1 _13681_ (.A(net6541),
    .B(net1028),
    .Y(_00005_));
 sg13g2_nor4_1 _13682_ (.A(net6543),
    .B(net6505),
    .C(_07875_),
    .D(_08652_),
    .Y(_00004_));
 sg13g2_nor3_1 _13683_ (.A(net6541),
    .B(_07877_),
    .C(_08658_),
    .Y(_00003_));
 sg13g2_nor3_1 _13684_ (.A(net227),
    .B(_08418_),
    .C(_08421_),
    .Y(_00002_));
 sg13g2_nor3_1 _13685_ (.A(_07784_),
    .B(_08907_),
    .C(_09300_),
    .Y(_00172_));
 sg13g2_and2_1 _13686_ (.A(_08667_),
    .B(net5564),
    .X(_09367_));
 sg13g2_nand2_1 _13687_ (.Y(_09368_),
    .A(_08908_),
    .B(net5336));
 sg13g2_mux2_1 _13688_ (.A0(net6470),
    .A1(net2247),
    .S(net5140),
    .X(_00321_));
 sg13g2_mux2_1 _13689_ (.A0(net6468),
    .A1(net2173),
    .S(net5140),
    .X(_00322_));
 sg13g2_nor2_1 _13690_ (.A(net6465),
    .B(net5140),
    .Y(_09369_));
 sg13g2_a21oi_1 _13691_ (.A1(_07955_),
    .A2(net5140),
    .Y(_00323_),
    .B1(_09369_));
 sg13g2_nor2_1 _13692_ (.A(net6463),
    .B(net5141),
    .Y(_09370_));
 sg13g2_a21oi_1 _13693_ (.A1(_07957_),
    .A2(net5140),
    .Y(_00324_),
    .B1(_09370_));
 sg13g2_nor2_1 _13694_ (.A(net6461),
    .B(net5140),
    .Y(_09371_));
 sg13g2_a21oi_1 _13695_ (.A1(_07959_),
    .A2(net5140),
    .Y(_00325_),
    .B1(_09371_));
 sg13g2_mux2_1 _13696_ (.A0(net6459),
    .A1(net2849),
    .S(net5141),
    .X(_00326_));
 sg13g2_mux2_1 _13697_ (.A0(net6457),
    .A1(net2844),
    .S(net5141),
    .X(_00327_));
 sg13g2_mux2_1 _13698_ (.A0(net6455),
    .A1(net2425),
    .S(net5140),
    .X(_00328_));
 sg13g2_mux2_1 _13699_ (.A0(net6454),
    .A1(net2568),
    .S(net5138),
    .X(_00329_));
 sg13g2_mux2_1 _13700_ (.A0(net6453),
    .A1(net2749),
    .S(net5138),
    .X(_00330_));
 sg13g2_mux2_1 _13701_ (.A0(net1533),
    .A1(net2824),
    .S(net5138),
    .X(_00331_));
 sg13g2_mux2_1 _13702_ (.A0(\soc_inst.core_mem_wdata[11] ),
    .A1(net2551),
    .S(net5138),
    .X(_00332_));
 sg13g2_nor2_1 _13703_ (.A(net1825),
    .B(net5139),
    .Y(_09372_));
 sg13g2_a21oi_1 _13704_ (.A1(_07964_),
    .A2(net5138),
    .Y(_00333_),
    .B1(_09372_));
 sg13g2_nor2_1 _13705_ (.A(net1321),
    .B(net5139),
    .Y(_09373_));
 sg13g2_a21oi_1 _13706_ (.A1(_07965_),
    .A2(net5138),
    .Y(_00334_),
    .B1(_09373_));
 sg13g2_nor2_1 _13707_ (.A(net1503),
    .B(net5139),
    .Y(_09374_));
 sg13g2_a21oi_1 _13708_ (.A1(_07966_),
    .A2(net5138),
    .Y(_00335_),
    .B1(_09374_));
 sg13g2_mux2_1 _13709_ (.A0(\soc_inst.core_mem_wdata[15] ),
    .A1(net2580),
    .S(net5138),
    .X(_00336_));
 sg13g2_a21oi_1 _13710_ (.A1(\soc_inst.spi_inst.cpha ),
    .A2(_08697_),
    .Y(_09375_),
    .B1(_08423_));
 sg13g2_o21ai_1 _13711_ (.B1(_09375_),
    .Y(_09376_),
    .A1(\soc_inst.spi_inst.cpha ),
    .A2(_08700_));
 sg13g2_nand2_1 _13712_ (.Y(_09377_),
    .A(\soc_inst.spi_inst.state[0] ),
    .B(\soc_inst.spi_inst.cpha ));
 sg13g2_nand4_1 _13713_ (.B(_00127_),
    .C(_09376_),
    .A(net1442),
    .Y(_09378_),
    .D(_09377_));
 sg13g2_o21ai_1 _13714_ (.B1(net1443),
    .Y(_00337_),
    .A1(_08186_),
    .A2(_09376_));
 sg13g2_xnor2_1 _13715_ (.Y(_09379_),
    .A(net2843),
    .B(net5017));
 sg13g2_nor2_1 _13716_ (.A(net6110),
    .B(_09379_),
    .Y(_00338_));
 sg13g2_a21oi_1 _13717_ (.A1(\soc_inst.spi_inst.bit_counter[0] ),
    .A2(net5016),
    .Y(_09380_),
    .B1(net2083));
 sg13g2_and3_1 _13718_ (.X(_09381_),
    .A(\soc_inst.spi_inst.bit_counter[0] ),
    .B(net2083),
    .C(net5017));
 sg13g2_nor3_1 _13719_ (.A(net6110),
    .B(net2084),
    .C(_09381_),
    .Y(_00339_));
 sg13g2_and4_1 _13720_ (.A(net2843),
    .B(net2083),
    .C(net2606),
    .D(_08702_),
    .X(_09382_));
 sg13g2_xnor2_1 _13721_ (.Y(_09383_),
    .A(net2606),
    .B(_09381_));
 sg13g2_nor2_1 _13722_ (.A(net6110),
    .B(net2607),
    .Y(_00340_));
 sg13g2_nor2_1 _13723_ (.A(net2428),
    .B(_09382_),
    .Y(_09384_));
 sg13g2_and2_1 _13724_ (.A(net2428),
    .B(_09382_),
    .X(_09385_));
 sg13g2_nor3_1 _13725_ (.A(net6110),
    .B(net2429),
    .C(_09385_),
    .Y(_00341_));
 sg13g2_nor2_1 _13726_ (.A(net2897),
    .B(_09385_),
    .Y(_09386_));
 sg13g2_and2_1 _13727_ (.A(net2897),
    .B(_09385_),
    .X(_09387_));
 sg13g2_nor3_1 _13728_ (.A(net6110),
    .B(_09386_),
    .C(_09387_),
    .Y(_00342_));
 sg13g2_a21oi_1 _13729_ (.A1(net2918),
    .A2(_09387_),
    .Y(_09388_),
    .B1(net6110));
 sg13g2_o21ai_1 _13730_ (.B1(_09388_),
    .Y(_09389_),
    .A1(net2918),
    .A2(_09387_));
 sg13g2_inv_1 _13731_ (.Y(_00343_),
    .A(_09389_));
 sg13g2_a21oi_1 _13732_ (.A1(_07804_),
    .A2(\soc_inst.spi_inst.state[0] ),
    .Y(_09390_),
    .B1(_08702_));
 sg13g2_a22oi_1 _13733_ (.Y(_09391_),
    .B1(net4920),
    .B2(net2730),
    .A2(net5016),
    .A1(net1));
 sg13g2_inv_1 _13734_ (.Y(_00344_),
    .A(_09391_));
 sg13g2_a22oi_1 _13735_ (.Y(_09392_),
    .B1(net4922),
    .B2(net2756),
    .A2(net5018),
    .A1(net2730));
 sg13g2_inv_1 _13736_ (.Y(_00345_),
    .A(_09392_));
 sg13g2_a22oi_1 _13737_ (.Y(_09393_),
    .B1(net4922),
    .B2(net2689),
    .A2(net5020),
    .A1(\soc_inst.spi_inst.rx_shift_reg[1] ));
 sg13g2_inv_1 _13738_ (.Y(_00346_),
    .A(net2690));
 sg13g2_a22oi_1 _13739_ (.Y(_09394_),
    .B1(net4923),
    .B2(net2850),
    .A2(net5021),
    .A1(net2689));
 sg13g2_inv_1 _13740_ (.Y(_00347_),
    .A(_09394_));
 sg13g2_a22oi_1 _13741_ (.Y(_09395_),
    .B1(net4922),
    .B2(net2327),
    .A2(net5021),
    .A1(\soc_inst.spi_inst.rx_shift_reg[3] ));
 sg13g2_inv_1 _13742_ (.Y(_00348_),
    .A(net2328));
 sg13g2_a22oi_1 _13743_ (.Y(_09396_),
    .B1(net4923),
    .B2(net2547),
    .A2(net5021),
    .A1(net2327));
 sg13g2_inv_1 _13744_ (.Y(_00349_),
    .A(_09396_));
 sg13g2_a22oi_1 _13745_ (.Y(_09397_),
    .B1(net4923),
    .B2(net2438),
    .A2(net5021),
    .A1(\soc_inst.spi_inst.rx_shift_reg[5] ));
 sg13g2_inv_1 _13746_ (.Y(_00350_),
    .A(net2439));
 sg13g2_a22oi_1 _13747_ (.Y(_09398_),
    .B1(net4923),
    .B2(net2600),
    .A2(net5021),
    .A1(net2438));
 sg13g2_inv_1 _13748_ (.Y(_00351_),
    .A(_09398_));
 sg13g2_a22oi_1 _13749_ (.Y(_09399_),
    .B1(net4923),
    .B2(net2554),
    .A2(net5022),
    .A1(\soc_inst.spi_inst.rx_shift_reg[7] ));
 sg13g2_inv_1 _13750_ (.Y(_00352_),
    .A(net2555));
 sg13g2_a22oi_1 _13751_ (.Y(_09400_),
    .B1(net4922),
    .B2(net2397),
    .A2(net5022),
    .A1(\soc_inst.spi_inst.rx_shift_reg[8] ));
 sg13g2_inv_1 _13752_ (.Y(_00353_),
    .A(net2398));
 sg13g2_a22oi_1 _13753_ (.Y(_09401_),
    .B1(net4922),
    .B2(net2229),
    .A2(net5018),
    .A1(\soc_inst.spi_inst.rx_shift_reg[9] ));
 sg13g2_inv_1 _13754_ (.Y(_00354_),
    .A(net2230));
 sg13g2_a22oi_1 _13755_ (.Y(_09402_),
    .B1(net4922),
    .B2(net2515),
    .A2(net5018),
    .A1(net2229));
 sg13g2_inv_1 _13756_ (.Y(_00355_),
    .A(_09402_));
 sg13g2_a22oi_1 _13757_ (.Y(_09403_),
    .B1(net4922),
    .B2(net2156),
    .A2(net5018),
    .A1(\soc_inst.spi_inst.rx_shift_reg[11] ));
 sg13g2_inv_1 _13758_ (.Y(_00356_),
    .A(net2157));
 sg13g2_a22oi_1 _13759_ (.Y(_09404_),
    .B1(net4923),
    .B2(net2922),
    .A2(net5018),
    .A1(net2156));
 sg13g2_inv_1 _13760_ (.Y(_00357_),
    .A(_09404_));
 sg13g2_a22oi_1 _13761_ (.Y(_09405_),
    .B1(net4923),
    .B2(net2485),
    .A2(net5021),
    .A1(\soc_inst.spi_inst.rx_shift_reg[13] ));
 sg13g2_inv_1 _13762_ (.Y(_00358_),
    .A(net2486));
 sg13g2_a22oi_1 _13763_ (.Y(_09406_),
    .B1(net4922),
    .B2(net2481),
    .A2(net5021),
    .A1(\soc_inst.spi_inst.rx_shift_reg[14] ));
 sg13g2_inv_1 _13764_ (.Y(_00359_),
    .A(net2482));
 sg13g2_a22oi_1 _13765_ (.Y(_09407_),
    .B1(net4921),
    .B2(net1557),
    .A2(net5018),
    .A1(\soc_inst.spi_inst.rx_shift_reg[15] ));
 sg13g2_inv_1 _13766_ (.Y(_00360_),
    .A(net1558));
 sg13g2_a22oi_1 _13767_ (.Y(_09408_),
    .B1(net4921),
    .B2(net1723),
    .A2(net5018),
    .A1(net1557));
 sg13g2_inv_1 _13768_ (.Y(_00361_),
    .A(_09408_));
 sg13g2_a22oi_1 _13769_ (.Y(_09409_),
    .B1(net4921),
    .B2(net1365),
    .A2(net5018),
    .A1(\soc_inst.spi_inst.rx_shift_reg[17] ));
 sg13g2_inv_1 _13770_ (.Y(_00362_),
    .A(net1366));
 sg13g2_a22oi_1 _13771_ (.Y(_09410_),
    .B1(net4921),
    .B2(net1622),
    .A2(net5019),
    .A1(net1365));
 sg13g2_inv_1 _13772_ (.Y(_00363_),
    .A(_09410_));
 sg13g2_a22oi_1 _13773_ (.Y(_09411_),
    .B1(net4920),
    .B2(net1361),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[19] ));
 sg13g2_inv_1 _13774_ (.Y(_00364_),
    .A(net1362));
 sg13g2_a22oi_1 _13775_ (.Y(_09412_),
    .B1(net4924),
    .B2(net1162),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[20] ));
 sg13g2_inv_1 _13776_ (.Y(_00365_),
    .A(net1163));
 sg13g2_a22oi_1 _13777_ (.Y(_09413_),
    .B1(net4924),
    .B2(net1845),
    .A2(net5020),
    .A1(net1162));
 sg13g2_inv_1 _13778_ (.Y(_00366_),
    .A(_09413_));
 sg13g2_a22oi_1 _13779_ (.Y(_09414_),
    .B1(net4921),
    .B2(net2391),
    .A2(net5020),
    .A1(net1845));
 sg13g2_inv_1 _13780_ (.Y(_00367_),
    .A(_09414_));
 sg13g2_a22oi_1 _13781_ (.Y(_09415_),
    .B1(net4920),
    .B2(net1125),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[23] ));
 sg13g2_inv_1 _13782_ (.Y(_00368_),
    .A(net1126));
 sg13g2_a22oi_1 _13783_ (.Y(_09416_),
    .B1(net4920),
    .B2(net1542),
    .A2(net5019),
    .A1(net1125));
 sg13g2_inv_1 _13784_ (.Y(_00369_),
    .A(_09416_));
 sg13g2_a22oi_1 _13785_ (.Y(_09417_),
    .B1(net4920),
    .B2(net1467),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[25] ));
 sg13g2_inv_1 _13786_ (.Y(_00370_),
    .A(net1468));
 sg13g2_a22oi_1 _13787_ (.Y(_09418_),
    .B1(net4921),
    .B2(net1301),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[26] ));
 sg13g2_inv_1 _13788_ (.Y(_00371_),
    .A(net1302));
 sg13g2_a22oi_1 _13789_ (.Y(_09419_),
    .B1(net4921),
    .B2(net1160),
    .A2(net5016),
    .A1(\soc_inst.spi_inst.rx_shift_reg[27] ));
 sg13g2_inv_1 _13790_ (.Y(_00372_),
    .A(net1161));
 sg13g2_a22oi_1 _13791_ (.Y(_09420_),
    .B1(net4920),
    .B2(net1146),
    .A2(net5016),
    .A1(\soc_inst.spi_inst.rx_shift_reg[28] ));
 sg13g2_inv_1 _13792_ (.Y(_00373_),
    .A(net1147));
 sg13g2_a22oi_1 _13793_ (.Y(_09421_),
    .B1(net4920),
    .B2(net1054),
    .A2(net5016),
    .A1(\soc_inst.spi_inst.rx_shift_reg[29] ));
 sg13g2_inv_1 _13794_ (.Y(_00374_),
    .A(net1055));
 sg13g2_a22oi_1 _13795_ (.Y(_09422_),
    .B1(net4920),
    .B2(net457),
    .A2(net5019),
    .A1(\soc_inst.spi_inst.rx_shift_reg[30] ));
 sg13g2_inv_1 _13796_ (.Y(_00375_),
    .A(net458));
 sg13g2_nand4_1 _13797_ (.B(_07890_),
    .C(_07891_),
    .A(\soc_inst.pwm_inst.channel_idx [0]),
    .Y(_09423_),
    .D(_07892_));
 sg13g2_nor2_2 _13798_ (.A(net6047),
    .B(_09423_),
    .Y(_09424_));
 sg13g2_nand2b_1 _13799_ (.Y(_09425_),
    .B(net5530),
    .A_N(_08677_));
 sg13g2_mux2_1 _13800_ (.A0(net6454),
    .A1(net3158),
    .S(net5137),
    .X(_00376_));
 sg13g2_and2_1 _13801_ (.A(_08667_),
    .B(net6056),
    .X(_09426_));
 sg13g2_nand2b_1 _13802_ (.Y(_09427_),
    .B(_09426_),
    .A_N(_08677_));
 sg13g2_nor2_1 _13803_ (.A(net6470),
    .B(_09427_),
    .Y(_09428_));
 sg13g2_a21oi_1 _13804_ (.A1(_07899_),
    .A2(_09427_),
    .Y(_00377_),
    .B1(_09428_));
 sg13g2_nand2_1 _13805_ (.Y(_09429_),
    .A(net2095),
    .B(net5135));
 sg13g2_o21ai_1 _13806_ (.B1(_09429_),
    .Y(_00378_),
    .A1(net6471),
    .A2(net5135));
 sg13g2_nor2_1 _13807_ (.A(_07784_),
    .B(net5136),
    .Y(_09430_));
 sg13g2_a21oi_1 _13808_ (.A1(_07798_),
    .A2(net5136),
    .Y(_00379_),
    .B1(_09430_));
 sg13g2_nand2_1 _13809_ (.Y(_09431_),
    .A(net1205),
    .B(net5135));
 sg13g2_o21ai_1 _13810_ (.B1(_09431_),
    .Y(_00380_),
    .A1(net6466),
    .A2(net5135));
 sg13g2_nand2_1 _13811_ (.Y(_09432_),
    .A(net2065),
    .B(net5135));
 sg13g2_o21ai_1 _13812_ (.B1(_09432_),
    .Y(_00381_),
    .A1(net6464),
    .A2(net5136));
 sg13g2_nand2_1 _13813_ (.Y(_09433_),
    .A(net1496),
    .B(net5135));
 sg13g2_o21ai_1 _13814_ (.B1(_09433_),
    .Y(_00382_),
    .A1(net6462),
    .A2(net5135));
 sg13g2_mux2_1 _13815_ (.A0(net6459),
    .A1(net2996),
    .S(net5137),
    .X(_00383_));
 sg13g2_mux2_1 _13816_ (.A0(net6458),
    .A1(net2913),
    .S(net5135),
    .X(_00384_));
 sg13g2_nor2_1 _13817_ (.A(net6456),
    .B(net5136),
    .Y(_09434_));
 sg13g2_a21oi_1 _13818_ (.A1(_07896_),
    .A2(net5136),
    .Y(_00385_),
    .B1(_09434_));
 sg13g2_a22oi_1 _13819_ (.Y(_09435_),
    .B1(net1480),
    .B2(_09312_),
    .A2(\soc_inst.spi_inst.state[0] ),
    .A1(net850));
 sg13g2_inv_1 _13820_ (.Y(_00386_),
    .A(net1481));
 sg13g2_mux2_1 _13821_ (.A0(net6453),
    .A1(net3185),
    .S(net5137),
    .X(_00387_));
 sg13g2_nor2b_1 _13822_ (.A(\soc_inst.gpio_inst.gpio_sync2[0] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[0] ),
    .Y(_09436_));
 sg13g2_a21oi_1 _13823_ (.A1(net93),
    .A2(_09436_),
    .Y(_09437_),
    .B1(net978));
 sg13g2_nor3_1 _13824_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(_08228_),
    .C(_08676_),
    .Y(_09438_));
 sg13g2_nand3_1 _13825_ (.B(_08237_),
    .C(_09438_),
    .A(net6205),
    .Y(_09439_));
 sg13g2_nor3_2 _13826_ (.A(net6051),
    .B(_09423_),
    .C(_09439_),
    .Y(_09440_));
 sg13g2_nor3_2 _13827_ (.A(\soc_inst.core_mem_addr[13] ),
    .B(_08231_),
    .C(_08676_),
    .Y(_09441_));
 sg13g2_a21oi_1 _13828_ (.A1(net6471),
    .A2(_09440_),
    .Y(_00388_),
    .B1(net979));
 sg13g2_mux2_1 _13829_ (.A0(net6546),
    .A1(net6465),
    .S(_08795_),
    .X(_00389_));
 sg13g2_mux2_1 _13830_ (.A0(net2192),
    .A1(net6463),
    .S(_08795_),
    .X(_00390_));
 sg13g2_mux2_1 _13831_ (.A0(net1677),
    .A1(net6461),
    .S(_08795_),
    .X(_00391_));
 sg13g2_nor4_1 _13832_ (.A(net111),
    .B(net13),
    .C(net6546),
    .D(_09273_),
    .Y(_09442_));
 sg13g2_a21o_1 _13833_ (.A2(net112),
    .A1(_09272_),
    .B1(net90),
    .X(_00392_));
 sg13g2_nor2_1 _13834_ (.A(_08672_),
    .B(_08794_),
    .Y(_09443_));
 sg13g2_nor2_1 _13835_ (.A(net1934),
    .B(net5134),
    .Y(_09444_));
 sg13g2_a21oi_1 _13836_ (.A1(net6470),
    .A2(net5134),
    .Y(_00393_),
    .B1(_09444_));
 sg13g2_nor2_1 _13837_ (.A(net2306),
    .B(net5133),
    .Y(_09445_));
 sg13g2_a21oi_1 _13838_ (.A1(net6468),
    .A2(net5133),
    .Y(_00394_),
    .B1(_09445_));
 sg13g2_nor2_1 _13839_ (.A(net2030),
    .B(net5133),
    .Y(_09446_));
 sg13g2_a21oi_1 _13840_ (.A1(net6465),
    .A2(net5133),
    .Y(_00395_),
    .B1(_09446_));
 sg13g2_nor2_1 _13841_ (.A(net2593),
    .B(net5133),
    .Y(_09447_));
 sg13g2_a21oi_1 _13842_ (.A1(net6463),
    .A2(net5133),
    .Y(_00396_),
    .B1(_09447_));
 sg13g2_nor2_1 _13843_ (.A(net2598),
    .B(net5134),
    .Y(_09448_));
 sg13g2_a21oi_1 _13844_ (.A1(net6461),
    .A2(net5134),
    .Y(_00397_),
    .B1(_09448_));
 sg13g2_mux2_1 _13845_ (.A0(net2635),
    .A1(net6460),
    .S(net5134),
    .X(_00398_));
 sg13g2_mux2_1 _13846_ (.A0(net2563),
    .A1(net6457),
    .S(net5134),
    .X(_00399_));
 sg13g2_nor2_1 _13847_ (.A(net2158),
    .B(net5133),
    .Y(_09449_));
 sg13g2_a21oi_1 _13848_ (.A1(net6455),
    .A2(net5133),
    .Y(_00400_),
    .B1(_09449_));
 sg13g2_o21ai_1 _13849_ (.B1(_09225_),
    .Y(_09450_),
    .A1(net6539),
    .A2(_08826_));
 sg13g2_nor2_1 _13850_ (.A(_08404_),
    .B(_09450_),
    .Y(_09451_));
 sg13g2_a21oi_1 _13851_ (.A1(net5565),
    .A2(_09450_),
    .Y(_09452_),
    .B1(_09451_));
 sg13g2_o21ai_1 _13852_ (.B1(_09452_),
    .Y(_09453_),
    .A1(net5565),
    .A2(_09231_));
 sg13g2_nor4_1 _13853_ (.A(net6540),
    .B(net6538),
    .C(_08828_),
    .D(_09453_),
    .Y(_09454_));
 sg13g2_mux2_1 _13854_ (.A0(_09454_),
    .A1(_09453_),
    .S(net3121),
    .X(_00401_));
 sg13g2_nand2_1 _13855_ (.Y(_09455_),
    .A(\soc_inst.i2c_inst.bit_cnt[0] ),
    .B(\soc_inst.i2c_inst.bit_cnt[1] ));
 sg13g2_xor2_1 _13856_ (.B(net2965),
    .A(\soc_inst.i2c_inst.bit_cnt[0] ),
    .X(_09456_));
 sg13g2_a22oi_1 _13857_ (.Y(_09457_),
    .B1(_09454_),
    .B2(_09456_),
    .A2(_09453_),
    .A1(net2965));
 sg13g2_inv_1 _13858_ (.Y(_00402_),
    .A(net2966));
 sg13g2_nand3_1 _13859_ (.B(net2965),
    .C(net1013),
    .A(net3121),
    .Y(_09458_));
 sg13g2_a21oi_1 _13860_ (.A1(_09266_),
    .A2(_09458_),
    .Y(_09459_),
    .B1(_09453_));
 sg13g2_nor2_1 _13861_ (.A(_09453_),
    .B(_09455_),
    .Y(_09460_));
 sg13g2_nor2_1 _13862_ (.A(net1013),
    .B(_09460_),
    .Y(_09461_));
 sg13g2_nor2_1 _13863_ (.A(_09459_),
    .B(net1014),
    .Y(_00403_));
 sg13g2_nor2b_1 _13864_ (.A(_09459_),
    .B_N(net3186),
    .Y(_09462_));
 sg13g2_nor2_1 _13865_ (.A(net3186),
    .B(_09458_),
    .Y(_09463_));
 sg13g2_a21oi_1 _13866_ (.A1(_09454_),
    .A2(_09463_),
    .Y(_09464_),
    .B1(_09462_));
 sg13g2_inv_1 _13867_ (.Y(_00404_),
    .A(net3187));
 sg13g2_nor2_1 _13868_ (.A(_08831_),
    .B(_09274_),
    .Y(_09465_));
 sg13g2_nor2_2 _13869_ (.A(net6539),
    .B(_09228_),
    .Y(_09466_));
 sg13g2_nand2_1 _13870_ (.Y(_09467_),
    .A(net6537),
    .B(_09466_));
 sg13g2_nand3b_1 _13871_ (.B(_09465_),
    .C(_09467_),
    .Y(_09468_),
    .A_N(_08798_));
 sg13g2_o21ai_1 _13872_ (.B1(_08818_),
    .Y(_09469_),
    .A1(_09226_),
    .A2(_09468_));
 sg13g2_nor2_1 _13873_ (.A(_08798_),
    .B(_09265_),
    .Y(_09470_));
 sg13g2_nor3_1 _13874_ (.A(_08405_),
    .B(_08798_),
    .C(_09265_),
    .Y(_09471_));
 sg13g2_a21oi_1 _13875_ (.A1(net6540),
    .A2(net6538),
    .Y(_09472_),
    .B1(_08402_));
 sg13g2_a21o_1 _13876_ (.A2(_09228_),
    .A1(_08828_),
    .B1(_09472_),
    .X(_09473_));
 sg13g2_o21ai_1 _13877_ (.B1(_09471_),
    .Y(_09474_),
    .A1(net5565),
    .A2(_09473_));
 sg13g2_nand2b_1 _13878_ (.Y(_09475_),
    .B(_09265_),
    .A_N(_09272_));
 sg13g2_nand3_1 _13879_ (.B(_09474_),
    .C(_09475_),
    .A(_09469_),
    .Y(_09476_));
 sg13g2_nand2_1 _13880_ (.Y(_09477_),
    .A(net6539),
    .B(_09265_));
 sg13g2_a21oi_1 _13881_ (.A1(net6546),
    .A2(net2192),
    .Y(_09478_),
    .B1(_09477_));
 sg13g2_o21ai_1 _13882_ (.B1(_09266_),
    .Y(_09479_),
    .A1(net6546),
    .A2(net2049));
 sg13g2_inv_1 _13883_ (.Y(_09480_),
    .A(_09479_));
 sg13g2_nor3_1 _13884_ (.A(_09470_),
    .B(_09478_),
    .C(_09480_),
    .Y(_09481_));
 sg13g2_mux2_1 _13885_ (.A0(_09481_),
    .A1(net111),
    .S(_09476_),
    .X(_00405_));
 sg13g2_nor3_1 _13886_ (.A(_08401_),
    .B(_08403_),
    .C(_08827_),
    .Y(_09482_));
 sg13g2_a22oi_1 _13887_ (.Y(_09483_),
    .B1(_08830_),
    .B2(net6540),
    .A2(_08825_),
    .A1(_08401_));
 sg13g2_nand2b_1 _13888_ (.Y(_09484_),
    .B(_09483_),
    .A_N(_09466_));
 sg13g2_a22oi_1 _13889_ (.Y(_09485_),
    .B1(_09484_),
    .B2(_08814_),
    .A2(_09482_),
    .A1(_09273_));
 sg13g2_a221oi_1 _13890_ (.B2(_08814_),
    .C1(_08831_),
    .B1(_09482_),
    .A1(_08401_),
    .Y(_09486_),
    .A2(_08826_));
 sg13g2_mux2_1 _13891_ (.A0(net1615),
    .A1(_09486_),
    .S(_09485_),
    .X(_00406_));
 sg13g2_mux2_1 _13892_ (.A0(net6),
    .A1(net2538),
    .S(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_latched ),
    .X(_00407_));
 sg13g2_mux2_1 _13893_ (.A0(net7),
    .A1(net2322),
    .S(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_latched ),
    .X(_00408_));
 sg13g2_nor2_1 _13894_ (.A(net2143),
    .B(net5174),
    .Y(_09487_));
 sg13g2_a21oi_1 _13895_ (.A1(net6470),
    .A2(net5174),
    .Y(_00409_),
    .B1(_09487_));
 sg13g2_nor2_1 _13896_ (.A(net2181),
    .B(net5174),
    .Y(_09488_));
 sg13g2_a21oi_1 _13897_ (.A1(net6468),
    .A2(net5174),
    .Y(_00410_),
    .B1(_09488_));
 sg13g2_nor2_1 _13898_ (.A(net2595),
    .B(net5174),
    .Y(_09489_));
 sg13g2_a21oi_1 _13899_ (.A1(net6465),
    .A2(net5174),
    .Y(_00411_),
    .B1(_09489_));
 sg13g2_nor2_1 _13900_ (.A(net2062),
    .B(net5174),
    .Y(_09490_));
 sg13g2_a21oi_1 _13901_ (.A1(net6463),
    .A2(net5174),
    .Y(_00412_),
    .B1(_09490_));
 sg13g2_nor2_1 _13902_ (.A(net2122),
    .B(net5173),
    .Y(_09491_));
 sg13g2_a21oi_1 _13903_ (.A1(net6461),
    .A2(net5173),
    .Y(_00413_),
    .B1(_09491_));
 sg13g2_nor2_1 _13904_ (.A(net1910),
    .B(net5173),
    .Y(_09492_));
 sg13g2_a21oi_1 _13905_ (.A1(net6459),
    .A2(net5173),
    .Y(_00414_),
    .B1(_09492_));
 sg13g2_nor2_1 _13906_ (.A(net1829),
    .B(net5173),
    .Y(_09493_));
 sg13g2_a21oi_1 _13907_ (.A1(net6458),
    .A2(net5173),
    .Y(_00415_),
    .B1(_09493_));
 sg13g2_nor2_1 _13908_ (.A(net1760),
    .B(net5173),
    .Y(_09494_));
 sg13g2_a21oi_1 _13909_ (.A1(net6455),
    .A2(net5173),
    .Y(_00416_),
    .B1(_09494_));
 sg13g2_nor2_1 _13910_ (.A(net2651),
    .B(net5172),
    .Y(_09495_));
 sg13g2_a21oi_1 _13911_ (.A1(net6454),
    .A2(net5172),
    .Y(_00417_),
    .B1(_09495_));
 sg13g2_nor2_1 _13912_ (.A(net2625),
    .B(net5172),
    .Y(_09496_));
 sg13g2_a21oi_1 _13913_ (.A1(net6453),
    .A2(net5172),
    .Y(_00418_),
    .B1(_09496_));
 sg13g2_nor2_1 _13914_ (.A(net1777),
    .B(net5170),
    .Y(_09497_));
 sg13g2_a21oi_1 _13915_ (.A1(net1533),
    .A2(net5170),
    .Y(_00419_),
    .B1(_09497_));
 sg13g2_nor2_1 _13916_ (.A(net1678),
    .B(net5170),
    .Y(_09498_));
 sg13g2_a21oi_1 _13917_ (.A1(\soc_inst.core_mem_wdata[11] ),
    .A2(net5170),
    .Y(_00420_),
    .B1(_09498_));
 sg13g2_nor2_1 _13918_ (.A(net2039),
    .B(net5170),
    .Y(_09499_));
 sg13g2_a21oi_1 _13919_ (.A1(net1825),
    .A2(net5171),
    .Y(_00421_),
    .B1(_09499_));
 sg13g2_nor2_1 _13920_ (.A(net2036),
    .B(net5170),
    .Y(_09500_));
 sg13g2_a21oi_1 _13921_ (.A1(net1321),
    .A2(net5171),
    .Y(_00422_),
    .B1(_09500_));
 sg13g2_nor2_1 _13922_ (.A(net2317),
    .B(net5171),
    .Y(_09501_));
 sg13g2_a21oi_1 _13923_ (.A1(net1503),
    .A2(net5171),
    .Y(_00423_),
    .B1(_09501_));
 sg13g2_nor2_1 _13924_ (.A(net2055),
    .B(net5170),
    .Y(_09502_));
 sg13g2_a21oi_1 _13925_ (.A1(\soc_inst.core_mem_wdata[15] ),
    .A2(net5171),
    .Y(_00424_),
    .B1(_09502_));
 sg13g2_nor2_1 _13926_ (.A(net2024),
    .B(net722),
    .Y(_09503_));
 sg13g2_a21oi_1 _13927_ (.A1(_07784_),
    .A2(net722),
    .Y(_00425_),
    .B1(_09503_));
 sg13g2_mux2_1 _13928_ (.A0(net6545),
    .A1(net6466),
    .S(net722),
    .X(_00426_));
 sg13g2_and2_1 _13929_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[4] ),
    .B(\soc_inst.cpu_core.mem_reg_we ),
    .X(_09504_));
 sg13g2_nand2_2 _13930_ (.Y(_09505_),
    .A(\soc_inst.cpu_core._unused_mem_rd_addr[4] ),
    .B(\soc_inst.cpu_core.mem_reg_we ));
 sg13g2_nand2_2 _13931_ (.Y(_09506_),
    .A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ));
 sg13g2_inv_2 _13932_ (.Y(_09507_),
    .A(_09506_));
 sg13g2_nand2_1 _13933_ (.Y(_09508_),
    .A(net6214),
    .B(net6217));
 sg13g2_nor3_2 _13934_ (.A(_09505_),
    .B(_09506_),
    .C(_09508_),
    .Y(_09509_));
 sg13g2_nor2_1 _13935_ (.A(\soc_inst.cpu_core.mem_instr[5] ),
    .B(\soc_inst.cpu_core.mem_instr[6] ),
    .Y(_09510_));
 sg13g2_and3_1 _13936_ (.X(_09511_),
    .A(_00260_),
    .B(_08985_),
    .C(_09510_));
 sg13g2_nand3_1 _13937_ (.B(_08985_),
    .C(_09510_),
    .A(_00260_),
    .Y(_09512_));
 sg13g2_nor2_2 _13938_ (.A(net6172),
    .B(net6168),
    .Y(_09513_));
 sg13g2_nand2_2 _13939_ (.Y(_09514_),
    .A(net6301),
    .B(net6294));
 sg13g2_nor3_2 _13940_ (.A(net6105),
    .B(net6031),
    .C(_09513_),
    .Y(_09515_));
 sg13g2_nor2_2 _13941_ (.A(_08982_),
    .B(_09003_),
    .Y(_09516_));
 sg13g2_a22oi_1 _13942_ (.Y(_09517_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .A2(net5348),
    .A1(\soc_inst.cpu_core.csr_file.mepc[0] ));
 sg13g2_a22oi_1 _13943_ (.Y(_09518_),
    .B1(net5156),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[0] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[0] ));
 sg13g2_a22oi_1 _13944_ (.Y(_09519_),
    .B1(net5536),
    .B2(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .A2(net5542),
    .A1(\soc_inst.cpu_core.csr_file.mtime[32] ));
 sg13g2_nand2_1 _13945_ (.Y(_09520_),
    .A(net5553),
    .B(_09519_));
 sg13g2_a221oi_1 _13946_ (.B2(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .C1(_09520_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .Y(_09521_),
    .A2(net5342));
 sg13g2_nand3_1 _13947_ (.B(_09518_),
    .C(_09521_),
    .A(_09517_),
    .Y(_09522_));
 sg13g2_a21oi_1 _13948_ (.A1(_07886_),
    .A2(net5547),
    .Y(_09523_),
    .B1(net6032));
 sg13g2_a22oi_1 _13949_ (.Y(_09524_),
    .B1(_09522_),
    .B2(_09523_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[0] ));
 sg13g2_nor2_1 _13950_ (.A(net1640),
    .B(net6036),
    .Y(_09525_));
 sg13g2_a21oi_1 _13951_ (.A1(net6036),
    .A2(net4997),
    .Y(_00427_),
    .B1(_09525_));
 sg13g2_a22oi_1 _13952_ (.Y(_09526_),
    .B1(net5155),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[1] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[1] ));
 sg13g2_a22oi_1 _13953_ (.Y(_09527_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .A2(net5348),
    .A1(\soc_inst.cpu_core.csr_file.mepc[1] ));
 sg13g2_a22oi_1 _13954_ (.Y(_09528_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[33] ));
 sg13g2_nand2_1 _13955_ (.Y(_09529_),
    .A(net5555),
    .B(_09528_));
 sg13g2_a221oi_1 _13956_ (.B2(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .C1(_09529_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .Y(_09530_),
    .A2(net5342));
 sg13g2_nand3_1 _13957_ (.B(_09527_),
    .C(_09530_),
    .A(_09526_),
    .Y(_09531_));
 sg13g2_a21oi_1 _13958_ (.A1(_07885_),
    .A2(net5547),
    .Y(_09532_),
    .B1(net6032));
 sg13g2_a22oi_1 _13959_ (.Y(_09533_),
    .B1(_09531_),
    .B2(_09532_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[1] ));
 sg13g2_nor2_1 _13960_ (.A(net1916),
    .B(net6036),
    .Y(_09534_));
 sg13g2_a21oi_1 _13961_ (.A1(net6036),
    .A2(net4990),
    .Y(_00428_),
    .B1(_09534_));
 sg13g2_a22oi_1 _13962_ (.Y(_09535_),
    .B1(net5155),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[2] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[2] ));
 sg13g2_nand2_2 _13963_ (.Y(_09536_),
    .A(net5552),
    .B(_09021_));
 sg13g2_a221oi_1 _13964_ (.B2(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .C1(_09536_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .Y(_09537_),
    .A2(net5544));
 sg13g2_a22oi_1 _13965_ (.Y(_09538_),
    .B1(net5341),
    .B2(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .A2(net5540),
    .A1(\soc_inst.cpu_core.csr_file.mtime[2] ));
 sg13g2_a22oi_1 _13966_ (.Y(_09539_),
    .B1(net5335),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .A2(net5347),
    .A1(\soc_inst.cpu_core.csr_file.mepc[2] ));
 sg13g2_nand4_1 _13967_ (.B(_09537_),
    .C(_09538_),
    .A(_09535_),
    .Y(_09540_),
    .D(_09539_));
 sg13g2_a21oi_1 _13968_ (.A1(_07887_),
    .A2(net5548),
    .Y(_09541_),
    .B1(net6032));
 sg13g2_a22oi_1 _13969_ (.Y(_09542_),
    .B1(_09540_),
    .B2(_09541_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[2] ));
 sg13g2_nor2_1 _13970_ (.A(net1662),
    .B(net6036),
    .Y(_09543_));
 sg13g2_a21oi_1 _13971_ (.A1(net6036),
    .A2(net4984),
    .Y(_00429_),
    .B1(_09543_));
 sg13g2_a22oi_1 _13972_ (.Y(_09544_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[35] ));
 sg13g2_nand2_1 _13973_ (.Y(_09545_),
    .A(net5554),
    .B(_09544_));
 sg13g2_a221oi_1 _13974_ (.B2(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .C1(_09545_),
    .B1(net5150),
    .A1(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .Y(_09546_),
    .A2(net5342));
 sg13g2_a22oi_1 _13975_ (.Y(_09547_),
    .B1(net5348),
    .B2(\soc_inst.cpu_core.csr_file.mepc[3] ),
    .A2(net5155),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[3] ));
 sg13g2_a22oi_1 _13976_ (.Y(_09548_),
    .B1(net5335),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .A2(net5353),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[3] ));
 sg13g2_nand3_1 _13977_ (.B(_09547_),
    .C(_09548_),
    .A(_09546_),
    .Y(_09549_));
 sg13g2_a21oi_1 _13978_ (.A1(_07888_),
    .A2(net5547),
    .Y(_09550_),
    .B1(net6032));
 sg13g2_a22oi_1 _13979_ (.Y(_09551_),
    .B1(_09549_),
    .B2(_09550_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[3] ));
 sg13g2_nor2_1 _13980_ (.A(net1915),
    .B(net6035),
    .Y(_09552_));
 sg13g2_a21oi_1 _13981_ (.A1(net6035),
    .A2(net4982),
    .Y(_00430_),
    .B1(_09552_));
 sg13g2_a22oi_1 _13982_ (.Y(_09553_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[36] ));
 sg13g2_nand2_1 _13983_ (.Y(_09554_),
    .A(net5555),
    .B(_09553_));
 sg13g2_a221oi_1 _13984_ (.B2(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .C1(_09554_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .Y(_09555_),
    .A2(net5341));
 sg13g2_a22oi_1 _13985_ (.Y(_09556_),
    .B1(net5156),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[4] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[4] ));
 sg13g2_a22oi_1 _13986_ (.Y(_09557_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .A2(net5348),
    .A1(\soc_inst.cpu_core.csr_file.mepc[4] ));
 sg13g2_nand3_1 _13987_ (.B(_09556_),
    .C(_09557_),
    .A(_09555_),
    .Y(_09558_));
 sg13g2_a21oi_1 _13988_ (.A1(_07889_),
    .A2(net5547),
    .Y(_09559_),
    .B1(net6033));
 sg13g2_a22oi_1 _13989_ (.Y(_09560_),
    .B1(_09558_),
    .B2(_09559_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[4] ));
 sg13g2_nor2_1 _13990_ (.A(net2033),
    .B(net6041),
    .Y(_09561_));
 sg13g2_a21oi_1 _13991_ (.A1(net6041),
    .A2(net4975),
    .Y(_00431_),
    .B1(_09561_));
 sg13g2_a22oi_1 _13992_ (.Y(_09562_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[37] ));
 sg13g2_nand2_1 _13993_ (.Y(_09563_),
    .A(net5554),
    .B(_09562_));
 sg13g2_a221oi_1 _13994_ (.B2(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .C1(_09563_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .Y(_09564_),
    .A2(net5341));
 sg13g2_a22oi_1 _13995_ (.Y(_09565_),
    .B1(net5347),
    .B2(\soc_inst.cpu_core.csr_file.mepc[5] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[5] ));
 sg13g2_a22oi_1 _13996_ (.Y(_09566_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .A2(net5155),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[5] ));
 sg13g2_nand3_1 _13997_ (.B(_09565_),
    .C(_09566_),
    .A(_09564_),
    .Y(_09567_));
 sg13g2_a21oi_1 _13998_ (.A1(_07890_),
    .A2(net5547),
    .Y(_09568_),
    .B1(net6033));
 sg13g2_a22oi_1 _13999_ (.Y(_09569_),
    .B1(_09567_),
    .B2(_09568_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[5] ));
 sg13g2_nor2_1 _14000_ (.A(net2245),
    .B(net6042),
    .Y(_09570_));
 sg13g2_a21oi_1 _14001_ (.A1(net6042),
    .A2(net4973),
    .Y(_00432_),
    .B1(_09570_));
 sg13g2_a22oi_1 _14002_ (.Y(_09571_),
    .B1(net5347),
    .B2(\soc_inst.cpu_core.csr_file.mepc[6] ),
    .A2(net5353),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[6] ));
 sg13g2_a22oi_1 _14003_ (.Y(_09572_),
    .B1(net5335),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .A2(net5157),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[6] ));
 sg13g2_a22oi_1 _14004_ (.Y(_09573_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[38] ));
 sg13g2_nand2_1 _14005_ (.Y(_09574_),
    .A(net5554),
    .B(_09573_));
 sg13g2_a221oi_1 _14006_ (.B2(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .C1(_09574_),
    .B1(net5150),
    .A1(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .Y(_09575_),
    .A2(net5343));
 sg13g2_nand3_1 _14007_ (.B(_09572_),
    .C(_09575_),
    .A(_09571_),
    .Y(_09576_));
 sg13g2_a21oi_1 _14008_ (.A1(_07892_),
    .A2(net5547),
    .Y(_09577_),
    .B1(net6032));
 sg13g2_a22oi_1 _14009_ (.Y(_09578_),
    .B1(_09576_),
    .B2(_09577_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[6] ));
 sg13g2_nor2_1 _14010_ (.A(net1694),
    .B(net6036),
    .Y(_09579_));
 sg13g2_a21oi_1 _14011_ (.A1(net6037),
    .A2(net4964),
    .Y(_00433_),
    .B1(_09579_));
 sg13g2_a22oi_1 _14012_ (.Y(_09580_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .A2(net5156),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[7] ));
 sg13g2_nor2_1 _14013_ (.A(_09001_),
    .B(_09003_),
    .Y(_09581_));
 sg13g2_a22oi_1 _14014_ (.Y(_09582_),
    .B1(_09581_),
    .B2(\soc_inst.cpu_core.csr_file.mip_tip ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[7] ));
 sg13g2_a22oi_1 _14015_ (.Y(_09583_),
    .B1(net5537),
    .B2(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .A2(net5543),
    .A1(\soc_inst.cpu_core.csr_file.mtime[39] ));
 sg13g2_a22oi_1 _14016_ (.Y(_09584_),
    .B1(net5348),
    .B2(\soc_inst.cpu_core.csr_file.mepc[7] ),
    .A2(_09025_),
    .A1(\soc_inst.cpu_core.csr_file.mie[7] ));
 sg13g2_nand3_1 _14017_ (.B(_09583_),
    .C(_09584_),
    .A(net5553),
    .Y(_09585_));
 sg13g2_a221oi_1 _14018_ (.B2(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .C1(_09585_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mcause[7] ),
    .Y(_09586_),
    .A2(net5342));
 sg13g2_nand3_1 _14019_ (.B(_09582_),
    .C(_09586_),
    .A(_09580_),
    .Y(_09587_));
 sg13g2_a21oi_1 _14020_ (.A1(_07891_),
    .A2(net5547),
    .Y(_09588_),
    .B1(net6033));
 sg13g2_a22oi_1 _14021_ (.Y(_09589_),
    .B1(_09587_),
    .B2(_09588_),
    .A2(_09515_),
    .A1(\soc_inst.core_mem_rdata[7] ));
 sg13g2_nor2_1 _14022_ (.A(net2185),
    .B(net6040),
    .Y(_09590_));
 sg13g2_a21oi_1 _14023_ (.A1(net6040),
    .A2(net4918),
    .Y(_00434_),
    .B1(_09590_));
 sg13g2_and2_1 _14024_ (.A(\soc_inst.core_mem_rdata[7] ),
    .B(_08988_),
    .X(_09591_));
 sg13g2_nor2_1 _14025_ (.A(net6290),
    .B(_09064_),
    .Y(_09592_));
 sg13g2_nand2b_1 _14026_ (.Y(_09593_),
    .B(net6168),
    .A_N(_09064_));
 sg13g2_nand2_2 _14027_ (.Y(_09594_),
    .A(net6045),
    .B(net6024));
 sg13g2_a21o_1 _14028_ (.A2(net5528),
    .A1(\soc_inst.core_mem_rdata[8] ),
    .B1(net5529),
    .X(_09595_));
 sg13g2_a22oi_1 _14029_ (.Y(_09596_),
    .B1(net5335),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .A2(net5155),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[8] ));
 sg13g2_a22oi_1 _14030_ (.Y(_09597_),
    .B1(net5347),
    .B2(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .A2(net5353),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[8] ));
 sg13g2_a221oi_1 _14031_ (.B2(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .C1(_09536_),
    .B1(net5149),
    .A1(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .Y(_09598_),
    .A2(net5544));
 sg13g2_nand3_1 _14032_ (.B(_09597_),
    .C(_09598_),
    .A(_09596_),
    .Y(_09599_));
 sg13g2_a221oi_1 _14033_ (.B2(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .C1(_09599_),
    .B1(net5341),
    .A1(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .Y(_09600_),
    .A2(net5540));
 sg13g2_o21ai_1 _14034_ (.B1(net6031),
    .Y(_09601_),
    .A1(\soc_inst.core_mem_addr[8] ),
    .A2(net5553));
 sg13g2_nor2_1 _14035_ (.A(_09600_),
    .B(_09601_),
    .Y(_09602_));
 sg13g2_a21oi_2 _14036_ (.B1(_09602_),
    .Y(_09603_),
    .A2(_09595_),
    .A1(net6032));
 sg13g2_nor2_1 _14037_ (.A(net1811),
    .B(net6037),
    .Y(_09604_));
 sg13g2_a21oi_1 _14038_ (.A1(net6037),
    .A2(net4779),
    .Y(_00435_),
    .B1(_09604_));
 sg13g2_a21oi_1 _14039_ (.A1(\soc_inst.core_mem_rdata[9] ),
    .A2(net5528),
    .Y(_09605_),
    .B1(_09591_));
 sg13g2_a22oi_1 _14040_ (.Y(_09606_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .A2(net5157),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[9] ));
 sg13g2_a22oi_1 _14041_ (.Y(_09607_),
    .B1(net5349),
    .B2(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[9] ));
 sg13g2_a221oi_1 _14042_ (.B2(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .C1(net5549),
    .B1(net5536),
    .A1(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .Y(_09608_),
    .A2(net5542));
 sg13g2_a22oi_1 _14043_ (.Y(_09609_),
    .B1(net5150),
    .B2(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .A2(net5343),
    .A1(\soc_inst.cpu_core.csr_file.mcause[9] ));
 sg13g2_nand4_1 _14044_ (.B(_09607_),
    .C(_09608_),
    .A(_09606_),
    .Y(_09610_),
    .D(_09609_));
 sg13g2_o21ai_1 _14045_ (.B1(_09610_),
    .Y(_09611_),
    .A1(\soc_inst.core_mem_addr[9] ),
    .A2(net5553));
 sg13g2_mux2_1 _14046_ (.A0(_09605_),
    .A1(_09611_),
    .S(net6030),
    .X(_09612_));
 sg13g2_nor2_1 _14047_ (.A(net1740),
    .B(net6042),
    .Y(_09613_));
 sg13g2_a21oi_1 _14048_ (.A1(net6042),
    .A2(net4915),
    .Y(_00436_),
    .B1(_09613_));
 sg13g2_a21oi_1 _14049_ (.A1(\soc_inst.core_mem_rdata[10] ),
    .A2(net5528),
    .Y(_09614_),
    .B1(net5529));
 sg13g2_a22oi_1 _14050_ (.Y(_09615_),
    .B1(net5347),
    .B2(\soc_inst.cpu_core.csr_file.mepc[10] ),
    .A2(net5155),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[10] ));
 sg13g2_a22oi_1 _14051_ (.Y(_09616_),
    .B1(net5334),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .A2(net5353),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[10] ));
 sg13g2_a221oi_1 _14052_ (.B2(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .C1(net5549),
    .B1(net5536),
    .A1(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .Y(_09617_),
    .A2(net5542));
 sg13g2_a22oi_1 _14053_ (.Y(_09618_),
    .B1(net5148),
    .B2(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .A2(net5343),
    .A1(\soc_inst.cpu_core.csr_file.mcause[10] ));
 sg13g2_nand4_1 _14054_ (.B(_09616_),
    .C(_09617_),
    .A(_09615_),
    .Y(_09619_),
    .D(_09618_));
 sg13g2_o21ai_1 _14055_ (.B1(_09619_),
    .Y(_09620_),
    .A1(\soc_inst.core_mem_addr[10] ),
    .A2(net5553));
 sg13g2_mux2_1 _14056_ (.A0(_09614_),
    .A1(_09620_),
    .S(net6029),
    .X(_09621_));
 sg13g2_nor2_1 _14057_ (.A(net1688),
    .B(net6043),
    .Y(_09622_));
 sg13g2_a21oi_1 _14058_ (.A1(net6043),
    .A2(net4906),
    .Y(_00437_),
    .B1(_09622_));
 sg13g2_a21o_1 _14059_ (.A2(net5528),
    .A1(\soc_inst.core_mem_rdata[11] ),
    .B1(net5529),
    .X(_09623_));
 sg13g2_a22oi_1 _14060_ (.Y(_09624_),
    .B1(_09581_),
    .B2(\soc_inst.cpu_core.csr_file.mip_eip ),
    .A2(net5334),
    .A1(\soc_inst.cpu_core.csr_file.mscratch[11] ));
 sg13g2_a22oi_1 _14061_ (.Y(_09625_),
    .B1(net5348),
    .B2(\soc_inst.cpu_core.csr_file.mepc[11] ),
    .A2(_09025_),
    .A1(\soc_inst.cpu_core.csr_file.mie[11] ));
 sg13g2_a22oi_1 _14062_ (.Y(_09626_),
    .B1(net5536),
    .B2(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .A2(net5542),
    .A1(\soc_inst.cpu_core.csr_file.mtime[43] ));
 sg13g2_a22oi_1 _14063_ (.Y(_09627_),
    .B1(net5155),
    .B2(_07790_),
    .A2(net5352),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[11] ));
 sg13g2_nand3_1 _14064_ (.B(_09626_),
    .C(_09627_),
    .A(net5553),
    .Y(_09628_));
 sg13g2_a221oi_1 _14065_ (.B2(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .C1(_09628_),
    .B1(net5148),
    .A1(\soc_inst.cpu_core.csr_file.mcause[11] ),
    .Y(_09629_),
    .A2(net5342));
 sg13g2_nand3_1 _14066_ (.B(_09625_),
    .C(_09629_),
    .A(_09624_),
    .Y(_09630_));
 sg13g2_a21oi_1 _14067_ (.A1(_07812_),
    .A2(net5547),
    .Y(_09631_),
    .B1(net6032));
 sg13g2_a22oi_1 _14068_ (.Y(_09632_),
    .B1(_09630_),
    .B2(_09631_),
    .A2(_09623_),
    .A1(net6032));
 sg13g2_nor2_1 _14069_ (.A(net1430),
    .B(net6037),
    .Y(_09633_));
 sg13g2_a21oi_1 _14070_ (.A1(net6036),
    .A2(net4777),
    .Y(_00438_),
    .B1(_09633_));
 sg13g2_a21oi_1 _14071_ (.A1(\soc_inst.core_mem_rdata[12] ),
    .A2(net5528),
    .Y(_09634_),
    .B1(net5529));
 sg13g2_a22oi_1 _14072_ (.Y(_09635_),
    .B1(net5154),
    .B2(_07789_),
    .A2(net5351),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[12] ));
 sg13g2_a22oi_1 _14073_ (.Y(_09636_),
    .B1(net5332),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .A2(net5345),
    .A1(\soc_inst.cpu_core.csr_file.mepc[12] ));
 sg13g2_a221oi_1 _14074_ (.B2(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .C1(net5549),
    .B1(net5536),
    .A1(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .Y(_09637_),
    .A2(net5542));
 sg13g2_a22oi_1 _14075_ (.Y(_09638_),
    .B1(net5147),
    .B2(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .A2(net5344),
    .A1(\soc_inst.cpu_core.csr_file.mcause[12] ));
 sg13g2_nand4_1 _14076_ (.B(_09636_),
    .C(_09637_),
    .A(_09635_),
    .Y(_09639_),
    .D(_09638_));
 sg13g2_o21ai_1 _14077_ (.B1(_09639_),
    .Y(_09640_),
    .A1(\soc_inst.core_mem_addr[12] ),
    .A2(net5551));
 sg13g2_mux2_1 _14078_ (.A0(_09634_),
    .A1(_09640_),
    .S(net6029),
    .X(_09641_));
 sg13g2_nor2_1 _14079_ (.A(net2166),
    .B(net6040),
    .Y(_09642_));
 sg13g2_a21oi_1 _14080_ (.A1(net6040),
    .A2(net4900),
    .Y(_00439_),
    .B1(_09642_));
 sg13g2_a21o_1 _14081_ (.A2(net5528),
    .A1(\soc_inst.core_mem_rdata[13] ),
    .B1(net5529),
    .X(_09643_));
 sg13g2_a22oi_1 _14082_ (.Y(_09644_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[13] ));
 sg13g2_a22oi_1 _14083_ (.Y(_09645_),
    .B1(net5345),
    .B2(\soc_inst.cpu_core.csr_file.mepc[13] ),
    .A2(net5351),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[13] ));
 sg13g2_a221oi_1 _14084_ (.B2(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .C1(net5549),
    .B1(net5536),
    .A1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .Y(_09646_),
    .A2(net5542));
 sg13g2_a22oi_1 _14085_ (.Y(_09647_),
    .B1(net5143),
    .B2(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .A2(net5338),
    .A1(\soc_inst.cpu_core.csr_file.mcause[13] ));
 sg13g2_nand4_1 _14086_ (.B(_09645_),
    .C(_09646_),
    .A(_09644_),
    .Y(_09648_),
    .D(_09647_));
 sg13g2_a21oi_1 _14087_ (.A1(_07813_),
    .A2(net5545),
    .Y(_09649_),
    .B1(net6033));
 sg13g2_a22oi_1 _14088_ (.Y(_09650_),
    .B1(_09648_),
    .B2(_09649_),
    .A2(_09643_),
    .A1(net6033));
 sg13g2_nor2_1 _14089_ (.A(net2364),
    .B(net6039),
    .Y(_09651_));
 sg13g2_a21oi_1 _14090_ (.A1(net6039),
    .A2(net4963),
    .Y(_00440_),
    .B1(_09651_));
 sg13g2_a21o_1 _14091_ (.A2(net5528),
    .A1(\soc_inst.core_mem_rdata[14] ),
    .B1(net5529),
    .X(_09652_));
 sg13g2_a22oi_1 _14092_ (.Y(_09653_),
    .B1(net5345),
    .B2(\soc_inst.cpu_core.csr_file.mepc[14] ),
    .A2(net5152),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[14] ));
 sg13g2_a22oi_1 _14093_ (.Y(_09654_),
    .B1(net5333),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .A2(net5351),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[14] ));
 sg13g2_a221oi_1 _14094_ (.B2(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .C1(net5549),
    .B1(net5536),
    .A1(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .Y(_09655_),
    .A2(net5542));
 sg13g2_a22oi_1 _14095_ (.Y(_09656_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .A2(net5339),
    .A1(\soc_inst.cpu_core.csr_file.mcause[14] ));
 sg13g2_nand4_1 _14096_ (.B(_09654_),
    .C(_09655_),
    .A(_09653_),
    .Y(_09657_),
    .D(_09656_));
 sg13g2_a21oi_1 _14097_ (.A1(_07815_),
    .A2(net5548),
    .Y(_09658_),
    .B1(net6033));
 sg13g2_a22oi_1 _14098_ (.Y(_09659_),
    .B1(_09657_),
    .B2(_09658_),
    .A2(_09652_),
    .A1(net6033));
 sg13g2_nor2_1 _14099_ (.A(net2146),
    .B(net6034),
    .Y(_09660_));
 sg13g2_a21oi_1 _14100_ (.A1(net6034),
    .A2(net4955),
    .Y(_00441_),
    .B1(_09660_));
 sg13g2_a21oi_1 _14101_ (.A1(\soc_inst.core_mem_rdata[15] ),
    .A2(net5528),
    .Y(_09661_),
    .B1(net5529));
 sg13g2_a22oi_1 _14102_ (.Y(_09662_),
    .B1(net5536),
    .B2(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .A2(net5542),
    .A1(\soc_inst.cpu_core.csr_file.mtime[47] ));
 sg13g2_nand2_1 _14103_ (.Y(_09663_),
    .A(net5550),
    .B(_09662_));
 sg13g2_a221oi_1 _14104_ (.B2(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .C1(_09663_),
    .B1(net5142),
    .A1(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .Y(_09664_),
    .A2(net5338));
 sg13g2_a22oi_1 _14105_ (.Y(_09665_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .A2(net5345),
    .A1(\soc_inst.cpu_core.csr_file.mepc[15] ));
 sg13g2_a22oi_1 _14106_ (.Y(_09666_),
    .B1(net5154),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[15] ),
    .A2(net5350),
    .A1(\soc_inst.cpu_core.csr_file.mtvec[15] ));
 sg13g2_nand3_1 _14107_ (.B(_09665_),
    .C(_09666_),
    .A(_09664_),
    .Y(_09667_));
 sg13g2_o21ai_1 _14108_ (.B1(_09667_),
    .Y(_09668_),
    .A1(\soc_inst.core_mem_addr[15] ),
    .A2(net5552));
 sg13g2_mux2_1 _14109_ (.A0(_09661_),
    .A1(_09668_),
    .S(net6029),
    .X(_09669_));
 sg13g2_nor2_1 _14110_ (.A(net1346),
    .B(net6039),
    .Y(_09670_));
 sg13g2_a21oi_1 _14111_ (.A1(net6039),
    .A2(net4898),
    .Y(_00442_),
    .B1(_09670_));
 sg13g2_nor2_2 _14112_ (.A(net6290),
    .B(net6045),
    .Y(_09671_));
 sg13g2_a21o_1 _14113_ (.A2(_09671_),
    .A1(\soc_inst.core_mem_rdata[15] ),
    .B1(net5529),
    .X(_09672_));
 sg13g2_a21oi_1 _14114_ (.A1(\soc_inst.core_mem_rdata[16] ),
    .A2(net6025),
    .Y(_09673_),
    .B1(net5330));
 sg13g2_nand2_1 _14115_ (.Y(_09674_),
    .A(\soc_inst.cpu_core.csr_file.mtvec[16] ),
    .B(net5351));
 sg13g2_a22oi_1 _14116_ (.Y(_09675_),
    .B1(net5147),
    .B2(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .A2(net5344),
    .A1(\soc_inst.cpu_core.csr_file.mcause[16] ));
 sg13g2_a22oi_1 _14117_ (.Y(_09676_),
    .B1(net5333),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .A2(net5346),
    .A1(\soc_inst.cpu_core.csr_file.mepc[16] ));
 sg13g2_a221oi_1 _14118_ (.B2(\soc_inst.cpu_core.csr_file.mstatus[16] ),
    .C1(net5545),
    .B1(net5152),
    .A1(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .Y(_09677_),
    .A2(net5539));
 sg13g2_nand4_1 _14119_ (.B(_09675_),
    .C(_09676_),
    .A(_09674_),
    .Y(_09678_),
    .D(_09677_));
 sg13g2_o21ai_1 _14120_ (.B1(_09678_),
    .Y(_09679_),
    .A1(\soc_inst.core_mem_addr[16] ),
    .A2(net5551));
 sg13g2_mux2_1 _14121_ (.A0(_09673_),
    .A1(_09679_),
    .S(net6031),
    .X(_09680_));
 sg13g2_nor2_1 _14122_ (.A(net2266),
    .B(net6039),
    .Y(_09681_));
 sg13g2_a21oi_1 _14123_ (.A1(net6039),
    .A2(net4892),
    .Y(_00443_),
    .B1(_09681_));
 sg13g2_a21oi_1 _14124_ (.A1(\soc_inst.core_mem_rdata[17] ),
    .A2(net6025),
    .Y(_09682_),
    .B1(net5330));
 sg13g2_and2_1 _14125_ (.A(\soc_inst.cpu_core.csr_file.mtvec[17] ),
    .B(net5351),
    .X(_09683_));
 sg13g2_a221oi_1 _14126_ (.B2(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .C1(_09683_),
    .B1(net5346),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .Y(_09684_),
    .A2(net5154));
 sg13g2_a221oi_1 _14127_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .C1(net5545),
    .B1(net5331),
    .A1(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .Y(_09685_),
    .A2(net5538));
 sg13g2_a22oi_1 _14128_ (.Y(_09686_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .A2(net5340),
    .A1(\soc_inst.cpu_core.csr_file.mcause[17] ));
 sg13g2_nand3_1 _14129_ (.B(_09685_),
    .C(_09686_),
    .A(_09684_),
    .Y(_09687_));
 sg13g2_o21ai_1 _14130_ (.B1(_09687_),
    .Y(_09688_),
    .A1(\soc_inst.core_mem_addr[17] ),
    .A2(net5550));
 sg13g2_mux2_1 _14131_ (.A0(_09682_),
    .A1(_09688_),
    .S(net6029),
    .X(_09689_));
 sg13g2_nor2_1 _14132_ (.A(net1616),
    .B(net6035),
    .Y(_09690_));
 sg13g2_a21oi_1 _14133_ (.A1(net6035),
    .A2(net4888),
    .Y(_00444_),
    .B1(_09690_));
 sg13g2_a21oi_1 _14134_ (.A1(\soc_inst.core_mem_rdata[18] ),
    .A2(net6025),
    .Y(_09691_),
    .B1(net5330));
 sg13g2_nor2_1 _14135_ (.A(_08018_),
    .B(_09058_),
    .Y(_09692_));
 sg13g2_a221oi_1 _14136_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .C1(_09692_),
    .B1(net5333),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[18] ),
    .Y(_09693_),
    .A2(net5154));
 sg13g2_a221oi_1 _14137_ (.B2(\soc_inst.cpu_core.csr_file.mtvec[18] ),
    .C1(net5545),
    .B1(net5350),
    .A1(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .Y(_09694_),
    .A2(net5538));
 sg13g2_a22oi_1 _14138_ (.Y(_09695_),
    .B1(net5147),
    .B2(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .A2(net5344),
    .A1(\soc_inst.cpu_core.csr_file.mcause[18] ));
 sg13g2_nand3_1 _14139_ (.B(_09694_),
    .C(_09695_),
    .A(_09693_),
    .Y(_09696_));
 sg13g2_o21ai_1 _14140_ (.B1(_09696_),
    .Y(_09697_),
    .A1(\soc_inst.core_mem_addr[18] ),
    .A2(net5552));
 sg13g2_mux2_1 _14141_ (.A0(_09691_),
    .A1(_09697_),
    .S(net6029),
    .X(_09698_));
 sg13g2_nor2_1 _14142_ (.A(net1816),
    .B(net6039),
    .Y(_09699_));
 sg13g2_a21oi_1 _14143_ (.A1(net6039),
    .A2(net4769),
    .Y(_00445_),
    .B1(_09699_));
 sg13g2_a21oi_1 _14144_ (.A1(\soc_inst.core_mem_rdata[19] ),
    .A2(net6025),
    .Y(_09700_),
    .B1(net5330));
 sg13g2_and2_1 _14145_ (.A(\soc_inst.cpu_core.csr_file.mtvec[19] ),
    .B(net5351),
    .X(_09701_));
 sg13g2_a22oi_1 _14146_ (.Y(_09702_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .A2(net5338),
    .A1(\soc_inst.cpu_core.csr_file.mcause[19] ));
 sg13g2_a221oi_1 _14147_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .C1(_09701_),
    .B1(net5333),
    .A1(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .Y(_09703_),
    .A2(net5346));
 sg13g2_a22oi_1 _14148_ (.Y(_09704_),
    .B1(net5151),
    .B2(\soc_inst.cpu_core.csr_file.mstatus[19] ),
    .A2(net5538),
    .A1(\soc_inst.cpu_core.csr_file.mtime[19] ));
 sg13g2_nand4_1 _14149_ (.B(_09702_),
    .C(_09703_),
    .A(net5550),
    .Y(_09705_),
    .D(_09704_));
 sg13g2_o21ai_1 _14150_ (.B1(_09705_),
    .Y(_09706_),
    .A1(\soc_inst.core_mem_addr[19] ),
    .A2(net5550));
 sg13g2_mux2_1 _14151_ (.A0(_09700_),
    .A1(_09706_),
    .S(net6029),
    .X(_09707_));
 sg13g2_nor2_1 _14152_ (.A(net2352),
    .B(net6041),
    .Y(_09708_));
 sg13g2_a21oi_1 _14153_ (.A1(net6041),
    .A2(net4881),
    .Y(_00446_),
    .B1(_09708_));
 sg13g2_a21oi_1 _14154_ (.A1(\soc_inst.core_mem_rdata[20] ),
    .A2(net6027),
    .Y(_09709_),
    .B1(net5329));
 sg13g2_and2_1 _14155_ (.A(\soc_inst.cpu_core.csr_file.mtvec[20] ),
    .B(net5351),
    .X(_09710_));
 sg13g2_a221oi_1 _14156_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[20] ),
    .C1(_09710_),
    .B1(net5333),
    .A1(\soc_inst.cpu_core.csr_file.mepc[20] ),
    .Y(_09711_),
    .A2(net5346));
 sg13g2_a221oi_1 _14157_ (.B2(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .C1(net5545),
    .B1(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .Y(_09712_),
    .A2(net5538));
 sg13g2_a22oi_1 _14158_ (.Y(_09713_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .A2(net5338),
    .A1(\soc_inst.cpu_core.csr_file.mcause[20] ));
 sg13g2_nand3_1 _14159_ (.B(_09712_),
    .C(_09713_),
    .A(_09711_),
    .Y(_09714_));
 sg13g2_o21ai_1 _14160_ (.B1(_09714_),
    .Y(_09715_),
    .A1(\soc_inst.core_mem_addr[20] ),
    .A2(net5551));
 sg13g2_mux2_1 _14161_ (.A0(_09709_),
    .A1(_09715_),
    .S(net6031),
    .X(_09716_));
 sg13g2_nor2_1 _14162_ (.A(net2196),
    .B(net6043),
    .Y(_09717_));
 sg13g2_a21oi_1 _14163_ (.A1(net6043),
    .A2(net4876),
    .Y(_00447_),
    .B1(_09717_));
 sg13g2_a21oi_1 _14164_ (.A1(\soc_inst.core_mem_rdata[21] ),
    .A2(net6027),
    .Y(_09718_),
    .B1(net5329));
 sg13g2_nor2_1 _14165_ (.A(_08021_),
    .B(_09058_),
    .Y(_09719_));
 sg13g2_a221oi_1 _14166_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .C1(_09719_),
    .B1(net5332),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[21] ),
    .Y(_09720_),
    .A2(net5152));
 sg13g2_a221oi_1 _14167_ (.B2(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .C1(net5545),
    .B1(net5350),
    .A1(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .Y(_09721_),
    .A2(net5539));
 sg13g2_a22oi_1 _14168_ (.Y(_09722_),
    .B1(net5147),
    .B2(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .A2(net5344),
    .A1(\soc_inst.cpu_core.csr_file.mcause[21] ));
 sg13g2_nand3_1 _14169_ (.B(_09721_),
    .C(_09722_),
    .A(_09720_),
    .Y(_09723_));
 sg13g2_o21ai_1 _14170_ (.B1(_09723_),
    .Y(_09724_),
    .A1(\soc_inst.core_mem_addr[21] ),
    .A2(net5551));
 sg13g2_mux2_1 _14171_ (.A0(_09718_),
    .A1(_09724_),
    .S(net6030),
    .X(_09725_));
 sg13g2_nor2_1 _14172_ (.A(net1297),
    .B(net6042),
    .Y(_09726_));
 sg13g2_a21oi_1 _14173_ (.A1(net6042),
    .A2(net4765),
    .Y(_00448_),
    .B1(_09726_));
 sg13g2_a21oi_1 _14174_ (.A1(\soc_inst.core_mem_rdata[22] ),
    .A2(net6025),
    .Y(_09727_),
    .B1(net5330));
 sg13g2_nand2_1 _14175_ (.Y(_09728_),
    .A(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .B(net5345));
 sg13g2_a22oi_1 _14176_ (.Y(_09729_),
    .B1(net5332),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .A2(net5152),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[22] ));
 sg13g2_a221oi_1 _14177_ (.B2(\soc_inst.cpu_core.csr_file.mtvec[22] ),
    .C1(net5545),
    .B1(net5350),
    .A1(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .Y(_09730_),
    .A2(net5539));
 sg13g2_a22oi_1 _14178_ (.Y(_09731_),
    .B1(net5144),
    .B2(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .A2(net5340),
    .A1(\soc_inst.cpu_core.csr_file.mcause[22] ));
 sg13g2_nand4_1 _14179_ (.B(_09729_),
    .C(_09730_),
    .A(_09728_),
    .Y(_09732_),
    .D(_09731_));
 sg13g2_o21ai_1 _14180_ (.B1(_09732_),
    .Y(_09733_),
    .A1(\soc_inst.core_mem_addr[22] ),
    .A2(net5550));
 sg13g2_mux2_1 _14181_ (.A0(_09727_),
    .A1(_09733_),
    .S(net6029),
    .X(_09734_));
 sg13g2_nor2_1 _14182_ (.A(net1478),
    .B(net6034),
    .Y(_09735_));
 sg13g2_a21oi_1 _14183_ (.A1(net6034),
    .A2(net4867),
    .Y(_00449_),
    .B1(_09735_));
 sg13g2_a21oi_1 _14184_ (.A1(\soc_inst.core_mem_rdata[23] ),
    .A2(net6027),
    .Y(_09736_),
    .B1(net5329));
 sg13g2_and2_1 _14185_ (.A(\soc_inst.cpu_core.csr_file.mtvec[23] ),
    .B(net5350),
    .X(_09737_));
 sg13g2_a221oi_1 _14186_ (.B2(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .C1(_09737_),
    .B1(net5333),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[23] ),
    .Y(_09738_),
    .A2(net5154));
 sg13g2_a22oi_1 _14187_ (.Y(_09739_),
    .B1(net5340),
    .B2(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .A2(net5539),
    .A1(\soc_inst.cpu_core.csr_file.mtime[23] ));
 sg13g2_a221oi_1 _14188_ (.B2(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .C1(net5545),
    .B1(net5144),
    .A1(\soc_inst.cpu_core.csr_file.mepc[23] ),
    .Y(_09740_),
    .A2(net5345));
 sg13g2_nand3_1 _14189_ (.B(_09739_),
    .C(_09740_),
    .A(_09738_),
    .Y(_09741_));
 sg13g2_o21ai_1 _14190_ (.B1(_09741_),
    .Y(_09742_),
    .A1(\soc_inst.core_mem_addr[23] ),
    .A2(net5551));
 sg13g2_mux2_1 _14191_ (.A0(_09736_),
    .A1(_09742_),
    .S(net6030),
    .X(_09743_));
 sg13g2_nor2_1 _14192_ (.A(net2448),
    .B(net6043),
    .Y(_09744_));
 sg13g2_a21oi_1 _14193_ (.A1(net6043),
    .A2(net4863),
    .Y(_00450_),
    .B1(_09744_));
 sg13g2_a21oi_1 _14194_ (.A1(\soc_inst.core_mem_rdata[24] ),
    .A2(net6027),
    .Y(_09745_),
    .B1(net5329));
 sg13g2_nand2_1 _14195_ (.Y(_09746_),
    .A(\soc_inst.cpu_core.csr_file.mcause[24] ),
    .B(net5338));
 sg13g2_a22oi_1 _14196_ (.Y(_09747_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[24] ));
 sg13g2_a22oi_1 _14197_ (.Y(_09748_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .A2(net5538),
    .A1(\soc_inst.cpu_core.csr_file.mtime[24] ));
 sg13g2_nand4_1 _14198_ (.B(_09746_),
    .C(_09747_),
    .A(net5550),
    .Y(_09749_),
    .D(_09748_));
 sg13g2_o21ai_1 _14199_ (.B1(_09749_),
    .Y(_09750_),
    .A1(\soc_inst.core_mem_addr[24] ),
    .A2(net5554));
 sg13g2_mux2_1 _14200_ (.A0(_09745_),
    .A1(_09750_),
    .S(net6030),
    .X(_09751_));
 sg13g2_nor2_1 _14201_ (.A(net1583),
    .B(net6035),
    .Y(_09752_));
 sg13g2_a21oi_1 _14202_ (.A1(net6035),
    .A2(net4858),
    .Y(_00451_),
    .B1(_09752_));
 sg13g2_a21oi_1 _14203_ (.A1(\soc_inst.core_mem_rdata[25] ),
    .A2(net6025),
    .Y(_09753_),
    .B1(net5330));
 sg13g2_nand2_1 _14204_ (.Y(_09754_),
    .A(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .B(net5145));
 sg13g2_a22oi_1 _14205_ (.Y(_09755_),
    .B1(net5332),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[25] ),
    .A2(net5153),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[25] ));
 sg13g2_a22oi_1 _14206_ (.Y(_09756_),
    .B1(net5339),
    .B2(\soc_inst.cpu_core.csr_file.mcause[25] ),
    .A2(net5541),
    .A1(\soc_inst.cpu_core.csr_file.mtime[25] ));
 sg13g2_nand4_1 _14207_ (.B(_09754_),
    .C(_09755_),
    .A(net5552),
    .Y(_09757_),
    .D(_09756_));
 sg13g2_o21ai_1 _14208_ (.B1(_09757_),
    .Y(_09758_),
    .A1(\soc_inst.core_mem_addr[25] ),
    .A2(net5554));
 sg13g2_mux2_1 _14209_ (.A0(_09753_),
    .A1(_09758_),
    .S(net6029),
    .X(_09759_));
 sg13g2_nor2_1 _14210_ (.A(net1751),
    .B(net6034),
    .Y(_09760_));
 sg13g2_a21oi_1 _14211_ (.A1(net6034),
    .A2(net4852),
    .Y(_00452_),
    .B1(_09760_));
 sg13g2_a21oi_1 _14212_ (.A1(\soc_inst.core_mem_rdata[26] ),
    .A2(net6027),
    .Y(_09761_),
    .B1(net5329));
 sg13g2_nand2_1 _14213_ (.Y(_09762_),
    .A(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .B(net5338));
 sg13g2_a22oi_1 _14214_ (.Y(_09763_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[26] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[26] ));
 sg13g2_a22oi_1 _14215_ (.Y(_09764_),
    .B1(net5142),
    .B2(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .A2(net5538),
    .A1(\soc_inst.cpu_core.csr_file.mtime[26] ));
 sg13g2_nand4_1 _14216_ (.B(_09762_),
    .C(_09763_),
    .A(net5550),
    .Y(_09765_),
    .D(_09764_));
 sg13g2_o21ai_1 _14217_ (.B1(_09765_),
    .Y(_09766_),
    .A1(\soc_inst.core_mem_addr[26] ),
    .A2(net5554));
 sg13g2_mux2_1 _14218_ (.A0(_09761_),
    .A1(_09766_),
    .S(net6030),
    .X(_09767_));
 sg13g2_nor2_1 _14219_ (.A(net2233),
    .B(net6041),
    .Y(_09768_));
 sg13g2_a21oi_1 _14220_ (.A1(net6041),
    .A2(net4847),
    .Y(_00453_),
    .B1(_09768_));
 sg13g2_a21oi_1 _14221_ (.A1(\soc_inst.core_mem_rdata[27] ),
    .A2(net6027),
    .Y(_09769_),
    .B1(net5329));
 sg13g2_nand2_1 _14222_ (.Y(_09770_),
    .A(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .B(net5145));
 sg13g2_a22oi_1 _14223_ (.Y(_09771_),
    .B1(net5332),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .A2(net5153),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[27] ));
 sg13g2_a22oi_1 _14224_ (.Y(_09772_),
    .B1(net5339),
    .B2(\soc_inst.cpu_core.csr_file.mcause[27] ),
    .A2(net5541),
    .A1(\soc_inst.cpu_core.csr_file.mtime[27] ));
 sg13g2_nand4_1 _14225_ (.B(_09770_),
    .C(_09771_),
    .A(net5550),
    .Y(_09773_),
    .D(_09772_));
 sg13g2_o21ai_1 _14226_ (.B1(_09773_),
    .Y(_09774_),
    .A1(\soc_inst.core_mem_addr[27] ),
    .A2(net5554));
 sg13g2_mux2_1 _14227_ (.A0(_09769_),
    .A1(_09774_),
    .S(net6030),
    .X(_09775_));
 sg13g2_nor2_1 _14228_ (.A(net1939),
    .B(net6034),
    .Y(_09776_));
 sg13g2_a21oi_1 _14229_ (.A1(net6034),
    .A2(net4844),
    .Y(_00454_),
    .B1(_09776_));
 sg13g2_a21oi_1 _14230_ (.A1(\soc_inst.core_mem_rdata[28] ),
    .A2(net6027),
    .Y(_09777_),
    .B1(_09672_));
 sg13g2_nand2_1 _14231_ (.Y(_09778_),
    .A(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .B(net5144));
 sg13g2_a22oi_1 _14232_ (.Y(_09779_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[28] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[28] ));
 sg13g2_a22oi_1 _14233_ (.Y(_09780_),
    .B1(net5338),
    .B2(\soc_inst.cpu_core.csr_file.mcause[28] ),
    .A2(net5539),
    .A1(\soc_inst.cpu_core.csr_file.mtime[28] ));
 sg13g2_nand4_1 _14234_ (.B(_09778_),
    .C(_09779_),
    .A(net5551),
    .Y(_09781_),
    .D(_09780_));
 sg13g2_o21ai_1 _14235_ (.B1(_09781_),
    .Y(_09782_),
    .A1(\soc_inst.core_mem_addr[28] ),
    .A2(net5553));
 sg13g2_mux2_1 _14236_ (.A0(_09777_),
    .A1(_09782_),
    .S(net6031),
    .X(_09783_));
 sg13g2_nor2_1 _14237_ (.A(net1961),
    .B(net6041),
    .Y(_09784_));
 sg13g2_a21oi_1 _14238_ (.A1(net6041),
    .A2(net4840),
    .Y(_00455_),
    .B1(_09784_));
 sg13g2_a21oi_1 _14239_ (.A1(\soc_inst.core_mem_rdata[29] ),
    .A2(net6028),
    .Y(_09785_),
    .B1(net5330));
 sg13g2_nand2_1 _14240_ (.Y(_09786_),
    .A(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .B(net5143));
 sg13g2_a22oi_1 _14241_ (.Y(_09787_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[29] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[29] ));
 sg13g2_a22oi_1 _14242_ (.Y(_09788_),
    .B1(net5338),
    .B2(\soc_inst.cpu_core.csr_file.mcause[29] ),
    .A2(net5538),
    .A1(\soc_inst.cpu_core.csr_file.mtime[29] ));
 sg13g2_nand4_1 _14243_ (.B(_09786_),
    .C(_09787_),
    .A(net5551),
    .Y(_09789_),
    .D(_09788_));
 sg13g2_o21ai_1 _14244_ (.B1(_09789_),
    .Y(_09790_),
    .A1(\soc_inst.core_mem_addr[29] ),
    .A2(net5553));
 sg13g2_mux2_1 _14245_ (.A0(_09785_),
    .A1(_09790_),
    .S(net6030),
    .X(_09791_));
 sg13g2_nor2_1 _14246_ (.A(net2125),
    .B(net6035),
    .Y(_09792_));
 sg13g2_a21oi_1 _14247_ (.A1(net6035),
    .A2(net4833),
    .Y(_00456_),
    .B1(_09792_));
 sg13g2_a21oi_1 _14248_ (.A1(\soc_inst.core_mem_rdata[30] ),
    .A2(net6027),
    .Y(_09793_),
    .B1(net5329));
 sg13g2_a22oi_1 _14249_ (.Y(_09794_),
    .B1(net5331),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .A2(net5151),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[30] ));
 sg13g2_a21oi_1 _14250_ (.A1(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .A2(net5538),
    .Y(_09795_),
    .B1(_09536_));
 sg13g2_a22oi_1 _14251_ (.Y(_09796_),
    .B1(net5143),
    .B2(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .A2(net5340),
    .A1(\soc_inst.cpu_core.csr_file.mcause[30] ));
 sg13g2_nand3_1 _14252_ (.B(_09795_),
    .C(_09796_),
    .A(_09794_),
    .Y(_09797_));
 sg13g2_o21ai_1 _14253_ (.B1(_09797_),
    .Y(_09798_),
    .A1(\soc_inst.core_mem_addr[30] ),
    .A2(net5554));
 sg13g2_mux2_1 _14254_ (.A0(_09793_),
    .A1(_09798_),
    .S(net6030),
    .X(_09799_));
 sg13g2_nor2_1 _14255_ (.A(net2109),
    .B(net6043),
    .Y(_09800_));
 sg13g2_a21oi_1 _14256_ (.A1(net6043),
    .A2(net4829),
    .Y(_00457_),
    .B1(_09800_));
 sg13g2_a21oi_1 _14257_ (.A1(\soc_inst.core_mem_rdata[31] ),
    .A2(net6028),
    .Y(_09801_),
    .B1(net5329));
 sg13g2_nand2_1 _14258_ (.Y(_09802_),
    .A(net3070),
    .B(net5341));
 sg13g2_a22oi_1 _14259_ (.Y(_09803_),
    .B1(net5332),
    .B2(\soc_inst.cpu_core.csr_file.mscratch[31] ),
    .A2(net5156),
    .A1(\soc_inst.cpu_core.csr_file.mstatus[31] ));
 sg13g2_a22oi_1 _14260_ (.Y(_09804_),
    .B1(net5145),
    .B2(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .A2(net5540),
    .A1(\soc_inst.cpu_core.csr_file.mtime[31] ));
 sg13g2_nand4_1 _14261_ (.B(_09802_),
    .C(_09803_),
    .A(net5552),
    .Y(_09805_),
    .D(_09804_));
 sg13g2_o21ai_1 _14262_ (.B1(_09805_),
    .Y(_09806_),
    .A1(\soc_inst.core_mem_addr[31] ),
    .A2(net5555));
 sg13g2_mux2_1 _14263_ (.A0(_09801_),
    .A1(_09806_),
    .S(net6031),
    .X(_09807_));
 sg13g2_nor2_1 _14264_ (.A(net1484),
    .B(net6042),
    .Y(_09808_));
 sg13g2_a21oi_1 _14265_ (.A1(net6042),
    .A2(net4826),
    .Y(_00458_),
    .B1(_09808_));
 sg13g2_nand3_1 _14266_ (.B(_09426_),
    .C(_09441_),
    .A(net6204),
    .Y(_09809_));
 sg13g2_nand2_1 _14267_ (.Y(_09810_),
    .A(net814),
    .B(_09809_));
 sg13g2_o21ai_1 _14268_ (.B1(_09810_),
    .Y(_00459_),
    .A1(_07785_),
    .A2(_09809_));
 sg13g2_nand3_1 _14269_ (.B(net5362),
    .C(_09441_),
    .A(net6204),
    .Y(_09811_));
 sg13g2_nand2_1 _14270_ (.Y(_09812_),
    .A(net445),
    .B(net5070));
 sg13g2_o21ai_1 _14271_ (.B1(_09812_),
    .Y(_00460_),
    .A1(_07785_),
    .A2(net5069));
 sg13g2_mux2_1 _14272_ (.A0(net6468),
    .A1(net2297),
    .S(net5069),
    .X(_00461_));
 sg13g2_mux2_1 _14273_ (.A0(net6466),
    .A1(net1987),
    .S(net5070),
    .X(_00462_));
 sg13g2_nor2_1 _14274_ (.A(net6464),
    .B(net5069),
    .Y(_09813_));
 sg13g2_a21oi_1 _14275_ (.A1(_07956_),
    .A2(net5069),
    .Y(_00463_),
    .B1(_09813_));
 sg13g2_nor2_1 _14276_ (.A(net6462),
    .B(net5069),
    .Y(_09814_));
 sg13g2_a21oi_1 _14277_ (.A1(_07958_),
    .A2(net5069),
    .Y(_00464_),
    .B1(_09814_));
 sg13g2_nor2_1 _14278_ (.A(net6460),
    .B(net5069),
    .Y(_09815_));
 sg13g2_a21oi_1 _14279_ (.A1(_07960_),
    .A2(net5069),
    .Y(_00465_),
    .B1(_09815_));
 sg13g2_nor2_1 _14280_ (.A(net6457),
    .B(net5070),
    .Y(_09816_));
 sg13g2_a21oi_1 _14281_ (.A1(_07961_),
    .A2(net5070),
    .Y(_00466_),
    .B1(_09816_));
 sg13g2_and3_2 _14282_ (.X(_09817_),
    .A(net6205),
    .B(net5566),
    .C(_09441_));
 sg13g2_mux2_1 _14283_ (.A0(net2783),
    .A1(net6471),
    .S(_09817_),
    .X(_00467_));
 sg13g2_nor2_1 _14284_ (.A(net2466),
    .B(_09817_),
    .Y(_09818_));
 sg13g2_a21oi_1 _14285_ (.A1(_07784_),
    .A2(_09817_),
    .Y(_00468_),
    .B1(_09818_));
 sg13g2_mux2_1 _14286_ (.A0(net2898),
    .A1(net6466),
    .S(_09817_),
    .X(_00469_));
 sg13g2_mux2_1 _14287_ (.A0(net2782),
    .A1(net6464),
    .S(_09817_),
    .X(_00470_));
 sg13g2_mux2_1 _14288_ (.A0(net2536),
    .A1(net245),
    .S(_09817_),
    .X(_00471_));
 sg13g2_mux2_1 _14289_ (.A0(net2499),
    .A1(net6460),
    .S(_09817_),
    .X(_00472_));
 sg13g2_mux2_1 _14290_ (.A0(net2505),
    .A1(net6457),
    .S(_09817_),
    .X(_00473_));
 sg13g2_nor2_2 _14291_ (.A(_08250_),
    .B(_08293_),
    .Y(_09819_));
 sg13g2_nand2b_2 _14292_ (.Y(_09820_),
    .B(net3402),
    .A_N(\soc_inst.mem_ctrl.access_state[4] ));
 sg13g2_nand2_1 _14293_ (.Y(_09821_),
    .A(_09819_),
    .B(_09820_));
 sg13g2_a21oi_2 _14294_ (.B1(\soc_inst.mem_ctrl.access_state[4] ),
    .Y(_09822_),
    .A2(_08245_),
    .A1(_08244_));
 sg13g2_nand2b_2 _14295_ (.Y(_09823_),
    .B(_08246_),
    .A_N(net2751));
 sg13g2_nor3_1 _14296_ (.A(net6106),
    .B(net4820),
    .C(_09823_),
    .Y(_09824_));
 sg13g2_a21o_1 _14297_ (.A2(net4820),
    .A1(net2779),
    .B1(_09824_),
    .X(_00474_));
 sg13g2_nor3_1 _14298_ (.A(net6045),
    .B(net4820),
    .C(_09823_),
    .Y(_09825_));
 sg13g2_a21o_1 _14299_ (.A2(net4820),
    .A1(net2917),
    .B1(_09825_),
    .X(_00475_));
 sg13g2_nor3_1 _14300_ (.A(net6024),
    .B(net4820),
    .C(_09823_),
    .Y(_09826_));
 sg13g2_a21o_1 _14301_ (.A2(net4820),
    .A1(net2851),
    .B1(_09826_),
    .X(_00476_));
 sg13g2_a21oi_1 _14302_ (.A1(net6504),
    .A2(\soc_inst.mem_ctrl.spi_done ),
    .Y(_09827_),
    .B1(_07867_));
 sg13g2_a21oi_1 _14303_ (.A1(net6181),
    .A2(_08289_),
    .Y(_09828_),
    .B1(_09827_));
 sg13g2_nand2_1 _14304_ (.Y(_09829_),
    .A(_09819_),
    .B(_09828_));
 sg13g2_nand2b_2 _14305_ (.Y(_09830_),
    .B(_07866_),
    .A_N(_09820_));
 sg13g2_nor2_1 _14306_ (.A(net6179),
    .B(_09830_),
    .Y(_09831_));
 sg13g2_nor3_1 _14307_ (.A(net6194),
    .B(net6179),
    .C(_09830_),
    .Y(_09832_));
 sg13g2_nor4_1 _14308_ (.A(_08386_),
    .B(_08389_),
    .C(_09829_),
    .D(_09832_),
    .Y(_09833_));
 sg13g2_nand3_1 _14309_ (.B(_08394_),
    .C(_09833_),
    .A(_08385_),
    .Y(_09834_));
 sg13g2_a22oi_1 _14310_ (.Y(_00477_),
    .B1(_09834_),
    .B2(_07883_),
    .A2(_09833_),
    .A1(_07865_));
 sg13g2_nor2_2 _14311_ (.A(_08988_),
    .B(_09823_),
    .Y(_09835_));
 sg13g2_nor2_2 _14312_ (.A(_08987_),
    .B(_09823_),
    .Y(_09836_));
 sg13g2_a21oi_1 _14313_ (.A1(net268),
    .A2(net5328),
    .Y(_09837_),
    .B1(net4816));
 sg13g2_a21oi_1 _14314_ (.A1(_08212_),
    .A2(net4817),
    .Y(_00478_),
    .B1(_09837_));
 sg13g2_nand2_1 _14315_ (.Y(_09838_),
    .A(net233),
    .B(net5328));
 sg13g2_nand2_1 _14316_ (.Y(_09839_),
    .A(net341),
    .B(net4817));
 sg13g2_o21ai_1 _14317_ (.B1(_09839_),
    .Y(_00479_),
    .A1(net4817),
    .A2(_09838_));
 sg13g2_nand2_1 _14318_ (.Y(_09840_),
    .A(\soc_inst.core_mem_wdata[26] ),
    .B(net5328));
 sg13g2_nand2_1 _14319_ (.Y(_09841_),
    .A(net318),
    .B(net4817));
 sg13g2_o21ai_1 _14320_ (.B1(_09841_),
    .Y(_00480_),
    .A1(net4816),
    .A2(_09840_));
 sg13g2_nand2_1 _14321_ (.Y(_09842_),
    .A(net712),
    .B(net5328));
 sg13g2_nand2_1 _14322_ (.Y(_09843_),
    .A(net745),
    .B(net4816));
 sg13g2_o21ai_1 _14323_ (.B1(_09843_),
    .Y(_00481_),
    .A1(net4816),
    .A2(_09842_));
 sg13g2_nand2_1 _14324_ (.Y(_09844_),
    .A(net369),
    .B(net5327));
 sg13g2_nand2_1 _14325_ (.Y(_09845_),
    .A(net802),
    .B(net4810));
 sg13g2_o21ai_1 _14326_ (.B1(_09845_),
    .Y(_00482_),
    .A1(net4810),
    .A2(_09844_));
 sg13g2_nand2_1 _14327_ (.Y(_09846_),
    .A(net313),
    .B(net5327));
 sg13g2_nand2_1 _14328_ (.Y(_09847_),
    .A(net415),
    .B(net4810));
 sg13g2_o21ai_1 _14329_ (.B1(_09847_),
    .Y(_00483_),
    .A1(net4810),
    .A2(_09846_));
 sg13g2_nand2_1 _14330_ (.Y(_09848_),
    .A(\soc_inst.core_mem_wdata[30] ),
    .B(net5328));
 sg13g2_nand2_1 _14331_ (.Y(_09849_),
    .A(net418),
    .B(net4817));
 sg13g2_o21ai_1 _14332_ (.B1(_09849_),
    .Y(_00484_),
    .A1(net4817),
    .A2(_09848_));
 sg13g2_nand2_1 _14333_ (.Y(_09850_),
    .A(\soc_inst.core_mem_wdata[31] ),
    .B(net5327));
 sg13g2_nand2_1 _14334_ (.Y(_09851_),
    .A(net266),
    .B(net4817));
 sg13g2_o21ai_1 _14335_ (.B1(_09851_),
    .Y(_00485_),
    .A1(net4812),
    .A2(_09850_));
 sg13g2_nand2_1 _14336_ (.Y(_09852_),
    .A(net225),
    .B(net5328));
 sg13g2_nand2_1 _14337_ (.Y(_09853_),
    .A(net853),
    .B(net4815));
 sg13g2_o21ai_1 _14338_ (.B1(_09853_),
    .Y(_00486_),
    .A1(net4815),
    .A2(_09852_));
 sg13g2_nand2_1 _14339_ (.Y(_09854_),
    .A(net160),
    .B(net5328));
 sg13g2_nand2_1 _14340_ (.Y(_09855_),
    .A(net1086),
    .B(net4815));
 sg13g2_o21ai_1 _14341_ (.B1(_09855_),
    .Y(_00487_),
    .A1(net4815),
    .A2(_09854_));
 sg13g2_nand2_1 _14342_ (.Y(_09856_),
    .A(\soc_inst.core_mem_wdata[18] ),
    .B(net5327));
 sg13g2_nand2_1 _14343_ (.Y(_09857_),
    .A(net1099),
    .B(net4816));
 sg13g2_o21ai_1 _14344_ (.B1(_09857_),
    .Y(_00488_),
    .A1(net4816),
    .A2(_09856_));
 sg13g2_nand2_1 _14345_ (.Y(_09858_),
    .A(net295),
    .B(net5327));
 sg13g2_nand2_1 _14346_ (.Y(_09859_),
    .A(net841),
    .B(net4815));
 sg13g2_o21ai_1 _14347_ (.B1(_09859_),
    .Y(_00489_),
    .A1(net4815),
    .A2(_09858_));
 sg13g2_nand2_1 _14348_ (.Y(_09860_),
    .A(net548),
    .B(net5328));
 sg13g2_nand2_1 _14349_ (.Y(_09861_),
    .A(net931),
    .B(net4815));
 sg13g2_o21ai_1 _14350_ (.B1(_09861_),
    .Y(_00490_),
    .A1(net4815),
    .A2(_09860_));
 sg13g2_nand2_1 _14351_ (.Y(_09862_),
    .A(net571),
    .B(net5327));
 sg13g2_nand2_1 _14352_ (.Y(_09863_),
    .A(net590),
    .B(net4810));
 sg13g2_o21ai_1 _14353_ (.B1(_09863_),
    .Y(_00491_),
    .A1(net4810),
    .A2(_09862_));
 sg13g2_nand2_1 _14354_ (.Y(_09864_),
    .A(\soc_inst.core_mem_wdata[22] ),
    .B(net5327));
 sg13g2_nand2_1 _14355_ (.Y(_09865_),
    .A(net964),
    .B(net4811));
 sg13g2_o21ai_1 _14356_ (.B1(_09865_),
    .Y(_00492_),
    .A1(net4810),
    .A2(_09864_));
 sg13g2_nand2_1 _14357_ (.Y(_09866_),
    .A(\soc_inst.core_mem_wdata[23] ),
    .B(net5327));
 sg13g2_nand2_1 _14358_ (.Y(_09867_),
    .A(net866),
    .B(net4816));
 sg13g2_o21ai_1 _14359_ (.B1(_09867_),
    .Y(_00493_),
    .A1(net4810),
    .A2(_09866_));
 sg13g2_a21oi_1 _14360_ (.A1(net6454),
    .A2(_09835_),
    .Y(_09868_),
    .B1(net4813));
 sg13g2_a21oi_1 _14361_ (.A1(_08213_),
    .A2(net4812),
    .Y(_00494_),
    .B1(_09868_));
 sg13g2_a21oi_1 _14362_ (.A1(net6453),
    .A2(_09835_),
    .Y(_09869_),
    .B1(net4813));
 sg13g2_a21oi_1 _14363_ (.A1(_08214_),
    .A2(net4813),
    .Y(_00495_),
    .B1(_09869_));
 sg13g2_a21oi_1 _14364_ (.A1(\soc_inst.core_mem_wdata[10] ),
    .A2(_09835_),
    .Y(_09870_),
    .B1(net4813));
 sg13g2_a21oi_1 _14365_ (.A1(_08215_),
    .A2(net4812),
    .Y(_00496_),
    .B1(_09870_));
 sg13g2_a21oi_1 _14366_ (.A1(\soc_inst.core_mem_wdata[11] ),
    .A2(_09835_),
    .Y(_09871_),
    .B1(net4812));
 sg13g2_a21oi_1 _14367_ (.A1(_08216_),
    .A2(net4812),
    .Y(_00497_),
    .B1(_09871_));
 sg13g2_a21oi_1 _14368_ (.A1(\soc_inst.core_mem_wdata[12] ),
    .A2(_09835_),
    .Y(_09872_),
    .B1(net4811));
 sg13g2_a21oi_1 _14369_ (.A1(_08217_),
    .A2(net4812),
    .Y(_00498_),
    .B1(_09872_));
 sg13g2_a21oi_1 _14370_ (.A1(\soc_inst.core_mem_wdata[13] ),
    .A2(_09835_),
    .Y(_09873_),
    .B1(net4811));
 sg13g2_a21oi_1 _14371_ (.A1(_08218_),
    .A2(net4814),
    .Y(_00499_),
    .B1(_09873_));
 sg13g2_a21oi_1 _14372_ (.A1(\soc_inst.core_mem_wdata[14] ),
    .A2(_09835_),
    .Y(_09874_),
    .B1(net4811));
 sg13g2_a21oi_1 _14373_ (.A1(_08219_),
    .A2(net4814),
    .Y(_00500_),
    .B1(_09874_));
 sg13g2_a21oi_1 _14374_ (.A1(\soc_inst.core_mem_wdata[15] ),
    .A2(_09835_),
    .Y(_09875_),
    .B1(net4812));
 sg13g2_a21oi_1 _14375_ (.A1(_08220_),
    .A2(net4812),
    .Y(_00501_),
    .B1(_09875_));
 sg13g2_nand2_1 _14376_ (.Y(_09876_),
    .A(net6471),
    .B(_09822_));
 sg13g2_nand2_1 _14377_ (.Y(_09877_),
    .A(net305),
    .B(net4818));
 sg13g2_o21ai_1 _14378_ (.B1(_09877_),
    .Y(_00502_),
    .A1(net4818),
    .A2(_09876_));
 sg13g2_nand2_1 _14379_ (.Y(_09878_),
    .A(net6469),
    .B(_09822_));
 sg13g2_nand2_1 _14380_ (.Y(_09879_),
    .A(net383),
    .B(net4818));
 sg13g2_o21ai_1 _14381_ (.B1(_09879_),
    .Y(_00503_),
    .A1(net4819),
    .A2(_09878_));
 sg13g2_nand2_1 _14382_ (.Y(_09880_),
    .A(net6467),
    .B(_09822_));
 sg13g2_nand2_1 _14383_ (.Y(_09881_),
    .A(net202),
    .B(net4821));
 sg13g2_o21ai_1 _14384_ (.B1(_09881_),
    .Y(_00504_),
    .A1(net4820),
    .A2(_09880_));
 sg13g2_nand2_1 _14385_ (.Y(_09882_),
    .A(net6464),
    .B(_09822_));
 sg13g2_nand2_1 _14386_ (.Y(_09883_),
    .A(net332),
    .B(net4819));
 sg13g2_o21ai_1 _14387_ (.B1(_09883_),
    .Y(_00505_),
    .A1(net4818),
    .A2(_09882_));
 sg13g2_nand2_1 _14388_ (.Y(_09884_),
    .A(net6462),
    .B(_09822_));
 sg13g2_nand2_1 _14389_ (.Y(_09885_),
    .A(net356),
    .B(net4818));
 sg13g2_o21ai_1 _14390_ (.B1(_09885_),
    .Y(_00506_),
    .A1(net4818),
    .A2(_09884_));
 sg13g2_nand2_1 _14391_ (.Y(_09886_),
    .A(net6460),
    .B(_09822_));
 sg13g2_nand2_1 _14392_ (.Y(_09887_),
    .A(net350),
    .B(net4818));
 sg13g2_o21ai_1 _14393_ (.B1(_09887_),
    .Y(_00507_),
    .A1(net4818),
    .A2(_09886_));
 sg13g2_nand2_1 _14394_ (.Y(_09888_),
    .A(net6458),
    .B(_09822_));
 sg13g2_nand2_1 _14395_ (.Y(_09889_),
    .A(net181),
    .B(net4819));
 sg13g2_o21ai_1 _14396_ (.B1(_09889_),
    .Y(_00508_),
    .A1(net4819),
    .A2(_09888_));
 sg13g2_nand2_1 _14397_ (.Y(_09890_),
    .A(net6455),
    .B(_09822_));
 sg13g2_nand2_1 _14398_ (.Y(_09891_),
    .A(net165),
    .B(net4819));
 sg13g2_o21ai_1 _14399_ (.B1(_09891_),
    .Y(_00509_),
    .A1(net4819),
    .A2(_09890_));
 sg13g2_nand2_1 _14400_ (.Y(_09892_),
    .A(net6168),
    .B(net6105));
 sg13g2_nand2_2 _14401_ (.Y(_09893_),
    .A(net6301),
    .B(net6169));
 sg13g2_inv_1 _14402_ (.Y(_09894_),
    .A(_09893_));
 sg13g2_a21oi_2 _14403_ (.B1(_09893_),
    .Y(_09895_),
    .A2(net6023),
    .A1(\soc_inst.cpu_core.mem_rs1_data[5] ));
 sg13g2_nand2_2 _14404_ (.Y(_09896_),
    .A(net4792),
    .B(_09514_));
 sg13g2_o21ai_1 _14405_ (.B1(net619),
    .Y(_09897_),
    .A1(_09895_),
    .A2(_09896_));
 sg13g2_nor2b_2 _14406_ (.A(net6293),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .Y(_09898_));
 sg13g2_nor2_2 _14407_ (.A(net6294),
    .B(_09067_),
    .Y(_09899_));
 sg13g2_nand2_1 _14408_ (.Y(_09900_),
    .A(net5534),
    .B(_09898_));
 sg13g2_o21ai_1 _14409_ (.B1(net620),
    .Y(_00510_),
    .A1(net4760),
    .A2(_09900_));
 sg13g2_a21oi_2 _14410_ (.B1(_09893_),
    .Y(_09901_),
    .A2(net6023),
    .A1(\soc_inst.cpu_core.mem_rs1_data[6] ));
 sg13g2_o21ai_1 _14411_ (.B1(net573),
    .Y(_09902_),
    .A1(net4760),
    .A2(_09901_));
 sg13g2_nor2b_1 _14412_ (.A(net6294),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .Y(_09903_));
 sg13g2_nand2_1 _14413_ (.Y(_09904_),
    .A(net5533),
    .B(_09903_));
 sg13g2_o21ai_1 _14414_ (.B1(net574),
    .Y(_00511_),
    .A1(net4760),
    .A2(_09904_));
 sg13g2_a21oi_2 _14415_ (.B1(_09893_),
    .Y(_09905_),
    .A2(net6023),
    .A1(net1413));
 sg13g2_o21ai_1 _14416_ (.B1(net440),
    .Y(_09906_),
    .A1(net4760),
    .A2(_09905_));
 sg13g2_nor2b_2 _14417_ (.A(net6293),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .Y(_09907_));
 sg13g2_nand2_1 _14418_ (.Y(_09908_),
    .A(net5534),
    .B(_09907_));
 sg13g2_o21ai_1 _14419_ (.B1(net441),
    .Y(_00512_),
    .A1(_09896_),
    .A2(_09908_));
 sg13g2_a21oi_2 _14420_ (.B1(_09893_),
    .Y(_09909_),
    .A2(net6023),
    .A1(net1456));
 sg13g2_o21ai_1 _14421_ (.B1(net785),
    .Y(_09910_),
    .A1(net4760),
    .A2(_09909_));
 sg13g2_nor2b_2 _14422_ (.A(net6294),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .Y(_09911_));
 sg13g2_nand2_1 _14423_ (.Y(_09912_),
    .A(net5534),
    .B(_09911_));
 sg13g2_o21ai_1 _14424_ (.B1(net786),
    .Y(_00513_),
    .A1(net4760),
    .A2(_09912_));
 sg13g2_a21oi_1 _14425_ (.A1(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .A2(net6024),
    .Y(_09913_),
    .B1(_09893_));
 sg13g2_o21ai_1 _14426_ (.B1(net476),
    .Y(_09914_),
    .A1(net4760),
    .A2(_09913_));
 sg13g2_nor2b_2 _14427_ (.A(net6293),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .Y(_09915_));
 sg13g2_nand2_1 _14428_ (.Y(_09916_),
    .A(net5534),
    .B(_09915_));
 sg13g2_o21ai_1 _14429_ (.B1(net477),
    .Y(_00514_),
    .A1(net4760),
    .A2(_09916_));
 sg13g2_o21ai_1 _14430_ (.B1(_09268_),
    .Y(_09917_),
    .A1(net5368),
    .A2(_09280_));
 sg13g2_nor2_1 _14431_ (.A(\soc_inst.i2c_inst.start_pending ),
    .B(_08831_),
    .Y(_09918_));
 sg13g2_o21ai_1 _14432_ (.B1(net92),
    .Y(_09919_),
    .A1(_09917_),
    .A2(_09918_));
 sg13g2_o21ai_1 _14433_ (.B1(_08831_),
    .Y(_09920_),
    .A1(_07895_),
    .A2(net241));
 sg13g2_o21ai_1 _14434_ (.B1(_09919_),
    .Y(_00515_),
    .A1(_09917_),
    .A2(_09920_));
 sg13g2_a21oi_2 _14435_ (.B1(net6105),
    .Y(_09921_),
    .A2(_08984_),
    .A1(net6290));
 sg13g2_o21ai_1 _14436_ (.B1(_09016_),
    .Y(_09922_),
    .A1(_08977_),
    .A2(net6016));
 sg13g2_nand2b_1 _14437_ (.Y(_09923_),
    .B(_09037_),
    .A_N(_09922_));
 sg13g2_nor2_2 _14438_ (.A(_09044_),
    .B(_09922_),
    .Y(_09924_));
 sg13g2_nor2_1 _14439_ (.A(net2544),
    .B(net4757),
    .Y(_09925_));
 sg13g2_nand2b_1 _14440_ (.Y(_09926_),
    .B(_09070_),
    .A_N(net2544));
 sg13g2_nor2_1 _14441_ (.A(net6301),
    .B(_09070_),
    .Y(_09927_));
 sg13g2_a21oi_1 _14442_ (.A1(_09073_),
    .A2(_09926_),
    .Y(_09928_),
    .B1(_09927_));
 sg13g2_a21oi_1 _14443_ (.A1(net4757),
    .A2(_09928_),
    .Y(_00516_),
    .B1(_09925_));
 sg13g2_nor2_1 _14444_ (.A(net2150),
    .B(net4757),
    .Y(_09929_));
 sg13g2_nand2_1 _14445_ (.Y(_09930_),
    .A(_08001_),
    .B(_09082_));
 sg13g2_nor2_1 _14446_ (.A(net6301),
    .B(_09082_),
    .Y(_09931_));
 sg13g2_a21oi_1 _14447_ (.A1(_09085_),
    .A2(_09930_),
    .Y(_09932_),
    .B1(_09931_));
 sg13g2_a21oi_1 _14448_ (.A1(net4757),
    .A2(_09932_),
    .Y(_00517_),
    .B1(_09929_));
 sg13g2_nor2_1 _14449_ (.A(net2744),
    .B(net4757),
    .Y(_09933_));
 sg13g2_nand2b_1 _14450_ (.Y(_09934_),
    .B(_09091_),
    .A_N(net2744));
 sg13g2_nor2_1 _14451_ (.A(net6302),
    .B(_09091_),
    .Y(_09935_));
 sg13g2_a21oi_1 _14452_ (.A1(_09093_),
    .A2(_09934_),
    .Y(_09936_),
    .B1(_09935_));
 sg13g2_a21oi_1 _14453_ (.A1(net4757),
    .A2(_09936_),
    .Y(_00518_),
    .B1(_09933_));
 sg13g2_a21oi_1 _14454_ (.A1(_09052_),
    .A2(net4758),
    .Y(_09937_),
    .B1(net718));
 sg13g2_a21oi_1 _14455_ (.A1(_09055_),
    .A2(net4758),
    .Y(_00519_),
    .B1(_09937_));
 sg13g2_nor2_1 _14456_ (.A(net2381),
    .B(net4757),
    .Y(_09938_));
 sg13g2_nand2b_1 _14457_ (.Y(_09939_),
    .B(_09108_),
    .A_N(net2381));
 sg13g2_nor2_1 _14458_ (.A(net6301),
    .B(_09108_),
    .Y(_09940_));
 sg13g2_a21oi_1 _14459_ (.A1(_09111_),
    .A2(_09939_),
    .Y(_09941_),
    .B1(_09940_));
 sg13g2_a21oi_1 _14460_ (.A1(net4757),
    .A2(_09941_),
    .Y(_00520_),
    .B1(_09938_));
 sg13g2_nand2_2 _14461_ (.Y(_09942_),
    .A(net5354),
    .B(net4948));
 sg13g2_nor2_1 _14462_ (.A(net6164),
    .B(net3021),
    .Y(_09943_));
 sg13g2_nor2_1 _14463_ (.A(net6475),
    .B(_09942_),
    .Y(_09944_));
 sg13g2_a21oi_2 _14464_ (.B1(net6328),
    .Y(_09945_),
    .A2(_09944_),
    .A1(_08290_));
 sg13g2_a21o_2 _14465_ (.A2(_09944_),
    .A1(_08290_),
    .B1(net6328),
    .X(_09946_));
 sg13g2_o21ai_1 _14466_ (.B1(_09945_),
    .Y(_09947_),
    .A1(_09942_),
    .A2(_09943_));
 sg13g2_a21oi_1 _14467_ (.A1(net2544),
    .A2(net4940),
    .Y(_09948_),
    .B1(net6475));
 sg13g2_nor3_1 _14468_ (.A(_09943_),
    .B(net4735),
    .C(_09948_),
    .Y(_09949_));
 sg13g2_a21o_1 _14469_ (.A2(_09947_),
    .A1(net2927),
    .B1(_09949_),
    .X(_00521_));
 sg13g2_nor2b_2 _14470_ (.A(net6533),
    .B_N(net6532),
    .Y(_09950_));
 sg13g2_nand2b_1 _14471_ (.Y(_09951_),
    .B(net6532),
    .A_N(net6533));
 sg13g2_nor4_2 _14472_ (.A(net6519),
    .B(net6525),
    .C(\soc_inst.core_instr_data[9] ),
    .Y(_09952_),
    .D(net6521));
 sg13g2_or4_1 _14473_ (.A(net6519),
    .B(net6524),
    .C(\soc_inst.core_instr_data[9] ),
    .D(net6521),
    .X(_09953_));
 sg13g2_nor4_1 _14474_ (.A(net6525),
    .B(net6523),
    .C(\soc_inst.core_instr_data[9] ),
    .D(net6520),
    .Y(_09954_));
 sg13g2_nor2_1 _14475_ (.A(net6522),
    .B(_09953_),
    .Y(_09955_));
 sg13g2_nor2_2 _14476_ (.A(net6513),
    .B(net6511),
    .Y(_09956_));
 sg13g2_and2_1 _14477_ (.A(net6509),
    .B(_09956_),
    .X(_09957_));
 sg13g2_nand2_2 _14478_ (.Y(_09958_),
    .A(net6509),
    .B(_09956_));
 sg13g2_or2_1 _14479_ (.X(_09959_),
    .B(net6527),
    .A(\soc_inst.core_instr_data[5] ));
 sg13g2_or2_1 _14480_ (.X(_09960_),
    .B(\soc_inst.core_instr_data[4] ),
    .A(\soc_inst.core_instr_data[3] ));
 sg13g2_nor3_2 _14481_ (.A(net6531),
    .B(_09959_),
    .C(_09960_),
    .Y(_09961_));
 sg13g2_nor4_2 _14482_ (.A(net6531),
    .B(net6517),
    .C(_09959_),
    .Y(_09962_),
    .D(_09960_));
 sg13g2_and3_1 _14483_ (.X(_09963_),
    .A(net6015),
    .B(net6014),
    .C(net6012));
 sg13g2_nand3_1 _14484_ (.B(net6013),
    .C(net6012),
    .A(net6015),
    .Y(_09964_));
 sg13g2_nor2b_2 _14485_ (.A(\soc_inst.core_instr_data[15] ),
    .B_N(\soc_inst.core_instr_data[14] ),
    .Y(_09965_));
 sg13g2_nor2b_2 _14486_ (.A(net6513),
    .B_N(\soc_inst.core_instr_data[14] ),
    .Y(_09966_));
 sg13g2_nor2b_2 _14487_ (.A(net6514),
    .B_N(_09965_),
    .Y(_09967_));
 sg13g2_a21oi_2 _14488_ (.B1(net6513),
    .Y(_09968_),
    .A2(_09965_),
    .A1(net6015));
 sg13g2_a21o_2 _14489_ (.A2(_09965_),
    .A1(net6015),
    .B1(net6513),
    .X(_09969_));
 sg13g2_nand2_2 _14490_ (.Y(_09970_),
    .A(_09964_),
    .B(_09968_));
 sg13g2_nor3_1 _14491_ (.A(net6093),
    .B(_09963_),
    .C(_09969_),
    .Y(_09971_));
 sg13g2_nor2b_2 _14492_ (.A(net6532),
    .B_N(net6533),
    .Y(_09972_));
 sg13g2_nand2b_2 _14493_ (.Y(_09973_),
    .B(\soc_inst.core_instr_data[0] ),
    .A_N(net6532));
 sg13g2_nand2_1 _14494_ (.Y(_09974_),
    .A(net6518),
    .B(net6013));
 sg13g2_and2_1 _14495_ (.A(net6519),
    .B(net6520),
    .X(_09975_));
 sg13g2_nand2_1 _14496_ (.Y(_09976_),
    .A(net6518),
    .B(net6520));
 sg13g2_nand2_1 _14497_ (.Y(_09977_),
    .A(net6520),
    .B(net6013));
 sg13g2_nand3_1 _14498_ (.B(net6013),
    .C(_09975_),
    .A(net6515),
    .Y(_09978_));
 sg13g2_nand2_1 _14499_ (.Y(_09979_),
    .A(net6514),
    .B(net6511));
 sg13g2_nor2_2 _14500_ (.A(net6509),
    .B(_09979_),
    .Y(_09980_));
 sg13g2_nand2_2 _14501_ (.Y(_09981_),
    .A(net6513),
    .B(_09965_));
 sg13g2_nand2_2 _14502_ (.Y(_09982_),
    .A(net6012),
    .B(_09980_));
 sg13g2_and2_1 _14503_ (.A(_09978_),
    .B(_09982_),
    .X(_09983_));
 sg13g2_nand2_2 _14504_ (.Y(_09984_),
    .A(_09978_),
    .B(_09982_));
 sg13g2_a21oi_1 _14505_ (.A1(net6091),
    .A2(_09983_),
    .Y(_09985_),
    .B1(_09971_));
 sg13g2_nor2_2 _14506_ (.A(\soc_inst.core_instr_data[1] ),
    .B(\soc_inst.core_instr_data[0] ),
    .Y(_09986_));
 sg13g2_or2_1 _14507_ (.X(_09987_),
    .B(net6533),
    .A(\soc_inst.core_instr_data[1] ));
 sg13g2_nor2_2 _14508_ (.A(net6512),
    .B(net6508),
    .Y(_09988_));
 sg13g2_nor3_2 _14509_ (.A(net6522),
    .B(net6517),
    .C(_09953_),
    .Y(_09989_));
 sg13g2_nand2b_2 _14510_ (.Y(_09990_),
    .B(_09989_),
    .A_N(_09959_));
 sg13g2_a21oi_2 _14511_ (.B1(_09966_),
    .Y(_09991_),
    .A2(_09990_),
    .A1(net6090));
 sg13g2_a21o_2 _14512_ (.A2(_09990_),
    .A1(net6090),
    .B1(_09966_),
    .X(_09992_));
 sg13g2_a221oi_1 _14513_ (.B2(_09992_),
    .C1(_09971_),
    .B1(_09986_),
    .A1(net6091),
    .Y(_09993_),
    .A2(_09983_));
 sg13g2_o21ai_1 _14514_ (.B1(_09985_),
    .Y(_09994_),
    .A1(_09987_),
    .A2(_09991_));
 sg13g2_xnor2_1 _14515_ (.Y(_09995_),
    .A(_07820_),
    .B(net5130));
 sg13g2_a21oi_1 _14516_ (.A1(net3012),
    .A2(net5361),
    .Y(_09996_),
    .B1(net4940));
 sg13g2_o21ai_1 _14517_ (.B1(_09996_),
    .Y(_09997_),
    .A1(net5361),
    .A2(_09995_));
 sg13g2_a21oi_1 _14518_ (.A1(_08001_),
    .A2(net4940),
    .Y(_09998_),
    .B1(net6475));
 sg13g2_a221oi_1 _14519_ (.B2(_09998_),
    .C1(net4735),
    .B1(_09997_),
    .A1(net6475),
    .Y(_09999_),
    .A2(net3149));
 sg13g2_a21oi_1 _14520_ (.A1(_07820_),
    .A2(net4735),
    .Y(_00522_),
    .B1(_09999_));
 sg13g2_o21ai_1 _14521_ (.B1(\soc_inst.core_instr_addr[2] ),
    .Y(_10000_),
    .A1(\soc_inst.core_instr_addr[1] ),
    .A2(net5131));
 sg13g2_inv_1 _14522_ (.Y(_10001_),
    .A(_10000_));
 sg13g2_nand3_1 _14523_ (.B(_07822_),
    .C(net5063),
    .A(_07820_),
    .Y(_10002_));
 sg13g2_a21oi_1 _14524_ (.A1(_10000_),
    .A2(_10002_),
    .Y(_10003_),
    .B1(net5361));
 sg13g2_o21ai_1 _14525_ (.B1(net4949),
    .Y(_10004_),
    .A1(net1784),
    .A2(net5354));
 sg13g2_a21oi_1 _14526_ (.A1(net2744),
    .A2(net4941),
    .Y(_10005_),
    .B1(net6475));
 sg13g2_o21ai_1 _14527_ (.B1(_10005_),
    .Y(_10006_),
    .A1(_10003_),
    .A2(_10004_));
 sg13g2_o21ai_1 _14528_ (.B1(_10006_),
    .Y(_10007_),
    .A1(net6164),
    .A2(net3246));
 sg13g2_nor2_1 _14529_ (.A(net3076),
    .B(_09945_),
    .Y(_10008_));
 sg13g2_a21oi_1 _14530_ (.A1(_09945_),
    .A2(_10007_),
    .Y(_00523_),
    .B1(_10008_));
 sg13g2_xnor2_1 _14531_ (.Y(_10009_),
    .A(_07824_),
    .B(_10000_));
 sg13g2_o21ai_1 _14532_ (.B1(net4948),
    .Y(_10010_),
    .A1(\soc_inst.cpu_core.ex_branch_target[3] ),
    .A2(net5354));
 sg13g2_a21o_1 _14533_ (.A2(_10009_),
    .A1(net5354),
    .B1(_10010_),
    .X(_10011_));
 sg13g2_a21oi_1 _14534_ (.A1(net718),
    .A2(net4940),
    .Y(_10012_),
    .B1(net6475));
 sg13g2_a21oi_1 _14535_ (.A1(_10011_),
    .A2(_10012_),
    .Y(_10013_),
    .B1(net4735));
 sg13g2_o21ai_1 _14536_ (.B1(_10013_),
    .Y(_10014_),
    .A1(net6164),
    .A2(net3245));
 sg13g2_o21ai_1 _14537_ (.B1(_10014_),
    .Y(_00524_),
    .A1(_07824_),
    .A2(_09945_));
 sg13g2_nand2_1 _14538_ (.Y(_10015_),
    .A(net2738),
    .B(net4735));
 sg13g2_nor3_2 _14539_ (.A(_07824_),
    .B(_07826_),
    .C(_10000_),
    .Y(_10016_));
 sg13g2_a21oi_1 _14540_ (.A1(\soc_inst.core_instr_addr[3] ),
    .A2(_10001_),
    .Y(_10017_),
    .B1(\soc_inst.core_instr_addr[4] ));
 sg13g2_o21ai_1 _14541_ (.B1(net5354),
    .Y(_10018_),
    .A1(_10016_),
    .A2(_10017_));
 sg13g2_a21oi_1 _14542_ (.A1(_08118_),
    .A2(net5360),
    .Y(_10019_),
    .B1(net4942));
 sg13g2_a221oi_1 _14543_ (.B2(_10019_),
    .C1(net6475),
    .B1(_10018_),
    .A1(net2381),
    .Y(_10020_),
    .A2(net4940));
 sg13g2_o21ai_1 _14544_ (.B1(_09945_),
    .Y(_10021_),
    .A1(net6164),
    .A2(net2959));
 sg13g2_o21ai_1 _14545_ (.B1(_10015_),
    .Y(_00525_),
    .A1(_10020_),
    .A2(_10021_));
 sg13g2_nand2_1 _14546_ (.Y(_10022_),
    .A(\soc_inst.core_instr_addr[5] ),
    .B(_10016_));
 sg13g2_nor2_1 _14547_ (.A(\soc_inst.core_instr_addr[5] ),
    .B(_10016_),
    .Y(_10023_));
 sg13g2_nor2_1 _14548_ (.A(net5360),
    .B(_10023_),
    .Y(_10024_));
 sg13g2_a22oi_1 _14549_ (.Y(_10025_),
    .B1(_10022_),
    .B2(_10024_),
    .A2(net5360),
    .A1(net3073));
 sg13g2_o21ai_1 _14550_ (.B1(net6163),
    .Y(_10026_),
    .A1(net776),
    .A2(net4950));
 sg13g2_a21o_1 _14551_ (.A2(_10025_),
    .A1(net4950),
    .B1(_10026_),
    .X(_10027_));
 sg13g2_a21oi_1 _14552_ (.A1(net6476),
    .A2(net2256),
    .Y(_10028_),
    .B1(net4734));
 sg13g2_a22oi_1 _14553_ (.Y(_00526_),
    .B1(_10027_),
    .B2(_10028_),
    .A2(net4734),
    .A1(_07828_));
 sg13g2_nor2_1 _14554_ (.A(_07830_),
    .B(_10022_),
    .Y(_10029_));
 sg13g2_a21oi_1 _14555_ (.A1(_07830_),
    .A2(_10022_),
    .Y(_10030_),
    .B1(net5360));
 sg13g2_nor2b_1 _14556_ (.A(_10029_),
    .B_N(_10030_),
    .Y(_10031_));
 sg13g2_a21oi_1 _14557_ (.A1(net3036),
    .A2(net5360),
    .Y(_10032_),
    .B1(_10031_));
 sg13g2_o21ai_1 _14558_ (.B1(net6163),
    .Y(_10033_),
    .A1(net715),
    .A2(net4949));
 sg13g2_a21o_1 _14559_ (.A2(_10032_),
    .A1(net4950),
    .B1(_10033_),
    .X(_10034_));
 sg13g2_a21oi_1 _14560_ (.A1(net6476),
    .A2(net1420),
    .Y(_10035_),
    .B1(net4734));
 sg13g2_a22oi_1 _14561_ (.Y(_00527_),
    .B1(_10034_),
    .B2(_10035_),
    .A2(net4734),
    .A1(_07830_));
 sg13g2_and4_1 _14562_ (.A(\soc_inst.core_instr_addr[5] ),
    .B(\soc_inst.core_instr_addr[6] ),
    .C(\soc_inst.core_instr_addr[7] ),
    .D(_10016_),
    .X(_10036_));
 sg13g2_nor2_1 _14563_ (.A(net5361),
    .B(_10036_),
    .Y(_10037_));
 sg13g2_o21ai_1 _14564_ (.B1(_10037_),
    .Y(_10038_),
    .A1(net2807),
    .A2(_10029_));
 sg13g2_a21oi_1 _14565_ (.A1(net2910),
    .A2(net5361),
    .Y(_10039_),
    .B1(net4942));
 sg13g2_o21ai_1 _14566_ (.B1(net6163),
    .Y(_10040_),
    .A1(net1193),
    .A2(net4948));
 sg13g2_a21o_1 _14567_ (.A2(_10039_),
    .A1(_10038_),
    .B1(_10040_),
    .X(_10041_));
 sg13g2_a21oi_1 _14568_ (.A1(net6476),
    .A2(net2706),
    .Y(_10042_),
    .B1(net4733));
 sg13g2_a22oi_1 _14569_ (.Y(_00528_),
    .B1(_10041_),
    .B2(_10042_),
    .A2(net4734),
    .A1(_07832_));
 sg13g2_or2_1 _14570_ (.X(_10043_),
    .B(_10036_),
    .A(\soc_inst.core_instr_addr[8] ));
 sg13g2_and2_1 _14571_ (.A(\soc_inst.core_instr_addr[8] ),
    .B(_10036_),
    .X(_10044_));
 sg13g2_nor2_1 _14572_ (.A(net5359),
    .B(_10044_),
    .Y(_10045_));
 sg13g2_a221oi_1 _14573_ (.B2(_10045_),
    .C1(net4942),
    .B1(_10043_),
    .A1(net2839),
    .Y(_10046_),
    .A2(net5359));
 sg13g2_o21ai_1 _14574_ (.B1(net6163),
    .Y(_10047_),
    .A1(net500),
    .A2(net4951));
 sg13g2_or2_1 _14575_ (.X(_10048_),
    .B(_10047_),
    .A(_10046_));
 sg13g2_a21oi_1 _14576_ (.A1(net6476),
    .A2(net1261),
    .Y(_10049_),
    .B1(net4733));
 sg13g2_a22oi_1 _14577_ (.Y(_00529_),
    .B1(_10048_),
    .B2(_10049_),
    .A2(net4733),
    .A1(_07834_));
 sg13g2_and3_2 _14578_ (.X(_10050_),
    .A(\soc_inst.core_instr_addr[8] ),
    .B(\soc_inst.core_instr_addr[9] ),
    .C(_10036_));
 sg13g2_o21ai_1 _14579_ (.B1(_08955_),
    .Y(_10051_),
    .A1(\soc_inst.core_instr_addr[9] ),
    .A2(_10044_));
 sg13g2_a21oi_1 _14580_ (.A1(net2780),
    .A2(net5359),
    .Y(_10052_),
    .B1(net4942));
 sg13g2_o21ai_1 _14581_ (.B1(_10052_),
    .Y(_10053_),
    .A1(_10050_),
    .A2(_10051_));
 sg13g2_o21ai_1 _14582_ (.B1(net6163),
    .Y(_10054_),
    .A1(net1068),
    .A2(net4950));
 sg13g2_nand2b_1 _14583_ (.Y(_10055_),
    .B(_10053_),
    .A_N(_10054_));
 sg13g2_a21oi_1 _14584_ (.A1(net6476),
    .A2(net1292),
    .Y(_10056_),
    .B1(net4733));
 sg13g2_a22oi_1 _14585_ (.Y(_00530_),
    .B1(_10055_),
    .B2(_10056_),
    .A2(net4733),
    .A1(_07836_));
 sg13g2_nand2_1 _14586_ (.Y(_10057_),
    .A(\soc_inst.core_instr_addr[10] ),
    .B(_10050_));
 sg13g2_nor2_1 _14587_ (.A(\soc_inst.core_instr_addr[10] ),
    .B(_10050_),
    .Y(_10058_));
 sg13g2_nor2_1 _14588_ (.A(net5359),
    .B(_10058_),
    .Y(_10059_));
 sg13g2_a221oi_1 _14589_ (.B2(_10059_),
    .C1(net4942),
    .B1(_10057_),
    .A1(net2721),
    .Y(_10060_),
    .A2(net5359));
 sg13g2_o21ai_1 _14590_ (.B1(net6163),
    .Y(_10061_),
    .A1(net1056),
    .A2(net4951));
 sg13g2_or2_1 _14591_ (.X(_10062_),
    .B(_10061_),
    .A(_10060_));
 sg13g2_a21oi_1 _14592_ (.A1(net6476),
    .A2(net1216),
    .Y(_10063_),
    .B1(net4733));
 sg13g2_a22oi_1 _14593_ (.Y(_00531_),
    .B1(_10062_),
    .B2(_10063_),
    .A2(net4734),
    .A1(_07838_));
 sg13g2_nand3_1 _14594_ (.B(\soc_inst.core_instr_addr[11] ),
    .C(_10050_),
    .A(\soc_inst.core_instr_addr[10] ),
    .Y(_10064_));
 sg13g2_a21oi_1 _14595_ (.A1(_07840_),
    .A2(_10057_),
    .Y(_10065_),
    .B1(net5359));
 sg13g2_a221oi_1 _14596_ (.B2(_10065_),
    .C1(net4942),
    .B1(_10064_),
    .A1(net1513),
    .Y(_10066_),
    .A2(net5359));
 sg13g2_o21ai_1 _14597_ (.B1(net6163),
    .Y(_10067_),
    .A1(net535),
    .A2(net4951));
 sg13g2_or2_1 _14598_ (.X(_10068_),
    .B(_10067_),
    .A(_10066_));
 sg13g2_a21oi_1 _14599_ (.A1(net6476),
    .A2(net3225),
    .Y(_10069_),
    .B1(net4733));
 sg13g2_a22oi_1 _14600_ (.Y(_00532_),
    .B1(_10068_),
    .B2(_10069_),
    .A2(net4733),
    .A1(_07840_));
 sg13g2_and4_1 _14601_ (.A(\soc_inst.core_instr_addr[10] ),
    .B(\soc_inst.core_instr_addr[11] ),
    .C(\soc_inst.core_instr_addr[12] ),
    .D(_10050_),
    .X(_10070_));
 sg13g2_xnor2_1 _14602_ (.Y(_10071_),
    .A(_07842_),
    .B(_10064_));
 sg13g2_a21oi_1 _14603_ (.A1(net2741),
    .A2(net5359),
    .Y(_10072_),
    .B1(_08971_));
 sg13g2_o21ai_1 _14604_ (.B1(_10072_),
    .Y(_10073_),
    .A1(net5357),
    .A2(_10071_));
 sg13g2_a21oi_1 _14605_ (.A1(_08010_),
    .A2(net4938),
    .Y(_10074_),
    .B1(net6474));
 sg13g2_a221oi_1 _14606_ (.B2(_10074_),
    .C1(net4731),
    .B1(_10073_),
    .A1(net6474),
    .Y(_10075_),
    .A2(net2077));
 sg13g2_a21oi_1 _14607_ (.A1(_07842_),
    .A2(net4731),
    .Y(_00533_),
    .B1(_10075_));
 sg13g2_and2_1 _14608_ (.A(\soc_inst.core_instr_addr[13] ),
    .B(_10070_),
    .X(_10076_));
 sg13g2_o21ai_1 _14609_ (.B1(net5354),
    .Y(_10077_),
    .A1(\soc_inst.core_instr_addr[13] ),
    .A2(_10070_));
 sg13g2_a21oi_1 _14610_ (.A1(net2446),
    .A2(net5357),
    .Y(_10078_),
    .B1(net4938));
 sg13g2_o21ai_1 _14611_ (.B1(_10078_),
    .Y(_10079_),
    .A1(_10076_),
    .A2(_10077_));
 sg13g2_a21oi_1 _14612_ (.A1(_08012_),
    .A2(net4938),
    .Y(_10080_),
    .B1(net6474));
 sg13g2_a221oi_1 _14613_ (.B2(_10080_),
    .C1(net4731),
    .B1(_10079_),
    .A1(net6474),
    .Y(_10081_),
    .A2(net2346));
 sg13g2_a21oi_1 _14614_ (.A1(_07844_),
    .A2(net4731),
    .Y(_00534_),
    .B1(_10081_));
 sg13g2_and2_1 _14615_ (.A(\soc_inst.core_instr_addr[14] ),
    .B(_10076_),
    .X(_10082_));
 sg13g2_o21ai_1 _14616_ (.B1(net5354),
    .Y(_10083_),
    .A1(\soc_inst.core_instr_addr[14] ),
    .A2(_10076_));
 sg13g2_a21oi_1 _14617_ (.A1(net2818),
    .A2(net5357),
    .Y(_10084_),
    .B1(net4938));
 sg13g2_o21ai_1 _14618_ (.B1(_10084_),
    .Y(_10085_),
    .A1(_10082_),
    .A2(_10083_));
 sg13g2_a21oi_1 _14619_ (.A1(_08014_),
    .A2(net4937),
    .Y(_10086_),
    .B1(net6474));
 sg13g2_a221oi_1 _14620_ (.B2(_10086_),
    .C1(net4730),
    .B1(_10085_),
    .A1(net6474),
    .Y(_10087_),
    .A2(net2510));
 sg13g2_a21oi_1 _14621_ (.A1(_07846_),
    .A2(net4731),
    .Y(_00535_),
    .B1(_10087_));
 sg13g2_and4_1 _14622_ (.A(\soc_inst.core_instr_addr[13] ),
    .B(\soc_inst.core_instr_addr[14] ),
    .C(\soc_inst.core_instr_addr[15] ),
    .D(_10070_),
    .X(_10088_));
 sg13g2_nor2_1 _14623_ (.A(net5355),
    .B(_10088_),
    .Y(_10089_));
 sg13g2_o21ai_1 _14624_ (.B1(_10089_),
    .Y(_10090_),
    .A1(\soc_inst.core_instr_addr[15] ),
    .A2(_10082_));
 sg13g2_a21oi_1 _14625_ (.A1(\soc_inst.cpu_core.ex_branch_target[15] ),
    .A2(net5356),
    .Y(_10091_),
    .B1(net4937));
 sg13g2_o21ai_1 _14626_ (.B1(net6162),
    .Y(_10092_),
    .A1(net503),
    .A2(net4946));
 sg13g2_a21oi_1 _14627_ (.A1(_10090_),
    .A2(_10091_),
    .Y(_10093_),
    .B1(_10092_));
 sg13g2_nand2_1 _14628_ (.Y(_10094_),
    .A(net6473),
    .B(net2449));
 sg13g2_nor2_1 _14629_ (.A(net4730),
    .B(_10093_),
    .Y(_10095_));
 sg13g2_a22oi_1 _14630_ (.Y(_00536_),
    .B1(_10094_),
    .B2(_10095_),
    .A2(net4731),
    .A1(_07848_));
 sg13g2_a21oi_1 _14631_ (.A1(\soc_inst.core_instr_addr[16] ),
    .A2(_10088_),
    .Y(_10096_),
    .B1(net5355));
 sg13g2_o21ai_1 _14632_ (.B1(_10096_),
    .Y(_10097_),
    .A1(\soc_inst.core_instr_addr[16] ),
    .A2(_10088_));
 sg13g2_a21oi_1 _14633_ (.A1(net2005),
    .A2(net5356),
    .Y(_10098_),
    .B1(net4938));
 sg13g2_o21ai_1 _14634_ (.B1(net6162),
    .Y(_10099_),
    .A1(net1143),
    .A2(net4946));
 sg13g2_a21o_1 _14635_ (.A2(_10098_),
    .A1(_10097_),
    .B1(_10099_),
    .X(_10100_));
 sg13g2_a21oi_1 _14636_ (.A1(net6473),
    .A2(net2114),
    .Y(_10101_),
    .B1(net4729));
 sg13g2_a22oi_1 _14637_ (.Y(_00537_),
    .B1(_10100_),
    .B2(_10101_),
    .A2(net4729),
    .A1(_07850_));
 sg13g2_a21oi_1 _14638_ (.A1(\soc_inst.core_instr_addr[16] ),
    .A2(_10088_),
    .Y(_10102_),
    .B1(\soc_inst.core_instr_addr[17] ));
 sg13g2_nand3_1 _14639_ (.B(\soc_inst.core_instr_addr[17] ),
    .C(_10088_),
    .A(\soc_inst.core_instr_addr[16] ),
    .Y(_10103_));
 sg13g2_nor2_1 _14640_ (.A(net5355),
    .B(_10102_),
    .Y(_10104_));
 sg13g2_a221oi_1 _14641_ (.B2(_10104_),
    .C1(net4937),
    .B1(_10103_),
    .A1(net3034),
    .Y(_10105_),
    .A2(net5355));
 sg13g2_o21ai_1 _14642_ (.B1(net6162),
    .Y(_10106_),
    .A1(net1024),
    .A2(net4946));
 sg13g2_or2_1 _14643_ (.X(_10107_),
    .B(_10106_),
    .A(_10105_));
 sg13g2_a21oi_1 _14644_ (.A1(net6473),
    .A2(net1966),
    .Y(_10108_),
    .B1(net4729));
 sg13g2_a22oi_1 _14645_ (.Y(_00538_),
    .B1(_10107_),
    .B2(_10108_),
    .A2(net4729),
    .A1(_07852_));
 sg13g2_nand2_1 _14646_ (.Y(_10109_),
    .A(_07854_),
    .B(_10103_));
 sg13g2_and4_1 _14647_ (.A(\soc_inst.core_instr_addr[16] ),
    .B(\soc_inst.core_instr_addr[17] ),
    .C(\soc_inst.core_instr_addr[18] ),
    .D(_10088_),
    .X(_10110_));
 sg13g2_nor2_1 _14648_ (.A(net5355),
    .B(_10110_),
    .Y(_10111_));
 sg13g2_a221oi_1 _14649_ (.B2(_10111_),
    .C1(net4937),
    .B1(_10109_),
    .A1(net2476),
    .Y(_10112_),
    .A2(net5355));
 sg13g2_o21ai_1 _14650_ (.B1(net6162),
    .Y(_10113_),
    .A1(net464),
    .A2(net4946));
 sg13g2_or2_1 _14651_ (.X(_10114_),
    .B(_10113_),
    .A(_10112_));
 sg13g2_a21oi_1 _14652_ (.A1(net6473),
    .A2(net2534),
    .Y(_10115_),
    .B1(net4730));
 sg13g2_a22oi_1 _14653_ (.Y(_00539_),
    .B1(_10114_),
    .B2(_10115_),
    .A2(net4730),
    .A1(_07854_));
 sg13g2_nor2_1 _14654_ (.A(\soc_inst.core_instr_addr[19] ),
    .B(_10110_),
    .Y(_10116_));
 sg13g2_nand2_1 _14655_ (.Y(_10117_),
    .A(\soc_inst.core_instr_addr[19] ),
    .B(_10110_));
 sg13g2_nor2_1 _14656_ (.A(net5355),
    .B(_10116_),
    .Y(_10118_));
 sg13g2_a221oi_1 _14657_ (.B2(_10118_),
    .C1(net4937),
    .B1(_10117_),
    .A1(net2441),
    .Y(_10119_),
    .A2(net5356));
 sg13g2_o21ai_1 _14658_ (.B1(net6162),
    .Y(_10120_),
    .A1(net611),
    .A2(net4946));
 sg13g2_or2_1 _14659_ (.X(_10121_),
    .B(_10120_),
    .A(_10119_));
 sg13g2_a21oi_1 _14660_ (.A1(net6473),
    .A2(net2796),
    .Y(_10122_),
    .B1(net4729));
 sg13g2_a22oi_1 _14661_ (.Y(_00540_),
    .B1(_10121_),
    .B2(_10122_),
    .A2(net4729),
    .A1(_07856_));
 sg13g2_nand3_1 _14662_ (.B(\soc_inst.core_instr_addr[20] ),
    .C(_10110_),
    .A(\soc_inst.core_instr_addr[19] ),
    .Y(_10123_));
 sg13g2_xnor2_1 _14663_ (.Y(_10124_),
    .A(_07858_),
    .B(_10117_));
 sg13g2_a21oi_1 _14664_ (.A1(net2719),
    .A2(net5355),
    .Y(_10125_),
    .B1(net4938));
 sg13g2_o21ai_1 _14665_ (.B1(_10125_),
    .Y(_10126_),
    .A1(net5356),
    .A2(_10124_));
 sg13g2_o21ai_1 _14666_ (.B1(net6162),
    .Y(_10127_),
    .A1(net344),
    .A2(net4946));
 sg13g2_nand2b_1 _14667_ (.Y(_10128_),
    .B(_10126_),
    .A_N(_10127_));
 sg13g2_a21oi_1 _14668_ (.A1(net6473),
    .A2(net1576),
    .Y(_10129_),
    .B1(net4729));
 sg13g2_a22oi_1 _14669_ (.Y(_00541_),
    .B1(_10128_),
    .B2(_10129_),
    .A2(net4729),
    .A1(_07858_));
 sg13g2_nor2_1 _14670_ (.A(_07860_),
    .B(_10123_),
    .Y(_10130_));
 sg13g2_xnor2_1 _14671_ (.Y(_10131_),
    .A(_07860_),
    .B(_10123_));
 sg13g2_a21oi_1 _14672_ (.A1(net2754),
    .A2(net5358),
    .Y(_10132_),
    .B1(net4937));
 sg13g2_o21ai_1 _14673_ (.B1(_10132_),
    .Y(_10133_),
    .A1(net5358),
    .A2(_10131_));
 sg13g2_a21oi_1 _14674_ (.A1(_08022_),
    .A2(net4939),
    .Y(_10134_),
    .B1(net6472));
 sg13g2_a221oi_1 _14675_ (.B2(_10134_),
    .C1(net4732),
    .B1(_10133_),
    .A1(net6472),
    .Y(_10135_),
    .A2(net2586));
 sg13g2_a21oi_1 _14676_ (.A1(_07860_),
    .A2(net4732),
    .Y(_00542_),
    .B1(_10135_));
 sg13g2_nand2_1 _14677_ (.Y(_10136_),
    .A(net3405),
    .B(_10130_));
 sg13g2_xnor2_1 _14678_ (.Y(_10137_),
    .A(\soc_inst.core_instr_addr[22] ),
    .B(_10130_));
 sg13g2_a21oi_1 _14679_ (.A1(net2830),
    .A2(net5358),
    .Y(_10138_),
    .B1(net4937));
 sg13g2_o21ai_1 _14680_ (.B1(_10138_),
    .Y(_10139_),
    .A1(net5358),
    .A2(_10137_));
 sg13g2_a21oi_1 _14681_ (.A1(_08024_),
    .A2(net4939),
    .Y(_10140_),
    .B1(net6472));
 sg13g2_a221oi_1 _14682_ (.B2(_10140_),
    .C1(net4732),
    .B1(_10139_),
    .A1(net6472),
    .Y(_10141_),
    .A2(net2133));
 sg13g2_a21oi_1 _14683_ (.A1(_07862_),
    .A2(net4732),
    .Y(_00543_),
    .B1(_10141_));
 sg13g2_xnor2_1 _14684_ (.Y(_10142_),
    .A(_07864_),
    .B(_10136_));
 sg13g2_a21oi_1 _14685_ (.A1(net2238),
    .A2(net5358),
    .Y(_10143_),
    .B1(net4937));
 sg13g2_o21ai_1 _14686_ (.B1(_10143_),
    .Y(_10144_),
    .A1(net5358),
    .A2(_10142_));
 sg13g2_o21ai_1 _14687_ (.B1(net6162),
    .Y(_10145_),
    .A1(net948),
    .A2(net4947));
 sg13g2_nand2b_1 _14688_ (.Y(_10146_),
    .B(_10144_),
    .A_N(_10145_));
 sg13g2_a21oi_1 _14689_ (.A1(net6473),
    .A2(net2460),
    .Y(_10147_),
    .B1(net4730));
 sg13g2_a22oi_1 _14690_ (.Y(_00544_),
    .B1(_10146_),
    .B2(_10147_),
    .A2(net4732),
    .A1(_07864_));
 sg13g2_a22oi_1 _14691_ (.Y(_10148_),
    .B1(_09265_),
    .B2(net6539),
    .A2(_08825_),
    .A1(_08401_));
 sg13g2_nand2_1 _14692_ (.Y(_10149_),
    .A(_09473_),
    .B(_10148_));
 sg13g2_nor3_1 _14693_ (.A(\soc_inst.i2c_inst.stop_pending ),
    .B(net5565),
    .C(_09231_),
    .Y(_10150_));
 sg13g2_a21oi_1 _14694_ (.A1(_08814_),
    .A2(_10149_),
    .Y(_10151_),
    .B1(_10150_));
 sg13g2_nand3_1 _14695_ (.B(_09469_),
    .C(_10151_),
    .A(_09267_),
    .Y(_10152_));
 sg13g2_nand2b_1 _14696_ (.Y(_10153_),
    .B(net3186),
    .A_N(net1013));
 sg13g2_nor4_1 _14697_ (.A(net3121),
    .B(net2965),
    .C(_09273_),
    .D(_10153_),
    .Y(_10154_));
 sg13g2_o21ai_1 _14698_ (.B1(_09226_),
    .Y(_10155_),
    .A1(net1565),
    .A2(net594));
 sg13g2_nor4_1 _14699_ (.A(_08404_),
    .B(_09466_),
    .C(_10152_),
    .D(_10154_),
    .Y(_10156_));
 sg13g2_a22oi_1 _14700_ (.Y(_00545_),
    .B1(_10155_),
    .B2(_10156_),
    .A2(_10152_),
    .A1(_07893_));
 sg13g2_nor2_1 _14701_ (.A(net1565),
    .B(_09227_),
    .Y(_10157_));
 sg13g2_nand2b_1 _14702_ (.Y(_10158_),
    .B(_09226_),
    .A_N(net1565));
 sg13g2_a22oi_1 _14703_ (.Y(_10159_),
    .B1(_10157_),
    .B2(net594),
    .A2(_09466_),
    .A1(net6537));
 sg13g2_a21oi_1 _14704_ (.A1(_09470_),
    .A2(_10159_),
    .Y(_10160_),
    .B1(_10152_));
 sg13g2_a21o_1 _14705_ (.A2(_10152_),
    .A1(net6538),
    .B1(_10160_),
    .X(_00546_));
 sg13g2_nand3_1 _14706_ (.B(_10148_),
    .C(_10158_),
    .A(_09465_),
    .Y(_10161_));
 sg13g2_mux2_1 _14707_ (.A0(_10161_),
    .A1(net6536),
    .S(_10152_),
    .X(_00547_));
 sg13g2_nand3_1 _14708_ (.B(_08829_),
    .C(_09467_),
    .A(_08799_),
    .Y(_10162_));
 sg13g2_a21oi_1 _14709_ (.A1(net1565),
    .A2(_09226_),
    .Y(_10163_),
    .B1(_10162_));
 sg13g2_nand2_1 _14710_ (.Y(_10164_),
    .A(net6534),
    .B(_10152_));
 sg13g2_o21ai_1 _14711_ (.B1(_10164_),
    .Y(_00548_),
    .A1(_10152_),
    .A2(_10163_));
 sg13g2_a21o_1 _14712_ (.A2(_08366_),
    .A1(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .B1(_07866_),
    .X(_10165_));
 sg13g2_nor3_1 _14713_ (.A(_07866_),
    .B(net3150),
    .C(_08383_),
    .Y(_10166_));
 sg13g2_nand3_1 _14714_ (.B(_09830_),
    .C(_10165_),
    .A(_09819_),
    .Y(_10167_));
 sg13g2_o21ai_1 _14715_ (.B1(_07866_),
    .Y(_10168_),
    .A1(\soc_inst.mem_ctrl.access_state[4] ),
    .A2(_08246_));
 sg13g2_nor2_1 _14716_ (.A(net6181),
    .B(_09823_),
    .Y(_10169_));
 sg13g2_a221oi_1 _14717_ (.B2(\soc_inst.core_mem_addr[0] ),
    .C1(net4712),
    .B1(net5324),
    .A1(net2927),
    .Y(_10170_),
    .A2(net5523));
 sg13g2_a21oi_1 _14718_ (.A1(_07817_),
    .A2(net4712),
    .Y(_00549_),
    .B1(_10170_));
 sg13g2_a221oi_1 _14719_ (.B2(\soc_inst.core_mem_addr[1] ),
    .C1(net4710),
    .B1(net5324),
    .A1(net2685),
    .Y(_10171_),
    .A2(net5523));
 sg13g2_a21oi_1 _14720_ (.A1(_07819_),
    .A2(net4712),
    .Y(_00550_),
    .B1(_10171_));
 sg13g2_a221oi_1 _14721_ (.B2(\soc_inst.core_mem_addr[2] ),
    .C1(net4710),
    .B1(net5325),
    .A1(\soc_inst.core_instr_addr[2] ),
    .Y(_10172_),
    .A2(net5524));
 sg13g2_a21oi_1 _14722_ (.A1(_07821_),
    .A2(net4709),
    .Y(_00551_),
    .B1(_10172_));
 sg13g2_a221oi_1 _14723_ (.B2(net6210),
    .C1(net4710),
    .B1(net5324),
    .A1(net2492),
    .Y(_10173_),
    .A2(net5523));
 sg13g2_a21oi_1 _14724_ (.A1(_07823_),
    .A2(net4710),
    .Y(_00552_),
    .B1(_10173_));
 sg13g2_a221oi_1 _14725_ (.B2(net2908),
    .C1(net4709),
    .B1(net5325),
    .A1(net2738),
    .Y(_10174_),
    .A2(net5524));
 sg13g2_a21oi_1 _14726_ (.A1(_07825_),
    .A2(net4709),
    .Y(_00553_),
    .B1(_10174_));
 sg13g2_a221oi_1 _14727_ (.B2(net3038),
    .C1(net4709),
    .B1(net5324),
    .A1(net2703),
    .Y(_10175_),
    .A2(net5523));
 sg13g2_a21oi_1 _14728_ (.A1(_07827_),
    .A2(net4709),
    .Y(_00554_),
    .B1(_10175_));
 sg13g2_a221oi_1 _14729_ (.B2(net2958),
    .C1(net4709),
    .B1(net5324),
    .A1(net2713),
    .Y(_10176_),
    .A2(net5523));
 sg13g2_a21oi_1 _14730_ (.A1(_07829_),
    .A2(net4709),
    .Y(_00555_),
    .B1(_10176_));
 sg13g2_a221oi_1 _14731_ (.B2(net3104),
    .C1(net4709),
    .B1(net5324),
    .A1(net2807),
    .Y(_10177_),
    .A2(net5523));
 sg13g2_a21oi_1 _14732_ (.A1(_07831_),
    .A2(net4711),
    .Y(_00556_),
    .B1(_10177_));
 sg13g2_a221oi_1 _14733_ (.B2(net1051),
    .C1(net4711),
    .B1(net5324),
    .A1(net2493),
    .Y(_10178_),
    .A2(net5523));
 sg13g2_a21oi_1 _14734_ (.A1(_07833_),
    .A2(net4708),
    .Y(_00557_),
    .B1(_10178_));
 sg13g2_a221oi_1 _14735_ (.B2(net1927),
    .C1(net4711),
    .B1(net5324),
    .A1(net3044),
    .Y(_10179_),
    .A2(net5523));
 sg13g2_a21oi_1 _14736_ (.A1(_07835_),
    .A2(net4712),
    .Y(_00558_),
    .B1(_10179_));
 sg13g2_a221oi_1 _14737_ (.B2(net1110),
    .C1(net4708),
    .B1(net5323),
    .A1(\soc_inst.core_instr_addr[10] ),
    .Y(_10180_),
    .A2(net5522));
 sg13g2_a21oi_1 _14738_ (.A1(_07837_),
    .A2(net4708),
    .Y(_00559_),
    .B1(_10180_));
 sg13g2_a221oi_1 _14739_ (.B2(net1538),
    .C1(net4708),
    .B1(net5323),
    .A1(\soc_inst.core_instr_addr[11] ),
    .Y(_10181_),
    .A2(net5522));
 sg13g2_a21oi_1 _14740_ (.A1(_07839_),
    .A2(net4707),
    .Y(_00560_),
    .B1(_10181_));
 sg13g2_a221oi_1 _14741_ (.B2(\soc_inst.core_mem_addr[12] ),
    .C1(net4707),
    .B1(net5322),
    .A1(\soc_inst.core_instr_addr[12] ),
    .Y(_10182_),
    .A2(net5521));
 sg13g2_a21oi_1 _14742_ (.A1(_07841_),
    .A2(net4712),
    .Y(_00561_),
    .B1(_10182_));
 sg13g2_a221oi_1 _14743_ (.B2(\soc_inst.core_mem_addr[13] ),
    .C1(net4707),
    .B1(net5322),
    .A1(\soc_inst.core_instr_addr[13] ),
    .Y(_10183_),
    .A2(net5521));
 sg13g2_a21oi_1 _14744_ (.A1(_07843_),
    .A2(net4707),
    .Y(_00562_),
    .B1(_10183_));
 sg13g2_a221oi_1 _14745_ (.B2(\soc_inst.core_mem_addr[14] ),
    .C1(net4705),
    .B1(net5321),
    .A1(\soc_inst.core_instr_addr[14] ),
    .Y(_10184_),
    .A2(net5520));
 sg13g2_a21oi_1 _14746_ (.A1(_07845_),
    .A2(net4705),
    .Y(_00563_),
    .B1(_10184_));
 sg13g2_a221oi_1 _14747_ (.B2(net2365),
    .C1(net4708),
    .B1(net5323),
    .A1(\soc_inst.core_instr_addr[15] ),
    .Y(_10185_),
    .A2(net5522));
 sg13g2_a21oi_1 _14748_ (.A1(_07847_),
    .A2(net4708),
    .Y(_00564_),
    .B1(_10185_));
 sg13g2_a221oi_1 _14749_ (.B2(net3105),
    .C1(net4705),
    .B1(net5321),
    .A1(net3138),
    .Y(_10186_),
    .A2(net5520));
 sg13g2_a21oi_1 _14750_ (.A1(_07849_),
    .A2(net4705),
    .Y(_00565_),
    .B1(_10186_));
 sg13g2_a221oi_1 _14751_ (.B2(net2856),
    .C1(net4705),
    .B1(net5321),
    .A1(net3092),
    .Y(_10187_),
    .A2(net5520));
 sg13g2_a21oi_1 _14752_ (.A1(_07851_),
    .A2(net4705),
    .Y(_00566_),
    .B1(_10187_));
 sg13g2_a221oi_1 _14753_ (.B2(net2836),
    .C1(net4706),
    .B1(net5321),
    .A1(net2925),
    .Y(_10188_),
    .A2(net5520));
 sg13g2_a21oi_1 _14754_ (.A1(_07853_),
    .A2(net4705),
    .Y(_00567_),
    .B1(_10188_));
 sg13g2_a221oi_1 _14755_ (.B2(net2687),
    .C1(net4706),
    .B1(net5321),
    .A1(\soc_inst.core_instr_addr[19] ),
    .Y(_10189_),
    .A2(net5520));
 sg13g2_a21oi_1 _14756_ (.A1(_07855_),
    .A2(net4705),
    .Y(_00568_),
    .B1(_10189_));
 sg13g2_a221oi_1 _14757_ (.B2(net2805),
    .C1(net4706),
    .B1(net5321),
    .A1(\soc_inst.core_instr_addr[20] ),
    .Y(_10190_),
    .A2(net5520));
 sg13g2_a21oi_1 _14758_ (.A1(_07857_),
    .A2(net4707),
    .Y(_00569_),
    .B1(_10190_));
 sg13g2_a221oi_1 _14759_ (.B2(net2889),
    .C1(net4706),
    .B1(net5321),
    .A1(net2693),
    .Y(_10191_),
    .A2(net5520));
 sg13g2_a21oi_1 _14760_ (.A1(_07859_),
    .A2(net4706),
    .Y(_00570_),
    .B1(_10191_));
 sg13g2_a221oi_1 _14761_ (.B2(net2694),
    .C1(net4706),
    .B1(net5321),
    .A1(\soc_inst.core_instr_addr[22] ),
    .Y(_10192_),
    .A2(net5520));
 sg13g2_a21oi_1 _14762_ (.A1(_07861_),
    .A2(net4707),
    .Y(_00571_),
    .B1(_10192_));
 sg13g2_a221oi_1 _14763_ (.B2(\soc_inst.core_mem_addr[23] ),
    .C1(net4706),
    .B1(net5322),
    .A1(\soc_inst.core_instr_addr[23] ),
    .Y(_10193_),
    .A2(net5521));
 sg13g2_a21oi_1 _14764_ (.A1(_07863_),
    .A2(net4707),
    .Y(_00572_),
    .B1(_10193_));
 sg13g2_o21ai_1 _14765_ (.B1(_09828_),
    .Y(_10194_),
    .A1(net6181),
    .A2(\soc_inst.mem_ctrl.access_state[3] ));
 sg13g2_or3_1 _14766_ (.A(_08387_),
    .B(_10166_),
    .C(_10194_),
    .X(_10195_));
 sg13g2_nor2_1 _14767_ (.A(net6183),
    .B(net2759),
    .Y(_10196_));
 sg13g2_a21oi_1 _14768_ (.A1(net6183),
    .A2(_07967_),
    .Y(_10197_),
    .B1(_10196_));
 sg13g2_mux2_1 _14769_ (.A0(_10197_),
    .A1(net6533),
    .S(net4700),
    .X(_00573_));
 sg13g2_nor2_1 _14770_ (.A(net6182),
    .B(net2602),
    .Y(_10198_));
 sg13g2_a21oi_1 _14771_ (.A1(net6183),
    .A2(_07968_),
    .Y(_10199_),
    .B1(_10198_));
 sg13g2_mux2_1 _14772_ (.A0(_10199_),
    .A1(net6532),
    .S(net4700),
    .X(_00574_));
 sg13g2_nor2_1 _14773_ (.A(net6185),
    .B(net2409),
    .Y(_10200_));
 sg13g2_a21oi_1 _14774_ (.A1(net6189),
    .A2(_07969_),
    .Y(_10201_),
    .B1(_10200_));
 sg13g2_mux2_1 _14775_ (.A0(_10201_),
    .A1(net2761),
    .S(net4701),
    .X(_00575_));
 sg13g2_nor2_1 _14776_ (.A(net6186),
    .B(net2507),
    .Y(_10202_));
 sg13g2_a21oi_1 _14777_ (.A1(net6189),
    .A2(_07970_),
    .Y(_10203_),
    .B1(_10202_));
 sg13g2_mux2_1 _14778_ (.A0(_10203_),
    .A1(net2799),
    .S(net4702),
    .X(_00576_));
 sg13g2_nor2_1 _14779_ (.A(net6183),
    .B(net2105),
    .Y(_10204_));
 sg13g2_a21oi_1 _14780_ (.A1(net6188),
    .A2(_07971_),
    .Y(_10205_),
    .B1(_10204_));
 sg13g2_mux2_1 _14781_ (.A0(_10205_),
    .A1(net6529),
    .S(net4700),
    .X(_00577_));
 sg13g2_nor2_1 _14782_ (.A(net6184),
    .B(net2410),
    .Y(_10206_));
 sg13g2_a21oi_1 _14783_ (.A1(net6185),
    .A2(_07972_),
    .Y(_10207_),
    .B1(_10206_));
 sg13g2_mux2_1 _14784_ (.A0(_10207_),
    .A1(net6528),
    .S(net4704),
    .X(_00578_));
 sg13g2_nor2_1 _14785_ (.A(net6187),
    .B(net2641),
    .Y(_10208_));
 sg13g2_a21oi_1 _14786_ (.A1(net6186),
    .A2(_07973_),
    .Y(_10209_),
    .B1(_10208_));
 sg13g2_mux2_1 _14787_ (.A0(_10209_),
    .A1(net6526),
    .S(net4702),
    .X(_00579_));
 sg13g2_nor2_1 _14788_ (.A(net6187),
    .B(net2619),
    .Y(_10210_));
 sg13g2_a21oi_1 _14789_ (.A1(net6189),
    .A2(_07974_),
    .Y(_10211_),
    .B1(_10210_));
 sg13g2_mux2_1 _14790_ (.A0(_10211_),
    .A1(net6525),
    .S(net4702),
    .X(_00580_));
 sg13g2_nor2_1 _14791_ (.A(net6184),
    .B(net2957),
    .Y(_10212_));
 sg13g2_a21oi_1 _14792_ (.A1(net6184),
    .A2(_07975_),
    .Y(_10213_),
    .B1(_10212_));
 sg13g2_mux2_1 _14793_ (.A0(_10213_),
    .A1(net6523),
    .S(net4701),
    .X(_00581_));
 sg13g2_nor2_1 _14794_ (.A(net6189),
    .B(net3006),
    .Y(_10214_));
 sg13g2_a21oi_1 _14795_ (.A1(net6189),
    .A2(_07976_),
    .Y(_10215_),
    .B1(_10214_));
 sg13g2_nor2_1 _14796_ (.A(net4701),
    .B(_10215_),
    .Y(_10216_));
 sg13g2_a21oi_1 _14797_ (.A1(_08026_),
    .A2(net4701),
    .Y(_00582_),
    .B1(_10216_));
 sg13g2_nor2_1 _14798_ (.A(net6187),
    .B(net2709),
    .Y(_10217_));
 sg13g2_a21oi_1 _14799_ (.A1(net6186),
    .A2(_07977_),
    .Y(_10218_),
    .B1(_10217_));
 sg13g2_nor2_1 _14800_ (.A(net4702),
    .B(_10218_),
    .Y(_10219_));
 sg13g2_a21oi_1 _14801_ (.A1(_08027_),
    .A2(net4701),
    .Y(_00583_),
    .B1(_10219_));
 sg13g2_nor2_1 _14802_ (.A(net6187),
    .B(net2916),
    .Y(_10220_));
 sg13g2_a21oi_1 _14803_ (.A1(net6187),
    .A2(_07978_),
    .Y(_10221_),
    .B1(_10220_));
 sg13g2_mux2_1 _14804_ (.A0(_10221_),
    .A1(net6518),
    .S(net4704),
    .X(_00584_));
 sg13g2_nor2_1 _14805_ (.A(net6190),
    .B(net2981),
    .Y(_10222_));
 sg13g2_a21oi_1 _14806_ (.A1(net6189),
    .A2(_07979_),
    .Y(_10223_),
    .B1(_10222_));
 sg13g2_nor2_1 _14807_ (.A(net4704),
    .B(_10223_),
    .Y(_10224_));
 sg13g2_a21oi_1 _14808_ (.A1(_08028_),
    .A2(net4703),
    .Y(_00585_),
    .B1(_10224_));
 sg13g2_nor2_1 _14809_ (.A(net6180),
    .B(net2776),
    .Y(_10225_));
 sg13g2_a21oi_1 _14810_ (.A1(net6180),
    .A2(_07980_),
    .Y(_10226_),
    .B1(_10225_));
 sg13g2_mux2_1 _14811_ (.A0(_10226_),
    .A1(net6512),
    .S(net4700),
    .X(_00586_));
 sg13g2_nor2_1 _14812_ (.A(net6180),
    .B(net2533),
    .Y(_10227_));
 sg13g2_a21oi_1 _14813_ (.A1(net6180),
    .A2(_07981_),
    .Y(_10228_),
    .B1(_10227_));
 sg13g2_mux2_1 _14814_ (.A0(_10228_),
    .A1(net6510),
    .S(net4701),
    .X(_00587_));
 sg13g2_nor2_1 _14815_ (.A(net6181),
    .B(net2722),
    .Y(_10229_));
 sg13g2_a21oi_1 _14816_ (.A1(net6180),
    .A2(_07982_),
    .Y(_10230_),
    .B1(_10229_));
 sg13g2_mux2_1 _14817_ (.A0(_10230_),
    .A1(net6508),
    .S(net4701),
    .X(_00588_));
 sg13g2_nor2_1 _14818_ (.A(net6184),
    .B(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .Y(_10231_));
 sg13g2_a21oi_1 _14819_ (.A1(net6188),
    .A2(_07983_),
    .Y(_10232_),
    .B1(_10231_));
 sg13g2_mux2_1 _14820_ (.A0(_10232_),
    .A1(net2667),
    .S(net4703),
    .X(_00589_));
 sg13g2_nor2_1 _14821_ (.A(net6185),
    .B(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .Y(_10233_));
 sg13g2_a21oi_1 _14822_ (.A1(net6188),
    .A2(_07984_),
    .Y(_10234_),
    .B1(_10233_));
 sg13g2_mux2_1 _14823_ (.A0(_10234_),
    .A1(net2696),
    .S(net4703),
    .X(_00590_));
 sg13g2_nor2_1 _14824_ (.A(net6182),
    .B(net2633),
    .Y(_10235_));
 sg13g2_a21oi_1 _14825_ (.A1(net6182),
    .A2(_07985_),
    .Y(_10236_),
    .B1(_10235_));
 sg13g2_mux2_1 _14826_ (.A0(_10236_),
    .A1(net2740),
    .S(net4703),
    .X(_00591_));
 sg13g2_nor2_1 _14827_ (.A(net6180),
    .B(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .Y(_10237_));
 sg13g2_a21oi_1 _14828_ (.A1(net6180),
    .A2(_07986_),
    .Y(_10238_),
    .B1(_10237_));
 sg13g2_mux2_1 _14829_ (.A0(_10238_),
    .A1(net2645),
    .S(net4703),
    .X(_00592_));
 sg13g2_nor2_1 _14830_ (.A(net6186),
    .B(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .Y(_10239_));
 sg13g2_a21oi_1 _14831_ (.A1(net6186),
    .A2(_07987_),
    .Y(_10240_),
    .B1(_10239_));
 sg13g2_mux2_1 _14832_ (.A0(_10240_),
    .A1(net2867),
    .S(net4702),
    .X(_00593_));
 sg13g2_nor2_1 _14833_ (.A(net6180),
    .B(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .Y(_10241_));
 sg13g2_a21oi_1 _14834_ (.A1(net6184),
    .A2(_07988_),
    .Y(_10242_),
    .B1(_10241_));
 sg13g2_mux2_1 _14835_ (.A0(_10242_),
    .A1(net2541),
    .S(net4702),
    .X(_00594_));
 sg13g2_nor2_1 _14836_ (.A(net6186),
    .B(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .Y(_10243_));
 sg13g2_a21oi_1 _14837_ (.A1(net6189),
    .A2(_07989_),
    .Y(_10244_),
    .B1(_10243_));
 sg13g2_mux2_1 _14838_ (.A0(_10244_),
    .A1(net2402),
    .S(net4701),
    .X(_00595_));
 sg13g2_nor2_1 _14839_ (.A(net6190),
    .B(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .Y(_10245_));
 sg13g2_a21oi_1 _14840_ (.A1(net6189),
    .A2(_07990_),
    .Y(_10246_),
    .B1(_10245_));
 sg13g2_mux2_1 _14841_ (.A0(_10246_),
    .A1(net2453),
    .S(net4704),
    .X(_00596_));
 sg13g2_nor2_1 _14842_ (.A(net6186),
    .B(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .Y(_10247_));
 sg13g2_a21oi_1 _14843_ (.A1(net6186),
    .A2(_07991_),
    .Y(_10248_),
    .B1(_10247_));
 sg13g2_mux2_1 _14844_ (.A0(_10248_),
    .A1(net2474),
    .S(net4702),
    .X(_00597_));
 sg13g2_nor2_1 _14845_ (.A(net6188),
    .B(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .Y(_10249_));
 sg13g2_a21oi_1 _14846_ (.A1(net6188),
    .A2(_07992_),
    .Y(_10250_),
    .B1(_10249_));
 sg13g2_mux2_1 _14847_ (.A0(_10250_),
    .A1(net2436),
    .S(net4703),
    .X(_00598_));
 sg13g2_nor2_1 _14848_ (.A(net6188),
    .B(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .Y(_10251_));
 sg13g2_a21oi_1 _14849_ (.A1(net6188),
    .A2(_07993_),
    .Y(_10252_),
    .B1(_10251_));
 sg13g2_mux2_1 _14850_ (.A0(_10252_),
    .A1(net2549),
    .S(net4703),
    .X(_00599_));
 sg13g2_nor2_1 _14851_ (.A(net6184),
    .B(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .Y(_10253_));
 sg13g2_a21oi_1 _14852_ (.A1(net6185),
    .A2(_07994_),
    .Y(_10254_),
    .B1(_10253_));
 sg13g2_mux2_1 _14853_ (.A0(_10254_),
    .A1(net2578),
    .S(net4703),
    .X(_00600_));
 sg13g2_nor2_1 _14854_ (.A(net6182),
    .B(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .Y(_10255_));
 sg13g2_a21oi_1 _14855_ (.A1(net6188),
    .A2(_07995_),
    .Y(_10256_),
    .B1(_10255_));
 sg13g2_mux2_1 _14856_ (.A0(_10256_),
    .A1(net2576),
    .S(net4700),
    .X(_00601_));
 sg13g2_nor2_1 _14857_ (.A(net6182),
    .B(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .Y(_10257_));
 sg13g2_a21oi_1 _14858_ (.A1(net6182),
    .A2(_07996_),
    .Y(_10258_),
    .B1(_10257_));
 sg13g2_mux2_1 _14859_ (.A0(_10258_),
    .A1(net2503),
    .S(net4700),
    .X(_00602_));
 sg13g2_nor2_1 _14860_ (.A(net6182),
    .B(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .Y(_10259_));
 sg13g2_a21oi_1 _14861_ (.A1(net6182),
    .A2(_07997_),
    .Y(_10260_),
    .B1(_10259_));
 sg13g2_mux2_1 _14862_ (.A0(_10260_),
    .A1(net1848),
    .S(net4700),
    .X(_00603_));
 sg13g2_nor2_1 _14863_ (.A(net6184),
    .B(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .Y(_10261_));
 sg13g2_a21oi_1 _14864_ (.A1(net6184),
    .A2(_07998_),
    .Y(_10262_),
    .B1(_10261_));
 sg13g2_mux2_1 _14865_ (.A0(_10262_),
    .A1(net1446),
    .S(net4700),
    .X(_00604_));
 sg13g2_nand2_1 _14866_ (.Y(_10263_),
    .A(_08248_),
    .B(_08391_));
 sg13g2_a21oi_1 _14867_ (.A1(net5190),
    .A2(_10263_),
    .Y(_10264_),
    .B1(_08399_));
 sg13g2_nor2_1 _14868_ (.A(net6507),
    .B(_07867_),
    .Y(_10265_));
 sg13g2_o21ai_1 _14869_ (.B1(_10264_),
    .Y(_10266_),
    .A1(_08250_),
    .A2(_10265_));
 sg13g2_nand2_2 _14870_ (.Y(_10267_),
    .A(net6290),
    .B(net6103));
 sg13g2_inv_1 _14871_ (.Y(_10268_),
    .A(_10267_));
 sg13g2_nand2_1 _14872_ (.Y(_10269_),
    .A(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .B(_10267_));
 sg13g2_a22oi_1 _14873_ (.Y(_10270_),
    .B1(_10268_),
    .B2(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .A2(net6107),
    .A1(net6290));
 sg13g2_nor2_2 _14874_ (.A(_08983_),
    .B(_08987_),
    .Y(_10271_));
 sg13g2_a221oi_1 _14875_ (.B2(_10270_),
    .C1(_08987_),
    .B1(_10269_),
    .A1(_07950_),
    .Y(_10272_),
    .A2(net6107));
 sg13g2_a221oi_1 _14876_ (.B2(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .C1(_10272_),
    .B1(_09671_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .Y(_10273_),
    .A2(_08988_));
 sg13g2_nor2_2 _14877_ (.A(net2919),
    .B(net6487),
    .Y(_10274_));
 sg13g2_nor2_2 _14878_ (.A(_08792_),
    .B(_09423_),
    .Y(_10275_));
 sg13g2_or2_1 _14879_ (.X(_10276_),
    .B(_09423_),
    .A(_08792_));
 sg13g2_a22oi_1 _14880_ (.Y(_10277_),
    .B1(_10275_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .A2(net5566),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ));
 sg13g2_a21oi_1 _14881_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ),
    .A2(net5336),
    .Y(_10278_),
    .B1(net5364));
 sg13g2_nand2b_1 _14882_ (.Y(_10279_),
    .B(net5530),
    .A_N(_00221_));
 sg13g2_or2_1 _14883_ (.X(_10280_),
    .B(net6097),
    .A(\soc_inst.spi_inst.rx_shift_reg[0] ));
 sg13g2_o21ai_1 _14884_ (.B1(_10280_),
    .Y(_10281_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .A2(_09244_));
 sg13g2_a21oi_1 _14885_ (.A1(_07939_),
    .A2(net6544),
    .Y(_10282_),
    .B1(_10281_));
 sg13g2_a221oi_1 _14886_ (.B2(_10282_),
    .C1(_09426_),
    .B1(_10275_),
    .A1(\soc_inst.spi_inst.busy ),
    .Y(_10283_),
    .A2(net5336));
 sg13g2_nand3_1 _14887_ (.B(_08229_),
    .C(_08675_),
    .A(net6212),
    .Y(_10284_));
 sg13g2_a221oi_1 _14888_ (.B2(_10283_),
    .C1(_10284_),
    .B1(_10279_),
    .A1(_07899_),
    .Y(_10285_),
    .A2(_09426_));
 sg13g2_a21oi_1 _14889_ (.A1(_07788_),
    .A2(net6068),
    .Y(_10286_),
    .B1(net6108));
 sg13g2_o21ai_1 _14890_ (.B1(_10286_),
    .Y(_10287_),
    .A1(_00283_),
    .A2(net6050));
 sg13g2_o21ai_1 _14891_ (.B1(_10287_),
    .Y(_10288_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .A2(net6048));
 sg13g2_a21oi_1 _14892_ (.A1(_00173_),
    .A2(net6056),
    .Y(_10289_),
    .B1(_10288_));
 sg13g2_nand2_1 _14893_ (.Y(_10290_),
    .A(net13),
    .B(net5336));
 sg13g2_a22oi_1 _14894_ (.Y(_10291_),
    .B1(net5530),
    .B2(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .A2(net5566),
    .A1(\soc_inst.gpio_inst.int_en_reg[0] ));
 sg13g2_a22oi_1 _14895_ (.Y(_10292_),
    .B1(_09426_),
    .B2(\soc_inst.gpio_bidir_oe [0]),
    .A2(net5363),
    .A1(\soc_inst.gpio_bidir_out [0]));
 sg13g2_nand3_1 _14896_ (.B(_10291_),
    .C(_10292_),
    .A(_10290_),
    .Y(_10293_));
 sg13g2_and2_1 _14897_ (.A(net6212),
    .B(_09441_),
    .X(_10294_));
 sg13g2_a221oi_1 _14898_ (.B2(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .C1(net6109),
    .B1(net5563),
    .A1(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .Y(_10295_),
    .A2(net6067));
 sg13g2_a221oi_1 _14899_ (.B2(_00234_),
    .C1(_10295_),
    .B1(net5559),
    .A1(_07949_),
    .Y(_10296_),
    .A2(net6056));
 sg13g2_nand2_1 _14900_ (.Y(_10297_),
    .A(net6212),
    .B(_08667_));
 sg13g2_nand3_1 _14901_ (.B(_08229_),
    .C(_08793_),
    .A(net6212),
    .Y(_10298_));
 sg13g2_inv_1 _14902_ (.Y(_10299_),
    .A(_10298_));
 sg13g2_nand2_1 _14903_ (.Y(_10300_),
    .A(_00226_),
    .B(net6206));
 sg13g2_a22oi_1 _14904_ (.Y(_10301_),
    .B1(_10300_),
    .B2(net6067),
    .A2(net5563),
    .A1(\soc_inst.i2c_inst.data_reg[0] ));
 sg13g2_nor2_1 _14905_ (.A(\soc_inst.i2c_inst.status_reg[0] ),
    .B(net6049),
    .Y(_10302_));
 sg13g2_nor3_1 _14906_ (.A(_10298_),
    .B(_10301_),
    .C(_10302_),
    .Y(_10303_));
 sg13g2_nand2_2 _14907_ (.Y(_10304_),
    .A(net6212),
    .B(_09308_));
 sg13g2_a221oi_1 _14908_ (.B2(_10278_),
    .C1(_10304_),
    .B1(_10277_),
    .A1(net5364),
    .Y(_10305_),
    .A2(_10274_));
 sg13g2_nor3_2 _14909_ (.A(net5193),
    .B(_10285_),
    .C(_10305_),
    .Y(_10306_));
 sg13g2_nor4_2 _14910_ (.A(_07813_),
    .B(_08231_),
    .C(_08676_),
    .Y(_10307_),
    .D(_10297_));
 sg13g2_a21o_1 _14911_ (.A2(net5128),
    .A1(_10296_),
    .B1(_10303_),
    .X(_10308_));
 sg13g2_nor3_2 _14912_ (.A(_07811_),
    .B(_07813_),
    .C(_09307_),
    .Y(_10309_));
 sg13g2_inv_1 _14913_ (.Y(_10310_),
    .A(net5127));
 sg13g2_a221oi_1 _14914_ (.B2(_10289_),
    .C1(_10308_),
    .B1(net5127),
    .A1(_10293_),
    .Y(_10311_),
    .A2(_10294_));
 sg13g2_a221oi_1 _14915_ (.B2(_10311_),
    .C1(net5041),
    .B1(_10306_),
    .A1(net5188),
    .Y(_10312_),
    .A2(_10273_));
 sg13g2_a21o_1 _14916_ (.A2(net5043),
    .A1(net1314),
    .B1(_10312_),
    .X(_00605_));
 sg13g2_nand2_1 _14917_ (.Y(_10313_),
    .A(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .B(net5128));
 sg13g2_o21ai_1 _14918_ (.B1(_10313_),
    .Y(_10314_),
    .A1(_00227_),
    .A2(_10298_));
 sg13g2_o21ai_1 _14919_ (.B1(net6067),
    .Y(_10315_),
    .A1(_07888_),
    .A2(_10314_));
 sg13g2_a22oi_1 _14920_ (.Y(_10316_),
    .B1(net5128),
    .B2(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .A2(_10299_),
    .A1(\soc_inst.i2c_inst.data_reg[1] ));
 sg13g2_nand2b_1 _14921_ (.Y(_10317_),
    .B(net5563),
    .A_N(_10316_));
 sg13g2_a22oi_1 _14922_ (.Y(_10318_),
    .B1(net5128),
    .B2(_07794_),
    .A2(_10299_),
    .A1(\soc_inst.i2c_inst.status_reg[1] ));
 sg13g2_a22oi_1 _14923_ (.Y(_10319_),
    .B1(_10318_),
    .B2(net5559),
    .A2(_10317_),
    .A1(_10315_));
 sg13g2_a22oi_1 _14924_ (.Y(_10320_),
    .B1(net5530),
    .B2(\soc_inst.gpio_inst.int_pend_reg[1] ),
    .A2(net5566),
    .A1(\soc_inst.gpio_inst.int_en_reg[1] ));
 sg13g2_nor2_2 _14925_ (.A(_10276_),
    .B(_10284_),
    .Y(_10321_));
 sg13g2_and2_1 _14926_ (.A(net6097),
    .B(net5123),
    .X(_10322_));
 sg13g2_nor2b_1 _14927_ (.A(\soc_inst.spi_inst.rx_shift_reg[25] ),
    .B_N(net6544),
    .Y(_10323_));
 sg13g2_nor2_1 _14928_ (.A(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .B(net6098),
    .Y(_10324_));
 sg13g2_nor3_2 _14929_ (.A(net6048),
    .B(_09423_),
    .C(_10284_),
    .Y(_10325_));
 sg13g2_nand2b_1 _14930_ (.Y(_10326_),
    .B(net6103),
    .A_N(\soc_inst.mem_ctrl.spi_data_out[9] ));
 sg13g2_o21ai_1 _14931_ (.B1(net6045),
    .Y(_10327_),
    .A1(net6168),
    .A2(net6106));
 sg13g2_o21ai_1 _14932_ (.B1(_10326_),
    .Y(_10328_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .A2(_10327_));
 sg13g2_a22oi_1 _14933_ (.Y(_10329_),
    .B1(net6046),
    .B2(_10328_),
    .A2(net6107),
    .A1(_07951_));
 sg13g2_nor2_1 _14934_ (.A(_00284_),
    .B(net6050),
    .Y(_10330_));
 sg13g2_nor2_1 _14935_ (.A(_00268_),
    .B(net6063),
    .Y(_10331_));
 sg13g2_nor3_1 _14936_ (.A(net6109),
    .B(_10330_),
    .C(_10331_),
    .Y(_10332_));
 sg13g2_nor2_1 _14937_ (.A(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .B(_08792_),
    .Y(_10333_));
 sg13g2_nor2_1 _14938_ (.A(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .B(net6048),
    .Y(_10334_));
 sg13g2_nor3_1 _14939_ (.A(_10332_),
    .B(_10333_),
    .C(_10334_),
    .Y(_10335_));
 sg13g2_nand2_1 _14940_ (.Y(_10336_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ),
    .B(net5336));
 sg13g2_a22oi_1 _14941_ (.Y(_10337_),
    .B1(_10275_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .A2(net5566),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ));
 sg13g2_a21oi_1 _14942_ (.A1(net2),
    .A2(net5337),
    .Y(_10338_),
    .B1(net5362));
 sg13g2_nor2_1 _14943_ (.A(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .B(_09248_),
    .Y(_10339_));
 sg13g2_a21oi_1 _14944_ (.A1(_10336_),
    .A2(_10337_),
    .Y(_10340_),
    .B1(_10304_));
 sg13g2_a21oi_1 _14945_ (.A1(net5127),
    .A2(_10335_),
    .Y(_10341_),
    .B1(_10340_));
 sg13g2_nor4_1 _14946_ (.A(_10276_),
    .B(_10323_),
    .C(_10324_),
    .D(_10339_),
    .Y(_10342_));
 sg13g2_a221oi_1 _14947_ (.B2(_07798_),
    .C1(_10342_),
    .B1(net5530),
    .A1(\soc_inst.spi_inst.done ),
    .Y(_10343_),
    .A2(net5336));
 sg13g2_o21ai_1 _14948_ (.B1(_10341_),
    .Y(_10344_),
    .A1(_10284_),
    .A2(_10343_));
 sg13g2_o21ai_1 _14949_ (.B1(_10294_),
    .Y(_10345_),
    .A1(\soc_inst.gpio_inst.gpio_out[0] ),
    .A2(_08907_));
 sg13g2_a21oi_1 _14950_ (.A1(_10320_),
    .A2(_10338_),
    .Y(_10346_),
    .B1(_10345_));
 sg13g2_nor3_2 _14951_ (.A(_10319_),
    .B(_10344_),
    .C(_10346_),
    .Y(_10347_));
 sg13g2_a21oi_1 _14952_ (.A1(net5190),
    .A2(_10329_),
    .Y(_10348_),
    .B1(net5038));
 sg13g2_a22oi_1 _14953_ (.Y(_00606_),
    .B1(_10347_),
    .B2(_10348_),
    .A2(net5038),
    .A1(_08000_));
 sg13g2_a21o_1 _14954_ (.A2(net6208),
    .A1(_00269_),
    .B1(net6063),
    .X(_10349_));
 sg13g2_o21ai_1 _14955_ (.B1(_10349_),
    .Y(_10350_),
    .A1(_00285_),
    .A2(net6050));
 sg13g2_nand2_1 _14956_ (.Y(_10351_),
    .A(_07906_),
    .B(net6108));
 sg13g2_a22oi_1 _14957_ (.Y(_10352_),
    .B1(_10350_),
    .B2(_10351_),
    .A2(net6061),
    .A1(\soc_inst.cpu_core.csr_file.mtime[2] ));
 sg13g2_nand2b_1 _14958_ (.Y(_10353_),
    .B(net6545),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[26] ));
 sg13g2_o21ai_1 _14959_ (.B1(_10353_),
    .Y(_10354_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .A2(net6097));
 sg13g2_a21oi_1 _14960_ (.A1(_07934_),
    .A2(_09243_),
    .Y(_10355_),
    .B1(_10354_));
 sg13g2_nor2_1 _14961_ (.A(_00315_),
    .B(_10276_),
    .Y(_10356_));
 sg13g2_a221oi_1 _14962_ (.B2(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .C1(net5559),
    .B1(net5563),
    .A1(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .Y(_10357_),
    .A2(net6067));
 sg13g2_a21oi_1 _14963_ (.A1(_00236_),
    .A2(net5560),
    .Y(_10358_),
    .B1(_10357_));
 sg13g2_a21oi_1 _14964_ (.A1(_00228_),
    .A2(net6206),
    .Y(_10359_),
    .B1(net6064));
 sg13g2_a21o_1 _14965_ (.A2(net5563),
    .A1(\soc_inst.i2c_inst.data_reg[2] ),
    .B1(_10359_),
    .X(_10360_));
 sg13g2_o21ai_1 _14966_ (.B1(_10360_),
    .Y(_10361_),
    .A1(\soc_inst.i2c_inst.status_reg[2] ),
    .A2(net6049));
 sg13g2_nand2_1 _14967_ (.Y(_10362_),
    .A(net6546),
    .B(net6056));
 sg13g2_a21oi_1 _14968_ (.A1(_10361_),
    .A2(_10362_),
    .Y(_10363_),
    .B1(_10298_));
 sg13g2_nand2b_1 _14969_ (.Y(_10364_),
    .B(net6104),
    .A_N(\soc_inst.mem_ctrl.spi_data_out[10] ));
 sg13g2_o21ai_1 _14970_ (.B1(_10364_),
    .Y(_10365_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .A2(_10327_));
 sg13g2_a22oi_1 _14971_ (.Y(_10366_),
    .B1(net6046),
    .B2(_10365_),
    .A2(net6107),
    .A1(_07952_));
 sg13g2_nand2_1 _14972_ (.Y(_10367_),
    .A(\soc_inst.gpio_inst.gpio_out[1] ),
    .B(net5363));
 sg13g2_nand2_1 _14973_ (.Y(_10368_),
    .A(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .B(net5530));
 sg13g2_a22oi_1 _14974_ (.Y(_10369_),
    .B1(net5337),
    .B2(net3),
    .A2(net5566),
    .A1(\soc_inst.gpio_inst.int_en_reg[2] ));
 sg13g2_nand3_1 _14975_ (.B(_10368_),
    .C(_10369_),
    .A(_10367_),
    .Y(_10370_));
 sg13g2_a221oi_1 _14976_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ),
    .C1(_10356_),
    .B1(net5336),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ),
    .Y(_10371_),
    .A2(net5566));
 sg13g2_nor2_1 _14977_ (.A(_10304_),
    .B(_10371_),
    .Y(_10372_));
 sg13g2_nor2_1 _14978_ (.A(_10310_),
    .B(_10352_),
    .Y(_10373_));
 sg13g2_nand2_1 _14979_ (.Y(_10374_),
    .A(net5128),
    .B(_10358_));
 sg13g2_a22oi_1 _14980_ (.Y(_10375_),
    .B1(_10275_),
    .B2(_10355_),
    .A2(net5530),
    .A1(_07797_));
 sg13g2_o21ai_1 _14981_ (.B1(_10374_),
    .Y(_10376_),
    .A1(_10284_),
    .A2(_10375_));
 sg13g2_or4_1 _14982_ (.A(_10363_),
    .B(_10372_),
    .C(_10373_),
    .D(_10376_),
    .X(_10377_));
 sg13g2_a21oi_2 _14983_ (.B1(_10377_),
    .Y(_10378_),
    .A2(_10370_),
    .A1(_10294_));
 sg13g2_a21oi_1 _14984_ (.A1(net5191),
    .A2(_10366_),
    .Y(_10379_),
    .B1(net5038));
 sg13g2_a22oi_1 _14985_ (.Y(_00607_),
    .B1(_10378_),
    .B2(_10379_),
    .A2(net5038),
    .A1(_08002_));
 sg13g2_nor2_1 _14986_ (.A(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .B(net6045),
    .Y(_10380_));
 sg13g2_nor2_1 _14987_ (.A(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .B(_10327_),
    .Y(_10381_));
 sg13g2_o21ai_1 _14988_ (.B1(net6046),
    .Y(_10382_),
    .A1(_10380_),
    .A2(_10381_));
 sg13g2_o21ai_1 _14989_ (.B1(_10382_),
    .Y(_10383_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .A2(net6106));
 sg13g2_a21oi_1 _14990_ (.A1(net5190),
    .A2(_10383_),
    .Y(_10384_),
    .B1(net5038));
 sg13g2_nand2b_1 _14991_ (.Y(_10385_),
    .B(net6544),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[27] ));
 sg13g2_o21ai_1 _14992_ (.B1(_10385_),
    .Y(_10386_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .A2(net6097));
 sg13g2_a21oi_1 _14993_ (.A1(_07935_),
    .A2(_09243_),
    .Y(_10387_),
    .B1(_10386_));
 sg13g2_nand2_1 _14994_ (.Y(_10388_),
    .A(net6206),
    .B(_07948_));
 sg13g2_a22oi_1 _14995_ (.Y(_10389_),
    .B1(_10388_),
    .B2(net6067),
    .A2(net5564),
    .A1(\soc_inst.pwm_inst.channel_duty[0][3] ));
 sg13g2_a21oi_1 _14996_ (.A1(_00237_),
    .A2(net5560),
    .Y(_10390_),
    .B1(_10389_));
 sg13g2_nor2_1 _14997_ (.A(_00286_),
    .B(net6050),
    .Y(_10391_));
 sg13g2_nor2_1 _14998_ (.A(_00270_),
    .B(net6063),
    .Y(_10392_));
 sg13g2_nor3_1 _14999_ (.A(net6108),
    .B(_10391_),
    .C(_10392_),
    .Y(_10393_));
 sg13g2_nor2_1 _15000_ (.A(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .B(net6048),
    .Y(_10394_));
 sg13g2_nor2_1 _15001_ (.A(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .B(_08792_),
    .Y(_10395_));
 sg13g2_nor3_1 _15002_ (.A(_10393_),
    .B(_10394_),
    .C(_10395_),
    .Y(_10396_));
 sg13g2_nand2_1 _15003_ (.Y(_10397_),
    .A(_00229_),
    .B(net6206));
 sg13g2_a22oi_1 _15004_ (.Y(_10398_),
    .B1(_10397_),
    .B2(net6067),
    .A2(net5563),
    .A1(\soc_inst.i2c_inst.data_reg[3] ));
 sg13g2_nor2_1 _15005_ (.A(\soc_inst.i2c_inst.status_reg[3] ),
    .B(net6049),
    .Y(_10399_));
 sg13g2_o21ai_1 _15006_ (.B1(_08792_),
    .Y(_10400_),
    .A1(_10398_),
    .A2(_10399_));
 sg13g2_a22oi_1 _15007_ (.Y(_10401_),
    .B1(net5530),
    .B2(\soc_inst.gpio_inst.int_pend_reg[3] ),
    .A2(net5567),
    .A1(\soc_inst.gpio_inst.int_en_reg[3] ));
 sg13g2_a21oi_1 _15008_ (.A1(net4),
    .A2(net5337),
    .Y(_10402_),
    .B1(net5363));
 sg13g2_a22oi_1 _15009_ (.Y(_10403_),
    .B1(_10401_),
    .B2(_10402_),
    .A2(net5362),
    .A1(_07956_));
 sg13g2_o21ai_1 _15010_ (.B1(_10400_),
    .Y(_10404_),
    .A1(\soc_inst.i2c_inst.ack_enable ),
    .A2(_08792_));
 sg13g2_nor2_1 _15011_ (.A(_10298_),
    .B(_10404_),
    .Y(_10405_));
 sg13g2_nor2_2 _15012_ (.A(_10276_),
    .B(_10304_),
    .Y(_10406_));
 sg13g2_a22oi_1 _15013_ (.Y(_10407_),
    .B1(_10406_),
    .B2(_07780_),
    .A2(_10403_),
    .A1(_10294_));
 sg13g2_and3_2 _15014_ (.X(_10408_),
    .A(net6212),
    .B(_09308_),
    .C(net5336));
 sg13g2_a221oi_1 _15015_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .C1(net5193),
    .B1(_10408_),
    .A1(_07796_),
    .Y(_10409_),
    .A2(_10325_));
 sg13g2_a21oi_1 _15016_ (.A1(net5128),
    .A2(_10390_),
    .Y(_10410_),
    .B1(_10405_));
 sg13g2_a22oi_1 _15017_ (.Y(_10411_),
    .B1(_10396_),
    .B2(net5127),
    .A2(_10387_),
    .A1(net5123));
 sg13g2_nand4_1 _15018_ (.B(_10409_),
    .C(_10410_),
    .A(_10407_),
    .Y(_10412_),
    .D(_10411_));
 sg13g2_a22oi_1 _15019_ (.Y(_10413_),
    .B1(_10384_),
    .B2(_10412_),
    .A2(net5040),
    .A1(net2462));
 sg13g2_inv_1 _15020_ (.Y(_00608_),
    .A(net2463));
 sg13g2_nor2_1 _15021_ (.A(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .B(net6045),
    .Y(_10414_));
 sg13g2_nor2_1 _15022_ (.A(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .B(_10327_),
    .Y(_10415_));
 sg13g2_o21ai_1 _15023_ (.B1(net6046),
    .Y(_10416_),
    .A1(_10414_),
    .A2(_10415_));
 sg13g2_o21ai_1 _15024_ (.B1(_10416_),
    .Y(_10417_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .A2(net6106));
 sg13g2_a21oi_1 _15025_ (.A1(net5190),
    .A2(_10417_),
    .Y(_10418_),
    .B1(net5042));
 sg13g2_a22oi_1 _15026_ (.Y(_10419_),
    .B1(_09424_),
    .B2(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .A2(net5567),
    .A1(\soc_inst.gpio_inst.int_en_reg[4] ));
 sg13g2_a21oi_1 _15027_ (.A1(net5),
    .A2(net5337),
    .Y(_10420_),
    .B1(net5363));
 sg13g2_a22oi_1 _15028_ (.Y(_10421_),
    .B1(_10419_),
    .B2(_10420_),
    .A2(net5362),
    .A1(_07958_));
 sg13g2_a22oi_1 _15029_ (.Y(_10422_),
    .B1(_10421_),
    .B2(_10294_),
    .A2(_10325_),
    .A1(_07795_));
 sg13g2_or2_1 _15030_ (.X(_10423_),
    .B(net6097),
    .A(\soc_inst.spi_inst.rx_shift_reg[4] ));
 sg13g2_o21ai_1 _15031_ (.B1(_10423_),
    .Y(_10424_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .A2(net6098));
 sg13g2_a21oi_1 _15032_ (.A1(_07940_),
    .A2(net6544),
    .Y(_10425_),
    .B1(_10424_));
 sg13g2_nand2_1 _15033_ (.Y(_10426_),
    .A(net6206),
    .B(_07947_));
 sg13g2_a22oi_1 _15034_ (.Y(_10427_),
    .B1(_10426_),
    .B2(net6067),
    .A2(net5564),
    .A1(\soc_inst.pwm_inst.channel_duty[0][4] ));
 sg13g2_a21oi_1 _15035_ (.A1(_00238_),
    .A2(net5559),
    .Y(_10428_),
    .B1(_10427_));
 sg13g2_a21oi_1 _15036_ (.A1(_07787_),
    .A2(net6068),
    .Y(_10429_),
    .B1(net6108));
 sg13g2_o21ai_1 _15037_ (.B1(_10429_),
    .Y(_10430_),
    .A1(_00287_),
    .A2(net6050));
 sg13g2_o21ai_1 _15038_ (.B1(_10430_),
    .Y(_10431_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .A2(net6048));
 sg13g2_a21oi_1 _15039_ (.A1(_07902_),
    .A2(net6056),
    .Y(_10432_),
    .B1(_10431_));
 sg13g2_nor2_1 _15040_ (.A(_00230_),
    .B(_08672_),
    .Y(_10433_));
 sg13g2_a221oi_1 _15041_ (.B2(\soc_inst.i2c_inst.data_reg[4] ),
    .C1(_10433_),
    .B1(net5563),
    .A1(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .Y(_10434_),
    .A2(net6056));
 sg13g2_a22oi_1 _15042_ (.Y(_10435_),
    .B1(_10432_),
    .B2(net5127),
    .A2(_10408_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ));
 sg13g2_nand2_1 _15043_ (.Y(_10436_),
    .A(net5128),
    .B(_10428_));
 sg13g2_o21ai_1 _15044_ (.B1(_10436_),
    .Y(_10437_),
    .A1(_10298_),
    .A2(_10434_));
 sg13g2_nor2_1 _15045_ (.A(net5193),
    .B(_10437_),
    .Y(_10438_));
 sg13g2_a22oi_1 _15046_ (.Y(_10439_),
    .B1(_10425_),
    .B2(net5123),
    .A2(_10406_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ));
 sg13g2_nand4_1 _15047_ (.B(_10435_),
    .C(_10438_),
    .A(_10422_),
    .Y(_10440_),
    .D(_10439_));
 sg13g2_a22oi_1 _15048_ (.Y(_10441_),
    .B1(_10418_),
    .B2(_10440_),
    .A2(net5042),
    .A1(net2636));
 sg13g2_inv_1 _15049_ (.Y(_00609_),
    .A(net2637));
 sg13g2_nand2_1 _15050_ (.Y(_10442_),
    .A(net315),
    .B(net5043));
 sg13g2_nand2b_1 _15051_ (.Y(_10443_),
    .B(net6104),
    .A_N(\soc_inst.mem_ctrl.spi_data_out[13] ));
 sg13g2_o21ai_1 _15052_ (.B1(_10443_),
    .Y(_10444_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .A2(_10327_));
 sg13g2_a22oi_1 _15053_ (.Y(_10445_),
    .B1(net6046),
    .B2(_10444_),
    .A2(net6107),
    .A1(_07953_));
 sg13g2_a22oi_1 _15054_ (.Y(_10446_),
    .B1(_09424_),
    .B2(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .A2(net5567),
    .A1(\soc_inst.gpio_inst.int_en_reg[5] ));
 sg13g2_a21oi_1 _15055_ (.A1(net6),
    .A2(net5337),
    .Y(_10447_),
    .B1(net5362));
 sg13g2_a22oi_1 _15056_ (.Y(_10448_),
    .B1(_10446_),
    .B2(_10447_),
    .A2(net5362),
    .A1(_07960_));
 sg13g2_or2_1 _15057_ (.X(_10449_),
    .B(net6050),
    .A(_00288_));
 sg13g2_o21ai_1 _15058_ (.B1(_10449_),
    .Y(_10450_),
    .A1(_00272_),
    .A2(_08672_));
 sg13g2_a221oi_1 _15059_ (.B2(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .C1(_10450_),
    .B1(net5560),
    .A1(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .Y(_10451_),
    .A2(net6056));
 sg13g2_inv_1 _15060_ (.Y(_10452_),
    .A(_10451_));
 sg13g2_nor2_1 _15061_ (.A(_08671_),
    .B(_10298_),
    .Y(_10453_));
 sg13g2_mux2_1 _15062_ (.A0(\soc_inst.i2c_inst.data_reg[5] ),
    .A1(\soc_inst.i2c_inst.prescale_reg[5] ),
    .S(net6211),
    .X(_10454_));
 sg13g2_nand2b_1 _15063_ (.Y(_10455_),
    .B(net6544),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[29] ));
 sg13g2_o21ai_1 _15064_ (.B1(_10455_),
    .Y(_10456_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .A2(net6097));
 sg13g2_a21oi_1 _15065_ (.A1(_07936_),
    .A2(_09243_),
    .Y(_10457_),
    .B1(_10456_));
 sg13g2_nand2_1 _15066_ (.Y(_10458_),
    .A(net6209),
    .B(_07946_));
 sg13g2_a22oi_1 _15067_ (.Y(_10459_),
    .B1(_10458_),
    .B2(net6066),
    .A2(net5562),
    .A1(\soc_inst.pwm_inst.channel_duty[0][5] ));
 sg13g2_a21oi_1 _15068_ (.A1(_00239_),
    .A2(net5559),
    .Y(_10460_),
    .B1(_10459_));
 sg13g2_a221oi_1 _15069_ (.B2(net5127),
    .C1(net5193),
    .B1(_10452_),
    .A1(_10294_),
    .Y(_10461_),
    .A2(_10448_));
 sg13g2_a22oi_1 _15070_ (.Y(_10462_),
    .B1(_10408_),
    .B2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ),
    .A2(_10406_),
    .A1(_07779_));
 sg13g2_a22oi_1 _15071_ (.Y(_10463_),
    .B1(_10457_),
    .B2(net5123),
    .A2(_10454_),
    .A1(_10453_));
 sg13g2_a22oi_1 _15072_ (.Y(_10464_),
    .B1(_10460_),
    .B2(net5128),
    .A2(_10325_),
    .A1(\soc_inst.spi_inst.clock_divider[5] ));
 sg13g2_nand4_1 _15073_ (.B(_10462_),
    .C(_10463_),
    .A(_10461_),
    .Y(_10465_),
    .D(_10464_));
 sg13g2_o21ai_1 _15074_ (.B1(_10465_),
    .Y(_10466_),
    .A1(_08240_),
    .A2(_10445_));
 sg13g2_o21ai_1 _15075_ (.B1(_10442_),
    .Y(_00610_),
    .A1(net5043),
    .A2(_10466_));
 sg13g2_nor2_1 _15076_ (.A(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .B(net6045),
    .Y(_10467_));
 sg13g2_nor2_1 _15077_ (.A(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .B(_10327_),
    .Y(_10468_));
 sg13g2_o21ai_1 _15078_ (.B1(net6046),
    .Y(_10469_),
    .A1(_10467_),
    .A2(_10468_));
 sg13g2_o21ai_1 _15079_ (.B1(_10469_),
    .Y(_10470_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .A2(net6106));
 sg13g2_a21oi_1 _15080_ (.A1(net5190),
    .A2(_10470_),
    .Y(_10471_),
    .B1(net5038));
 sg13g2_nor2_1 _15081_ (.A(_00289_),
    .B(net6050),
    .Y(_10472_));
 sg13g2_nor2_1 _15082_ (.A(_00273_),
    .B(net6063),
    .Y(_10473_));
 sg13g2_nor3_1 _15083_ (.A(net6108),
    .B(_10472_),
    .C(_10473_),
    .Y(_10474_));
 sg13g2_nor2_1 _15084_ (.A(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .B(net6048),
    .Y(_10475_));
 sg13g2_nor2_1 _15085_ (.A(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .B(_08792_),
    .Y(_10476_));
 sg13g2_nor3_1 _15086_ (.A(_10474_),
    .B(_10475_),
    .C(_10476_),
    .Y(_10477_));
 sg13g2_mux2_1 _15087_ (.A0(\soc_inst.i2c_inst.data_reg[6] ),
    .A1(\soc_inst.i2c_inst.prescale_reg[6] ),
    .S(net6211),
    .X(_10478_));
 sg13g2_a21oi_1 _15088_ (.A1(net7),
    .A2(net5337),
    .Y(_10479_),
    .B1(net5363));
 sg13g2_a22oi_1 _15089_ (.Y(_10480_),
    .B1(_09424_),
    .B2(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .A2(net5567),
    .A1(\soc_inst.gpio_inst.int_en_reg[6] ));
 sg13g2_a22oi_1 _15090_ (.Y(_10481_),
    .B1(_10479_),
    .B2(_10480_),
    .A2(net5362),
    .A1(_07961_));
 sg13g2_nand2b_1 _15091_ (.Y(_10482_),
    .B(net6544),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[30] ));
 sg13g2_o21ai_1 _15092_ (.B1(_10482_),
    .Y(_10483_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .A2(net6097));
 sg13g2_a21oi_1 _15093_ (.A1(_07937_),
    .A2(_09243_),
    .Y(_10484_),
    .B1(_10483_));
 sg13g2_nand2_1 _15094_ (.Y(_10485_),
    .A(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .B(net5562));
 sg13g2_o21ai_1 _15095_ (.B1(net6068),
    .Y(_10486_),
    .A1(_07888_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][6] ));
 sg13g2_a22oi_1 _15096_ (.Y(_10487_),
    .B1(_10485_),
    .B2(_10486_),
    .A2(net5558),
    .A1(_00240_));
 sg13g2_a22oi_1 _15097_ (.Y(_10488_),
    .B1(_10484_),
    .B2(net5123),
    .A2(_10478_),
    .A1(_10453_));
 sg13g2_a22oi_1 _15098_ (.Y(_10489_),
    .B1(_10477_),
    .B2(net5127),
    .A2(_10325_),
    .A1(\soc_inst.spi_inst.clock_divider[6] ));
 sg13g2_a22oi_1 _15099_ (.Y(_10490_),
    .B1(_10481_),
    .B2(_10294_),
    .A2(_10408_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ));
 sg13g2_a221oi_1 _15100_ (.B2(net5129),
    .C1(net5193),
    .B1(_10487_),
    .A1(net6175),
    .Y(_10491_),
    .A2(_10406_));
 sg13g2_nand4_1 _15101_ (.B(_10489_),
    .C(_10490_),
    .A(_10488_),
    .Y(_10492_),
    .D(_10491_));
 sg13g2_a22oi_1 _15102_ (.Y(_10493_),
    .B1(_10471_),
    .B2(_10492_),
    .A2(net5040),
    .A1(net2353));
 sg13g2_inv_1 _15103_ (.Y(_00611_),
    .A(net2354));
 sg13g2_nor2_1 _15104_ (.A(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .B(net6045),
    .Y(_10494_));
 sg13g2_nor2_1 _15105_ (.A(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .B(_10327_),
    .Y(_10495_));
 sg13g2_o21ai_1 _15106_ (.B1(net6046),
    .Y(_10496_),
    .A1(_10494_),
    .A2(_10495_));
 sg13g2_o21ai_1 _15107_ (.B1(_10496_),
    .Y(_10497_),
    .A1(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .A2(net6106));
 sg13g2_nor2b_1 _15108_ (.A(net6211),
    .B_N(\soc_inst.i2c_inst.data_reg[7] ),
    .Y(_10498_));
 sg13g2_nor2_1 _15109_ (.A(_00231_),
    .B(_07887_),
    .Y(_10499_));
 sg13g2_o21ai_1 _15110_ (.B1(_10453_),
    .Y(_10500_),
    .A1(_10498_),
    .A2(_10499_));
 sg13g2_nand2b_1 _15111_ (.Y(_10501_),
    .B(net6544),
    .A_N(\soc_inst.spi_inst.rx_shift_reg[31] ));
 sg13g2_o21ai_1 _15112_ (.B1(_10501_),
    .Y(_10502_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .A2(net6097));
 sg13g2_a21oi_1 _15113_ (.A1(_07938_),
    .A2(_09243_),
    .Y(_10503_),
    .B1(_10502_));
 sg13g2_nand2_1 _15114_ (.Y(_10504_),
    .A(\soc_inst.pwm_inst.channel_duty[0][7] ),
    .B(net5564));
 sg13g2_o21ai_1 _15115_ (.B1(net6066),
    .Y(_10505_),
    .A1(_07888_),
    .A2(\soc_inst.pwm_inst.channel_counter[0][7] ));
 sg13g2_a22oi_1 _15116_ (.Y(_10506_),
    .B1(_10504_),
    .B2(_10505_),
    .A2(net5559),
    .A1(_00241_));
 sg13g2_a221oi_1 _15117_ (.B2(_07783_),
    .C1(net6108),
    .B1(net5562),
    .A1(_07786_),
    .Y(_10507_),
    .A2(net6066));
 sg13g2_a221oi_1 _15118_ (.B2(_07905_),
    .C1(_10507_),
    .B1(net5557),
    .A1(_07901_),
    .Y(_10508_),
    .A2(net6061));
 sg13g2_a22oi_1 _15119_ (.Y(_10509_),
    .B1(_10506_),
    .B2(net5129),
    .A2(_10325_),
    .A1(\soc_inst.spi_inst.clock_divider[7] ));
 sg13g2_nand2_1 _15120_ (.Y(_10510_),
    .A(_10500_),
    .B(_10509_));
 sg13g2_a22oi_1 _15121_ (.Y(_10511_),
    .B1(_10503_),
    .B2(net5123),
    .A2(_10406_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ));
 sg13g2_a22oi_1 _15122_ (.Y(_10512_),
    .B1(_10508_),
    .B2(net5127),
    .A2(_10408_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ));
 sg13g2_nand2_1 _15123_ (.Y(_10513_),
    .A(_10511_),
    .B(_10512_));
 sg13g2_nor3_2 _15124_ (.A(net5193),
    .B(_10510_),
    .C(_10513_),
    .Y(_10514_));
 sg13g2_a21oi_1 _15125_ (.A1(net5191),
    .A2(_10497_),
    .Y(_10515_),
    .B1(_10514_));
 sg13g2_mux2_1 _15126_ (.A0(_10515_),
    .A1(net2589),
    .S(net5042),
    .X(_00612_));
 sg13g2_a22oi_1 _15127_ (.Y(_10516_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .A1(net6297));
 sg13g2_a221oi_1 _15128_ (.B2(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .C1(net5558),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .Y(_10517_),
    .A2(net6065));
 sg13g2_a21oi_2 _15129_ (.B1(_10517_),
    .Y(_10518_),
    .A2(net5558),
    .A1(_00242_));
 sg13g2_a21o_1 _15130_ (.A2(net6207),
    .A1(_00275_),
    .B1(net6062),
    .X(_10519_));
 sg13g2_o21ai_1 _15131_ (.B1(_10519_),
    .Y(_10520_),
    .A1(_00291_),
    .A2(net6051));
 sg13g2_o21ai_1 _15132_ (.B1(_10520_),
    .Y(_10521_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .A2(net6047));
 sg13g2_nand2_1 _15133_ (.Y(_10522_),
    .A(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .B(net6056));
 sg13g2_and2_1 _15134_ (.A(net6544),
    .B(net5123),
    .X(_10523_));
 sg13g2_and2_1 _15135_ (.A(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .B(_09243_),
    .X(_10524_));
 sg13g2_a21oi_1 _15136_ (.A1(_10521_),
    .A2(_10522_),
    .Y(_10525_),
    .B1(_10310_));
 sg13g2_a221oi_1 _15137_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .C1(_10525_),
    .B1(_10406_),
    .A1(\soc_inst.spi_inst.cpha ),
    .Y(_10526_),
    .A2(_10325_));
 sg13g2_a22oi_1 _15138_ (.Y(_10527_),
    .B1(_10524_),
    .B2(net5123),
    .A2(_10518_),
    .A1(net5129));
 sg13g2_nand2b_1 _15139_ (.Y(_10528_),
    .B(_10527_),
    .A_N(net5193));
 sg13g2_a21oi_1 _15140_ (.A1(net1557),
    .A2(net5061),
    .Y(_10529_),
    .B1(_10528_));
 sg13g2_a221oi_1 _15141_ (.B2(_10529_),
    .C1(net5041),
    .B1(_10526_),
    .A1(net5188),
    .Y(_10530_),
    .A2(_10516_));
 sg13g2_a21o_1 _15142_ (.A2(net5042),
    .A1(net2137),
    .B1(_10530_),
    .X(_00613_));
 sg13g2_a22oi_1 _15143_ (.Y(_10531_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .A1(net6298));
 sg13g2_a21o_1 _15144_ (.A2(net6207),
    .A1(_00276_),
    .B1(net6062),
    .X(_10532_));
 sg13g2_o21ai_1 _15145_ (.B1(_10532_),
    .Y(_10533_),
    .A1(_00292_),
    .A2(net6051));
 sg13g2_nand2b_1 _15146_ (.Y(_10534_),
    .B(net6108),
    .A_N(\soc_inst.cpu_core.csr_file.mtime[41] ));
 sg13g2_a22oi_1 _15147_ (.Y(_10535_),
    .B1(_10533_),
    .B2(_10534_),
    .A2(net6061),
    .A1(\soc_inst.cpu_core.csr_file.mtime[9] ));
 sg13g2_a221oi_1 _15148_ (.B2(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .C1(net5556),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .Y(_10536_),
    .A2(net6065));
 sg13g2_a21oi_2 _15149_ (.B1(_10536_),
    .Y(_10537_),
    .A2(net5557),
    .A1(_00243_));
 sg13g2_nand3_1 _15150_ (.B(_09243_),
    .C(_10321_),
    .A(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .Y(_10538_));
 sg13g2_nor2_1 _15151_ (.A(_10310_),
    .B(_10535_),
    .Y(_10539_));
 sg13g2_a221oi_1 _15152_ (.B2(_07778_),
    .C1(_10539_),
    .B1(_10406_),
    .A1(\soc_inst.spi_inst.cpol ),
    .Y(_10540_),
    .A2(_10325_));
 sg13g2_a221oi_1 _15153_ (.B2(net5129),
    .C1(net5193),
    .B1(_10537_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .Y(_10541_),
    .A2(net5061));
 sg13g2_and2_1 _15154_ (.A(_10538_),
    .B(_10541_),
    .X(_10542_));
 sg13g2_a22oi_1 _15155_ (.Y(_10543_),
    .B1(_10540_),
    .B2(_10542_),
    .A2(_10531_),
    .A1(net5188));
 sg13g2_mux2_1 _15156_ (.A0(_10543_),
    .A1(net2344),
    .S(net5042),
    .X(_00614_));
 sg13g2_a22oi_1 _15157_ (.Y(_10544_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .B2(net6104),
    .A2(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .A1(net6296));
 sg13g2_a21o_1 _15158_ (.A2(net6208),
    .A1(_00277_),
    .B1(net6062),
    .X(_10545_));
 sg13g2_o21ai_1 _15159_ (.B1(_10545_),
    .Y(_10546_),
    .A1(_00293_),
    .A2(net6055));
 sg13g2_o21ai_1 _15160_ (.B1(_10546_),
    .Y(_10547_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .A2(net6047));
 sg13g2_nand2_1 _15161_ (.Y(_10548_),
    .A(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .B(net6060));
 sg13g2_nand2_1 _15162_ (.Y(_10549_),
    .A(_10547_),
    .B(_10548_));
 sg13g2_a221oi_1 _15163_ (.B2(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .C1(net5558),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .Y(_10550_),
    .A2(net6065));
 sg13g2_a21oi_1 _15164_ (.A1(_00244_),
    .A2(net5556),
    .Y(_10551_),
    .B1(_10550_));
 sg13g2_mux2_1 _15165_ (.A0(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .S(net6098),
    .X(_10552_));
 sg13g2_nand2_1 _15166_ (.Y(_10553_),
    .A(_10322_),
    .B(_10552_));
 sg13g2_o21ai_1 _15167_ (.B1(_10553_),
    .Y(_10554_),
    .A1(net5197),
    .A2(_10544_));
 sg13g2_a221oi_1 _15168_ (.B2(net5129),
    .C1(_10554_),
    .B1(_10551_),
    .A1(net5126),
    .Y(_10555_),
    .A2(_10549_));
 sg13g2_nand2_1 _15169_ (.Y(_10556_),
    .A(net1165),
    .B(net5035));
 sg13g2_o21ai_1 _15170_ (.B1(_10556_),
    .Y(_00615_),
    .A1(net5035),
    .A2(_10555_));
 sg13g2_a22oi_1 _15171_ (.Y(_10557_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .A1(net6297));
 sg13g2_a21o_1 _15172_ (.A2(net6207),
    .A1(_00278_),
    .B1(net6062),
    .X(_10558_));
 sg13g2_o21ai_1 _15173_ (.B1(_10558_),
    .Y(_10559_),
    .A1(_00294_),
    .A2(net6055));
 sg13g2_o21ai_1 _15174_ (.B1(_10559_),
    .Y(_10560_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .A2(net6047));
 sg13g2_nand2_1 _15175_ (.Y(_10561_),
    .A(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .B(net6060));
 sg13g2_nand2_1 _15176_ (.Y(_10562_),
    .A(_10560_),
    .B(_10561_));
 sg13g2_a221oi_1 _15177_ (.B2(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .C1(net5558),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .Y(_10563_),
    .A2(net6065));
 sg13g2_a21oi_1 _15178_ (.A1(_00245_),
    .A2(net5556),
    .Y(_10564_),
    .B1(_10563_));
 sg13g2_mux2_1 _15179_ (.A0(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .S(net6098),
    .X(_10565_));
 sg13g2_nand2_1 _15180_ (.Y(_10566_),
    .A(_10322_),
    .B(_10565_));
 sg13g2_o21ai_1 _15181_ (.B1(_10566_),
    .Y(_10567_),
    .A1(net5197),
    .A2(_10557_));
 sg13g2_a221oi_1 _15182_ (.B2(net5129),
    .C1(_10567_),
    .B1(_10564_),
    .A1(net5126),
    .Y(_10568_),
    .A2(_10562_));
 sg13g2_nand2_1 _15183_ (.Y(_10569_),
    .A(net1310),
    .B(net5037));
 sg13g2_o21ai_1 _15184_ (.B1(_10569_),
    .Y(_00616_),
    .A1(net5037),
    .A2(_10568_));
 sg13g2_a22oi_1 _15185_ (.Y(_10570_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .A1(net6297));
 sg13g2_a21o_1 _15186_ (.A2(net6207),
    .A1(_00279_),
    .B1(net6062),
    .X(_10571_));
 sg13g2_o21ai_1 _15187_ (.B1(_10571_),
    .Y(_10572_),
    .A1(_00295_),
    .A2(net6055));
 sg13g2_o21ai_1 _15188_ (.B1(_10572_),
    .Y(_10573_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .A2(net6047));
 sg13g2_nand2_1 _15189_ (.Y(_10574_),
    .A(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .B(net6060));
 sg13g2_nand2_1 _15190_ (.Y(_10575_),
    .A(_10573_),
    .B(_10574_));
 sg13g2_nand2_1 _15191_ (.Y(_10576_),
    .A(net6207),
    .B(_07942_));
 sg13g2_a22oi_1 _15192_ (.Y(_10577_),
    .B1(_10576_),
    .B2(net6065),
    .A2(net5561),
    .A1(\soc_inst.pwm_inst.channel_duty[0][12] ));
 sg13g2_a21oi_1 _15193_ (.A1(_00246_),
    .A2(net5556),
    .Y(_10578_),
    .B1(_10577_));
 sg13g2_mux2_1 _15194_ (.A0(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .S(net6098),
    .X(_10579_));
 sg13g2_nand2_1 _15195_ (.Y(_10580_),
    .A(_10322_),
    .B(_10579_));
 sg13g2_o21ai_1 _15196_ (.B1(_10580_),
    .Y(_10581_),
    .A1(net5197),
    .A2(_10570_));
 sg13g2_a221oi_1 _15197_ (.B2(net5129),
    .C1(_10581_),
    .B1(_10578_),
    .A1(net5126),
    .Y(_10582_),
    .A2(_10575_));
 sg13g2_nand2_1 _15198_ (.Y(_10583_),
    .A(net773),
    .B(net5037));
 sg13g2_o21ai_1 _15199_ (.B1(_10583_),
    .Y(_00617_),
    .A1(net5037),
    .A2(_10582_));
 sg13g2_a22oi_1 _15200_ (.Y(_10584_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .A1(net6297));
 sg13g2_a21o_1 _15201_ (.A2(net6207),
    .A1(_00280_),
    .B1(net6062),
    .X(_10585_));
 sg13g2_o21ai_1 _15202_ (.B1(_10585_),
    .Y(_10586_),
    .A1(_00296_),
    .A2(net6055));
 sg13g2_o21ai_1 _15203_ (.B1(_10586_),
    .Y(_10587_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .A2(net6047));
 sg13g2_nand2_1 _15204_ (.Y(_10588_),
    .A(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .B(net6060));
 sg13g2_nand2_1 _15205_ (.Y(_10589_),
    .A(_10587_),
    .B(_10588_));
 sg13g2_a221oi_1 _15206_ (.B2(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .C1(net5558),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .Y(_10590_),
    .A2(net6065));
 sg13g2_a21oi_1 _15207_ (.A1(_00247_),
    .A2(net5556),
    .Y(_10591_),
    .B1(_10590_));
 sg13g2_mux2_1 _15208_ (.A0(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .S(net6098),
    .X(_10592_));
 sg13g2_nand2_1 _15209_ (.Y(_10593_),
    .A(_10322_),
    .B(_10592_));
 sg13g2_o21ai_1 _15210_ (.B1(_10593_),
    .Y(_10594_),
    .A1(net5197),
    .A2(_10584_));
 sg13g2_a221oi_1 _15211_ (.B2(_10307_),
    .C1(_10594_),
    .B1(_10591_),
    .A1(net5126),
    .Y(_10595_),
    .A2(_10589_));
 sg13g2_nand2_1 _15212_ (.Y(_10596_),
    .A(net683),
    .B(net5044));
 sg13g2_o21ai_1 _15213_ (.B1(_10596_),
    .Y(_00618_),
    .A1(net5035),
    .A2(_10595_));
 sg13g2_a22oi_1 _15214_ (.Y(_10597_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .B2(net6104),
    .A2(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .A1(net6299));
 sg13g2_a21o_1 _15215_ (.A2(net6207),
    .A1(_00281_),
    .B1(net6062),
    .X(_10598_));
 sg13g2_o21ai_1 _15216_ (.B1(_10598_),
    .Y(_10599_),
    .A1(_00297_),
    .A2(net6055));
 sg13g2_o21ai_1 _15217_ (.B1(_10599_),
    .Y(_10600_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .A2(net6047));
 sg13g2_nand2_1 _15218_ (.Y(_10601_),
    .A(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .B(net6060));
 sg13g2_nand2_1 _15219_ (.Y(_10602_),
    .A(_10600_),
    .B(_10601_));
 sg13g2_a221oi_1 _15220_ (.B2(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .C1(net5556),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .Y(_10603_),
    .A2(net6065));
 sg13g2_a21oi_1 _15221_ (.A1(_00248_),
    .A2(net5556),
    .Y(_10604_),
    .B1(_10603_));
 sg13g2_mux2_1 _15222_ (.A0(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .S(net6098),
    .X(_10605_));
 sg13g2_nand2_1 _15223_ (.Y(_10606_),
    .A(_10322_),
    .B(_10605_));
 sg13g2_o21ai_1 _15224_ (.B1(_10606_),
    .Y(_10607_),
    .A1(net5197),
    .A2(_10597_));
 sg13g2_a221oi_1 _15225_ (.B2(_10307_),
    .C1(_10607_),
    .B1(_10604_),
    .A1(net5126),
    .Y(_10608_),
    .A2(_10602_));
 sg13g2_nand2_1 _15226_ (.Y(_10609_),
    .A(net981),
    .B(net5044));
 sg13g2_o21ai_1 _15227_ (.B1(_10609_),
    .Y(_00619_),
    .A1(net5036),
    .A2(_10608_));
 sg13g2_a22oi_1 _15228_ (.Y(_10610_),
    .B1(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .B2(net6103),
    .A2(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .A1(net6297));
 sg13g2_a21o_1 _15229_ (.A2(net6207),
    .A1(_00282_),
    .B1(net6062),
    .X(_10611_));
 sg13g2_o21ai_1 _15230_ (.B1(_10611_),
    .Y(_10612_),
    .A1(_00298_),
    .A2(net6055));
 sg13g2_o21ai_1 _15231_ (.B1(_10612_),
    .Y(_10613_),
    .A1(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .A2(net6047));
 sg13g2_nand2_1 _15232_ (.Y(_10614_),
    .A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .B(net6060));
 sg13g2_nand2_1 _15233_ (.Y(_10615_),
    .A(_10613_),
    .B(_10614_));
 sg13g2_a221oi_1 _15234_ (.B2(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .C1(net5556),
    .B1(net5561),
    .A1(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .Y(_10616_),
    .A2(net6065));
 sg13g2_a21oi_1 _15235_ (.A1(_00249_),
    .A2(net5557),
    .Y(_10617_),
    .B1(_10616_));
 sg13g2_mux2_1 _15236_ (.A0(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .A1(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .S(net6098),
    .X(_10618_));
 sg13g2_nand2_1 _15237_ (.Y(_10619_),
    .A(_10322_),
    .B(_10618_));
 sg13g2_o21ai_1 _15238_ (.B1(_10619_),
    .Y(_10620_),
    .A1(net5197),
    .A2(_10610_));
 sg13g2_a221oi_1 _15239_ (.B2(_10307_),
    .C1(_10620_),
    .B1(_10617_),
    .A1(net5126),
    .Y(_10621_),
    .A2(_10615_));
 sg13g2_nand2_1 _15240_ (.Y(_10622_),
    .A(net1556),
    .B(net5044));
 sg13g2_o21ai_1 _15241_ (.B1(_10622_),
    .Y(_00620_),
    .A1(net5035),
    .A2(_10621_));
 sg13g2_nand2_1 _15242_ (.Y(_10623_),
    .A(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .B(net6057));
 sg13g2_o21ai_1 _15243_ (.B1(_10623_),
    .Y(_10624_),
    .A1(_00299_),
    .A2(net6052));
 sg13g2_a21oi_1 _15244_ (.A1(net6298),
    .A2(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .Y(_10625_),
    .B1(net5196));
 sg13g2_a221oi_1 _15245_ (.B2(net5125),
    .C1(net5189),
    .B1(_10624_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .Y(_10626_),
    .A2(net5059));
 sg13g2_nor3_1 _15246_ (.A(net5036),
    .B(_10625_),
    .C(_10626_),
    .Y(_10627_));
 sg13g2_a21o_1 _15247_ (.A2(net5035),
    .A1(net1998),
    .B1(_10627_),
    .X(_00621_));
 sg13g2_nand2_1 _15248_ (.Y(_10628_),
    .A(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .B(net6057));
 sg13g2_o21ai_1 _15249_ (.B1(_10628_),
    .Y(_10629_),
    .A1(_00300_),
    .A2(net6052));
 sg13g2_a21oi_1 _15250_ (.A1(net6298),
    .A2(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .Y(_10630_),
    .B1(net5196));
 sg13g2_a221oi_1 _15251_ (.B2(net5125),
    .C1(net5189),
    .B1(_10629_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .Y(_10631_),
    .A2(net5059));
 sg13g2_nor3_1 _15252_ (.A(net5036),
    .B(_10630_),
    .C(_10631_),
    .Y(_10632_));
 sg13g2_a21o_1 _15253_ (.A2(net5035),
    .A1(net2204),
    .B1(_10632_),
    .X(_00622_));
 sg13g2_nand2_1 _15254_ (.Y(_10633_),
    .A(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .B(net6057));
 sg13g2_o21ai_1 _15255_ (.B1(_10633_),
    .Y(_10634_),
    .A1(_00301_),
    .A2(net6052));
 sg13g2_a21oi_1 _15256_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .Y(_10635_),
    .B1(net5196));
 sg13g2_a221oi_1 _15257_ (.B2(net5125),
    .C1(net5189),
    .B1(_10634_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .Y(_10636_),
    .A2(net5059));
 sg13g2_nor3_1 _15258_ (.A(net5036),
    .B(_10635_),
    .C(_10636_),
    .Y(_10637_));
 sg13g2_a21o_1 _15259_ (.A2(net5044),
    .A1(net2212),
    .B1(_10637_),
    .X(_00623_));
 sg13g2_nand2_1 _15260_ (.Y(_10638_),
    .A(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .B(net6057));
 sg13g2_o21ai_1 _15261_ (.B1(_10638_),
    .Y(_10639_),
    .A1(_00302_),
    .A2(net6052));
 sg13g2_a21oi_1 _15262_ (.A1(net6298),
    .A2(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .Y(_10640_),
    .B1(net5196));
 sg13g2_a221oi_1 _15263_ (.B2(net5125),
    .C1(net5189),
    .B1(_10639_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .Y(_10641_),
    .A2(net5059));
 sg13g2_nor3_1 _15264_ (.A(net5036),
    .B(_10640_),
    .C(_10641_),
    .Y(_10642_));
 sg13g2_a21o_1 _15265_ (.A2(net5035),
    .A1(net2190),
    .B1(_10642_),
    .X(_00624_));
 sg13g2_nand2_1 _15266_ (.Y(_10643_),
    .A(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .B(net6057));
 sg13g2_o21ai_1 _15267_ (.B1(_10643_),
    .Y(_10644_),
    .A1(_00303_),
    .A2(net6052));
 sg13g2_a21oi_1 _15268_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .Y(_10645_),
    .B1(net5195));
 sg13g2_a221oi_1 _15269_ (.B2(net5124),
    .C1(net5189),
    .B1(_10644_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .Y(_10646_),
    .A2(net5059));
 sg13g2_nor3_1 _15270_ (.A(net5039),
    .B(_10645_),
    .C(_10646_),
    .Y(_10647_));
 sg13g2_a21o_1 _15271_ (.A2(net5042),
    .A1(net1380),
    .B1(_10647_),
    .X(_00625_));
 sg13g2_nand2_1 _15272_ (.Y(_10648_),
    .A(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .B(net6057));
 sg13g2_o21ai_1 _15273_ (.B1(_10648_),
    .Y(_10649_),
    .A1(_00304_),
    .A2(net6052));
 sg13g2_a21oi_1 _15274_ (.A1(net6300),
    .A2(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .Y(_10650_),
    .B1(net5195));
 sg13g2_a221oi_1 _15275_ (.B2(net5124),
    .C1(net5189),
    .B1(_10649_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .Y(_10651_),
    .A2(net5059));
 sg13g2_nor3_1 _15276_ (.A(net5042),
    .B(_10650_),
    .C(_10651_),
    .Y(_10652_));
 sg13g2_a21o_1 _15277_ (.A2(net5043),
    .A1(net1020),
    .B1(_10652_),
    .X(_00626_));
 sg13g2_nand2_1 _15278_ (.Y(_10653_),
    .A(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .B(net6057));
 sg13g2_o21ai_1 _15279_ (.B1(_10653_),
    .Y(_10654_),
    .A1(_00305_),
    .A2(net6052));
 sg13g2_a21oi_1 _15280_ (.A1(net6300),
    .A2(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .Y(_10655_),
    .B1(net5196));
 sg13g2_a221oi_1 _15281_ (.B2(net5125),
    .C1(net5189),
    .B1(_10654_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .Y(_10656_),
    .A2(net5059));
 sg13g2_nor3_1 _15282_ (.A(net5036),
    .B(_10655_),
    .C(_10656_),
    .Y(_10657_));
 sg13g2_a21o_1 _15283_ (.A2(net5035),
    .A1(net2060),
    .B1(_10657_),
    .X(_00627_));
 sg13g2_nand2_1 _15284_ (.Y(_10658_),
    .A(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .B(net6057));
 sg13g2_o21ai_1 _15285_ (.B1(_10658_),
    .Y(_10659_),
    .A1(_00306_),
    .A2(net6052));
 sg13g2_a21oi_1 _15286_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .Y(_10660_),
    .B1(net5195));
 sg13g2_a221oi_1 _15287_ (.B2(net5124),
    .C1(net5189),
    .B1(_10659_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .Y(_10661_),
    .A2(net5059));
 sg13g2_nor3_1 _15288_ (.A(net5039),
    .B(_10660_),
    .C(_10661_),
    .Y(_10662_));
 sg13g2_a21o_1 _15289_ (.A2(net5043),
    .A1(net1188),
    .B1(_10662_),
    .X(_00628_));
 sg13g2_nand2_1 _15290_ (.Y(_10663_),
    .A(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .B(net6058));
 sg13g2_o21ai_1 _15291_ (.B1(_10663_),
    .Y(_10664_),
    .A1(_00307_),
    .A2(net6053));
 sg13g2_a21oi_1 _15292_ (.A1(net6297),
    .A2(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .Y(_10665_),
    .B1(net5194));
 sg13g2_a221oi_1 _15293_ (.B2(net5124),
    .C1(net5188),
    .B1(_10664_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .Y(_10666_),
    .A2(net5060));
 sg13g2_nor3_1 _15294_ (.A(net5039),
    .B(_10665_),
    .C(_10666_),
    .Y(_10667_));
 sg13g2_a21o_1 _15295_ (.A2(net5038),
    .A1(net1224),
    .B1(_10667_),
    .X(_00629_));
 sg13g2_nand2_1 _15296_ (.Y(_10668_),
    .A(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .B(net6058));
 sg13g2_o21ai_1 _15297_ (.B1(_10668_),
    .Y(_10669_),
    .A1(_00308_),
    .A2(net6053));
 sg13g2_a21oi_1 _15298_ (.A1(net6298),
    .A2(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .Y(_10670_),
    .B1(net5196));
 sg13g2_a221oi_1 _15299_ (.B2(net5125),
    .C1(net5188),
    .B1(_10669_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .Y(_10671_),
    .A2(net5060));
 sg13g2_nor3_1 _15300_ (.A(net5040),
    .B(_10670_),
    .C(_10671_),
    .Y(_10672_));
 sg13g2_a21o_1 _15301_ (.A2(net5036),
    .A1(net1958),
    .B1(_10672_),
    .X(_00630_));
 sg13g2_nand2_1 _15302_ (.Y(_10673_),
    .A(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .B(net6058));
 sg13g2_o21ai_1 _15303_ (.B1(_10673_),
    .Y(_10674_),
    .A1(_00309_),
    .A2(net6053));
 sg13g2_a21oi_1 _15304_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .Y(_10675_),
    .B1(net5195));
 sg13g2_a221oi_1 _15305_ (.B2(net5126),
    .C1(net5191),
    .B1(_10674_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .Y(_10676_),
    .A2(net5061));
 sg13g2_nor3_1 _15306_ (.A(net5039),
    .B(_10675_),
    .C(_10676_),
    .Y(_10677_));
 sg13g2_a21o_1 _15307_ (.A2(net5040),
    .A1(net2333),
    .B1(_10677_),
    .X(_00631_));
 sg13g2_nand2_1 _15308_ (.Y(_10678_),
    .A(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .B(net6058));
 sg13g2_o21ai_1 _15309_ (.B1(_10678_),
    .Y(_10679_),
    .A1(_00310_),
    .A2(net6053));
 sg13g2_a21oi_1 _15310_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .Y(_10680_),
    .B1(net5194));
 sg13g2_a221oi_1 _15311_ (.B2(net5125),
    .C1(net5188),
    .B1(_10679_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .Y(_10681_),
    .A2(net5060));
 sg13g2_nor3_1 _15312_ (.A(net5039),
    .B(_10680_),
    .C(_10681_),
    .Y(_10682_));
 sg13g2_a21o_1 _15313_ (.A2(net5038),
    .A1(net2379),
    .B1(_10682_),
    .X(_00632_));
 sg13g2_nand2_1 _15314_ (.Y(_10683_),
    .A(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .B(net6058));
 sg13g2_o21ai_1 _15315_ (.B1(_10683_),
    .Y(_10684_),
    .A1(_00311_),
    .A2(net6053));
 sg13g2_a21oi_1 _15316_ (.A1(net6297),
    .A2(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .Y(_10685_),
    .B1(net5196));
 sg13g2_a221oi_1 _15317_ (.B2(net5124),
    .C1(net5188),
    .B1(_10684_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .Y(_10686_),
    .A2(net5060));
 sg13g2_nor3_1 _15318_ (.A(net5041),
    .B(_10685_),
    .C(_10686_),
    .Y(_10687_));
 sg13g2_a21o_1 _15319_ (.A2(net5040),
    .A1(net2315),
    .B1(_10687_),
    .X(_00633_));
 sg13g2_nand2_1 _15320_ (.Y(_10688_),
    .A(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .B(net6059));
 sg13g2_o21ai_1 _15321_ (.B1(_10688_),
    .Y(_10689_),
    .A1(_00312_),
    .A2(net6054));
 sg13g2_a21oi_1 _15322_ (.A1(net6296),
    .A2(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .Y(_10690_),
    .B1(net5194));
 sg13g2_a221oi_1 _15323_ (.B2(net5124),
    .C1(net5192),
    .B1(_10689_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .Y(_10691_),
    .A2(net5060));
 sg13g2_nor3_1 _15324_ (.A(net5039),
    .B(_10690_),
    .C(_10691_),
    .Y(_10692_));
 sg13g2_a21o_1 _15325_ (.A2(net5043),
    .A1(net1148),
    .B1(_10692_),
    .X(_00634_));
 sg13g2_nand2_1 _15326_ (.Y(_10693_),
    .A(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .B(net6059));
 sg13g2_o21ai_1 _15327_ (.B1(_10693_),
    .Y(_10694_),
    .A1(_00313_),
    .A2(net6054));
 sg13g2_a21oi_1 _15328_ (.A1(net6299),
    .A2(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .Y(_10695_),
    .B1(net5194));
 sg13g2_a221oi_1 _15329_ (.B2(net5124),
    .C1(net5192),
    .B1(_10694_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .Y(_10696_),
    .A2(net5060));
 sg13g2_nor3_1 _15330_ (.A(net5039),
    .B(_10695_),
    .C(_10696_),
    .Y(_10697_));
 sg13g2_a21o_1 _15331_ (.A2(net5042),
    .A1(net1508),
    .B1(_10697_),
    .X(_00635_));
 sg13g2_nand2_1 _15332_ (.Y(_10698_),
    .A(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .B(net6059));
 sg13g2_o21ai_1 _15333_ (.B1(_10698_),
    .Y(_10699_),
    .A1(_00314_),
    .A2(net6054));
 sg13g2_a21oi_1 _15334_ (.A1(net6297),
    .A2(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .Y(_10700_),
    .B1(net5194));
 sg13g2_a221oi_1 _15335_ (.B2(net5124),
    .C1(net5192),
    .B1(_10699_),
    .A1(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .Y(_10701_),
    .A2(net5060));
 sg13g2_nor3_1 _15336_ (.A(net5041),
    .B(_10700_),
    .C(_10701_),
    .Y(_10702_));
 sg13g2_a21o_1 _15337_ (.A2(net5043),
    .A1(net1119),
    .B1(_10702_),
    .X(_00636_));
 sg13g2_nor2_1 _15338_ (.A(net6193),
    .B(net6179),
    .Y(_10703_));
 sg13g2_nand2_1 _15339_ (.Y(_10704_),
    .A(_00266_),
    .B(_10703_));
 sg13g2_a21oi_1 _15340_ (.A1(_08398_),
    .A2(_10704_),
    .Y(_10705_),
    .B1(_08247_));
 sg13g2_nand3b_1 _15341_ (.B(net6193),
    .C(_08248_),
    .Y(_10706_),
    .A_N(_08384_));
 sg13g2_nor3_1 _15342_ (.A(net5197),
    .B(_08392_),
    .C(_10705_),
    .Y(_10707_));
 sg13g2_nand2_1 _15343_ (.Y(_10708_),
    .A(_10706_),
    .B(_10707_));
 sg13g2_o21ai_1 _15344_ (.B1(\soc_inst.core_mem_re ),
    .Y(_10709_),
    .A1(net6504),
    .A2(net6193));
 sg13g2_nand2_1 _15345_ (.Y(_10710_),
    .A(_07816_),
    .B(_10703_));
 sg13g2_and2_1 _15346_ (.A(_10709_),
    .B(_10710_),
    .X(_10711_));
 sg13g2_nor3_1 _15347_ (.A(_08244_),
    .B(_10708_),
    .C(_10711_),
    .Y(_10712_));
 sg13g2_a21o_1 _15348_ (.A2(_10708_),
    .A1(net1438),
    .B1(_10712_),
    .X(_00637_));
 sg13g2_nand2_1 _15349_ (.Y(_10713_),
    .A(_08249_),
    .B(_09831_));
 sg13g2_a21oi_1 _15350_ (.A1(_10264_),
    .A2(_10713_),
    .Y(_10714_),
    .B1(net421));
 sg13g2_nand3_1 _15351_ (.B(_09830_),
    .C(_10264_),
    .A(net5190),
    .Y(_10715_));
 sg13g2_nor2b_1 _15352_ (.A(_10714_),
    .B_N(_10715_),
    .Y(_00638_));
 sg13g2_nor3_1 _15353_ (.A(_09829_),
    .B(_09831_),
    .C(_10166_),
    .Y(_10716_));
 sg13g2_nand2_1 _15354_ (.Y(_10717_),
    .A(_07867_),
    .B(_08395_));
 sg13g2_mux2_1 _15355_ (.A0(net3148),
    .A1(_10717_),
    .S(_10716_),
    .X(_00639_));
 sg13g2_nor2_1 _15356_ (.A(net6194),
    .B(_09820_),
    .Y(_10718_));
 sg13g2_nor2_1 _15357_ (.A(_08389_),
    .B(_10718_),
    .Y(_10719_));
 sg13g2_and4_1 _15358_ (.A(_08385_),
    .B(_08394_),
    .C(_09819_),
    .D(_10719_),
    .X(_10720_));
 sg13g2_nand3_1 _15359_ (.B(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .C(net4691),
    .A(net6196),
    .Y(_10721_));
 sg13g2_o21ai_1 _15360_ (.B1(_10721_),
    .Y(_00640_),
    .A1(_07967_),
    .A2(net4691));
 sg13g2_nand3_1 _15361_ (.B(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .C(net4691),
    .A(net6196),
    .Y(_10722_));
 sg13g2_o21ai_1 _15362_ (.B1(_10722_),
    .Y(_00641_),
    .A1(_07968_),
    .A2(net4692));
 sg13g2_nand3_1 _15363_ (.B(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .C(net4696),
    .A(net6197),
    .Y(_10723_));
 sg13g2_o21ai_1 _15364_ (.B1(_10723_),
    .Y(_00642_),
    .A1(_07969_),
    .A2(net4696));
 sg13g2_nand3_1 _15365_ (.B(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .C(net4697),
    .A(net6197),
    .Y(_10724_));
 sg13g2_o21ai_1 _15366_ (.B1(_10724_),
    .Y(_00643_),
    .A1(_07970_),
    .A2(net4698));
 sg13g2_nand3_1 _15367_ (.B(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .C(net4691),
    .A(net6200),
    .Y(_10725_));
 sg13g2_o21ai_1 _15368_ (.B1(_10725_),
    .Y(_00644_),
    .A1(_07971_),
    .A2(net4692));
 sg13g2_nand3_1 _15369_ (.B(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .C(net4690),
    .A(net6196),
    .Y(_10726_));
 sg13g2_o21ai_1 _15370_ (.B1(_10726_),
    .Y(_00645_),
    .A1(_07972_),
    .A2(net4690));
 sg13g2_nand3_1 _15371_ (.B(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .C(net4694),
    .A(net6199),
    .Y(_10727_));
 sg13g2_o21ai_1 _15372_ (.B1(_10727_),
    .Y(_00646_),
    .A1(_07973_),
    .A2(net4694));
 sg13g2_nand3_1 _15373_ (.B(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .C(net4698),
    .A(net6197),
    .Y(_10728_));
 sg13g2_o21ai_1 _15374_ (.B1(_10728_),
    .Y(_00647_),
    .A1(_07974_),
    .A2(net4698));
 sg13g2_nand3_1 _15375_ (.B(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .C(net4693),
    .A(net6199),
    .Y(_10729_));
 sg13g2_o21ai_1 _15376_ (.B1(_10729_),
    .Y(_00648_),
    .A1(_07975_),
    .A2(net4693));
 sg13g2_nand3_1 _15377_ (.B(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .C(net4699),
    .A(net6198),
    .Y(_10730_));
 sg13g2_o21ai_1 _15378_ (.B1(_10730_),
    .Y(_00649_),
    .A1(_07976_),
    .A2(net4698));
 sg13g2_nand3_1 _15379_ (.B(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .C(net4695),
    .A(net6199),
    .Y(_10731_));
 sg13g2_o21ai_1 _15380_ (.B1(_10731_),
    .Y(_00650_),
    .A1(_07977_),
    .A2(net4695));
 sg13g2_nand3_1 _15381_ (.B(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .C(net4695),
    .A(net6199),
    .Y(_10732_));
 sg13g2_o21ai_1 _15382_ (.B1(_10732_),
    .Y(_00651_),
    .A1(_07978_),
    .A2(net4695));
 sg13g2_nand3_1 _15383_ (.B(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .C(net4697),
    .A(net6197),
    .Y(_10733_));
 sg13g2_o21ai_1 _15384_ (.B1(_10733_),
    .Y(_00652_),
    .A1(_07979_),
    .A2(net4697));
 sg13g2_nand3_1 _15385_ (.B(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .C(net4689),
    .A(net6196),
    .Y(_10734_));
 sg13g2_o21ai_1 _15386_ (.B1(_10734_),
    .Y(_00653_),
    .A1(_07980_),
    .A2(net4689));
 sg13g2_nand3_1 _15387_ (.B(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .C(net4694),
    .A(net6199),
    .Y(_10735_));
 sg13g2_o21ai_1 _15388_ (.B1(_10735_),
    .Y(_00654_),
    .A1(_07981_),
    .A2(net4694));
 sg13g2_nand3_1 _15389_ (.B(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .C(net4694),
    .A(net6195),
    .Y(_10736_));
 sg13g2_o21ai_1 _15390_ (.B1(_10736_),
    .Y(_00655_),
    .A1(_07982_),
    .A2(net4694));
 sg13g2_nand3_1 _15391_ (.B(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .C(net4691),
    .A(net6198),
    .Y(_10737_));
 sg13g2_o21ai_1 _15392_ (.B1(_10737_),
    .Y(_00656_),
    .A1(_07983_),
    .A2(net4692));
 sg13g2_nand3_1 _15393_ (.B(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .C(net4696),
    .A(net6198),
    .Y(_10738_));
 sg13g2_o21ai_1 _15394_ (.B1(_10738_),
    .Y(_00657_),
    .A1(_07984_),
    .A2(net4696));
 sg13g2_nand3_1 _15395_ (.B(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .C(net4689),
    .A(net6196),
    .Y(_10739_));
 sg13g2_o21ai_1 _15396_ (.B1(_10739_),
    .Y(_00658_),
    .A1(_07985_),
    .A2(net4689));
 sg13g2_nand3_1 _15397_ (.B(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .C(net4690),
    .A(net6195),
    .Y(_10740_));
 sg13g2_o21ai_1 _15398_ (.B1(_10740_),
    .Y(_00659_),
    .A1(_07986_),
    .A2(net4690));
 sg13g2_nand3_1 _15399_ (.B(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .C(net4696),
    .A(net6197),
    .Y(_10741_));
 sg13g2_o21ai_1 _15400_ (.B1(_10741_),
    .Y(_00660_),
    .A1(_07987_),
    .A2(net4696));
 sg13g2_nand3_1 _15401_ (.B(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .C(net4694),
    .A(net6199),
    .Y(_10742_));
 sg13g2_o21ai_1 _15402_ (.B1(_10742_),
    .Y(_00661_),
    .A1(_07988_),
    .A2(net4694));
 sg13g2_nand3_1 _15403_ (.B(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .C(net4698),
    .A(net6197),
    .Y(_10743_));
 sg13g2_o21ai_1 _15404_ (.B1(_10743_),
    .Y(_00662_),
    .A1(_07989_),
    .A2(net4698));
 sg13g2_nand3_1 _15405_ (.B(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .C(net4698),
    .A(net6197),
    .Y(_10744_));
 sg13g2_o21ai_1 _15406_ (.B1(_10744_),
    .Y(_00663_),
    .A1(_07990_),
    .A2(net4698));
 sg13g2_nand3_1 _15407_ (.B(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .C(net4696),
    .A(net6197),
    .Y(_10745_));
 sg13g2_o21ai_1 _15408_ (.B1(_10745_),
    .Y(_00664_),
    .A1(_07991_),
    .A2(net4696));
 sg13g2_nand3_1 _15409_ (.B(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .C(net4691),
    .A(net6200),
    .Y(_10746_));
 sg13g2_o21ai_1 _15410_ (.B1(_10746_),
    .Y(_00665_),
    .A1(_07992_),
    .A2(net4692));
 sg13g2_nand3_1 _15411_ (.B(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .C(net4692),
    .A(net6198),
    .Y(_10747_));
 sg13g2_o21ai_1 _15412_ (.B1(_10747_),
    .Y(_00666_),
    .A1(_07993_),
    .A2(net4692));
 sg13g2_nand3_1 _15413_ (.B(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .C(net4693),
    .A(net6199),
    .Y(_10748_));
 sg13g2_o21ai_1 _15414_ (.B1(_10748_),
    .Y(_00667_),
    .A1(_07994_),
    .A2(net4690));
 sg13g2_nand3_1 _15415_ (.B(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .C(net4691),
    .A(net6196),
    .Y(_10749_));
 sg13g2_o21ai_1 _15416_ (.B1(_10749_),
    .Y(_00668_),
    .A1(_07995_),
    .A2(net4691));
 sg13g2_nand3_1 _15417_ (.B(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .C(net4689),
    .A(net6196),
    .Y(_10750_));
 sg13g2_o21ai_1 _15418_ (.B1(_10750_),
    .Y(_00669_),
    .A1(_07996_),
    .A2(net4689));
 sg13g2_nand3_1 _15419_ (.B(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .C(net4689),
    .A(net6196),
    .Y(_10751_));
 sg13g2_o21ai_1 _15420_ (.B1(_10751_),
    .Y(_00670_),
    .A1(_07997_),
    .A2(net4689));
 sg13g2_nand3_1 _15421_ (.B(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .C(net4690),
    .A(net6199),
    .Y(_10752_));
 sg13g2_o21ai_1 _15422_ (.B1(_10752_),
    .Y(_00671_),
    .A1(_07998_),
    .A2(net4690));
 sg13g2_nor2_1 _15423_ (.A(_08293_),
    .B(_10708_),
    .Y(_10753_));
 sg13g2_o21ai_1 _15424_ (.B1(net6205),
    .Y(_10754_),
    .A1(net6504),
    .A2(net6193));
 sg13g2_a21oi_1 _15425_ (.A1(_10710_),
    .A2(_10754_),
    .Y(_10755_),
    .B1(_08245_));
 sg13g2_mux2_1 _15426_ (.A0(net6507),
    .A1(_10755_),
    .S(_10753_),
    .X(_00672_));
 sg13g2_nor2_1 _15427_ (.A(net6503),
    .B(_08419_),
    .Y(_10756_));
 sg13g2_nor2_2 _15428_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .Y(_10757_));
 sg13g2_or2_1 _15429_ (.X(_10758_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ));
 sg13g2_nand2_1 _15430_ (.Y(_10759_),
    .A(net6503),
    .B(_10757_));
 sg13g2_nand2b_1 _15431_ (.Y(_10760_),
    .B(_10759_),
    .A_N(_10756_));
 sg13g2_mux2_1 _15432_ (.A0(net6507),
    .A1(net6506),
    .S(_10760_),
    .X(_00673_));
 sg13g2_xor2_1 _15433_ (.B(net311),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .X(_00674_));
 sg13g2_nand3_1 _15434_ (.B(net3298),
    .C(net311),
    .A(net3222),
    .Y(_10761_));
 sg13g2_a21o_1 _15435_ (.A2(net311),
    .A1(net3222),
    .B1(net3298),
    .X(_10762_));
 sg13g2_and2_1 _15436_ (.A(_10761_),
    .B(_10762_),
    .X(_00675_));
 sg13g2_nand4_1 _15437_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .C(net363),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .Y(_10763_),
    .D(net311));
 sg13g2_xnor2_1 _15438_ (.Y(_00676_),
    .A(net363),
    .B(_10761_));
 sg13g2_nor2_1 _15439_ (.A(_07907_),
    .B(_10763_),
    .Y(_10764_));
 sg13g2_xnor2_1 _15440_ (.Y(_00677_),
    .A(net358),
    .B(_10763_));
 sg13g2_xor2_1 _15441_ (.B(_10764_),
    .A(net253),
    .X(_00678_));
 sg13g2_nand3_1 _15442_ (.B(net1638),
    .C(_10764_),
    .A(net253),
    .Y(_10765_));
 sg13g2_a21o_1 _15443_ (.A2(_10764_),
    .A1(net253),
    .B1(net1638),
    .X(_10766_));
 sg13g2_and2_1 _15444_ (.A(_10765_),
    .B(_10766_),
    .X(_00679_));
 sg13g2_nor2_1 _15445_ (.A(_07908_),
    .B(_10765_),
    .Y(_10767_));
 sg13g2_xnor2_1 _15446_ (.Y(_00680_),
    .A(net562),
    .B(_10765_));
 sg13g2_and2_1 _15447_ (.A(net338),
    .B(_10767_),
    .X(_10768_));
 sg13g2_xor2_1 _15448_ (.B(_10767_),
    .A(net338),
    .X(_00681_));
 sg13g2_xor2_1 _15449_ (.B(_10768_),
    .A(net354),
    .X(_00682_));
 sg13g2_nand3_1 _15450_ (.B(net354),
    .C(_10768_),
    .A(net3313),
    .Y(_10769_));
 sg13g2_a21o_1 _15451_ (.A2(_10768_),
    .A1(net354),
    .B1(net3313),
    .X(_10770_));
 sg13g2_and2_1 _15452_ (.A(_10769_),
    .B(_10770_),
    .X(_00683_));
 sg13g2_nand4_1 _15453_ (.B(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .Y(_10771_),
    .D(_10768_));
 sg13g2_xnor2_1 _15454_ (.Y(_00684_),
    .A(net388),
    .B(_10769_));
 sg13g2_xnor2_1 _15455_ (.Y(_00685_),
    .A(net144),
    .B(_10771_));
 sg13g2_nand2_2 _15456_ (.Y(_10772_),
    .A(net6484),
    .B(_08657_));
 sg13g2_nor4_1 _15457_ (.A(net6203),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .D(_10772_),
    .Y(_10773_));
 sg13g2_and3_2 _15458_ (.X(_10774_),
    .A(_08411_),
    .B(_08412_),
    .C(_08657_));
 sg13g2_nand3_1 _15459_ (.B(_08412_),
    .C(_08657_),
    .A(_08411_),
    .Y(_10775_));
 sg13g2_nor2_1 _15460_ (.A(net1745),
    .B(net5519),
    .Y(_10776_));
 sg13g2_nor2_1 _15461_ (.A(net1415),
    .B(net5519),
    .Y(_10777_));
 sg13g2_nor3_1 _15462_ (.A(_10773_),
    .B(_10776_),
    .C(_10777_),
    .Y(_10778_));
 sg13g2_nor3_2 _15463_ (.A(_07816_),
    .B(_07875_),
    .C(_10778_),
    .Y(_10779_));
 sg13g2_mux4_1 _15464_ (.S0(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[0] ),
    .A0(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger ),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d1 ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d2 ),
    .A3(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d3 ),
    .S1(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[1] ),
    .X(_10780_));
 sg13g2_a22oi_1 _15465_ (.Y(_10781_),
    .B1(_10780_),
    .B2(_08665_),
    .A2(_10759_),
    .A1(_07875_));
 sg13g2_or3_1 _15466_ (.A(_10756_),
    .B(_10779_),
    .C(_10781_),
    .X(_10782_));
 sg13g2_nand2_1 _15467_ (.Y(_10783_),
    .A(net6489),
    .B(net9));
 sg13g2_nand2_1 _15468_ (.Y(_10784_),
    .A(net1237),
    .B(net5025));
 sg13g2_o21ai_1 _15469_ (.B1(_10784_),
    .Y(_00686_),
    .A1(net5025),
    .A2(_10783_));
 sg13g2_nand2_1 _15470_ (.Y(_10785_),
    .A(net6495),
    .B(net10));
 sg13g2_nand2_1 _15471_ (.Y(_10786_),
    .A(net1357),
    .B(net5027));
 sg13g2_o21ai_1 _15472_ (.B1(_10786_),
    .Y(_00687_),
    .A1(net5027),
    .A2(_10785_));
 sg13g2_nand2_1 _15473_ (.Y(_10787_),
    .A(net6492),
    .B(net11));
 sg13g2_nand2_1 _15474_ (.Y(_10788_),
    .A(net1137),
    .B(net5034));
 sg13g2_o21ai_1 _15475_ (.B1(_10788_),
    .Y(_00688_),
    .A1(net5030),
    .A2(_10787_));
 sg13g2_nand2_1 _15476_ (.Y(_10789_),
    .A(net6494),
    .B(net12));
 sg13g2_nand2_1 _15477_ (.Y(_10790_),
    .A(net1039),
    .B(net5029));
 sg13g2_o21ai_1 _15478_ (.B1(_10790_),
    .Y(_00689_),
    .A1(net5028),
    .A2(_10789_));
 sg13g2_nand2_1 _15479_ (.Y(_10791_),
    .A(net6489),
    .B(net1237));
 sg13g2_nand2_1 _15480_ (.Y(_10792_),
    .A(net1415),
    .B(net5025));
 sg13g2_o21ai_1 _15481_ (.B1(_10792_),
    .Y(_00690_),
    .A1(net5025),
    .A2(_10791_));
 sg13g2_nand2_1 _15482_ (.Y(_10793_),
    .A(net6489),
    .B(net1357));
 sg13g2_nand2_1 _15483_ (.Y(_10794_),
    .A(net1745),
    .B(net5027));
 sg13g2_o21ai_1 _15484_ (.B1(_10794_),
    .Y(_00691_),
    .A1(net5027),
    .A2(_10793_));
 sg13g2_nand2_1 _15485_ (.Y(_10795_),
    .A(net6493),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ));
 sg13g2_nand2_1 _15486_ (.Y(_10796_),
    .A(net997),
    .B(net5030));
 sg13g2_o21ai_1 _15487_ (.B1(_10796_),
    .Y(_00692_),
    .A1(net5030),
    .A2(_10795_));
 sg13g2_nand2_1 _15488_ (.Y(_10797_),
    .A(net6491),
    .B(net1039));
 sg13g2_nand2_1 _15489_ (.Y(_10798_),
    .A(net1414),
    .B(net5031));
 sg13g2_o21ai_1 _15490_ (.B1(_10798_),
    .Y(_00693_),
    .A1(net5028),
    .A2(_10797_));
 sg13g2_nand2_1 _15491_ (.Y(_10799_),
    .A(net6491),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ));
 sg13g2_nand2_1 _15492_ (.Y(_10800_),
    .A(net1087),
    .B(net5026));
 sg13g2_o21ai_1 _15493_ (.B1(_10800_),
    .Y(_00694_),
    .A1(net5026),
    .A2(_10799_));
 sg13g2_nand2_1 _15494_ (.Y(_10801_),
    .A(net6495),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ));
 sg13g2_nand2_1 _15495_ (.Y(_10802_),
    .A(net1228),
    .B(net5028));
 sg13g2_o21ai_1 _15496_ (.B1(_10802_),
    .Y(_00695_),
    .A1(net5027),
    .A2(_10801_));
 sg13g2_nand2_1 _15497_ (.Y(_10803_),
    .A(net6493),
    .B(net997));
 sg13g2_nand2_1 _15498_ (.Y(_10804_),
    .A(net1093),
    .B(net5030));
 sg13g2_o21ai_1 _15499_ (.B1(_10804_),
    .Y(_00696_),
    .A1(net5030),
    .A2(_10803_));
 sg13g2_nand2_1 _15500_ (.Y(_10805_),
    .A(net6492),
    .B(net1414));
 sg13g2_nand2_1 _15501_ (.Y(_10806_),
    .A(net2023),
    .B(net5031));
 sg13g2_o21ai_1 _15502_ (.B1(_10806_),
    .Y(_00697_),
    .A1(net5031),
    .A2(_10805_));
 sg13g2_nand2_1 _15503_ (.Y(_10807_),
    .A(net6491),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ));
 sg13g2_nand2_1 _15504_ (.Y(_10808_),
    .A(net674),
    .B(net5026));
 sg13g2_o21ai_1 _15505_ (.B1(_10808_),
    .Y(_00698_),
    .A1(net5026),
    .A2(_10807_));
 sg13g2_nand2_1 _15506_ (.Y(_10809_),
    .A(net6491),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ));
 sg13g2_nand2_1 _15507_ (.Y(_10810_),
    .A(net1122),
    .B(net5028));
 sg13g2_o21ai_1 _15508_ (.B1(_10810_),
    .Y(_00699_),
    .A1(net5029),
    .A2(_10809_));
 sg13g2_nand2_1 _15509_ (.Y(_10811_),
    .A(net6493),
    .B(net1093));
 sg13g2_nand2_1 _15510_ (.Y(_10812_),
    .A(net1489),
    .B(net5032));
 sg13g2_o21ai_1 _15511_ (.B1(_10812_),
    .Y(_00700_),
    .A1(net5032),
    .A2(_10811_));
 sg13g2_nand2_1 _15512_ (.Y(_10813_),
    .A(net6492),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ));
 sg13g2_nand2_1 _15513_ (.Y(_10814_),
    .A(net1207),
    .B(net5031));
 sg13g2_o21ai_1 _15514_ (.B1(_10814_),
    .Y(_00701_),
    .A1(net5031),
    .A2(_10813_));
 sg13g2_nand2_1 _15515_ (.Y(_10815_),
    .A(net6491),
    .B(net674));
 sg13g2_nand2_1 _15516_ (.Y(_10816_),
    .A(net928),
    .B(net5025));
 sg13g2_o21ai_1 _15517_ (.B1(_10816_),
    .Y(_00702_),
    .A1(net5025),
    .A2(_10815_));
 sg13g2_nand2_1 _15518_ (.Y(_10817_),
    .A(net6489),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ));
 sg13g2_nand2_1 _15519_ (.Y(_10818_),
    .A(net937),
    .B(net5028));
 sg13g2_o21ai_1 _15520_ (.B1(_10818_),
    .Y(_00703_),
    .A1(net5027),
    .A2(_10817_));
 sg13g2_nand2_1 _15521_ (.Y(_10819_),
    .A(net6493),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ));
 sg13g2_nand2_1 _15522_ (.Y(_10820_),
    .A(net1063),
    .B(net5032));
 sg13g2_o21ai_1 _15523_ (.B1(_10820_),
    .Y(_00704_),
    .A1(net5032),
    .A2(_10819_));
 sg13g2_nand2_1 _15524_ (.Y(_10821_),
    .A(net6492),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ));
 sg13g2_nand2_1 _15525_ (.Y(_10822_),
    .A(net1060),
    .B(net5031));
 sg13g2_o21ai_1 _15526_ (.B1(_10822_),
    .Y(_00705_),
    .A1(net5034),
    .A2(_10821_));
 sg13g2_nand2_1 _15527_ (.Y(_10823_),
    .A(net6489),
    .B(net928));
 sg13g2_nand2_1 _15528_ (.Y(_10824_),
    .A(net943),
    .B(net5025));
 sg13g2_o21ai_1 _15529_ (.B1(_10824_),
    .Y(_00706_),
    .A1(net5026),
    .A2(_10823_));
 sg13g2_nand2_1 _15530_ (.Y(_10825_),
    .A(net6489),
    .B(net937));
 sg13g2_nand2_1 _15531_ (.Y(_10826_),
    .A(net1263),
    .B(net5027));
 sg13g2_o21ai_1 _15532_ (.B1(_10826_),
    .Y(_00707_),
    .A1(net5027),
    .A2(_10825_));
 sg13g2_nand2_1 _15533_ (.Y(_10827_),
    .A(net6493),
    .B(net1063));
 sg13g2_nand2_1 _15534_ (.Y(_10828_),
    .A(net1338),
    .B(net5033));
 sg13g2_o21ai_1 _15535_ (.B1(_10828_),
    .Y(_00708_),
    .A1(net5033),
    .A2(_10827_));
 sg13g2_nand2_1 _15536_ (.Y(_10829_),
    .A(net6492),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ));
 sg13g2_nand2_1 _15537_ (.Y(_10830_),
    .A(net915),
    .B(net5031));
 sg13g2_o21ai_1 _15538_ (.B1(_10830_),
    .Y(_00709_),
    .A1(net5031),
    .A2(_10829_));
 sg13g2_nand2_1 _15539_ (.Y(_10831_),
    .A(net6489),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ));
 sg13g2_nand2_1 _15540_ (.Y(_10832_),
    .A(net888),
    .B(net5026));
 sg13g2_o21ai_1 _15541_ (.B1(_10832_),
    .Y(_00710_),
    .A1(net5025),
    .A2(_10831_));
 sg13g2_nand2_1 _15542_ (.Y(_10833_),
    .A(net6491),
    .B(net1263));
 sg13g2_nand2_1 _15543_ (.Y(_10834_),
    .A(net1411),
    .B(net5028));
 sg13g2_o21ai_1 _15544_ (.B1(_10834_),
    .Y(_00711_),
    .A1(net5028),
    .A2(_10833_));
 sg13g2_nand2_1 _15545_ (.Y(_10835_),
    .A(net6493),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ));
 sg13g2_nand2_1 _15546_ (.Y(_10836_),
    .A(net1289),
    .B(net5033));
 sg13g2_o21ai_1 _15547_ (.B1(_10836_),
    .Y(_00712_),
    .A1(net5033),
    .A2(_10835_));
 sg13g2_nand2_1 _15548_ (.Y(_10837_),
    .A(net6492),
    .B(net915));
 sg13g2_nand2_1 _15549_ (.Y(_10838_),
    .A(net1174),
    .B(net5032));
 sg13g2_o21ai_1 _15550_ (.B1(_10838_),
    .Y(_00713_),
    .A1(net5032),
    .A2(_10837_));
 sg13g2_nand2_1 _15551_ (.Y(_10839_),
    .A(net6491),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ));
 sg13g2_nand2_1 _15552_ (.Y(_10840_),
    .A(net153),
    .B(net5030));
 sg13g2_o21ai_1 _15553_ (.B1(_10840_),
    .Y(_00714_),
    .A1(net5030),
    .A2(_10839_));
 sg13g2_nand2_1 _15554_ (.Y(_10841_),
    .A(net6491),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ));
 sg13g2_nand2_1 _15555_ (.Y(_10842_),
    .A(net247),
    .B(net5030));
 sg13g2_o21ai_1 _15556_ (.B1(_10842_),
    .Y(_00715_),
    .A1(net5026),
    .A2(_10841_));
 sg13g2_nand2_1 _15557_ (.Y(_10843_),
    .A(net6492),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ));
 sg13g2_nand2_1 _15558_ (.Y(_10844_),
    .A(net1117),
    .B(net5032));
 sg13g2_o21ai_1 _15559_ (.B1(_10844_),
    .Y(_00716_),
    .A1(net5032),
    .A2(_10843_));
 sg13g2_nand2_1 _15560_ (.Y(_10845_),
    .A(net6492),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ));
 sg13g2_nand2_1 _15561_ (.Y(_10846_),
    .A(net301),
    .B(net5033));
 sg13g2_o21ai_1 _15562_ (.B1(_10846_),
    .Y(_00717_),
    .A1(net5033),
    .A2(_10845_));
 sg13g2_nand2b_1 _15563_ (.Y(_00718_),
    .B(net1028),
    .A_N(net227));
 sg13g2_or2_1 _15564_ (.X(_10847_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .A(net6490));
 sg13g2_or2_1 _15565_ (.X(_10848_),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .A(net6501));
 sg13g2_nor3_2 _15566_ (.A(net6089),
    .B(_10847_),
    .C(_10848_),
    .Y(_10849_));
 sg13g2_or3_1 _15567_ (.A(_10758_),
    .B(_10847_),
    .C(_10848_),
    .X(_10850_));
 sg13g2_a21oi_1 _15568_ (.A1(net6142),
    .A2(net6501),
    .Y(_10851_),
    .B1(_10756_));
 sg13g2_nand2_2 _15569_ (.Y(_10852_),
    .A(_08666_),
    .B(_10851_));
 sg13g2_a21oi_2 _15570_ (.B1(_10852_),
    .Y(_10853_),
    .A2(_10849_),
    .A1(net6503));
 sg13g2_a21o_2 _15571_ (.A2(_10849_),
    .A1(net6503),
    .B1(_10852_),
    .X(_10854_));
 sg13g2_nand2_1 _15572_ (.Y(_10855_),
    .A(net1951),
    .B(net5118));
 sg13g2_nor2_2 _15573_ (.A(_08417_),
    .B(net6010),
    .Y(_10856_));
 sg13g2_nor2_2 _15574_ (.A(net5118),
    .B(_10856_),
    .Y(_10857_));
 sg13g2_o21ai_1 _15575_ (.B1(_10857_),
    .Y(_10858_),
    .A1(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .A2(net6009));
 sg13g2_nand2b_1 _15576_ (.Y(_10859_),
    .B(_08660_),
    .A_N(_10847_));
 sg13g2_and2_1 _15577_ (.A(net6142),
    .B(_10859_),
    .X(_10860_));
 sg13g2_nand2b_1 _15578_ (.Y(_10861_),
    .B(net5122),
    .A_N(net5116));
 sg13g2_nand2_1 _15579_ (.Y(_10862_),
    .A(net1951),
    .B(net5056));
 sg13g2_and2_1 _15580_ (.A(net6506),
    .B(_08634_),
    .X(_10863_));
 sg13g2_nand2_2 _15581_ (.Y(_10864_),
    .A(_10757_),
    .B(net6009));
 sg13g2_a22oi_1 _15582_ (.Y(_10865_),
    .B1(_10864_),
    .B2(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .A2(net5317),
    .A1(net605));
 sg13g2_a22oi_1 _15583_ (.Y(_00719_),
    .B1(_10862_),
    .B2(_10865_),
    .A2(_10858_),
    .A1(_10855_));
 sg13g2_nand2_2 _15584_ (.Y(_10866_),
    .A(_08417_),
    .B(net6011));
 sg13g2_nand2_1 _15585_ (.Y(_10867_),
    .A(_10757_),
    .B(_10866_));
 sg13g2_nand2_1 _15586_ (.Y(_10868_),
    .A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .B(net5115));
 sg13g2_a22oi_1 _15587_ (.Y(_10869_),
    .B1(net341),
    .B2(net5315),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .A1(net6497));
 sg13g2_a21oi_1 _15588_ (.A1(_10868_),
    .A2(_10869_),
    .Y(_10870_),
    .B1(net5118));
 sg13g2_a21o_1 _15589_ (.A2(net5057),
    .A1(net1929),
    .B1(_10870_),
    .X(_00720_));
 sg13g2_nand2_1 _15590_ (.Y(_10871_),
    .A(net318),
    .B(net5316));
 sg13g2_a22oi_1 _15591_ (.Y(_10872_),
    .B1(net5115),
    .B2(\soc_inst.mem_ctrl.spi_addr[2] ),
    .A2(net1929),
    .A1(net6498));
 sg13g2_a21oi_1 _15592_ (.A1(_10871_),
    .A2(_10872_),
    .Y(_10873_),
    .B1(net5117));
 sg13g2_a21o_1 _15593_ (.A2(net5057),
    .A1(net2295),
    .B1(_10873_),
    .X(_00721_));
 sg13g2_nand2_1 _15594_ (.Y(_10874_),
    .A(net745),
    .B(net5316));
 sg13g2_a22oi_1 _15595_ (.Y(_10875_),
    .B1(net5115),
    .B2(\soc_inst.mem_ctrl.spi_addr[3] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .A1(net6497));
 sg13g2_a21oi_1 _15596_ (.A1(_10874_),
    .A2(_10875_),
    .Y(_10876_),
    .B1(net5117));
 sg13g2_a21o_1 _15597_ (.A2(net5056),
    .A1(net2063),
    .B1(_10876_),
    .X(_00722_));
 sg13g2_nand2_1 _15598_ (.Y(_10877_),
    .A(net1391),
    .B(net5117));
 sg13g2_o21ai_1 _15599_ (.B1(_10857_),
    .Y(_10878_),
    .A1(\soc_inst.mem_ctrl.spi_addr[4] ),
    .A2(net6009));
 sg13g2_and2_1 _15600_ (.A(net6482),
    .B(_10859_),
    .X(_10879_));
 sg13g2_a22oi_1 _15601_ (.Y(_10880_),
    .B1(_10864_),
    .B2(\soc_inst.mem_ctrl.spi_addr[4] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .A1(net6498));
 sg13g2_inv_1 _15602_ (.Y(_10881_),
    .A(_10880_));
 sg13g2_a221oi_1 _15603_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .C1(_10881_),
    .B1(net5109),
    .A1(net802),
    .Y(_10882_),
    .A2(net5315));
 sg13g2_nand2_1 _15604_ (.Y(_10883_),
    .A(net1391),
    .B(net5056));
 sg13g2_a22oi_1 _15605_ (.Y(_00723_),
    .B1(_10882_),
    .B2(_10883_),
    .A2(_10878_),
    .A1(_10877_));
 sg13g2_o21ai_1 _15606_ (.B1(_10857_),
    .Y(_10884_),
    .A1(\soc_inst.mem_ctrl.spi_addr[5] ),
    .A2(net6009));
 sg13g2_and2_1 _15607_ (.A(net415),
    .B(net5314),
    .X(_10885_));
 sg13g2_a221oi_1 _15608_ (.B2(net5116),
    .C1(_10885_),
    .B1(net2360),
    .A1(net6497),
    .Y(_10886_),
    .A2(net1391));
 sg13g2_a22oi_1 _15609_ (.Y(_10887_),
    .B1(net5110),
    .B2(net1929),
    .A2(_10864_),
    .A1(\soc_inst.mem_ctrl.spi_addr[5] ));
 sg13g2_a21oi_1 _15610_ (.A1(_10886_),
    .A2(_10887_),
    .Y(_10888_),
    .B1(_10884_));
 sg13g2_a21o_1 _15611_ (.A2(net5117),
    .A1(net2360),
    .B1(_10888_),
    .X(_00724_));
 sg13g2_nand2_1 _15612_ (.Y(_10889_),
    .A(net908),
    .B(net5117));
 sg13g2_o21ai_1 _15613_ (.B1(_10857_),
    .Y(_10890_),
    .A1(\soc_inst.mem_ctrl.spi_addr[6] ),
    .A2(net6009));
 sg13g2_a22oi_1 _15614_ (.Y(_10891_),
    .B1(_10864_),
    .B2(\soc_inst.mem_ctrl.spi_addr[6] ),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .A1(net6497));
 sg13g2_inv_1 _15615_ (.Y(_10892_),
    .A(_10891_));
 sg13g2_a221oi_1 _15616_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .C1(_10892_),
    .B1(net5110),
    .A1(net418),
    .Y(_10893_),
    .A2(net5315));
 sg13g2_nand2_1 _15617_ (.Y(_10894_),
    .A(net908),
    .B(net5056));
 sg13g2_a22oi_1 _15618_ (.Y(_00725_),
    .B1(_10893_),
    .B2(_10894_),
    .A2(_10890_),
    .A1(_10889_));
 sg13g2_o21ai_1 _15619_ (.B1(_10857_),
    .Y(_10895_),
    .A1(\soc_inst.mem_ctrl.spi_addr[7] ),
    .A2(net6009));
 sg13g2_and2_1 _15620_ (.A(net266),
    .B(net5315),
    .X(_10896_));
 sg13g2_a221oi_1 _15621_ (.B2(net5116),
    .C1(_10896_),
    .B1(net2423),
    .A1(net6497),
    .Y(_10897_),
    .A2(net908));
 sg13g2_a22oi_1 _15622_ (.Y(_10898_),
    .B1(net5111),
    .B2(net2063),
    .A2(_10864_),
    .A1(\soc_inst.mem_ctrl.spi_addr[7] ));
 sg13g2_a21oi_1 _15623_ (.A1(_10897_),
    .A2(_10898_),
    .Y(_10899_),
    .B1(_10895_));
 sg13g2_a21o_1 _15624_ (.A2(net5117),
    .A1(net2423),
    .B1(_10899_),
    .X(_00726_));
 sg13g2_a221oi_1 _15625_ (.B2(\soc_inst.mem_ctrl.spi_addr[8] ),
    .C1(net6011),
    .B1(net6089),
    .A1(net6498),
    .Y(_10900_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ));
 sg13g2_a22oi_1 _15626_ (.Y(_10901_),
    .B1(net5109),
    .B2(net1391),
    .A2(net5316),
    .A1(net853));
 sg13g2_o21ai_1 _15627_ (.B1(net5122),
    .Y(_10902_),
    .A1(\soc_inst.mem_ctrl.spi_addr[8] ),
    .A2(_10866_));
 sg13g2_a221oi_1 _15628_ (.B2(_10901_),
    .C1(_10902_),
    .B1(_10900_),
    .A1(_07817_),
    .Y(_10903_),
    .A2(net5320));
 sg13g2_a21o_1 _15629_ (.A2(net5057),
    .A1(net2117),
    .B1(_10903_),
    .X(_00727_));
 sg13g2_a221oi_1 _15630_ (.B2(\soc_inst.mem_ctrl.spi_addr[9] ),
    .C1(net6011),
    .B1(net6089),
    .A1(net6498),
    .Y(_10904_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ));
 sg13g2_a22oi_1 _15631_ (.Y(_10905_),
    .B1(net5109),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .A2(net5316),
    .A1(net1086));
 sg13g2_o21ai_1 _15632_ (.B1(net5122),
    .Y(_10906_),
    .A1(\soc_inst.mem_ctrl.spi_addr[9] ),
    .A2(_10866_));
 sg13g2_a221oi_1 _15633_ (.B2(_10905_),
    .C1(_10906_),
    .B1(_10904_),
    .A1(_07819_),
    .Y(_10907_),
    .A2(_10856_));
 sg13g2_a21o_1 _15634_ (.A2(net5056),
    .A1(net2052),
    .B1(_10907_),
    .X(_00728_));
 sg13g2_nand2_1 _15635_ (.Y(_10908_),
    .A(net568),
    .B(net5056));
 sg13g2_nand2_1 _15636_ (.Y(_10909_),
    .A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .B(net5320));
 sg13g2_a22oi_1 _15637_ (.Y(_10910_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .B2(net5315),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .A1(net6497));
 sg13g2_nand2_1 _15638_ (.Y(_10911_),
    .A(_10909_),
    .B(_10910_));
 sg13g2_a221oi_1 _15639_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .C1(_10911_),
    .B1(net5109),
    .A1(\soc_inst.mem_ctrl.spi_addr[10] ),
    .Y(_10912_),
    .A2(net5115));
 sg13g2_o21ai_1 _15640_ (.B1(_10908_),
    .Y(_00729_),
    .A1(net5117),
    .A2(_10912_));
 sg13g2_nand2_1 _15641_ (.Y(_10913_),
    .A(net1075),
    .B(net5056));
 sg13g2_nand2_1 _15642_ (.Y(_10914_),
    .A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .B(net5320));
 sg13g2_a22oi_1 _15643_ (.Y(_10915_),
    .B1(net841),
    .B2(net5316),
    .A2(net568),
    .A1(net6497));
 sg13g2_nand2_1 _15644_ (.Y(_10916_),
    .A(_10914_),
    .B(_10915_));
 sg13g2_a221oi_1 _15645_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .C1(_10916_),
    .B1(net5110),
    .A1(\soc_inst.mem_ctrl.spi_addr[11] ),
    .Y(_10917_),
    .A2(net5115));
 sg13g2_o21ai_1 _15646_ (.B1(_10913_),
    .Y(_00730_),
    .A1(net5118),
    .A2(_10917_));
 sg13g2_o21ai_1 _15647_ (.B1(net6011),
    .Y(_10918_),
    .A1(_07841_),
    .A2(net5568));
 sg13g2_a21oi_1 _15648_ (.A1(\soc_inst.mem_ctrl.spi_addr[4] ),
    .A2(net5568),
    .Y(_10919_),
    .B1(_10918_));
 sg13g2_nand2_1 _15649_ (.Y(_10920_),
    .A(net2179),
    .B(net5057));
 sg13g2_a22oi_1 _15650_ (.Y(_10921_),
    .B1(net6089),
    .B2(\soc_inst.mem_ctrl.spi_addr[12] ),
    .A2(net1075),
    .A1(net6498));
 sg13g2_nand2_1 _15651_ (.Y(_10922_),
    .A(net6010),
    .B(_10921_));
 sg13g2_a221oi_1 _15652_ (.B2(net2117),
    .C1(_10922_),
    .B1(net5111),
    .A1(net931),
    .Y(_10923_),
    .A2(net5317));
 sg13g2_nor2_1 _15653_ (.A(net2179),
    .B(net5122),
    .Y(_10924_));
 sg13g2_a221oi_1 _15654_ (.B2(_10923_),
    .C1(_10924_),
    .B1(_10920_),
    .A1(net5122),
    .Y(_00731_),
    .A2(_10919_));
 sg13g2_nand2_1 _15655_ (.Y(_10925_),
    .A(net416),
    .B(net5055));
 sg13g2_nand2_1 _15656_ (.Y(_10926_),
    .A(\soc_inst.mem_ctrl.spi_addr[5] ),
    .B(net5320));
 sg13g2_a22oi_1 _15657_ (.Y(_10927_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[13] ),
    .B2(net5315),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .A1(net6496));
 sg13g2_nand2_1 _15658_ (.Y(_10928_),
    .A(_10926_),
    .B(_10927_));
 sg13g2_a221oi_1 _15659_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .C1(_10928_),
    .B1(net5109),
    .A1(\soc_inst.mem_ctrl.spi_addr[13] ),
    .Y(_10929_),
    .A2(net5114));
 sg13g2_o21ai_1 _15660_ (.B1(_10925_),
    .Y(_00732_),
    .A1(net5119),
    .A2(_10929_));
 sg13g2_nand2_1 _15661_ (.Y(_10930_),
    .A(net396),
    .B(net5056));
 sg13g2_nand2_1 _15662_ (.Y(_10931_),
    .A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .B(net5320));
 sg13g2_a22oi_1 _15663_ (.Y(_10932_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[14] ),
    .B2(net5315),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .A1(net6496));
 sg13g2_nand2_1 _15664_ (.Y(_10933_),
    .A(_10931_),
    .B(_10932_));
 sg13g2_a221oi_1 _15665_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ),
    .C1(_10933_),
    .B1(net5109),
    .A1(\soc_inst.mem_ctrl.spi_addr[14] ),
    .Y(_10934_),
    .A2(net5114));
 sg13g2_o21ai_1 _15666_ (.B1(_10930_),
    .Y(_00733_),
    .A1(net5117),
    .A2(_10934_));
 sg13g2_nand2_1 _15667_ (.Y(_10935_),
    .A(net601),
    .B(net5055));
 sg13g2_nand2_1 _15668_ (.Y(_10936_),
    .A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .B(net5320));
 sg13g2_a22oi_1 _15669_ (.Y(_10937_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[15] ),
    .B2(net5315),
    .A2(net396),
    .A1(net6497));
 sg13g2_nand2_1 _15670_ (.Y(_10938_),
    .A(_10936_),
    .B(_10937_));
 sg13g2_a221oi_1 _15671_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .C1(_10938_),
    .B1(net5110),
    .A1(\soc_inst.mem_ctrl.spi_addr[15] ),
    .Y(_10939_),
    .A2(net5114));
 sg13g2_o21ai_1 _15672_ (.B1(_10935_),
    .Y(_00734_),
    .A1(net5119),
    .A2(_10939_));
 sg13g2_nand2_1 _15673_ (.Y(_10940_),
    .A(net956),
    .B(net5055));
 sg13g2_nand2_1 _15674_ (.Y(_10941_),
    .A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .B(net5109));
 sg13g2_a22oi_1 _15675_ (.Y(_10942_),
    .B1(net352),
    .B2(net5314),
    .A2(net601),
    .A1(net6496));
 sg13g2_nand2_1 _15676_ (.Y(_10943_),
    .A(_10941_),
    .B(_10942_));
 sg13g2_a221oi_1 _15677_ (.B2(\soc_inst.mem_ctrl.spi_addr[16] ),
    .C1(_10943_),
    .B1(net5114),
    .A1(\soc_inst.mem_ctrl.spi_addr[8] ),
    .Y(_10944_),
    .A2(net5319));
 sg13g2_o21ai_1 _15678_ (.B1(_10940_),
    .Y(_00735_),
    .A1(net5119),
    .A2(_10944_));
 sg13g2_a221oi_1 _15679_ (.B2(\soc_inst.mem_ctrl.spi_addr[17] ),
    .C1(net6011),
    .B1(net6089),
    .A1(net6496),
    .Y(_10945_),
    .A2(net956));
 sg13g2_a22oi_1 _15680_ (.Y(_10946_),
    .B1(net5112),
    .B2(net416),
    .A2(net5314),
    .A1(net376));
 sg13g2_o21ai_1 _15681_ (.B1(net5122),
    .Y(_10947_),
    .A1(\soc_inst.mem_ctrl.spi_addr[17] ),
    .A2(_10866_));
 sg13g2_a221oi_1 _15682_ (.B2(_10946_),
    .C1(_10947_),
    .B1(_10945_),
    .A1(_07835_),
    .Y(_10948_),
    .A2(net5319));
 sg13g2_a21o_1 _15683_ (.A2(net5055),
    .A1(net1807),
    .B1(_10948_),
    .X(_00736_));
 sg13g2_nand2_1 _15684_ (.Y(_10949_),
    .A(net583),
    .B(net5058));
 sg13g2_nand2_1 _15685_ (.Y(_10950_),
    .A(net396),
    .B(net5109));
 sg13g2_a22oi_1 _15686_ (.Y(_10951_),
    .B1(net309),
    .B2(net5314),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .A1(net6496));
 sg13g2_nand2_1 _15687_ (.Y(_10952_),
    .A(_10950_),
    .B(_10951_));
 sg13g2_a221oi_1 _15688_ (.B2(\soc_inst.mem_ctrl.spi_addr[18] ),
    .C1(_10952_),
    .B1(net5114),
    .A1(\soc_inst.mem_ctrl.spi_addr[10] ),
    .Y(_10953_),
    .A2(net5319));
 sg13g2_o21ai_1 _15689_ (.B1(_10949_),
    .Y(_00737_),
    .A1(net5119),
    .A2(_10953_));
 sg13g2_a221oi_1 _15690_ (.B2(\soc_inst.mem_ctrl.spi_addr[19] ),
    .C1(net6011),
    .B1(net6089),
    .A1(net6499),
    .Y(_10954_),
    .A2(net583));
 sg13g2_a22oi_1 _15691_ (.Y(_10955_),
    .B1(net5112),
    .B2(net601),
    .A2(net5314),
    .A1(net379));
 sg13g2_o21ai_1 _15692_ (.B1(net5122),
    .Y(_10956_),
    .A1(\soc_inst.mem_ctrl.spi_addr[19] ),
    .A2(_10866_));
 sg13g2_a221oi_1 _15693_ (.B2(_10955_),
    .C1(_10956_),
    .B1(_10954_),
    .A1(_07839_),
    .Y(_10957_),
    .A2(net5319));
 sg13g2_a21o_1 _15694_ (.A2(net5055),
    .A1(net1670),
    .B1(_10957_),
    .X(_00738_));
 sg13g2_a221oi_1 _15695_ (.B2(\soc_inst.mem_ctrl.spi_addr[20] ),
    .C1(net6011),
    .B1(net6089),
    .A1(net6496),
    .Y(_10958_),
    .A2(net1670));
 sg13g2_a22oi_1 _15696_ (.Y(_10959_),
    .B1(net5112),
    .B2(net956),
    .A2(net5318),
    .A1(net701));
 sg13g2_o21ai_1 _15697_ (.B1(net5122),
    .Y(_10960_),
    .A1(\soc_inst.mem_ctrl.spi_addr[20] ),
    .A2(_10866_));
 sg13g2_a221oi_1 _15698_ (.B2(_10959_),
    .C1(_10960_),
    .B1(_10958_),
    .A1(_07841_),
    .Y(_10961_),
    .A2(net5319));
 sg13g2_a21o_1 _15699_ (.A2(net5055),
    .A1(net2335),
    .B1(_10961_),
    .X(_00739_));
 sg13g2_nand2_1 _15700_ (.Y(_10962_),
    .A(net1041),
    .B(net5055));
 sg13g2_nand2_1 _15701_ (.Y(_10963_),
    .A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .B(net5319));
 sg13g2_a22oi_1 _15702_ (.Y(_10964_),
    .B1(net431),
    .B2(net5314),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .A1(net6496));
 sg13g2_nand2_1 _15703_ (.Y(_10965_),
    .A(_10963_),
    .B(_10964_));
 sg13g2_a221oi_1 _15704_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .C1(_10965_),
    .B1(net5112),
    .A1(\soc_inst.mem_ctrl.spi_addr[21] ),
    .Y(_10966_),
    .A2(net5114));
 sg13g2_o21ai_1 _15705_ (.B1(_10962_),
    .Y(_00740_),
    .A1(net5119),
    .A2(_10966_));
 sg13g2_nand2_1 _15706_ (.Y(_10967_),
    .A(net994),
    .B(net5055));
 sg13g2_nand2_1 _15707_ (.Y(_10968_),
    .A(\soc_inst.mem_ctrl.spi_addr[14] ),
    .B(net5319));
 sg13g2_a22oi_1 _15708_ (.Y(_10969_),
    .B1(net898),
    .B2(net5314),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .A1(net6502));
 sg13g2_nand2_1 _15709_ (.Y(_10970_),
    .A(_10968_),
    .B(_10969_));
 sg13g2_a221oi_1 _15710_ (.B2(net583),
    .C1(_10970_),
    .B1(net5112),
    .A1(\soc_inst.mem_ctrl.spi_addr[22] ),
    .Y(_10971_),
    .A2(net5114));
 sg13g2_o21ai_1 _15711_ (.B1(_10967_),
    .Y(_00741_),
    .A1(net5119),
    .A2(_10971_));
 sg13g2_nand2_1 _15712_ (.Y(_10972_),
    .A(net1190),
    .B(net5058));
 sg13g2_nand2_1 _15713_ (.Y(_10973_),
    .A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .B(net5319));
 sg13g2_a22oi_1 _15714_ (.Y(_10974_),
    .B1(net342),
    .B2(net5314),
    .A2(net994),
    .A1(net6496));
 sg13g2_nand2_1 _15715_ (.Y(_10975_),
    .A(_10973_),
    .B(_10974_));
 sg13g2_a221oi_1 _15716_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .C1(_10975_),
    .B1(net5112),
    .A1(\soc_inst.mem_ctrl.spi_addr[23] ),
    .Y(_10976_),
    .A2(net5114));
 sg13g2_o21ai_1 _15717_ (.B1(_10972_),
    .Y(_00742_),
    .A1(net5121),
    .A2(_10976_));
 sg13g2_o21ai_1 _15718_ (.B1(net6011),
    .Y(_10977_),
    .A1(net6507),
    .A2(net5568));
 sg13g2_a21oi_1 _15719_ (.A1(\soc_inst.mem_ctrl.spi_addr[16] ),
    .A2(net5568),
    .Y(_10978_),
    .B1(_10977_));
 sg13g2_o21ai_1 _15720_ (.B1(net6010),
    .Y(_10979_),
    .A1(net6507),
    .A2(_10757_));
 sg13g2_a22oi_1 _15721_ (.Y(_10980_),
    .B1(net305),
    .B2(net5318),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .A1(net6500));
 sg13g2_nand2b_1 _15722_ (.Y(_10981_),
    .B(_10980_),
    .A_N(_10979_));
 sg13g2_a221oi_1 _15723_ (.B2(net2335),
    .C1(_10981_),
    .B1(net5113),
    .A1(net2519),
    .Y(_10982_),
    .A2(_10860_));
 sg13g2_nor3_1 _15724_ (.A(net5120),
    .B(_10978_),
    .C(_10982_),
    .Y(_10983_));
 sg13g2_a21o_1 _15725_ (.A2(net5120),
    .A1(net2519),
    .B1(_10983_),
    .X(_00743_));
 sg13g2_nand2_1 _15726_ (.Y(_10984_),
    .A(net880),
    .B(net5121));
 sg13g2_a21oi_1 _15727_ (.A1(\soc_inst.mem_ctrl.spi_addr[17] ),
    .A2(net5568),
    .Y(_10985_),
    .B1(_10977_));
 sg13g2_a21oi_1 _15728_ (.A1(net6500),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .Y(_10986_),
    .B1(_10979_));
 sg13g2_a22oi_1 _15729_ (.Y(_10987_),
    .B1(net5113),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .A2(net5318),
    .A1(net383));
 sg13g2_nand2_1 _15730_ (.Y(_10988_),
    .A(_10986_),
    .B(_10987_));
 sg13g2_a22oi_1 _15731_ (.Y(_10989_),
    .B1(_10988_),
    .B2(_10853_),
    .A2(net5116),
    .A1(net880));
 sg13g2_o21ai_1 _15732_ (.B1(_10984_),
    .Y(_00744_),
    .A1(_10985_),
    .A2(_10989_));
 sg13g2_nand2_1 _15733_ (.Y(_10990_),
    .A(net935),
    .B(net5058));
 sg13g2_a22oi_1 _15734_ (.Y(_10991_),
    .B1(net202),
    .B2(net5318),
    .A2(net880),
    .A1(net6502));
 sg13g2_inv_1 _15735_ (.Y(_10992_),
    .A(_10991_));
 sg13g2_a221oi_1 _15736_ (.B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .C1(_10992_),
    .B1(net5112),
    .A1(\soc_inst.mem_ctrl.spi_addr[18] ),
    .Y(_10993_),
    .A2(net5320));
 sg13g2_o21ai_1 _15737_ (.B1(_10990_),
    .Y(_00745_),
    .A1(net5121),
    .A2(_10993_));
 sg13g2_a21oi_1 _15738_ (.A1(net6502),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .Y(_10994_),
    .B1(_10864_));
 sg13g2_a22oi_1 _15739_ (.Y(_10995_),
    .B1(net5113),
    .B2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .A2(net5318),
    .A1(net332));
 sg13g2_nand2_1 _15740_ (.Y(_10996_),
    .A(_10994_),
    .B(_10995_));
 sg13g2_nand2_1 _15741_ (.Y(_10997_),
    .A(net788),
    .B(net5120));
 sg13g2_nor3_1 _15742_ (.A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .B(_08417_),
    .C(net6009),
    .Y(_10998_));
 sg13g2_a22oi_1 _15743_ (.Y(_10999_),
    .B1(_10996_),
    .B2(_10853_),
    .A2(net5116),
    .A1(net788));
 sg13g2_o21ai_1 _15744_ (.B1(_10997_),
    .Y(_00746_),
    .A1(_10998_),
    .A2(_10999_));
 sg13g2_nor2_1 _15745_ (.A(\soc_inst.mem_ctrl.spi_addr[20] ),
    .B(_08417_),
    .Y(_11000_));
 sg13g2_a22oi_1 _15746_ (.Y(_11001_),
    .B1(net6089),
    .B2(net6507),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ),
    .A1(net6500));
 sg13g2_inv_1 _15747_ (.Y(_11002_),
    .A(_11001_));
 sg13g2_a221oi_1 _15748_ (.B2(net2519),
    .C1(_11002_),
    .B1(net5113),
    .A1(net356),
    .Y(_11003_),
    .A2(net5318));
 sg13g2_o21ai_1 _15749_ (.B1(_11003_),
    .Y(_11004_),
    .A1(_10977_),
    .A2(_11000_));
 sg13g2_a22oi_1 _15750_ (.Y(_11005_),
    .B1(_11004_),
    .B2(_10853_),
    .A2(net5058),
    .A1(net2812));
 sg13g2_inv_1 _15751_ (.Y(_00747_),
    .A(net2813));
 sg13g2_a22oi_1 _15752_ (.Y(_11006_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[29] ),
    .B2(_10863_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .A1(net6500));
 sg13g2_nand2b_1 _15753_ (.Y(_11007_),
    .B(_11006_),
    .A_N(_10864_));
 sg13g2_a221oi_1 _15754_ (.B2(net880),
    .C1(_11007_),
    .B1(net5113),
    .A1(net2736),
    .Y(_11008_),
    .A2(net5116));
 sg13g2_nor3_1 _15755_ (.A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .B(_08417_),
    .C(net6009),
    .Y(_11009_));
 sg13g2_nor3_1 _15756_ (.A(net5120),
    .B(_11008_),
    .C(_11009_),
    .Y(_11010_));
 sg13g2_a21o_1 _15757_ (.A2(net5120),
    .A1(net2736),
    .B1(_11010_),
    .X(_00748_));
 sg13g2_a21oi_1 _15758_ (.A1(\soc_inst.mem_ctrl.spi_addr[22] ),
    .A2(net5568),
    .Y(_11011_),
    .B1(_10977_));
 sg13g2_a22oi_1 _15759_ (.Y(_11012_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[30] ),
    .B2(_10863_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .A1(net6500));
 sg13g2_nand2b_1 _15760_ (.Y(_11013_),
    .B(_11012_),
    .A_N(_10979_));
 sg13g2_a221oi_1 _15761_ (.B2(net935),
    .C1(_11013_),
    .B1(net5113),
    .A1(net2825),
    .Y(_11014_),
    .A2(net5116));
 sg13g2_nor3_1 _15762_ (.A(net5120),
    .B(_11011_),
    .C(_11014_),
    .Y(_11015_));
 sg13g2_a21o_1 _15763_ (.A2(net5120),
    .A1(net2825),
    .B1(_11015_),
    .X(_00749_));
 sg13g2_a21oi_1 _15764_ (.A1(\soc_inst.mem_ctrl.spi_addr[23] ),
    .A2(net5568),
    .Y(_11016_),
    .B1(_10977_));
 sg13g2_a22oi_1 _15765_ (.Y(_11017_),
    .B1(\soc_inst.mem_ctrl.spi_data_in[31] ),
    .B2(_10863_),
    .A2(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ),
    .A1(net6500));
 sg13g2_nand2b_1 _15766_ (.Y(_11018_),
    .B(_11017_),
    .A_N(_10979_));
 sg13g2_a221oi_1 _15767_ (.B2(net788),
    .C1(_11018_),
    .B1(net5113),
    .A1(net2663),
    .Y(_11019_),
    .A2(net5116));
 sg13g2_nor3_1 _15768_ (.A(net5120),
    .B(_11016_),
    .C(_11019_),
    .Y(_11020_));
 sg13g2_a21o_1 _15769_ (.A2(net5121),
    .A1(net2663),
    .B1(_11020_),
    .X(_00750_));
 sg13g2_nand3b_1 _15770_ (.B(_10779_),
    .C(_10780_),
    .Y(_11021_),
    .A_N(net6506));
 sg13g2_and2_1 _15771_ (.A(net6490),
    .B(_11021_),
    .X(_11022_));
 sg13g2_a21oi_1 _15772_ (.A1(net6167),
    .A2(_07875_),
    .Y(_11023_),
    .B1(_11022_));
 sg13g2_nor2_2 _15773_ (.A(net6167),
    .B(net97),
    .Y(_11024_));
 sg13g2_nor2_1 _15774_ (.A(net3399),
    .B(_10774_),
    .Y(_11025_));
 sg13g2_a22oi_1 _15775_ (.Y(_11026_),
    .B1(net5312),
    .B2(net9),
    .A2(net6004),
    .A1(net1237));
 sg13g2_nor2_1 _15776_ (.A(net3284),
    .B(net4802),
    .Y(_11027_));
 sg13g2_a21oi_1 _15777_ (.A1(net4802),
    .A2(_11026_),
    .Y(_00751_),
    .B1(_11027_));
 sg13g2_a22oi_1 _15778_ (.Y(_11028_),
    .B1(net5312),
    .B2(net10),
    .A2(net6004),
    .A1(net1357));
 sg13g2_nor2_1 _15779_ (.A(net3131),
    .B(net4798),
    .Y(_11029_));
 sg13g2_a21oi_1 _15780_ (.A1(net4798),
    .A2(_11028_),
    .Y(_00752_),
    .B1(_11029_));
 sg13g2_a22oi_1 _15781_ (.Y(_11030_),
    .B1(net5313),
    .B2(net11),
    .A2(net6008),
    .A1(net1137));
 sg13g2_nor2_1 _15782_ (.A(net3002),
    .B(net4803),
    .Y(_11031_));
 sg13g2_a21oi_1 _15783_ (.A1(net4803),
    .A2(_11030_),
    .Y(_00753_),
    .B1(_11031_));
 sg13g2_a22oi_1 _15784_ (.Y(_11032_),
    .B1(net5312),
    .B2(net12),
    .A2(net6006),
    .A1(net1039));
 sg13g2_nor2_1 _15785_ (.A(net3127),
    .B(net4800),
    .Y(_11033_));
 sg13g2_a21oi_1 _15786_ (.A1(net4801),
    .A2(_11032_),
    .Y(_00754_),
    .B1(_11033_));
 sg13g2_a22oi_1 _15787_ (.Y(_11034_),
    .B1(net5312),
    .B2(net1237),
    .A2(net6004),
    .A1(net1415));
 sg13g2_nor2_1 _15788_ (.A(net3147),
    .B(net4798),
    .Y(_11035_));
 sg13g2_a21oi_1 _15789_ (.A1(net4798),
    .A2(_11034_),
    .Y(_00755_),
    .B1(_11035_));
 sg13g2_a22oi_1 _15790_ (.Y(_11036_),
    .B1(net5312),
    .B2(net1357),
    .A2(net6004),
    .A1(net1745));
 sg13g2_nor2_1 _15791_ (.A(net3142),
    .B(net4798),
    .Y(_11037_));
 sg13g2_a21oi_1 _15792_ (.A1(net4798),
    .A2(_11036_),
    .Y(_00756_),
    .B1(_11037_));
 sg13g2_a22oi_1 _15793_ (.Y(_11038_),
    .B1(net5313),
    .B2(net1137),
    .A2(net6008),
    .A1(net997));
 sg13g2_nor2_1 _15794_ (.A(net3005),
    .B(net4803),
    .Y(_11039_));
 sg13g2_a21oi_1 _15795_ (.A1(net4803),
    .A2(_11038_),
    .Y(_00757_),
    .B1(_11039_));
 sg13g2_a22oi_1 _15796_ (.Y(_11040_),
    .B1(_11025_),
    .B2(net1039),
    .A2(net6006),
    .A1(net1414));
 sg13g2_nor2_1 _15797_ (.A(net3114),
    .B(net4800),
    .Y(_11041_));
 sg13g2_a21oi_1 _15798_ (.A1(net4801),
    .A2(_11040_),
    .Y(_00758_),
    .B1(_11041_));
 sg13g2_a22oi_1 _15799_ (.Y(_11042_),
    .B1(net5312),
    .B2(net1415),
    .A2(net6005),
    .A1(net1087));
 sg13g2_nor2_1 _15800_ (.A(net3084),
    .B(net4803),
    .Y(_11043_));
 sg13g2_a21oi_1 _15801_ (.A1(net4800),
    .A2(_11042_),
    .Y(_00759_),
    .B1(_11043_));
 sg13g2_a22oi_1 _15802_ (.Y(_11044_),
    .B1(net5312),
    .B2(net1745),
    .A2(net6005),
    .A1(net1228));
 sg13g2_nor2_1 _15803_ (.A(net3046),
    .B(net4803),
    .Y(_11045_));
 sg13g2_a21oi_1 _15804_ (.A1(net4800),
    .A2(_11044_),
    .Y(_00760_),
    .B1(_11045_));
 sg13g2_a22oi_1 _15805_ (.Y(_11046_),
    .B1(net5313),
    .B2(net997),
    .A2(net6008),
    .A1(net1093));
 sg13g2_nor2_1 _15806_ (.A(net2633),
    .B(net4804),
    .Y(_11047_));
 sg13g2_a21oi_1 _15807_ (.A1(net4803),
    .A2(_11046_),
    .Y(_00761_),
    .B1(_11047_));
 sg13g2_a22oi_1 _15808_ (.Y(_11048_),
    .B1(net5313),
    .B2(net1414),
    .A2(net6007),
    .A1(net2023));
 sg13g2_nor2_1 _15809_ (.A(net3069),
    .B(net4805),
    .Y(_11049_));
 sg13g2_a21oi_1 _15810_ (.A1(net4805),
    .A2(_11048_),
    .Y(_00762_),
    .B1(_11049_));
 sg13g2_a22oi_1 _15811_ (.Y(_11050_),
    .B1(net5312),
    .B2(net1087),
    .A2(net6005),
    .A1(net674));
 sg13g2_nor2_1 _15812_ (.A(net3057),
    .B(net4800),
    .Y(_11051_));
 sg13g2_a21oi_1 _15813_ (.A1(net4800),
    .A2(_11050_),
    .Y(_00763_),
    .B1(_11051_));
 sg13g2_a22oi_1 _15814_ (.Y(_11052_),
    .B1(net5313),
    .B2(net1228),
    .A2(net6006),
    .A1(net1122));
 sg13g2_nor2_1 _15815_ (.A(net2870),
    .B(net4804),
    .Y(_11053_));
 sg13g2_a21oi_1 _15816_ (.A1(net4808),
    .A2(_11052_),
    .Y(_00764_),
    .B1(_11053_));
 sg13g2_a22oi_1 _15817_ (.Y(_11054_),
    .B1(net5313),
    .B2(net1093),
    .A2(net6007),
    .A1(net1489));
 sg13g2_nor2_1 _15818_ (.A(net3087),
    .B(net4806),
    .Y(_11055_));
 sg13g2_a21oi_1 _15819_ (.A1(net4806),
    .A2(_11054_),
    .Y(_00765_),
    .B1(_11055_));
 sg13g2_a22oi_1 _15820_ (.Y(_11056_),
    .B1(net5313),
    .B2(net2023),
    .A2(net6007),
    .A1(net1207));
 sg13g2_nor2_1 _15821_ (.A(net3130),
    .B(net4808),
    .Y(_11057_));
 sg13g2_a21oi_1 _15822_ (.A1(net4808),
    .A2(_11056_),
    .Y(_00766_),
    .B1(_11057_));
 sg13g2_mux2_1 _15823_ (.A0(net9),
    .A1(net674),
    .S(net5519),
    .X(_11058_));
 sg13g2_a22oi_1 _15824_ (.Y(_11059_),
    .B1(_11058_),
    .B2(net6167),
    .A2(net6004),
    .A1(net928));
 sg13g2_nor2_1 _15825_ (.A(net2957),
    .B(net4798),
    .Y(_11060_));
 sg13g2_a21oi_1 _15826_ (.A1(net4799),
    .A2(_11059_),
    .Y(_00767_),
    .B1(_11060_));
 sg13g2_mux2_1 _15827_ (.A0(net10),
    .A1(net1122),
    .S(net5519),
    .X(_11061_));
 sg13g2_a22oi_1 _15828_ (.Y(_11062_),
    .B1(_11061_),
    .B2(net6167),
    .A2(net6006),
    .A1(net937));
 sg13g2_nor2_1 _15829_ (.A(net3006),
    .B(net4802),
    .Y(_11063_));
 sg13g2_a21oi_1 _15830_ (.A1(net4809),
    .A2(_11062_),
    .Y(_00768_),
    .B1(_11063_));
 sg13g2_mux2_1 _15831_ (.A0(net11),
    .A1(net1489),
    .S(net5518),
    .X(_11064_));
 sg13g2_a22oi_1 _15832_ (.Y(_11065_),
    .B1(_11064_),
    .B2(_07810_),
    .A2(net6008),
    .A1(net1063));
 sg13g2_nor2_1 _15833_ (.A(net2709),
    .B(net4806),
    .Y(_11066_));
 sg13g2_a21oi_1 _15834_ (.A1(net4806),
    .A2(_11065_),
    .Y(_00769_),
    .B1(_11066_));
 sg13g2_mux2_1 _15835_ (.A0(net12),
    .A1(net1207),
    .S(_10775_),
    .X(_11067_));
 sg13g2_a22oi_1 _15836_ (.Y(_11068_),
    .B1(_11067_),
    .B2(net6166),
    .A2(net6007),
    .A1(net1060));
 sg13g2_nor2_1 _15837_ (.A(net2916),
    .B(net4802),
    .Y(_11069_));
 sg13g2_a21oi_1 _15838_ (.A1(net4802),
    .A2(_11068_),
    .Y(_00770_),
    .B1(_11069_));
 sg13g2_mux2_1 _15839_ (.A0(net1237),
    .A1(net928),
    .S(net5519),
    .X(_11070_));
 sg13g2_a22oi_1 _15840_ (.Y(_11071_),
    .B1(_11070_),
    .B2(net6167),
    .A2(net6004),
    .A1(net943));
 sg13g2_nor2_1 _15841_ (.A(net2981),
    .B(net4799),
    .Y(_11072_));
 sg13g2_a21oi_1 _15842_ (.A1(net4799),
    .A2(_11071_),
    .Y(_00771_),
    .B1(_11072_));
 sg13g2_mux2_1 _15843_ (.A0(net1357),
    .A1(net937),
    .S(net5519),
    .X(_11073_));
 sg13g2_a22oi_1 _15844_ (.Y(_11074_),
    .B1(_11073_),
    .B2(net6167),
    .A2(net6004),
    .A1(net1263));
 sg13g2_nor2_1 _15845_ (.A(net2776),
    .B(net4798),
    .Y(_11075_));
 sg13g2_a21oi_1 _15846_ (.A1(net4799),
    .A2(_11074_),
    .Y(_00772_),
    .B1(_11075_));
 sg13g2_mux2_1 _15847_ (.A0(net1137),
    .A1(net1063),
    .S(net5518),
    .X(_11076_));
 sg13g2_a22oi_1 _15848_ (.Y(_11077_),
    .B1(_11076_),
    .B2(net6166),
    .A2(net6007),
    .A1(net1338));
 sg13g2_nor2_1 _15849_ (.A(net2533),
    .B(net4807),
    .Y(_11078_));
 sg13g2_a21oi_1 _15850_ (.A1(net4807),
    .A2(_11077_),
    .Y(_00773_),
    .B1(_11078_));
 sg13g2_mux2_1 _15851_ (.A0(net1039),
    .A1(net1060),
    .S(net5518),
    .X(_11079_));
 sg13g2_a22oi_1 _15852_ (.Y(_11080_),
    .B1(_11079_),
    .B2(net6166),
    .A2(net6007),
    .A1(net915));
 sg13g2_nor2_1 _15853_ (.A(net2722),
    .B(net4802),
    .Y(_11081_));
 sg13g2_a21oi_1 _15854_ (.A1(net4802),
    .A2(_11080_),
    .Y(_00774_),
    .B1(_11081_));
 sg13g2_nor2_1 _15855_ (.A(net943),
    .B(_10774_),
    .Y(_11082_));
 sg13g2_nor3_1 _15856_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(_10777_),
    .C(_11082_),
    .Y(_11083_));
 sg13g2_a21oi_1 _15857_ (.A1(net888),
    .A2(net6004),
    .Y(_11084_),
    .B1(_11083_));
 sg13g2_nor2_1 _15858_ (.A(net2759),
    .B(net4800),
    .Y(_11085_));
 sg13g2_a21oi_1 _15859_ (.A1(net4800),
    .A2(_11084_),
    .Y(_00775_),
    .B1(_11085_));
 sg13g2_nor2_1 _15860_ (.A(net1263),
    .B(_10774_),
    .Y(_11086_));
 sg13g2_nor3_1 _15861_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(_10776_),
    .C(_11086_),
    .Y(_11087_));
 sg13g2_a21oi_1 _15862_ (.A1(net1411),
    .A2(net6005),
    .Y(_11088_),
    .B1(_11087_));
 sg13g2_nor2_1 _15863_ (.A(net2602),
    .B(net4804),
    .Y(_11089_));
 sg13g2_a21oi_1 _15864_ (.A1(net4804),
    .A2(_11088_),
    .Y(_00776_),
    .B1(_11089_));
 sg13g2_mux2_1 _15865_ (.A0(net997),
    .A1(net1338),
    .S(net5518),
    .X(_11090_));
 sg13g2_a22oi_1 _15866_ (.Y(_11091_),
    .B1(_11090_),
    .B2(net6166),
    .A2(net6008),
    .A1(net1289));
 sg13g2_nor2_1 _15867_ (.A(net2409),
    .B(net4804),
    .Y(_11092_));
 sg13g2_a21oi_1 _15868_ (.A1(net4805),
    .A2(_11091_),
    .Y(_00777_),
    .B1(_11092_));
 sg13g2_mux2_1 _15869_ (.A0(net1414),
    .A1(net915),
    .S(net5518),
    .X(_11093_));
 sg13g2_a22oi_1 _15870_ (.Y(_11094_),
    .B1(_11093_),
    .B2(net6166),
    .A2(net6007),
    .A1(net1174));
 sg13g2_nor2_1 _15871_ (.A(net2507),
    .B(net4806),
    .Y(_11095_));
 sg13g2_a21oi_1 _15872_ (.A1(net4806),
    .A2(_11094_),
    .Y(_00778_),
    .B1(_11095_));
 sg13g2_mux2_1 _15873_ (.A0(net1087),
    .A1(net888),
    .S(net5518),
    .X(_11096_));
 sg13g2_a22oi_1 _15874_ (.Y(_11097_),
    .B1(_11096_),
    .B2(net6166),
    .A2(net6008),
    .A1(net153));
 sg13g2_nor2_1 _15875_ (.A(net2105),
    .B(net4804),
    .Y(_11098_));
 sg13g2_a21oi_1 _15876_ (.A1(net4804),
    .A2(_11097_),
    .Y(_00779_),
    .B1(_11098_));
 sg13g2_mux2_1 _15877_ (.A0(net1228),
    .A1(net1411),
    .S(net5519),
    .X(_11099_));
 sg13g2_a22oi_1 _15878_ (.Y(_11100_),
    .B1(_11099_),
    .B2(net6166),
    .A2(net6008),
    .A1(net247));
 sg13g2_nor2_1 _15879_ (.A(net2410),
    .B(net4804),
    .Y(_11101_));
 sg13g2_a21oi_1 _15880_ (.A1(net4803),
    .A2(_11100_),
    .Y(_00780_),
    .B1(_11101_));
 sg13g2_mux2_1 _15881_ (.A0(net1093),
    .A1(net1289),
    .S(net5518),
    .X(_11102_));
 sg13g2_a22oi_1 _15882_ (.Y(_11103_),
    .B1(_11102_),
    .B2(_07810_),
    .A2(_11024_),
    .A1(net1117));
 sg13g2_nor2_1 _15883_ (.A(net2641),
    .B(net4806),
    .Y(_11104_));
 sg13g2_a21oi_1 _15884_ (.A1(net4807),
    .A2(_11103_),
    .Y(_00781_),
    .B1(_11104_));
 sg13g2_mux2_1 _15885_ (.A0(net2023),
    .A1(net1174),
    .S(net5518),
    .X(_11105_));
 sg13g2_a22oi_1 _15886_ (.Y(_11106_),
    .B1(_11105_),
    .B2(net6166),
    .A2(net6007),
    .A1(net301));
 sg13g2_nor2_1 _15887_ (.A(net2619),
    .B(net4806),
    .Y(_11107_));
 sg13g2_a21oi_1 _15888_ (.A1(net4807),
    .A2(_11106_),
    .Y(_00782_),
    .B1(_11107_));
 sg13g2_nor3_1 _15889_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(net1027),
    .C(net405),
    .Y(_11108_));
 sg13g2_nor2_1 _15890_ (.A(net6142),
    .B(_08414_),
    .Y(_11109_));
 sg13g2_nor3_1 _15891_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ),
    .C(_11109_),
    .Y(_11110_));
 sg13g2_nand2_1 _15892_ (.Y(_11111_),
    .A(_08647_),
    .B(_11110_));
 sg13g2_inv_1 _15893_ (.Y(_11112_),
    .A(_11111_));
 sg13g2_nor3_1 _15894_ (.A(net1134),
    .B(net2659),
    .C(_10758_),
    .Y(_11113_));
 sg13g2_nand2_1 _15895_ (.Y(_11114_),
    .A(net6503),
    .B(_11113_));
 sg13g2_nor4_2 _15896_ (.A(net2273),
    .B(net1077),
    .C(_10847_),
    .Y(_11115_),
    .D(_10848_));
 sg13g2_nor2_1 _15897_ (.A(net6542),
    .B(_11114_),
    .Y(_11116_));
 sg13g2_and3_2 _15898_ (.X(_11117_),
    .A(_11108_),
    .B(_11115_),
    .C(_11116_));
 sg13g2_or2_1 _15899_ (.X(_11118_),
    .B(_11117_),
    .A(net6542));
 sg13g2_nor3_1 _15900_ (.A(net1134),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .C(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .Y(_11119_));
 sg13g2_nor3_1 _15901_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .C(_08419_),
    .Y(_11120_));
 sg13g2_nand4_1 _15902_ (.B(_11108_),
    .C(_11119_),
    .A(_10849_),
    .Y(_11121_),
    .D(_11120_));
 sg13g2_o21ai_1 _15903_ (.B1(_11121_),
    .Y(_11122_),
    .A1(_11108_),
    .A2(_11112_));
 sg13g2_nand2_1 _15904_ (.Y(_11123_),
    .A(net2141),
    .B(_11117_));
 sg13g2_o21ai_1 _15905_ (.B1(_11123_),
    .Y(_00783_),
    .A1(_11118_),
    .A2(_11122_));
 sg13g2_nand3_1 _15906_ (.B(_07875_),
    .C(net6503),
    .A(net3281),
    .Y(_11124_));
 sg13g2_nand3_1 _15907_ (.B(_11021_),
    .C(_11124_),
    .A(net6167),
    .Y(_00784_));
 sg13g2_o21ai_1 _15908_ (.B1(_11115_),
    .Y(_11125_),
    .A1(_11111_),
    .A2(_11114_));
 sg13g2_nor2b_1 _15909_ (.A(_11118_),
    .B_N(_11125_),
    .Y(_11126_));
 sg13g2_a21o_1 _15910_ (.A2(_11117_),
    .A1(net2874),
    .B1(_11126_),
    .X(_00785_));
 sg13g2_a21oi_1 _15911_ (.A1(_08974_),
    .A2(_09594_),
    .Y(_11127_),
    .B1(_09002_));
 sg13g2_and3_1 _15912_ (.X(_11128_),
    .A(_08981_),
    .B(_09030_),
    .C(_11127_));
 sg13g2_nor2b_1 _15913_ (.A(net5332),
    .B_N(_09594_),
    .Y(_11129_));
 sg13g2_or4_1 _15914_ (.A(_08982_),
    .B(_09002_),
    .C(_09044_),
    .D(_11129_),
    .X(_11130_));
 sg13g2_a21oi_1 _15915_ (.A1(_09898_),
    .A2(net4796),
    .Y(_11131_),
    .B1(net270));
 sg13g2_a21oi_1 _15916_ (.A1(net6173),
    .A2(_09898_),
    .Y(_11132_),
    .B1(_09895_));
 sg13g2_nor2_1 _15917_ (.A(_09513_),
    .B(_11130_),
    .Y(_11133_));
 sg13g2_nand2b_2 _15918_ (.Y(_11134_),
    .B(_09514_),
    .A_N(_11130_));
 sg13g2_a21oi_1 _15919_ (.A1(_11132_),
    .A2(net4727),
    .Y(_00786_),
    .B1(net271));
 sg13g2_a21oi_1 _15920_ (.A1(_09903_),
    .A2(net4795),
    .Y(_11135_),
    .B1(net140));
 sg13g2_a21oi_1 _15921_ (.A1(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .A2(_08987_),
    .Y(_11136_),
    .B1(_09901_));
 sg13g2_a21oi_1 _15922_ (.A1(net4727),
    .A2(_11136_),
    .Y(_00787_),
    .B1(net141));
 sg13g2_nor2b_2 _15923_ (.A(net6294),
    .B_N(net2390),
    .Y(_11137_));
 sg13g2_a21oi_1 _15924_ (.A1(net4795),
    .A2(_11137_),
    .Y(_11138_),
    .B1(net194));
 sg13g2_o21ai_1 _15925_ (.B1(net6023),
    .Y(_11139_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .A2(net6019));
 sg13g2_a21oi_1 _15926_ (.A1(net6172),
    .A2(_11137_),
    .Y(_11140_),
    .B1(_11139_));
 sg13g2_a21oi_1 _15927_ (.A1(net4728),
    .A2(_11140_),
    .Y(_00788_),
    .B1(net195));
 sg13g2_a21oi_1 _15928_ (.A1(_09907_),
    .A2(net4796),
    .Y(_11141_),
    .B1(net222));
 sg13g2_a21oi_1 _15929_ (.A1(net6173),
    .A2(_09907_),
    .Y(_11142_),
    .B1(_09905_));
 sg13g2_a21oi_1 _15930_ (.A1(net4727),
    .A2(_11142_),
    .Y(_00789_),
    .B1(net223));
 sg13g2_a21oi_1 _15931_ (.A1(_09911_),
    .A2(net4797),
    .Y(_11143_),
    .B1(net131));
 sg13g2_a21oi_1 _15932_ (.A1(net6173),
    .A2(_09911_),
    .Y(_11144_),
    .B1(_09909_));
 sg13g2_a21oi_1 _15933_ (.A1(net4728),
    .A2(_11144_),
    .Y(_00790_),
    .B1(net132));
 sg13g2_a21oi_1 _15934_ (.A1(_09915_),
    .A2(net4797),
    .Y(_11145_),
    .B1(net134));
 sg13g2_a21oi_1 _15935_ (.A1(net6173),
    .A2(_09915_),
    .Y(_11146_),
    .B1(_09913_));
 sg13g2_a21oi_1 _15936_ (.A1(net4728),
    .A2(_11146_),
    .Y(_00791_),
    .B1(net135));
 sg13g2_nor2b_2 _15937_ (.A(net6294),
    .B_N(net1582),
    .Y(_11147_));
 sg13g2_a21oi_1 _15938_ (.A1(net4795),
    .A2(_11147_),
    .Y(_11148_),
    .B1(net280));
 sg13g2_o21ai_1 _15939_ (.B1(net6023),
    .Y(_11149_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .A2(net6019));
 sg13g2_a21oi_1 _15940_ (.A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .A2(_08987_),
    .Y(_11150_),
    .B1(_11149_));
 sg13g2_a21oi_1 _15941_ (.A1(net4727),
    .A2(_11150_),
    .Y(_00792_),
    .B1(net281));
 sg13g2_nor2b_2 _15942_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .Y(_11151_));
 sg13g2_a21oi_1 _15943_ (.A1(net4793),
    .A2(_11151_),
    .Y(_11152_),
    .B1(net137));
 sg13g2_o21ai_1 _15944_ (.B1(net6021),
    .Y(_11153_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .A2(net6019));
 sg13g2_a21oi_1 _15945_ (.A1(net6170),
    .A2(_11151_),
    .Y(_11154_),
    .B1(_11153_));
 sg13g2_a21oi_1 _15946_ (.A1(net4728),
    .A2(_11154_),
    .Y(_00793_),
    .B1(net138));
 sg13g2_nor2b_2 _15947_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .Y(_11155_));
 sg13g2_a21oi_1 _15948_ (.A1(net4793),
    .A2(_11155_),
    .Y(_11156_),
    .B1(net423));
 sg13g2_o21ai_1 _15949_ (.B1(net6021),
    .Y(_11157_),
    .A1(net1452),
    .A2(net6018));
 sg13g2_a21oi_1 _15950_ (.A1(net6170),
    .A2(_11155_),
    .Y(_11158_),
    .B1(_11157_));
 sg13g2_a21oi_1 _15951_ (.A1(net4726),
    .A2(_11158_),
    .Y(_00794_),
    .B1(net424));
 sg13g2_nor2b_2 _15952_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .Y(_11159_));
 sg13g2_a21oi_1 _15953_ (.A1(net4794),
    .A2(_11159_),
    .Y(_11160_),
    .B1(net235));
 sg13g2_o21ai_1 _15954_ (.B1(net6022),
    .Y(_11161_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15955_ (.A1(net6170),
    .A2(_11159_),
    .Y(_11162_),
    .B1(_11161_));
 sg13g2_a21oi_1 _15956_ (.A1(net4727),
    .A2(_11162_),
    .Y(_00795_),
    .B1(net236));
 sg13g2_nor2b_2 _15957_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .Y(_11163_));
 sg13g2_a21oi_1 _15958_ (.A1(net4793),
    .A2(_11163_),
    .Y(_11164_),
    .B1(net126));
 sg13g2_o21ai_1 _15959_ (.B1(net6021),
    .Y(_11165_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .A2(net6018));
 sg13g2_a21oi_1 _15960_ (.A1(net6170),
    .A2(_11163_),
    .Y(_11166_),
    .B1(_11165_));
 sg13g2_a21oi_1 _15961_ (.A1(net4726),
    .A2(_11166_),
    .Y(_00796_),
    .B1(net127));
 sg13g2_nor2b_2 _15962_ (.A(net6292),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .Y(_11167_));
 sg13g2_a21oi_1 _15963_ (.A1(net4794),
    .A2(_11167_),
    .Y(_11168_),
    .B1(net283));
 sg13g2_o21ai_1 _15964_ (.B1(net6021),
    .Y(_11169_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15965_ (.A1(net6171),
    .A2(_11167_),
    .Y(_11170_),
    .B1(_11169_));
 sg13g2_a21oi_1 _15966_ (.A1(net4726),
    .A2(_11170_),
    .Y(_00797_),
    .B1(net284));
 sg13g2_nor2b_2 _15967_ (.A(net6292),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .Y(_11171_));
 sg13g2_a21oi_1 _15968_ (.A1(net4793),
    .A2(_11171_),
    .Y(_11172_),
    .B1(net726));
 sg13g2_o21ai_1 _15969_ (.B1(net6022),
    .Y(_11173_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15970_ (.A1(net6171),
    .A2(_11171_),
    .Y(_11174_),
    .B1(_11173_));
 sg13g2_a21oi_1 _15971_ (.A1(net4726),
    .A2(_11174_),
    .Y(_00798_),
    .B1(net727));
 sg13g2_nor2b_2 _15972_ (.A(net6292),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .Y(_11175_));
 sg13g2_a21oi_1 _15973_ (.A1(net4794),
    .A2(_11175_),
    .Y(_11176_),
    .B1(net148));
 sg13g2_o21ai_1 _15974_ (.B1(net6022),
    .Y(_11177_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15975_ (.A1(net6171),
    .A2(_11175_),
    .Y(_11178_),
    .B1(_11177_));
 sg13g2_a21oi_1 _15976_ (.A1(net4727),
    .A2(_11178_),
    .Y(_00799_),
    .B1(net149));
 sg13g2_nor2b_2 _15977_ (.A(net6292),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .Y(_11179_));
 sg13g2_a21oi_1 _15978_ (.A1(net4793),
    .A2(_11179_),
    .Y(_11180_),
    .B1(net191));
 sg13g2_o21ai_1 _15979_ (.B1(net6022),
    .Y(_11181_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15980_ (.A1(net6171),
    .A2(_11179_),
    .Y(_11182_),
    .B1(_11181_));
 sg13g2_a21oi_1 _15981_ (.A1(net4726),
    .A2(_11182_),
    .Y(_00800_),
    .B1(net192));
 sg13g2_nor2b_2 _15982_ (.A(net6292),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .Y(_11183_));
 sg13g2_a21oi_1 _15983_ (.A1(net4794),
    .A2(_11183_),
    .Y(_11184_),
    .B1(net169));
 sg13g2_o21ai_1 _15984_ (.B1(net6021),
    .Y(_11185_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .A2(net6020));
 sg13g2_a21oi_1 _15985_ (.A1(net6170),
    .A2(_11183_),
    .Y(_11186_),
    .B1(_11185_));
 sg13g2_a21oi_1 _15986_ (.A1(net4727),
    .A2(_11186_),
    .Y(_00801_),
    .B1(net170));
 sg13g2_nor2b_2 _15987_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .Y(_11187_));
 sg13g2_a21oi_1 _15988_ (.A1(net4793),
    .A2(_11187_),
    .Y(_11188_),
    .B1(net197));
 sg13g2_o21ai_1 _15989_ (.B1(net6021),
    .Y(_11189_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .A2(net6018));
 sg13g2_a21oi_1 _15990_ (.A1(net6170),
    .A2(_11187_),
    .Y(_11190_),
    .B1(_11189_));
 sg13g2_a21oi_1 _15991_ (.A1(net4726),
    .A2(_11190_),
    .Y(_00802_),
    .B1(net198));
 sg13g2_nor2b_2 _15992_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .Y(_11191_));
 sg13g2_a21oi_1 _15993_ (.A1(net4793),
    .A2(_11191_),
    .Y(_11192_),
    .B1(net176));
 sg13g2_o21ai_1 _15994_ (.B1(net6021),
    .Y(_11193_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .A2(net6017));
 sg13g2_a21oi_1 _15995_ (.A1(net6170),
    .A2(_11191_),
    .Y(_11194_),
    .B1(_11193_));
 sg13g2_a21oi_1 _15996_ (.A1(net4726),
    .A2(_11194_),
    .Y(_00803_),
    .B1(net177));
 sg13g2_nor2b_2 _15997_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .Y(_11195_));
 sg13g2_a21oi_1 _15998_ (.A1(net4793),
    .A2(_11195_),
    .Y(_11196_),
    .B1(net277));
 sg13g2_o21ai_1 _15999_ (.B1(net6021),
    .Y(_11197_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .A2(net6018));
 sg13g2_a21oi_1 _16000_ (.A1(net6170),
    .A2(_11195_),
    .Y(_11198_),
    .B1(_11197_));
 sg13g2_a21oi_1 _16001_ (.A1(net4726),
    .A2(_11198_),
    .Y(_00804_),
    .B1(net278));
 sg13g2_nand2_1 _16002_ (.Y(_11199_),
    .A(net749),
    .B(net4723));
 sg13g2_nor2b_1 _16003_ (.A(net6289),
    .B_N(net2674),
    .Y(_11200_));
 sg13g2_a21o_1 _16004_ (.A2(_10271_),
    .A1(net749),
    .B1(_11200_),
    .X(_11201_));
 sg13g2_nor2_1 _16005_ (.A(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .B(net6017),
    .Y(_11202_));
 sg13g2_o21ai_1 _16006_ (.B1(_11201_),
    .Y(_11203_),
    .A1(net6016),
    .A2(_11202_));
 sg13g2_o21ai_1 _16007_ (.B1(_11199_),
    .Y(_00805_),
    .A1(net4723),
    .A2(_11203_));
 sg13g2_nand2_1 _16008_ (.Y(_11204_),
    .A(net580),
    .B(net4725));
 sg13g2_nor2b_1 _16009_ (.A(net6289),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .Y(_11205_));
 sg13g2_a21o_1 _16010_ (.A2(_10271_),
    .A1(net580),
    .B1(_11205_),
    .X(_11206_));
 sg13g2_nor2_1 _16011_ (.A(net2145),
    .B(net6017),
    .Y(_11207_));
 sg13g2_o21ai_1 _16012_ (.B1(_11206_),
    .Y(_11208_),
    .A1(_09921_),
    .A2(_11207_));
 sg13g2_o21ai_1 _16013_ (.B1(_11204_),
    .Y(_00806_),
    .A1(net4725),
    .A2(_11208_));
 sg13g2_nand2_1 _16014_ (.Y(_11209_),
    .A(net553),
    .B(net4723));
 sg13g2_nor2b_1 _16015_ (.A(net6289),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .Y(_11210_));
 sg13g2_a21o_1 _16016_ (.A2(_10271_),
    .A1(net553),
    .B1(_11210_),
    .X(_11211_));
 sg13g2_nor2_1 _16017_ (.A(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .B(net6017),
    .Y(_11212_));
 sg13g2_o21ai_1 _16018_ (.B1(_11211_),
    .Y(_11213_),
    .A1(net6016),
    .A2(_11212_));
 sg13g2_o21ai_1 _16019_ (.B1(_11209_),
    .Y(_00807_),
    .A1(net4723),
    .A2(_11213_));
 sg13g2_nand2_1 _16020_ (.Y(_11214_),
    .A(net385),
    .B(net4724));
 sg13g2_nor2b_1 _16021_ (.A(net6289),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .Y(_11215_));
 sg13g2_a21o_1 _16022_ (.A2(_10271_),
    .A1(net385),
    .B1(_11215_),
    .X(_11216_));
 sg13g2_nor2_1 _16023_ (.A(net1591),
    .B(net6017),
    .Y(_11217_));
 sg13g2_o21ai_1 _16024_ (.B1(_11216_),
    .Y(_11218_),
    .A1(net6016),
    .A2(_11217_));
 sg13g2_o21ai_1 _16025_ (.B1(_11214_),
    .Y(_00808_),
    .A1(net4724),
    .A2(_11218_));
 sg13g2_nand2_1 _16026_ (.Y(_11219_),
    .A(net1152),
    .B(net4723));
 sg13g2_nor2b_1 _16027_ (.A(net6291),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .Y(_11220_));
 sg13g2_a21o_1 _16028_ (.A2(_10271_),
    .A1(net1152),
    .B1(_11220_),
    .X(_11221_));
 sg13g2_nor2_1 _16029_ (.A(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .B(net6017),
    .Y(_11222_));
 sg13g2_o21ai_1 _16030_ (.B1(_11221_),
    .Y(_11223_),
    .A1(net6016),
    .A2(_11222_));
 sg13g2_o21ai_1 _16031_ (.B1(_11219_),
    .Y(_00809_),
    .A1(net4723),
    .A2(_11223_));
 sg13g2_nand2_1 _16032_ (.Y(_11224_),
    .A(net482),
    .B(net4723));
 sg13g2_nor2b_1 _16033_ (.A(net6289),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .Y(_11225_));
 sg13g2_a21o_1 _16034_ (.A2(_10271_),
    .A1(net482),
    .B1(_11225_),
    .X(_11226_));
 sg13g2_nor2_1 _16035_ (.A(net2672),
    .B(net6017),
    .Y(_11227_));
 sg13g2_o21ai_1 _16036_ (.B1(_11226_),
    .Y(_11228_),
    .A1(net6016),
    .A2(_11227_));
 sg13g2_o21ai_1 _16037_ (.B1(_11224_),
    .Y(_00810_),
    .A1(net4723),
    .A2(_11228_));
 sg13g2_nand2_1 _16038_ (.Y(_11229_),
    .A(net541),
    .B(net4724));
 sg13g2_nor2b_1 _16039_ (.A(net6289),
    .B_N(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .Y(_11230_));
 sg13g2_a21o_1 _16040_ (.A2(_10271_),
    .A1(net541),
    .B1(_11230_),
    .X(_11231_));
 sg13g2_nor2_1 _16041_ (.A(net1348),
    .B(net6017),
    .Y(_11232_));
 sg13g2_o21ai_1 _16042_ (.B1(_11231_),
    .Y(_11233_),
    .A1(net6016),
    .A2(_11232_));
 sg13g2_o21ai_1 _16043_ (.B1(_11229_),
    .Y(_00811_),
    .A1(net4724),
    .A2(_11233_));
 sg13g2_a22oi_1 _16044_ (.Y(_11234_),
    .B1(_10271_),
    .B2(net1709),
    .A2(net1398),
    .A1(net6168));
 sg13g2_o21ai_1 _16045_ (.B1(net6024),
    .Y(_11235_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .A2(net6019));
 sg13g2_nor2_1 _16046_ (.A(net6016),
    .B(_11235_),
    .Y(_11236_));
 sg13g2_nor3_1 _16047_ (.A(net4725),
    .B(_11234_),
    .C(_11236_),
    .Y(_11237_));
 sg13g2_a21o_1 _16048_ (.A2(net4725),
    .A1(net1709),
    .B1(_11237_),
    .X(_00812_));
 sg13g2_nand2_1 _16049_ (.Y(_11238_),
    .A(net6488),
    .B(net6142));
 sg13g2_nor4_1 _16050_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .B(net6488),
    .C(net6490),
    .D(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .Y(_11239_));
 sg13g2_nand3_1 _16051_ (.B(_11113_),
    .C(_11239_),
    .A(net6503),
    .Y(_11240_));
 sg13g2_o21ai_1 _16052_ (.B1(_11238_),
    .Y(_11241_),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .A2(_11240_));
 sg13g2_nand4_1 _16053_ (.B(_07879_),
    .C(_08412_),
    .A(net6488),
    .Y(_11242_),
    .D(_08413_));
 sg13g2_nand2_1 _16054_ (.Y(_11243_),
    .A(_08419_),
    .B(_11239_));
 sg13g2_nand2_1 _16055_ (.Y(_11244_),
    .A(net6490),
    .B(net6506));
 sg13g2_nor2b_1 _16056_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .B_N(_11113_),
    .Y(_11245_));
 sg13g2_nand4_1 _16057_ (.B(_11243_),
    .C(_11244_),
    .A(_11242_),
    .Y(_11246_),
    .D(_11245_));
 sg13g2_mux2_1 _16058_ (.A0(_11246_),
    .A1(net3382),
    .S(_11241_),
    .X(_11247_));
 sg13g2_nor2b_1 _16059_ (.A(net6541),
    .B_N(net3383),
    .Y(_00813_));
 sg13g2_or2_1 _16060_ (.X(_00814_),
    .B(net405),
    .A(net1309));
 sg13g2_nor2_1 _16061_ (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .B(net6500),
    .Y(_11248_));
 sg13g2_a21oi_1 _16062_ (.A1(_08648_),
    .A2(_11248_),
    .Y(_11249_),
    .B1(net6482));
 sg13g2_nand4_1 _16063_ (.B(_07876_),
    .C(net6503),
    .A(net6167),
    .Y(_11250_),
    .D(_10757_));
 sg13g2_or4_1 _16064_ (.A(net6488),
    .B(_10847_),
    .C(_10848_),
    .D(_11250_),
    .X(_11251_));
 sg13g2_nor4_1 _16065_ (.A(net1134),
    .B(net2882),
    .C(net2273),
    .D(_11251_),
    .Y(_11252_));
 sg13g2_nor2_1 _16066_ (.A(net6488),
    .B(net1027),
    .Y(_11253_));
 sg13g2_a21o_2 _16067_ (.A2(_11253_),
    .A1(_11252_),
    .B1(_11249_),
    .X(_11254_));
 sg13g2_mux2_1 _16068_ (.A0(net6201),
    .A1(net6202),
    .S(net6486),
    .X(_11255_));
 sg13g2_nand2_1 _16069_ (.Y(_11256_),
    .A(_11252_),
    .B(_11255_));
 sg13g2_a21oi_1 _16070_ (.A1(net6490),
    .A2(net6506),
    .Y(_11257_),
    .B1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ));
 sg13g2_and2_1 _16071_ (.A(_07882_),
    .B(_11257_),
    .X(_11258_));
 sg13g2_nand2_2 _16072_ (.Y(_11259_),
    .A(_07882_),
    .B(_11257_));
 sg13g2_mux2_1 _16073_ (.A0(uio_out[1]),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .S(net6483),
    .X(_11260_));
 sg13g2_a22oi_1 _16074_ (.Y(_11261_),
    .B1(_11259_),
    .B2(_11260_),
    .A2(net2663),
    .A1(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ));
 sg13g2_a21oi_1 _16075_ (.A1(_11256_),
    .A2(_11261_),
    .Y(_11262_),
    .B1(_11254_));
 sg13g2_a21o_1 _16076_ (.A2(_11254_),
    .A1(net2988),
    .B1(_11262_),
    .X(_00815_));
 sg13g2_and2_1 _16077_ (.A(_11242_),
    .B(_11256_),
    .X(_11263_));
 sg13g2_mux2_1 _16078_ (.A0(net2991),
    .A1(net2736),
    .S(net6483),
    .X(_11264_));
 sg13g2_a21oi_1 _16079_ (.A1(_11259_),
    .A2(_11264_),
    .Y(_11265_),
    .B1(_11254_));
 sg13g2_a22oi_1 _16080_ (.Y(_00816_),
    .B1(_11263_),
    .B2(_11265_),
    .A2(_11254_),
    .A1(_08221_));
 sg13g2_nor2_1 _16081_ (.A(net6483),
    .B(net3066),
    .Y(_11266_));
 sg13g2_o21ai_1 _16082_ (.B1(_11259_),
    .Y(_11267_),
    .A1(net6142),
    .A2(net2825));
 sg13g2_o21ai_1 _16083_ (.B1(_11256_),
    .Y(_11268_),
    .A1(_11266_),
    .A2(_11267_));
 sg13g2_mux2_1 _16084_ (.A0(_11268_),
    .A1(net3066),
    .S(_11254_),
    .X(_00817_));
 sg13g2_mux2_1 _16085_ (.A0(net2862),
    .A1(net2663),
    .S(net6483),
    .X(_11269_));
 sg13g2_a21oi_1 _16086_ (.A1(_11259_),
    .A2(_11269_),
    .Y(_11270_),
    .B1(_11254_));
 sg13g2_a22oi_1 _16087_ (.Y(_00818_),
    .B1(_11263_),
    .B2(_11270_),
    .A2(_11254_),
    .A1(_08222_));
 sg13g2_nor3_1 _16088_ (.A(net6193),
    .B(_08247_),
    .C(_09820_),
    .Y(_11271_));
 sg13g2_nor3_1 _16089_ (.A(net5195),
    .B(_08293_),
    .C(_11271_),
    .Y(_11272_));
 sg13g2_nand2_1 _16090_ (.Y(_11273_),
    .A(_10706_),
    .B(_11272_));
 sg13g2_nor4_1 _16091_ (.A(net2751),
    .B(net6193),
    .C(_08246_),
    .D(_11273_),
    .Y(_11274_));
 sg13g2_a21o_1 _16092_ (.A2(_11273_),
    .A1(net6504),
    .B1(_11274_),
    .X(_00819_));
 sg13g2_a21oi_1 _16093_ (.A1(net6302),
    .A2(net2723),
    .Y(_11275_),
    .B1(_09071_));
 sg13g2_nand4_1 _16094_ (.B(net5156),
    .C(net6105),
    .A(net2723),
    .Y(_11276_),
    .D(_09070_));
 sg13g2_o21ai_1 _16095_ (.B1(_11276_),
    .Y(_11277_),
    .A1(_09067_),
    .A2(_11275_));
 sg13g2_mux2_1 _16096_ (.A0(net2723),
    .A1(_11277_),
    .S(net4792),
    .X(_00820_));
 sg13g2_a21oi_1 _16097_ (.A1(net6301),
    .A2(net2745),
    .Y(_11278_),
    .B1(_09083_));
 sg13g2_nand4_1 _16098_ (.B(net5155),
    .C(net6105),
    .A(net2745),
    .Y(_11279_),
    .D(_09082_));
 sg13g2_o21ai_1 _16099_ (.B1(_11279_),
    .Y(_11280_),
    .A1(_09067_),
    .A2(_11278_));
 sg13g2_mux2_1 _16100_ (.A0(net2745),
    .A1(_11280_),
    .S(net4792),
    .X(_00821_));
 sg13g2_nand4_1 _16101_ (.B(net5157),
    .C(net6105),
    .A(net2773),
    .Y(_11281_),
    .D(_09091_));
 sg13g2_a21oi_1 _16102_ (.A1(net6302),
    .A2(net2773),
    .Y(_11282_),
    .B1(_09092_));
 sg13g2_o21ai_1 _16103_ (.B1(_11281_),
    .Y(_11283_),
    .A1(_09067_),
    .A2(_11282_));
 sg13g2_mux2_1 _16104_ (.A0(net2773),
    .A1(_11283_),
    .S(net4792),
    .X(_00822_));
 sg13g2_a21oi_1 _16105_ (.A1(net6302),
    .A2(net2784),
    .Y(_11284_),
    .B1(_09109_));
 sg13g2_nand4_1 _16106_ (.B(net5156),
    .C(_09049_),
    .A(net2784),
    .Y(_11285_),
    .D(_09108_));
 sg13g2_o21ai_1 _16107_ (.B1(_11285_),
    .Y(_11286_),
    .A1(_09067_),
    .A2(_11284_));
 sg13g2_mux2_1 _16108_ (.A0(net2784),
    .A1(_11286_),
    .S(_09038_),
    .X(_00823_));
 sg13g2_nor2_1 _16109_ (.A(net2432),
    .B(net1860),
    .Y(_11287_));
 sg13g2_nand3b_1 _16110_ (.B(net2406),
    .C(_11287_),
    .Y(_11288_),
    .A_N(net2746));
 sg13g2_nand3_1 _16111_ (.B(net6487),
    .C(_11288_),
    .A(net2919),
    .Y(_11289_));
 sg13g2_and2_1 _16112_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .B(_10274_),
    .X(_11290_));
 sg13g2_nand2_1 _16113_ (.Y(_11291_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .B(_10274_));
 sg13g2_nand4_1 _16114_ (.B(_07782_),
    .C(net6487),
    .A(net2746),
    .Y(_11292_),
    .D(_11287_));
 sg13g2_nand3_1 _16115_ (.B(net6003),
    .C(_11292_),
    .A(_11289_),
    .Y(_11293_));
 sg13g2_nand2_1 _16116_ (.Y(_11294_),
    .A(net6549),
    .B(_11293_));
 sg13g2_nor2_1 _16117_ (.A(_07799_),
    .B(net6487),
    .Y(_11295_));
 sg13g2_nand2b_1 _16118_ (.Y(_11296_),
    .B(net2919),
    .A_N(net6487));
 sg13g2_xnor2_1 _16119_ (.Y(_11297_),
    .A(_00317_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ));
 sg13g2_xor2_1 _16120_ (.B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .X(_11298_));
 sg13g2_xor2_1 _16121_ (.B(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .X(_11299_));
 sg13g2_nand2b_1 _16122_ (.Y(_11300_),
    .B(net6175),
    .A_N(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ));
 sg13g2_nand2b_1 _16123_ (.Y(_11301_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .A_N(net6175));
 sg13g2_or2_1 _16124_ (.X(_11302_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ),
    .A(_00316_));
 sg13g2_o21ai_1 _16125_ (.B1(_11300_),
    .Y(_11303_),
    .A1(_00315_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ));
 sg13g2_a221oi_1 _16126_ (.B2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .C1(_11303_),
    .B1(_07803_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .Y(_11304_),
    .A2(_07801_));
 sg13g2_o21ai_1 _16127_ (.B1(_11301_),
    .Y(_11305_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .A2(_07800_));
 sg13g2_a221oi_1 _16128_ (.B2(_07781_),
    .C1(_11305_),
    .B1(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .A1(_00316_),
    .Y(_11306_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ));
 sg13g2_xnor2_1 _16129_ (.Y(_11307_),
    .A(_00318_),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ));
 sg13g2_nor4_1 _16130_ (.A(_11297_),
    .B(_11298_),
    .C(_11299_),
    .D(_11307_),
    .Y(_11308_));
 sg13g2_o21ai_1 _16131_ (.B1(_11302_),
    .Y(_11309_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .A2(_07801_));
 sg13g2_a221oi_1 _16132_ (.B2(_07800_),
    .C1(_11309_),
    .B1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .A1(_00315_),
    .Y(_11310_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ));
 sg13g2_and4_1 _16133_ (.A(_11304_),
    .B(_11306_),
    .C(_11308_),
    .D(_11310_),
    .X(_11311_));
 sg13g2_nand2b_1 _16134_ (.Y(_11312_),
    .B(net6553),
    .A_N(_11311_));
 sg13g2_o21ai_1 _16135_ (.B1(_11294_),
    .Y(_00824_),
    .A1(net2920),
    .A2(net5108));
 sg13g2_nor2b_2 _16136_ (.A(net2919),
    .B_N(net6487),
    .Y(_11313_));
 sg13g2_a21oi_1 _16137_ (.A1(_11295_),
    .A2(_11311_),
    .Y(_11314_),
    .B1(_11313_));
 sg13g2_a21oi_1 _16138_ (.A1(_11289_),
    .A2(_11314_),
    .Y(_00825_),
    .B1(_07884_));
 sg13g2_nor2_1 _16139_ (.A(net1488),
    .B(net4795),
    .Y(_11315_));
 sg13g2_nand2b_1 _16140_ (.Y(_11316_),
    .B(_09070_),
    .A_N(net1488));
 sg13g2_a21oi_1 _16141_ (.A1(_09073_),
    .A2(_11316_),
    .Y(_11317_),
    .B1(_09927_));
 sg13g2_a21oi_1 _16142_ (.A1(net4795),
    .A2(_11317_),
    .Y(_00826_),
    .B1(_11315_));
 sg13g2_nor2_1 _16143_ (.A(net1805),
    .B(net4795),
    .Y(_11318_));
 sg13g2_nand2b_1 _16144_ (.Y(_11319_),
    .B(_09082_),
    .A_N(net1805));
 sg13g2_a21oi_1 _16145_ (.A1(_09085_),
    .A2(_11319_),
    .Y(_11320_),
    .B1(_09931_));
 sg13g2_a21oi_1 _16146_ (.A1(net4795),
    .A2(_11320_),
    .Y(_00827_),
    .B1(_11318_));
 sg13g2_nor2_1 _16147_ (.A(net1783),
    .B(net4796),
    .Y(_11321_));
 sg13g2_nand2b_1 _16148_ (.Y(_11322_),
    .B(_09091_),
    .A_N(net1783));
 sg13g2_a21oi_1 _16149_ (.A1(_09093_),
    .A2(_11322_),
    .Y(_11323_),
    .B1(_09935_));
 sg13g2_a21oi_1 _16150_ (.A1(net4796),
    .A2(_11323_),
    .Y(_00828_),
    .B1(_11321_));
 sg13g2_a21oi_1 _16151_ (.A1(_09052_),
    .A2(net4796),
    .Y(_11324_),
    .B1(net162));
 sg13g2_a21oi_1 _16152_ (.A1(_09055_),
    .A2(net4796),
    .Y(_00829_),
    .B1(_11324_));
 sg13g2_nor2_1 _16153_ (.A(net1731),
    .B(net4796),
    .Y(_11325_));
 sg13g2_nand2b_1 _16154_ (.Y(_11326_),
    .B(_09108_),
    .A_N(net1731));
 sg13g2_a21oi_1 _16155_ (.A1(_09111_),
    .A2(_11326_),
    .Y(_11327_),
    .B1(_09940_));
 sg13g2_a21oi_1 _16156_ (.A1(net4795),
    .A2(_11327_),
    .Y(_00830_),
    .B1(_11325_));
 sg13g2_nand2_1 _16157_ (.Y(_11328_),
    .A(_11115_),
    .B(_11253_));
 sg13g2_o21ai_1 _16158_ (.B1(_09366_),
    .Y(_11329_),
    .A1(_11250_),
    .A2(_11328_));
 sg13g2_inv_1 _16159_ (.Y(_11330_),
    .A(_11329_));
 sg13g2_o21ai_1 _16160_ (.B1(_11330_),
    .Y(_11331_),
    .A1(_08666_),
    .A2(_10780_));
 sg13g2_nand2_2 _16161_ (.Y(_11332_),
    .A(_08627_),
    .B(_08660_));
 sg13g2_o21ai_1 _16162_ (.B1(_07874_),
    .Y(_11333_),
    .A1(net6506),
    .A2(_11332_));
 sg13g2_nor2_1 _16163_ (.A(net6490),
    .B(_11332_),
    .Y(_11334_));
 sg13g2_nor2_1 _16164_ (.A(net6486),
    .B(_08665_),
    .Y(_11335_));
 sg13g2_a221oi_1 _16165_ (.B2(net6142),
    .C1(_11334_),
    .B1(_11335_),
    .A1(net6486),
    .Y(_11336_),
    .A2(_11333_));
 sg13g2_inv_1 _16166_ (.Y(_11337_),
    .A(_11336_));
 sg13g2_nand2_1 _16167_ (.Y(_11338_),
    .A(_08632_),
    .B(_11251_));
 sg13g2_or2_1 _16168_ (.X(_11339_),
    .B(_11338_),
    .A(net6500));
 sg13g2_and2_1 _16169_ (.A(net6482),
    .B(net6202),
    .X(_11340_));
 sg13g2_and2_1 _16170_ (.A(net6203),
    .B(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .X(_11341_));
 sg13g2_nand2_1 _16171_ (.Y(_11342_),
    .A(net6201),
    .B(_11340_));
 sg13g2_nand3_1 _16172_ (.B(net6486),
    .C(_11340_),
    .A(net6201),
    .Y(_11343_));
 sg13g2_xnor2_1 _16173_ (.Y(_11344_),
    .A(net6486),
    .B(_11342_));
 sg13g2_a21oi_1 _16174_ (.A1(_11339_),
    .A2(_11344_),
    .Y(_11345_),
    .B1(_11331_));
 sg13g2_a22oi_1 _16175_ (.Y(_00831_),
    .B1(_11337_),
    .B2(_11345_),
    .A2(_11331_),
    .A1(_07878_));
 sg13g2_xnor2_1 _16176_ (.Y(_11346_),
    .A(net6486),
    .B(net6485));
 sg13g2_a21oi_1 _16177_ (.A1(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .A2(_08665_),
    .Y(_11347_),
    .B1(net6485));
 sg13g2_a221oi_1 _16178_ (.B2(net6142),
    .C1(_11334_),
    .B1(_11347_),
    .A1(_11333_),
    .Y(_11348_),
    .A2(_11346_));
 sg13g2_a21oi_1 _16179_ (.A1(net6501),
    .A2(_08414_),
    .Y(_11349_),
    .B1(net6488));
 sg13g2_xnor2_1 _16180_ (.Y(_11350_),
    .A(_07879_),
    .B(_11343_));
 sg13g2_a21oi_1 _16181_ (.A1(_11251_),
    .A2(_11349_),
    .Y(_11351_),
    .B1(_11350_));
 sg13g2_nor3_1 _16182_ (.A(_11331_),
    .B(_11348_),
    .C(_11351_),
    .Y(_11352_));
 sg13g2_a21oi_1 _16183_ (.A1(_07879_),
    .A2(_11331_),
    .Y(_00832_),
    .B1(_11352_));
 sg13g2_and2_1 _16184_ (.A(_11248_),
    .B(_11251_),
    .X(_11353_));
 sg13g2_nand3_1 _16185_ (.B(_08657_),
    .C(_11341_),
    .A(net6484),
    .Y(_11354_));
 sg13g2_nand2b_1 _16186_ (.Y(_11355_),
    .B(_11354_),
    .A_N(_11353_));
 sg13g2_a21oi_1 _16187_ (.A1(_08657_),
    .A2(_11341_),
    .Y(_11356_),
    .B1(net6484));
 sg13g2_o21ai_1 _16188_ (.B1(_11251_),
    .Y(_11357_),
    .A1(net6484),
    .A2(_08657_));
 sg13g2_nor2b_1 _16189_ (.A(_11357_),
    .B_N(_10772_),
    .Y(_11358_));
 sg13g2_and2_1 _16190_ (.A(_08660_),
    .B(_11257_),
    .X(_11359_));
 sg13g2_o21ai_1 _16191_ (.B1(_11359_),
    .Y(_11360_),
    .A1(net6482),
    .A2(_11353_));
 sg13g2_o21ai_1 _16192_ (.B1(_11360_),
    .Y(_11361_),
    .A1(_07874_),
    .A2(_11358_));
 sg13g2_o21ai_1 _16193_ (.B1(_11361_),
    .Y(_11362_),
    .A1(_11355_),
    .A2(_11356_));
 sg13g2_o21ai_1 _16194_ (.B1(_11362_),
    .Y(_11363_),
    .A1(net6483),
    .A2(net3261));
 sg13g2_nor2_1 _16195_ (.A(_08666_),
    .B(_10779_),
    .Y(_11364_));
 sg13g2_a21oi_1 _16196_ (.A1(_11358_),
    .A2(_11364_),
    .Y(_11365_),
    .B1(_11331_));
 sg13g2_a22oi_1 _16197_ (.Y(_00833_),
    .B1(net3262),
    .B2(_11365_),
    .A2(_11331_),
    .A1(_07881_));
 sg13g2_a21oi_1 _16198_ (.A1(_11258_),
    .A2(_11353_),
    .Y(_11366_),
    .B1(net6482));
 sg13g2_nor2_1 _16199_ (.A(_11331_),
    .B(_11366_),
    .Y(_11367_));
 sg13g2_and2_1 _16200_ (.A(_11355_),
    .B(_11367_),
    .X(_11368_));
 sg13g2_nor4_1 _16201_ (.A(net3334),
    .B(_10772_),
    .C(_11342_),
    .D(_11353_),
    .Y(_11369_));
 sg13g2_o21ai_1 _16202_ (.B1(_11259_),
    .Y(_11370_),
    .A1(net6482),
    .A2(net3334));
 sg13g2_o21ai_1 _16203_ (.B1(_11370_),
    .Y(_11371_),
    .A1(_08666_),
    .A2(_10779_));
 sg13g2_xnor2_1 _16204_ (.Y(_11372_),
    .A(_07880_),
    .B(_10772_));
 sg13g2_nor2_1 _16205_ (.A(_11331_),
    .B(_11372_),
    .Y(_11373_));
 sg13g2_o21ai_1 _16206_ (.B1(_11373_),
    .Y(_11374_),
    .A1(_11369_),
    .A2(_11371_));
 sg13g2_o21ai_1 _16207_ (.B1(_11374_),
    .Y(_00834_),
    .A1(_07880_),
    .A2(_11368_));
 sg13g2_or2_1 _16208_ (.X(_00835_),
    .B(net1776),
    .A(net436));
 sg13g2_o21ai_1 _16209_ (.B1(_09366_),
    .Y(_11375_),
    .A1(_11114_),
    .A2(_11328_));
 sg13g2_a21oi_1 _16210_ (.A1(_11115_),
    .A2(_11253_),
    .Y(_11376_),
    .B1(net6482));
 sg13g2_nand3_1 _16211_ (.B(_11115_),
    .C(_11253_),
    .A(_08419_),
    .Y(_11377_));
 sg13g2_nand2_1 _16212_ (.Y(_11378_),
    .A(_11113_),
    .B(_11377_));
 sg13g2_nor3_1 _16213_ (.A(_11375_),
    .B(_11376_),
    .C(_11378_),
    .Y(_11379_));
 sg13g2_a21oi_1 _16214_ (.A1(net6142),
    .A2(_11375_),
    .Y(_00836_),
    .B1(_11379_));
 sg13g2_and2_1 _16215_ (.A(\soc_inst.cpu_core.csr_file.mie[11] ),
    .B(\soc_inst.cpu_core.csr_file.mip_eip ),
    .X(_11380_));
 sg13g2_o21ai_1 _16216_ (.B1(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .Y(_11381_),
    .A1(_09130_),
    .A2(_11380_));
 sg13g2_nand4_1 _16217_ (.B(\soc_inst.cpu_core.if_pc[5] ),
    .C(\soc_inst.cpu_core.if_pc[6] ),
    .A(\soc_inst.cpu_core.if_pc[4] ),
    .Y(_11382_),
    .D(\soc_inst.cpu_core.if_pc[7] ));
 sg13g2_nand3_1 _16218_ (.B(\soc_inst.cpu_core.if_pc[0] ),
    .C(\soc_inst.cpu_core.if_pc[3] ),
    .A(\soc_inst.cpu_core.if_pc[1] ),
    .Y(_11383_));
 sg13g2_nor3_2 _16219_ (.A(_07912_),
    .B(_11382_),
    .C(_11383_),
    .Y(_11384_));
 sg13g2_nand4_1 _16220_ (.B(\soc_inst.cpu_core.if_pc[13] ),
    .C(\soc_inst.cpu_core.if_pc[14] ),
    .A(\soc_inst.cpu_core.if_pc[12] ),
    .Y(_11385_),
    .D(\soc_inst.cpu_core.if_pc[15] ));
 sg13g2_nand4_1 _16221_ (.B(\soc_inst.cpu_core.if_pc[9] ),
    .C(\soc_inst.cpu_core.if_pc[10] ),
    .A(\soc_inst.cpu_core.if_pc[8] ),
    .Y(_11386_),
    .D(\soc_inst.cpu_core.if_pc[11] ));
 sg13g2_nand4_1 _16222_ (.B(\soc_inst.cpu_core.if_pc[17] ),
    .C(\soc_inst.cpu_core.if_pc[18] ),
    .A(\soc_inst.cpu_core.if_pc[16] ),
    .Y(_11387_),
    .D(\soc_inst.cpu_core.if_pc[19] ));
 sg13g2_nand4_1 _16223_ (.B(\soc_inst.cpu_core.if_pc[21] ),
    .C(\soc_inst.cpu_core.if_pc[22] ),
    .A(\soc_inst.cpu_core.if_pc[20] ),
    .Y(_11388_),
    .D(\soc_inst.cpu_core.if_pc[23] ));
 sg13g2_nor4_1 _16224_ (.A(_11385_),
    .B(_11386_),
    .C(_11387_),
    .D(_11388_),
    .Y(_11389_));
 sg13g2_a21oi_2 _16225_ (.B1(_11381_),
    .Y(_11390_),
    .A2(_11389_),
    .A1(_11384_));
 sg13g2_nor2_1 _16226_ (.A(net6391),
    .B(_11390_),
    .Y(_11391_));
 sg13g2_a21oi_1 _16227_ (.A1(_07871_),
    .A2(net6369),
    .Y(_00837_),
    .B1(net5307));
 sg13g2_or3_1 _16228_ (.A(_00256_),
    .B(_00255_),
    .C(\soc_inst.cpu_core.id_instr[3] ),
    .X(_11392_));
 sg13g2_nor2_2 _16229_ (.A(\soc_inst.cpu_core.id_instr[2] ),
    .B(_11392_),
    .Y(_11393_));
 sg13g2_nor3_1 _16230_ (.A(_07792_),
    .B(\soc_inst.cpu_core.id_instr[5] ),
    .C(net6306),
    .Y(_11394_));
 sg13g2_a21oi_1 _16231_ (.A1(_11393_),
    .A2(_11394_),
    .Y(_11395_),
    .B1(net6413));
 sg13g2_nand4_1 _16232_ (.B(\soc_inst.cpu_core.id_instr[5] ),
    .C(net6306),
    .A(_07792_),
    .Y(_11396_),
    .D(_11393_));
 sg13g2_nor2_1 _16233_ (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_11397_));
 sg13g2_nor3_1 _16234_ (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[0] ),
    .C(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_11398_));
 sg13g2_nand2b_2 _16235_ (.Y(_11399_),
    .B(_11397_),
    .A_N(\soc_inst.cpu_core.id_funct3[0] ));
 sg13g2_nor4_1 _16236_ (.A(\soc_inst.cpu_core.id_instr[8] ),
    .B(\soc_inst.cpu_core.id_instr[7] ),
    .C(\soc_inst.cpu_core.id_instr[10] ),
    .D(\soc_inst.cpu_core.id_instr[11] ),
    .Y(_11400_));
 sg13g2_nor2b_1 _16237_ (.A(\soc_inst.cpu_core.id_instr[9] ),
    .B_N(_11400_),
    .Y(_11401_));
 sg13g2_nor3_1 _16238_ (.A(_11396_),
    .B(_11398_),
    .C(_11401_),
    .Y(_11402_));
 sg13g2_nand2_1 _16239_ (.Y(_11403_),
    .A(_00257_),
    .B(\soc_inst.cpu_core.id_instr[5] ));
 sg13g2_nand4_1 _16240_ (.B(\soc_inst.cpu_core.id_instr[2] ),
    .C(\soc_inst.cpu_core.id_instr[5] ),
    .A(_00257_),
    .Y(_11404_),
    .D(net6306));
 sg13g2_nor3_1 _16241_ (.A(_00256_),
    .B(_00255_),
    .C(_11404_),
    .Y(_11405_));
 sg13g2_nor3_1 _16242_ (.A(_00257_),
    .B(net6306),
    .C(_11392_),
    .Y(_11406_));
 sg13g2_nor3_1 _16243_ (.A(_11402_),
    .B(_11405_),
    .C(_11406_),
    .Y(_11407_));
 sg13g2_and2_1 _16244_ (.A(\soc_inst.cpu_core.id_instr[3] ),
    .B(_11405_),
    .X(_11408_));
 sg13g2_nand2_2 _16245_ (.Y(_11409_),
    .A(\soc_inst.cpu_core.id_instr[3] ),
    .B(_11405_));
 sg13g2_nor2_1 _16246_ (.A(_11392_),
    .B(_11404_),
    .Y(_11410_));
 sg13g2_or2_1 _16247_ (.X(_11411_),
    .B(_11404_),
    .A(_11392_));
 sg13g2_a22oi_1 _16248_ (.Y(_00838_),
    .B1(_11395_),
    .B2(_11407_),
    .A2(_07933_),
    .A1(net6413));
 sg13g2_or3_1 _16249_ (.A(net2885),
    .B(_11396_),
    .C(_11399_),
    .X(_11412_));
 sg13g2_nor2_1 _16250_ (.A(net6352),
    .B(net2556),
    .Y(_11413_));
 sg13g2_nor2_1 _16251_ (.A(net2726),
    .B(net2566),
    .Y(_11414_));
 sg13g2_nor4_1 _16252_ (.A(net1121),
    .B(net2286),
    .C(net2613),
    .D(net2698),
    .Y(_11415_));
 sg13g2_and4_1 _16253_ (.A(net2501),
    .B(net2893),
    .C(net2609),
    .D(_11414_),
    .X(_11416_));
 sg13g2_nor4_1 _16254_ (.A(net6355),
    .B(net630),
    .C(net2556),
    .D(_11412_),
    .Y(_11417_));
 sg13g2_nand3_1 _16255_ (.B(_11416_),
    .C(_11417_),
    .A(_11415_),
    .Y(_11418_));
 sg13g2_o21ai_1 _16256_ (.B1(_11418_),
    .Y(_00839_),
    .A1(net6163),
    .A2(net6145));
 sg13g2_nor3_1 _16257_ (.A(net2501),
    .B(\soc_inst.cpu_core.id_imm12[8] ),
    .C(net2609),
    .Y(_11419_));
 sg13g2_nand3_1 _16258_ (.B(_11415_),
    .C(net2610),
    .A(_11414_),
    .Y(_11420_));
 sg13g2_nor4_1 _16259_ (.A(net6356),
    .B(net2556),
    .C(_11412_),
    .D(net2611),
    .Y(_11421_));
 sg13g2_a22oi_1 _16260_ (.Y(_11422_),
    .B1(net630),
    .B2(net2612),
    .A2(net6356),
    .A1(net2562));
 sg13g2_inv_1 _16261_ (.Y(_00840_),
    .A(_11422_));
 sg13g2_nor2_1 _16262_ (.A(net6312),
    .B(net377),
    .Y(_11423_));
 sg13g2_a21oi_1 _16263_ (.A1(_07785_),
    .A2(net6312),
    .Y(_00841_),
    .B1(_11423_));
 sg13g2_nor2_1 _16264_ (.A(net6311),
    .B(net299),
    .Y(_11424_));
 sg13g2_a21oi_1 _16265_ (.A1(_07784_),
    .A2(net6310),
    .Y(_00842_),
    .B1(_11424_));
 sg13g2_mux2_1 _16266_ (.A0(net791),
    .A1(net6467),
    .S(net6331),
    .X(_00843_));
 sg13g2_mux2_1 _16267_ (.A0(net398),
    .A1(net6463),
    .S(net6312),
    .X(_00844_));
 sg13g2_mux2_1 _16268_ (.A0(net251),
    .A1(net6462),
    .S(net6310),
    .X(_00845_));
 sg13g2_mux2_1 _16269_ (.A0(net638),
    .A1(net6460),
    .S(net6311),
    .X(_00846_));
 sg13g2_mux2_1 _16270_ (.A0(net297),
    .A1(net6458),
    .S(net6310),
    .X(_00847_));
 sg13g2_mux2_1 _16271_ (.A0(net856),
    .A1(net6456),
    .S(net6313),
    .X(_00848_));
 sg13g2_mux2_1 _16272_ (.A0(net255),
    .A1(net1497),
    .S(net6321),
    .X(_00849_));
 sg13g2_mux2_1 _16273_ (.A0(net926),
    .A1(net6453),
    .S(net6308),
    .X(_00850_));
 sg13g2_mux2_1 _16274_ (.A0(net293),
    .A1(net1533),
    .S(net6320),
    .X(_00851_));
 sg13g2_mux2_1 _16275_ (.A0(net1396),
    .A1(\soc_inst.core_mem_wdata[11] ),
    .S(net6307),
    .X(_00852_));
 sg13g2_mux2_1 _16276_ (.A0(net1799),
    .A1(net1825),
    .S(net6308),
    .X(_00853_));
 sg13g2_mux2_1 _16277_ (.A0(net238),
    .A1(net1321),
    .S(net6309),
    .X(_00854_));
 sg13g2_mux2_1 _16278_ (.A0(net335),
    .A1(net1503),
    .S(net6309),
    .X(_00855_));
 sg13g2_mux2_1 _16279_ (.A0(net1548),
    .A1(net2861),
    .S(net6307),
    .X(_00856_));
 sg13g2_mux2_1 _16280_ (.A0(net324),
    .A1(net225),
    .S(net6314),
    .X(_00857_));
 sg13g2_mux2_1 _16281_ (.A0(net566),
    .A1(net160),
    .S(net6314),
    .X(_00858_));
 sg13g2_mux2_1 _16282_ (.A0(net510),
    .A1(net1272),
    .S(net6316),
    .X(_00859_));
 sg13g2_mux2_1 _16283_ (.A0(net687),
    .A1(net295),
    .S(net6314),
    .X(_00860_));
 sg13g2_mux2_1 _16284_ (.A0(net1976),
    .A1(net548),
    .S(net6314),
    .X(_00861_));
 sg13g2_mux2_1 _16285_ (.A0(net522),
    .A1(net571),
    .S(net6316),
    .X(_00862_));
 sg13g2_mux2_1 _16286_ (.A0(net586),
    .A1(net1311),
    .S(net6315),
    .X(_00863_));
 sg13g2_mux2_1 _16287_ (.A0(net273),
    .A1(net1329),
    .S(net6322),
    .X(_00864_));
 sg13g2_mux2_1 _16288_ (.A0(net347),
    .A1(net268),
    .S(net6314),
    .X(_00865_));
 sg13g2_mux2_1 _16289_ (.A0(net2573),
    .A1(net233),
    .S(net6307),
    .X(_00866_));
 sg13g2_mux2_1 _16290_ (.A0(net208),
    .A1(net1016),
    .S(net6317),
    .X(_00867_));
 sg13g2_mux2_1 _16291_ (.A0(net472),
    .A1(net712),
    .S(net6315),
    .X(_00868_));
 sg13g2_mux2_1 _16292_ (.A0(net1089),
    .A1(net369),
    .S(net6307),
    .X(_00869_));
 sg13g2_mux2_1 _16293_ (.A0(net852),
    .A1(net313),
    .S(net6307),
    .X(_00870_));
 sg13g2_mux2_1 _16294_ (.A0(net1795),
    .A1(net734),
    .S(net6315),
    .X(_00871_));
 sg13g2_mux2_1 _16295_ (.A0(net426),
    .A1(net854),
    .S(net6317),
    .X(_00872_));
 sg13g2_nor2b_1 _16296_ (.A(net630),
    .B_N(_11421_),
    .Y(_11425_));
 sg13g2_a21o_1 _16297_ (.A2(net6351),
    .A1(net2455),
    .B1(_11425_),
    .X(_00873_));
 sg13g2_a21o_1 _16298_ (.A2(_08962_),
    .A1(net6158),
    .B1(net896),
    .X(_00874_));
 sg13g2_nand2_1 _16299_ (.Y(_11426_),
    .A(net1886),
    .B(net6373));
 sg13g2_nor4_2 _16300_ (.A(net6475),
    .B(net6328),
    .C(_08290_),
    .Y(_11427_),
    .D(_09942_));
 sg13g2_nand4_1 _16301_ (.B(net6158),
    .C(_08289_),
    .A(net3148),
    .Y(_11428_),
    .D(_09944_));
 sg13g2_nand2_1 _16302_ (.Y(_11429_),
    .A(net5132),
    .B(net4754));
 sg13g2_o21ai_1 _16303_ (.B1(_11426_),
    .Y(_00875_),
    .A1(\soc_inst.core_instr_data[0] ),
    .A2(_11429_));
 sg13g2_nand2_1 _16304_ (.Y(_11430_),
    .A(net2013),
    .B(net6373));
 sg13g2_o21ai_1 _16305_ (.B1(_11430_),
    .Y(_00876_),
    .A1(\soc_inst.core_instr_data[1] ),
    .A2(_11429_));
 sg13g2_nand2_1 _16306_ (.Y(_11431_),
    .A(net6373),
    .B(net2936));
 sg13g2_nand2_1 _16307_ (.Y(_11432_),
    .A(net6522),
    .B(_09952_));
 sg13g2_nor2_1 _16308_ (.A(net6012),
    .B(net5997),
    .Y(_11433_));
 sg13g2_nor2_1 _16309_ (.A(_09981_),
    .B(_11433_),
    .Y(_11434_));
 sg13g2_o21ai_1 _16310_ (.B1(_09980_),
    .Y(_11435_),
    .A1(net6012),
    .A2(net5997));
 sg13g2_nor2b_2 _16311_ (.A(net6510),
    .B_N(net6512),
    .Y(_11436_));
 sg13g2_nand2b_2 _16312_ (.Y(_11437_),
    .B(net6514),
    .A_N(net6510));
 sg13g2_nand3_1 _16313_ (.B(_11435_),
    .C(_11437_),
    .A(_09978_),
    .Y(_11438_));
 sg13g2_nor2_1 _16314_ (.A(net6092),
    .B(_09968_),
    .Y(_11439_));
 sg13g2_and3_1 _16315_ (.X(_11440_),
    .A(net6095),
    .B(net6014),
    .C(_09961_));
 sg13g2_nor2_1 _16316_ (.A(_11439_),
    .B(_11440_),
    .Y(_11441_));
 sg13g2_inv_1 _16317_ (.Y(_11442_),
    .A(_11441_));
 sg13g2_nand3_1 _16318_ (.B(net6015),
    .C(_09968_),
    .A(net6517),
    .Y(_11443_));
 sg13g2_a22oi_1 _16319_ (.Y(_11444_),
    .B1(_11442_),
    .B2(_11443_),
    .A2(_11438_),
    .A1(net6091));
 sg13g2_nand2_1 _16320_ (.Y(_11445_),
    .A(net5067),
    .B(_11444_));
 sg13g2_o21ai_1 _16321_ (.B1(_11445_),
    .Y(_11446_),
    .A1(net6531),
    .A2(net5067));
 sg13g2_o21ai_1 _16322_ (.B1(_11431_),
    .Y(_00877_),
    .A1(net4719),
    .A2(_11446_));
 sg13g2_nand2_1 _16323_ (.Y(_11447_),
    .A(net6376),
    .B(net3065));
 sg13g2_nor2_1 _16324_ (.A(net5131),
    .B(_11437_),
    .Y(_11448_));
 sg13g2_a21oi_1 _16325_ (.A1(net6530),
    .A2(net5130),
    .Y(_11449_),
    .B1(_11448_));
 sg13g2_o21ai_1 _16326_ (.B1(_11447_),
    .Y(_00878_),
    .A1(net4720),
    .A2(_11449_));
 sg13g2_nand2_1 _16327_ (.Y(_11450_),
    .A(net2877),
    .B(net6416));
 sg13g2_nand2b_1 _16328_ (.Y(_11451_),
    .B(_09961_),
    .A_N(_09955_));
 sg13g2_nand2_1 _16329_ (.Y(_11452_),
    .A(net6014),
    .B(_11451_));
 sg13g2_nor2_2 _16330_ (.A(net6511),
    .B(net6508),
    .Y(_11453_));
 sg13g2_or2_1 _16331_ (.X(_11454_),
    .B(net6508),
    .A(net6510));
 sg13g2_nor3_1 _16332_ (.A(net6512),
    .B(net6510),
    .C(net6508),
    .Y(_11455_));
 sg13g2_nand2b_2 _16333_ (.Y(_11456_),
    .B(_09956_),
    .A_N(net6509));
 sg13g2_nand3_1 _16334_ (.B(_11452_),
    .C(_11456_),
    .A(_09968_),
    .Y(_11457_));
 sg13g2_nor2_2 _16335_ (.A(_09966_),
    .B(_09987_),
    .Y(_11458_));
 sg13g2_and2_1 _16336_ (.A(net6511),
    .B(net6508),
    .X(_11459_));
 sg13g2_nand2_2 _16337_ (.Y(_11460_),
    .A(net6510),
    .B(net6509));
 sg13g2_nand2_2 _16338_ (.Y(_11461_),
    .A(_11437_),
    .B(_11460_));
 sg13g2_a21oi_1 _16339_ (.A1(net6095),
    .A2(_11457_),
    .Y(_11462_),
    .B1(_11458_));
 sg13g2_o21ai_1 _16340_ (.B1(_11462_),
    .Y(_11463_),
    .A1(_09973_),
    .A2(_11461_));
 sg13g2_mux2_1 _16341_ (.A0(\soc_inst.core_instr_data[4] ),
    .A1(_11463_),
    .S(net5066),
    .X(_11464_));
 sg13g2_o21ai_1 _16342_ (.B1(_11450_),
    .Y(_00879_),
    .A1(net4720),
    .A2(_11464_));
 sg13g2_nand2_1 _16343_ (.Y(_11465_),
    .A(net6415),
    .B(net3174));
 sg13g2_nand2_1 _16344_ (.Y(_11466_),
    .A(net6092),
    .B(_09976_));
 sg13g2_a221oi_1 _16345_ (.B2(net6508),
    .C1(_11461_),
    .B1(_11466_),
    .A1(net6094),
    .Y(_11467_),
    .A2(_09969_));
 sg13g2_nand3_1 _16346_ (.B(_11435_),
    .C(_11467_),
    .A(net5065),
    .Y(_11468_));
 sg13g2_o21ai_1 _16347_ (.B1(_11468_),
    .Y(_11469_),
    .A1(net6528),
    .A2(net5065));
 sg13g2_o21ai_1 _16348_ (.B1(_11465_),
    .Y(_00880_),
    .A1(net4720),
    .A2(_11469_));
 sg13g2_nand2_1 _16349_ (.Y(_11470_),
    .A(net6415),
    .B(net6451));
 sg13g2_o21ai_1 _16350_ (.B1(net6091),
    .Y(_11471_),
    .A1(_09984_),
    .A2(_11461_));
 sg13g2_nand3_1 _16351_ (.B(_11441_),
    .C(_11471_),
    .A(net5067),
    .Y(_11472_));
 sg13g2_o21ai_1 _16352_ (.B1(_11472_),
    .Y(_11473_),
    .A1(net6526),
    .A2(net5067));
 sg13g2_o21ai_1 _16353_ (.B1(_11470_),
    .Y(_00881_),
    .A1(net4721),
    .A2(_11473_));
 sg13g2_nand2_1 _16354_ (.Y(_11474_),
    .A(net6378),
    .B(net1906));
 sg13g2_nor2b_2 _16355_ (.A(net6514),
    .B_N(\soc_inst.core_instr_data[2] ),
    .Y(_11475_));
 sg13g2_and2_1 _16356_ (.A(net6531),
    .B(_09988_),
    .X(_11476_));
 sg13g2_o21ai_1 _16357_ (.B1(_09986_),
    .Y(_11477_),
    .A1(_09991_),
    .A2(_11476_));
 sg13g2_nand2_1 _16358_ (.Y(_11478_),
    .A(net6517),
    .B(net6013));
 sg13g2_nor2_1 _16359_ (.A(_09958_),
    .B(_09961_),
    .Y(_11479_));
 sg13g2_o21ai_1 _16360_ (.B1(net6524),
    .Y(_11480_),
    .A1(net6090),
    .A2(_11479_));
 sg13g2_o21ai_1 _16361_ (.B1(_11480_),
    .Y(_11481_),
    .A1(_11451_),
    .A2(_11478_));
 sg13g2_a21oi_1 _16362_ (.A1(net6525),
    .A2(net6088),
    .Y(_11482_),
    .B1(_09969_));
 sg13g2_o21ai_1 _16363_ (.B1(net6094),
    .Y(_11483_),
    .A1(_09970_),
    .A2(_11481_));
 sg13g2_nor2_2 _16364_ (.A(_09973_),
    .B(net6088),
    .Y(_11484_));
 sg13g2_a21o_1 _16365_ (.A2(_09972_),
    .A1(net6524),
    .B1(_11484_),
    .X(_11485_));
 sg13g2_nand2_1 _16366_ (.Y(_11486_),
    .A(net6515),
    .B(net6086));
 sg13g2_nand4_1 _16367_ (.B(_11437_),
    .C(_11454_),
    .A(net6525),
    .Y(_11487_),
    .D(_11460_));
 sg13g2_nand3_1 _16368_ (.B(_11486_),
    .C(_11487_),
    .A(_11454_),
    .Y(_11488_));
 sg13g2_o21ai_1 _16369_ (.B1(_11485_),
    .Y(_11489_),
    .A1(_09984_),
    .A2(_11488_));
 sg13g2_nand4_1 _16370_ (.B(_11477_),
    .C(_11483_),
    .A(net5068),
    .Y(_11490_),
    .D(_11489_));
 sg13g2_o21ai_1 _16371_ (.B1(_11490_),
    .Y(_11491_),
    .A1(net6524),
    .A2(net5067));
 sg13g2_o21ai_1 _16372_ (.B1(_11474_),
    .Y(_00882_),
    .A1(net4719),
    .A2(_11491_));
 sg13g2_nand2_1 _16373_ (.Y(_11492_),
    .A(net6374),
    .B(net1270));
 sg13g2_o21ai_1 _16374_ (.B1(net6094),
    .Y(_11493_),
    .A1(net6090),
    .A2(_11479_));
 sg13g2_nand2_1 _16375_ (.Y(_11494_),
    .A(net5066),
    .B(_11493_));
 sg13g2_nand2_1 _16376_ (.Y(_11495_),
    .A(net6530),
    .B(_09988_));
 sg13g2_a21oi_1 _16377_ (.A1(_09992_),
    .A2(_11495_),
    .Y(_11496_),
    .B1(_09987_));
 sg13g2_nand2_1 _16378_ (.Y(_11497_),
    .A(net6523),
    .B(_11454_));
 sg13g2_a21oi_1 _16379_ (.A1(net6530),
    .A2(net6086),
    .Y(_11498_),
    .B1(net6088));
 sg13g2_o21ai_1 _16380_ (.B1(_11498_),
    .Y(_11499_),
    .A1(_11461_),
    .A2(_11497_));
 sg13g2_nor2_1 _16381_ (.A(_09984_),
    .B(_11499_),
    .Y(_11500_));
 sg13g2_o21ai_1 _16382_ (.B1(_09972_),
    .Y(_11501_),
    .A1(net6522),
    .A2(_11456_));
 sg13g2_nand2_1 _16383_ (.Y(_11502_),
    .A(net6094),
    .B(_09970_));
 sg13g2_o21ai_1 _16384_ (.B1(_11502_),
    .Y(_11503_),
    .A1(_11500_),
    .A2(_11501_));
 sg13g2_or2_1 _16385_ (.X(_11504_),
    .B(_11503_),
    .A(_11496_));
 sg13g2_a22oi_1 _16386_ (.Y(_11505_),
    .B1(_11504_),
    .B2(net5066),
    .A2(_11494_),
    .A1(net6522));
 sg13g2_o21ai_1 _16387_ (.B1(_11492_),
    .Y(_00883_),
    .A1(net4719),
    .A2(_11505_));
 sg13g2_nand2_1 _16388_ (.Y(_11506_),
    .A(net6374),
    .B(net1265));
 sg13g2_nor2_2 _16389_ (.A(net6514),
    .B(_11460_),
    .Y(_11507_));
 sg13g2_a221oi_1 _16390_ (.B2(net6527),
    .C1(_09991_),
    .B1(_11507_),
    .A1(net6529),
    .Y(_11508_),
    .A2(_09988_));
 sg13g2_nand2_1 _16391_ (.Y(_11509_),
    .A(net6529),
    .B(_11459_));
 sg13g2_nor2_1 _16392_ (.A(\soc_inst.core_instr_data[9] ),
    .B(_11453_),
    .Y(_11510_));
 sg13g2_o21ai_1 _16393_ (.B1(_11509_),
    .Y(_11511_),
    .A1(_11461_),
    .A2(_11510_));
 sg13g2_a21oi_1 _16394_ (.A1(_08026_),
    .A2(net6088),
    .Y(_11512_),
    .B1(_09973_));
 sg13g2_o21ai_1 _16395_ (.B1(_11512_),
    .Y(_11513_),
    .A1(_09984_),
    .A2(_11511_));
 sg13g2_o21ai_1 _16396_ (.B1(_11502_),
    .Y(_11514_),
    .A1(_09987_),
    .A2(_11508_));
 sg13g2_nand2b_1 _16397_ (.Y(_11515_),
    .B(_11513_),
    .A_N(_11514_));
 sg13g2_a21o_1 _16398_ (.A2(net6086),
    .A1(net6095),
    .B1(_11494_),
    .X(_11516_));
 sg13g2_a22oi_1 _16399_ (.Y(_11517_),
    .B1(_11516_),
    .B2(\soc_inst.core_instr_data[9] ),
    .A2(_11515_),
    .A1(net5065));
 sg13g2_o21ai_1 _16400_ (.B1(_11506_),
    .Y(_00884_),
    .A1(net4719),
    .A2(_11517_));
 sg13g2_nand2_1 _16401_ (.Y(_11518_),
    .A(net6374),
    .B(net873));
 sg13g2_o21ai_1 _16402_ (.B1(_08027_),
    .Y(_11519_),
    .A1(net6522),
    .A2(_09953_));
 sg13g2_o21ai_1 _16403_ (.B1(_11519_),
    .Y(_11520_),
    .A1(_09963_),
    .A2(_09967_));
 sg13g2_or3_1 _16404_ (.A(net6088),
    .B(net6086),
    .C(_11479_),
    .X(_11521_));
 sg13g2_a21oi_1 _16405_ (.A1(\soc_inst.core_instr_data[10] ),
    .A2(_11521_),
    .Y(_11522_),
    .B1(net6513));
 sg13g2_a21oi_1 _16406_ (.A1(_11520_),
    .A2(_11522_),
    .Y(_11523_),
    .B1(net6093));
 sg13g2_a21oi_1 _16407_ (.A1(_08027_),
    .A2(_11507_),
    .Y(_11524_),
    .B1(_09987_));
 sg13g2_a21oi_1 _16408_ (.A1(net6511),
    .A2(net6521),
    .Y(_11525_),
    .B1(_09956_));
 sg13g2_o21ai_1 _16409_ (.B1(_09972_),
    .Y(_11526_),
    .A1(net6521),
    .A2(_11456_));
 sg13g2_a21oi_1 _16410_ (.A1(_09982_),
    .A2(_11525_),
    .Y(_11527_),
    .B1(_11526_));
 sg13g2_or4_1 _16411_ (.A(net5131),
    .B(_11523_),
    .C(_11524_),
    .D(_11527_),
    .X(_11528_));
 sg13g2_o21ai_1 _16412_ (.B1(_11528_),
    .Y(_11529_),
    .A1(net6521),
    .A2(net5065));
 sg13g2_o21ai_1 _16413_ (.B1(_11518_),
    .Y(_00885_),
    .A1(net4719),
    .A2(_11529_));
 sg13g2_nand2_1 _16414_ (.Y(_11530_),
    .A(net6378),
    .B(net1248));
 sg13g2_o21ai_1 _16415_ (.B1(_09967_),
    .Y(_11531_),
    .A1(net6518),
    .A2(_09954_));
 sg13g2_nand2_1 _16416_ (.Y(_11532_),
    .A(net6519),
    .B(_11453_));
 sg13g2_o21ai_1 _16417_ (.B1(_11532_),
    .Y(_11533_),
    .A1(_09961_),
    .A2(_09974_));
 sg13g2_nor2_1 _16418_ (.A(net6512),
    .B(_11533_),
    .Y(_11534_));
 sg13g2_and3_1 _16419_ (.X(_11535_),
    .A(_09964_),
    .B(_11531_),
    .C(_11534_));
 sg13g2_nand2_1 _16420_ (.Y(_11536_),
    .A(net6519),
    .B(_09967_));
 sg13g2_nand2_1 _16421_ (.Y(_11537_),
    .A(_09982_),
    .B(_11536_));
 sg13g2_nand2_1 _16422_ (.Y(_11538_),
    .A(_11484_),
    .B(_11537_));
 sg13g2_o21ai_1 _16423_ (.B1(_11538_),
    .Y(_11539_),
    .A1(net6092),
    .A2(_11535_));
 sg13g2_o21ai_1 _16424_ (.B1(net6013),
    .Y(_11540_),
    .A1(net6515),
    .A2(_09976_));
 sg13g2_nor2b_1 _16425_ (.A(net6520),
    .B_N(net6518),
    .Y(_11541_));
 sg13g2_a21oi_1 _16426_ (.A1(net6512),
    .A2(net6510),
    .Y(_11542_),
    .B1(net6087));
 sg13g2_o21ai_1 _16427_ (.B1(_11542_),
    .Y(_11543_),
    .A1(_11540_),
    .A2(_11541_));
 sg13g2_a21oi_1 _16428_ (.A1(net6091),
    .A2(_11543_),
    .Y(_11544_),
    .B1(_11507_));
 sg13g2_nand2_1 _16429_ (.Y(_11545_),
    .A(net5063),
    .B(_11544_));
 sg13g2_a22oi_1 _16430_ (.Y(_11546_),
    .B1(_11545_),
    .B2(net6519),
    .A2(_11539_),
    .A1(net5063));
 sg13g2_o21ai_1 _16431_ (.B1(_11530_),
    .Y(_00886_),
    .A1(net4721),
    .A2(_11546_));
 sg13g2_nand2_1 _16432_ (.Y(_11547_),
    .A(net6415),
    .B(net3014));
 sg13g2_nor2_1 _16433_ (.A(net6531),
    .B(net6012),
    .Y(_11548_));
 sg13g2_nand2_1 _16434_ (.Y(_11549_),
    .A(net6515),
    .B(_11436_));
 sg13g2_nand2_1 _16435_ (.Y(_11550_),
    .A(_11540_),
    .B(_11549_));
 sg13g2_and2_1 _16436_ (.A(net6528),
    .B(net6527),
    .X(_11551_));
 sg13g2_a221oi_1 _16437_ (.B2(net6014),
    .C1(_11550_),
    .B1(_11551_),
    .A1(net6513),
    .Y(_11552_),
    .A2(_11459_));
 sg13g2_o21ai_1 _16438_ (.B1(_11552_),
    .Y(_11553_),
    .A1(_11435_),
    .A2(_11548_));
 sg13g2_nand2_1 _16439_ (.Y(_11554_),
    .A(net6091),
    .B(_11553_));
 sg13g2_o21ai_1 _16440_ (.B1(net6095),
    .Y(_11555_),
    .A1(_09970_),
    .A2(net6088));
 sg13g2_a21oi_1 _16441_ (.A1(_11554_),
    .A2(_11555_),
    .Y(_11556_),
    .B1(net5132));
 sg13g2_a21oi_1 _16442_ (.A1(net6517),
    .A2(net5132),
    .Y(_11557_),
    .B1(_11556_));
 sg13g2_o21ai_1 _16443_ (.B1(_11547_),
    .Y(_00887_),
    .A1(net4720),
    .A2(_11557_));
 sg13g2_nand2_1 _16444_ (.Y(_11558_),
    .A(net6376),
    .B(net2924));
 sg13g2_a22oi_1 _16445_ (.Y(_11559_),
    .B1(net5065),
    .B2(net6093),
    .A2(_09964_),
    .A1(_09956_));
 sg13g2_nand2_2 _16446_ (.Y(_11560_),
    .A(_09990_),
    .B(net6087));
 sg13g2_nand2_1 _16447_ (.Y(_11561_),
    .A(_09986_),
    .B(_11560_));
 sg13g2_nor2_1 _16448_ (.A(net6530),
    .B(net6012),
    .Y(_11562_));
 sg13g2_nand2b_1 _16449_ (.Y(_11563_),
    .B(net6521),
    .A_N(net6527));
 sg13g2_nand2_1 _16450_ (.Y(_11564_),
    .A(_09974_),
    .B(_11549_));
 sg13g2_o21ai_1 _16451_ (.B1(_11564_),
    .Y(_11565_),
    .A1(net6516),
    .A2(_11563_));
 sg13g2_o21ai_1 _16452_ (.B1(_11565_),
    .Y(_11566_),
    .A1(_11435_),
    .A2(_11562_));
 sg13g2_a21oi_1 _16453_ (.A1(net6091),
    .A2(_11566_),
    .Y(_11567_),
    .B1(_11559_));
 sg13g2_nand2_1 _16454_ (.Y(_11568_),
    .A(_11561_),
    .B(_11567_));
 sg13g2_o21ai_1 _16455_ (.B1(_11568_),
    .Y(_11569_),
    .A1(net6513),
    .A2(net5065));
 sg13g2_o21ai_1 _16456_ (.B1(_11558_),
    .Y(_00888_),
    .A1(net4719),
    .A2(_11569_));
 sg13g2_nand2_1 _16457_ (.Y(_11570_),
    .A(net6416),
    .B(net2945));
 sg13g2_or2_1 _16458_ (.X(_11571_),
    .B(net6012),
    .A(net6529));
 sg13g2_a221oi_1 _16459_ (.B2(_11571_),
    .C1(_11550_),
    .B1(_11434_),
    .A1(net6014),
    .Y(_11572_),
    .A2(_09959_));
 sg13g2_o21ai_1 _16460_ (.B1(net5066),
    .Y(_11573_),
    .A1(_09973_),
    .A2(_11572_));
 sg13g2_o21ai_1 _16461_ (.B1(_11573_),
    .Y(_11574_),
    .A1(net6511),
    .A2(net5067));
 sg13g2_o21ai_1 _16462_ (.B1(_11570_),
    .Y(_00889_),
    .A1(net4720),
    .A2(_11574_));
 sg13g2_nand2_1 _16463_ (.Y(_11575_),
    .A(net6375),
    .B(net6450));
 sg13g2_a21o_1 _16464_ (.A2(_09966_),
    .A1(net6524),
    .B1(_09991_),
    .X(_11576_));
 sg13g2_nor2_2 _16465_ (.A(net6517),
    .B(_09961_),
    .Y(_11577_));
 sg13g2_nor2_2 _16466_ (.A(_09958_),
    .B(_11577_),
    .Y(_11578_));
 sg13g2_inv_1 _16467_ (.Y(_11579_),
    .A(_11578_));
 sg13g2_o21ai_1 _16468_ (.B1(_11578_),
    .Y(_11580_),
    .A1(net6525),
    .A2(_09989_));
 sg13g2_a21oi_1 _16469_ (.A1(_11482_),
    .A2(_11580_),
    .Y(_11581_),
    .B1(net6093));
 sg13g2_or2_1 _16470_ (.X(_11582_),
    .B(_09962_),
    .A(\soc_inst.core_instr_data[5] ));
 sg13g2_nand2_1 _16471_ (.Y(_11583_),
    .A(_11434_),
    .B(_11582_));
 sg13g2_a21oi_2 _16472_ (.B1(net6087),
    .Y(_11584_),
    .A2(_11436_),
    .A1(net6515));
 sg13g2_nand2_1 _16473_ (.Y(_11585_),
    .A(_09978_),
    .B(_11584_));
 sg13g2_and2_1 _16474_ (.A(net6509),
    .B(_11437_),
    .X(_11586_));
 sg13g2_a21oi_1 _16475_ (.A1(net6524),
    .A2(_11586_),
    .Y(_11587_),
    .B1(_11585_));
 sg13g2_nand2_1 _16476_ (.Y(_11588_),
    .A(_11583_),
    .B(_11587_));
 sg13g2_a221oi_1 _16477_ (.B2(_11485_),
    .C1(_11581_),
    .B1(_11588_),
    .A1(_09986_),
    .Y(_11589_),
    .A2(_11576_));
 sg13g2_nand2_1 _16478_ (.Y(_11590_),
    .A(net5067),
    .B(_11589_));
 sg13g2_o21ai_1 _16479_ (.B1(_11590_),
    .Y(_11591_),
    .A1(net6509),
    .A2(net5067));
 sg13g2_o21ai_1 _16480_ (.B1(_11575_),
    .Y(_00890_),
    .A1(net4719),
    .A2(_11591_));
 sg13g2_or2_1 _16481_ (.X(_11592_),
    .B(_09962_),
    .A(net6527));
 sg13g2_nand2b_1 _16482_ (.Y(_11593_),
    .B(_11432_),
    .A_N(_11592_));
 sg13g2_a221oi_1 _16483_ (.B2(_09980_),
    .C1(_11585_),
    .B1(_11593_),
    .A1(net6522),
    .Y(_11594_),
    .A2(_11586_));
 sg13g2_nand2_2 _16484_ (.Y(_11595_),
    .A(_11456_),
    .B(_11579_));
 sg13g2_nand3_1 _16485_ (.B(_09952_),
    .C(_11578_),
    .A(_08028_),
    .Y(_11596_));
 sg13g2_nand2_1 _16486_ (.Y(_11597_),
    .A(net6522),
    .B(_11595_));
 sg13g2_nand3_1 _16487_ (.B(_11596_),
    .C(_11597_),
    .A(_09956_),
    .Y(_11598_));
 sg13g2_a221oi_1 _16488_ (.B2(net6095),
    .C1(_11458_),
    .B1(_11598_),
    .A1(net6523),
    .Y(_11599_),
    .A2(_09986_));
 sg13g2_o21ai_1 _16489_ (.B1(_11599_),
    .Y(_11600_),
    .A1(_11501_),
    .A2(_11594_));
 sg13g2_mux2_1 _16490_ (.A0(net2667),
    .A1(_11600_),
    .S(net5068),
    .X(_11601_));
 sg13g2_a22oi_1 _16491_ (.Y(_11602_),
    .B1(net4754),
    .B2(_11601_),
    .A2(net6448),
    .A1(net6363));
 sg13g2_inv_1 _16492_ (.Y(_00891_),
    .A(_11602_));
 sg13g2_nand2_1 _16493_ (.Y(_11603_),
    .A(net6375),
    .B(net6445));
 sg13g2_a22oi_1 _16494_ (.Y(_11604_),
    .B1(_11512_),
    .B2(_11586_),
    .A2(_09985_),
    .A1(_09966_));
 sg13g2_nor2_1 _16495_ (.A(_08026_),
    .B(net6092),
    .Y(_11605_));
 sg13g2_nor2_1 _16496_ (.A(_09981_),
    .B(_11577_),
    .Y(_11606_));
 sg13g2_a21oi_2 _16497_ (.B1(_09981_),
    .Y(_11607_),
    .A2(_11577_),
    .A1(net5997));
 sg13g2_nand2b_2 _16498_ (.Y(_11608_),
    .B(_11607_),
    .A_N(_11433_));
 sg13g2_and2_1 _16499_ (.A(_09978_),
    .B(_11608_),
    .X(_11609_));
 sg13g2_nand2_2 _16500_ (.Y(_11610_),
    .A(_11584_),
    .B(_11609_));
 sg13g2_a221oi_1 _16501_ (.B2(_11512_),
    .C1(net5131),
    .B1(_11610_),
    .A1(_11595_),
    .Y(_11611_),
    .A2(_11605_));
 sg13g2_o21ai_1 _16502_ (.B1(_11611_),
    .Y(_11612_),
    .A1(_08026_),
    .A2(_11604_));
 sg13g2_o21ai_1 _16503_ (.B1(_11612_),
    .Y(_11613_),
    .A1(net2696),
    .A2(net5063));
 sg13g2_o21ai_1 _16504_ (.B1(_11603_),
    .Y(_00892_),
    .A1(net4721),
    .A2(_11613_));
 sg13g2_nand2_1 _16505_ (.Y(_11614_),
    .A(net6362),
    .B(net6444));
 sg13g2_o21ai_1 _16506_ (.B1(_11578_),
    .Y(_11615_),
    .A1(\soc_inst.core_instr_data[10] ),
    .A2(_09989_));
 sg13g2_a21oi_1 _16507_ (.A1(\soc_inst.core_instr_data[10] ),
    .A2(_11453_),
    .Y(_11616_),
    .B1(_09969_));
 sg13g2_a21o_1 _16508_ (.A2(_11616_),
    .A1(_11615_),
    .B1(net6092),
    .X(_11617_));
 sg13g2_nor2b_1 _16509_ (.A(_11586_),
    .B_N(_11584_),
    .Y(_11618_));
 sg13g2_a21o_1 _16510_ (.A2(_11618_),
    .A1(_11608_),
    .B1(_11526_),
    .X(_11619_));
 sg13g2_nand4_1 _16511_ (.B(_11561_),
    .C(_11617_),
    .A(net5063),
    .Y(_11620_),
    .D(_11619_));
 sg13g2_o21ai_1 _16512_ (.B1(_11620_),
    .Y(_11621_),
    .A1(net2740),
    .A2(net5063));
 sg13g2_o21ai_1 _16513_ (.B1(_11614_),
    .Y(_00893_),
    .A1(net4722),
    .A2(_11621_));
 sg13g2_nand2_1 _16514_ (.Y(_11622_),
    .A(net6362),
    .B(net6443));
 sg13g2_o21ai_1 _16515_ (.B1(net6091),
    .Y(_11623_),
    .A1(net6519),
    .A2(_11456_));
 sg13g2_nand2b_1 _16516_ (.Y(_11624_),
    .B(_11610_),
    .A_N(_11623_));
 sg13g2_a21oi_1 _16517_ (.A1(_08028_),
    .A2(_09954_),
    .Y(_11625_),
    .B1(net6518));
 sg13g2_o21ai_1 _16518_ (.B1(_11532_),
    .Y(_11626_),
    .A1(_11579_),
    .A2(_11625_));
 sg13g2_o21ai_1 _16519_ (.B1(net6094),
    .Y(_11627_),
    .A1(_09969_),
    .A2(_11626_));
 sg13g2_nand3_1 _16520_ (.B(_11624_),
    .C(_11627_),
    .A(net5064),
    .Y(_11628_));
 sg13g2_o21ai_1 _16521_ (.B1(_11628_),
    .Y(_11629_),
    .A1(net2645),
    .A2(net5063));
 sg13g2_o21ai_1 _16522_ (.B1(_11622_),
    .Y(_00894_),
    .A1(net4722),
    .A2(_11629_));
 sg13g2_nand2_1 _16523_ (.Y(_11630_),
    .A(net6415),
    .B(net6438));
 sg13g2_and2_1 _16524_ (.A(_11459_),
    .B(_11475_),
    .X(_11631_));
 sg13g2_o21ai_1 _16525_ (.B1(_09986_),
    .Y(_11632_),
    .A1(_09991_),
    .A2(_11631_));
 sg13g2_nor2_2 _16526_ (.A(net6015),
    .B(_09973_),
    .Y(_11633_));
 sg13g2_a21oi_1 _16527_ (.A1(net6531),
    .A2(_11633_),
    .Y(_11634_),
    .B1(_11484_));
 sg13g2_a221oi_1 _16528_ (.B2(_11475_),
    .C1(_11610_),
    .B1(_09965_),
    .A1(net6531),
    .Y(_11635_),
    .A2(net6013));
 sg13g2_or2_1 _16529_ (.X(_11636_),
    .B(_11635_),
    .A(_11634_));
 sg13g2_nor2_2 _16530_ (.A(net6093),
    .B(_09965_),
    .Y(_11637_));
 sg13g2_a221oi_1 _16531_ (.B2(_11637_),
    .C1(_11439_),
    .B1(_11475_),
    .A1(net6015),
    .Y(_11638_),
    .A2(_11440_));
 sg13g2_nand4_1 _16532_ (.B(_11632_),
    .C(_11636_),
    .A(net5065),
    .Y(_11639_),
    .D(_11638_));
 sg13g2_o21ai_1 _16533_ (.B1(_11639_),
    .Y(_11640_),
    .A1(net2867),
    .A2(net5065));
 sg13g2_o21ai_1 _16534_ (.B1(_11630_),
    .Y(_00895_),
    .A1(net4720),
    .A2(_11640_));
 sg13g2_nand2_1 _16535_ (.Y(_11641_),
    .A(net6376),
    .B(net6436));
 sg13g2_a22oi_1 _16536_ (.Y(_11642_),
    .B1(_11637_),
    .B2(_09979_),
    .A2(_11507_),
    .A1(_09985_));
 sg13g2_nand2b_1 _16537_ (.Y(_11643_),
    .B(net6530),
    .A_N(_11642_));
 sg13g2_o21ai_1 _16538_ (.B1(net6511),
    .Y(_11644_),
    .A1(net6512),
    .A2(net6508));
 sg13g2_o21ai_1 _16539_ (.B1(_11644_),
    .Y(_11645_),
    .A1(net6530),
    .A2(net6087));
 sg13g2_a21oi_1 _16540_ (.A1(net6530),
    .A2(_11633_),
    .Y(_11646_),
    .B1(_11484_));
 sg13g2_a21o_1 _16541_ (.A2(_11645_),
    .A1(_11609_),
    .B1(_11646_),
    .X(_11647_));
 sg13g2_nand3_1 _16542_ (.B(_11643_),
    .C(_11647_),
    .A(net5064),
    .Y(_11648_));
 sg13g2_o21ai_1 _16543_ (.B1(_11648_),
    .Y(_11649_),
    .A1(net2541),
    .A2(net5064));
 sg13g2_o21ai_1 _16544_ (.B1(_11641_),
    .Y(_00896_),
    .A1(net4721),
    .A2(_11649_));
 sg13g2_nand2_1 _16545_ (.Y(_11650_),
    .A(net6415),
    .B(net6435));
 sg13g2_a21oi_1 _16546_ (.A1(net6529),
    .A2(_11633_),
    .Y(_11651_),
    .B1(_11484_));
 sg13g2_a21oi_1 _16547_ (.A1(net6529),
    .A2(_11644_),
    .Y(_11652_),
    .B1(net6087));
 sg13g2_a21oi_1 _16548_ (.A1(_11609_),
    .A2(_11652_),
    .Y(_11653_),
    .B1(_11651_));
 sg13g2_a221oi_1 _16549_ (.B2(net6529),
    .C1(_09991_),
    .B1(_11507_),
    .A1(net6526),
    .Y(_11654_),
    .A2(net6090));
 sg13g2_o21ai_1 _16550_ (.B1(net6094),
    .Y(_11655_),
    .A1(net6529),
    .A2(_09970_));
 sg13g2_o21ai_1 _16551_ (.B1(_11655_),
    .Y(_11656_),
    .A1(_09987_),
    .A2(_11654_));
 sg13g2_or3_1 _16552_ (.A(net5130),
    .B(_11653_),
    .C(_11656_),
    .X(_11657_));
 sg13g2_o21ai_1 _16553_ (.B1(_11657_),
    .Y(_11658_),
    .A1(net2402),
    .A2(net5064));
 sg13g2_o21ai_1 _16554_ (.B1(_11650_),
    .Y(_00897_),
    .A1(net4720),
    .A2(_11658_));
 sg13g2_nand2_1 _16555_ (.Y(_11659_),
    .A(net6415),
    .B(net6433));
 sg13g2_nand2b_1 _16556_ (.Y(_11660_),
    .B(_09990_),
    .A_N(net6528));
 sg13g2_a22oi_1 _16557_ (.Y(_11661_),
    .B1(net6087),
    .B2(_11660_),
    .A2(net6521),
    .A1(net6510));
 sg13g2_a21o_1 _16558_ (.A2(_11661_),
    .A1(net6090),
    .B1(_09987_),
    .X(_11662_));
 sg13g2_a21oi_1 _16559_ (.A1(net6528),
    .A2(_11633_),
    .Y(_11663_),
    .B1(_11484_));
 sg13g2_a221oi_1 _16560_ (.B2(net6528),
    .C1(net6087),
    .B1(_11644_),
    .A1(net6013),
    .Y(_11664_),
    .A2(_09975_));
 sg13g2_a21o_1 _16561_ (.A2(_11664_),
    .A1(_11608_),
    .B1(_11663_),
    .X(_11665_));
 sg13g2_o21ai_1 _16562_ (.B1(net6094),
    .Y(_11666_),
    .A1(net6528),
    .A2(_09970_));
 sg13g2_nand4_1 _16563_ (.B(_11662_),
    .C(_11665_),
    .A(net5062),
    .Y(_11667_),
    .D(_11666_));
 sg13g2_o21ai_1 _16564_ (.B1(_11667_),
    .Y(_11668_),
    .A1(net2453),
    .A2(net5064));
 sg13g2_o21ai_1 _16565_ (.B1(_11659_),
    .Y(_00898_),
    .A1(net4720),
    .A2(_11668_));
 sg13g2_a21o_1 _16566_ (.A2(_11633_),
    .A1(net6526),
    .B1(_11484_),
    .X(_11669_));
 sg13g2_o21ai_1 _16567_ (.B1(_11607_),
    .Y(_11670_),
    .A1(net5997),
    .A2(_11592_));
 sg13g2_a221oi_1 _16568_ (.B2(net6518),
    .C1(net6087),
    .B1(_11436_),
    .A1(net6526),
    .Y(_11671_),
    .A2(net6090));
 sg13g2_nor2_1 _16569_ (.A(net6526),
    .B(_09975_),
    .Y(_11672_));
 sg13g2_o21ai_1 _16570_ (.B1(_11671_),
    .Y(_11673_),
    .A1(_11540_),
    .A2(_11672_));
 sg13g2_nand2b_1 _16571_ (.Y(_11674_),
    .B(_11670_),
    .A_N(_11673_));
 sg13g2_a21oi_1 _16572_ (.A1(net6015),
    .A2(_09967_),
    .Y(_11675_),
    .B1(net6526));
 sg13g2_nand2_1 _16573_ (.Y(_11676_),
    .A(_09964_),
    .B(_11675_));
 sg13g2_a221oi_1 _16574_ (.B2(_11676_),
    .C1(net6512),
    .B1(_11644_),
    .A1(net6526),
    .Y(_11677_),
    .A2(net6086));
 sg13g2_a21o_1 _16575_ (.A2(net6090),
    .A1(net6519),
    .B1(_09991_),
    .X(_11678_));
 sg13g2_a22oi_1 _16576_ (.Y(_11679_),
    .B1(_11678_),
    .B2(_09986_),
    .A2(_11674_),
    .A1(_11669_));
 sg13g2_o21ai_1 _16577_ (.B1(_11679_),
    .Y(_11680_),
    .A1(net6092),
    .A2(_11677_));
 sg13g2_mux2_1 _16578_ (.A0(net2474),
    .A1(_11680_),
    .S(net5064),
    .X(_11681_));
 sg13g2_a22oi_1 _16579_ (.Y(_11682_),
    .B1(net4754),
    .B2(_11681_),
    .A2(net6431),
    .A1(net6373));
 sg13g2_inv_1 _16580_ (.Y(_00899_),
    .A(_11682_));
 sg13g2_nand2_1 _16581_ (.Y(_11683_),
    .A(net6363),
    .B(net2838));
 sg13g2_o21ai_1 _16582_ (.B1(_09986_),
    .Y(_11684_),
    .A1(net6515),
    .A2(_09991_));
 sg13g2_o21ai_1 _16583_ (.B1(net6516),
    .Y(_11685_),
    .A1(_09967_),
    .A2(net6086));
 sg13g2_a21oi_2 _16584_ (.B1(_11484_),
    .Y(_11686_),
    .A2(_11633_),
    .A1(net6516));
 sg13g2_nand2b_1 _16585_ (.Y(_11687_),
    .B(_11548_),
    .A_N(net5997));
 sg13g2_o21ai_1 _16586_ (.B1(_11456_),
    .Y(_11688_),
    .A1(_08028_),
    .A2(_09974_));
 sg13g2_a21oi_2 _16587_ (.B1(_11688_),
    .Y(_11689_),
    .A2(_09967_),
    .A1(net6515));
 sg13g2_a22oi_1 _16588_ (.Y(_11690_),
    .B1(_11607_),
    .B2(_11687_),
    .A2(_11461_),
    .A1(net6531));
 sg13g2_a21oi_1 _16589_ (.A1(_11689_),
    .A2(_11690_),
    .Y(_11691_),
    .B1(_11686_));
 sg13g2_o21ai_1 _16590_ (.B1(_11684_),
    .Y(_11692_),
    .A1(net6092),
    .A2(_11685_));
 sg13g2_or3_1 _16591_ (.A(net5130),
    .B(_11691_),
    .C(_11692_),
    .X(_11693_));
 sg13g2_o21ai_1 _16592_ (.B1(_11693_),
    .Y(_11694_),
    .A1(net2436),
    .A2(net5062));
 sg13g2_o21ai_1 _16593_ (.B1(_11683_),
    .Y(_00900_),
    .A1(net4722),
    .A2(_11694_));
 sg13g2_nand2_1 _16594_ (.Y(_11695_),
    .A(net6362),
    .B(net3209));
 sg13g2_a22oi_1 _16595_ (.Y(_11696_),
    .B1(net6088),
    .B2(net6524),
    .A2(_09966_),
    .A1(\soc_inst.core_instr_data[5] ));
 sg13g2_a21oi_1 _16596_ (.A1(_09992_),
    .A2(_11696_),
    .Y(_11697_),
    .B1(_09987_));
 sg13g2_a22oi_1 _16597_ (.Y(_11698_),
    .B1(_11507_),
    .B2(net6524),
    .A2(_11475_),
    .A1(_09965_));
 sg13g2_o21ai_1 _16598_ (.B1(_11607_),
    .Y(_11699_),
    .A1(net5997),
    .A2(_11582_));
 sg13g2_a22oi_1 _16599_ (.Y(_11700_),
    .B1(net6086),
    .B2(net6528),
    .A2(_11436_),
    .A1(net6525));
 sg13g2_nand3_1 _16600_ (.B(_11699_),
    .C(_11700_),
    .A(_11689_),
    .Y(_11701_));
 sg13g2_nand2b_1 _16601_ (.Y(_11702_),
    .B(_11701_),
    .A_N(_11686_));
 sg13g2_o21ai_1 _16602_ (.B1(_11702_),
    .Y(_11703_),
    .A1(net6092),
    .A2(_11698_));
 sg13g2_or3_1 _16603_ (.A(net5131),
    .B(_11697_),
    .C(_11703_),
    .X(_11704_));
 sg13g2_o21ai_1 _16604_ (.B1(_11704_),
    .Y(_11705_),
    .A1(net2549),
    .A2(net5063));
 sg13g2_o21ai_1 _16605_ (.B1(_11695_),
    .Y(_00901_),
    .A1(net4722),
    .A2(_11705_));
 sg13g2_nand2_1 _16606_ (.Y(_11706_),
    .A(net6363),
    .B(net2649));
 sg13g2_o21ai_1 _16607_ (.B1(_11458_),
    .Y(_11707_),
    .A1(net6523),
    .A2(_11560_));
 sg13g2_nand2b_1 _16608_ (.Y(_11708_),
    .B(_11562_),
    .A_N(net5997));
 sg13g2_a22oi_1 _16609_ (.Y(_11709_),
    .B1(_11607_),
    .B2(_11708_),
    .A2(_11461_),
    .A1(net6527));
 sg13g2_a21o_1 _16610_ (.A2(_11709_),
    .A1(_11689_),
    .B1(_11686_),
    .X(_11710_));
 sg13g2_a22oi_1 _16611_ (.Y(_11711_),
    .B1(net6086),
    .B2(net6523),
    .A2(_09967_),
    .A1(net6530));
 sg13g2_nand2b_1 _16612_ (.Y(_11712_),
    .B(net6094),
    .A_N(_11711_));
 sg13g2_nand4_1 _16613_ (.B(_11707_),
    .C(_11710_),
    .A(net5062),
    .Y(_11713_),
    .D(_11712_));
 sg13g2_o21ai_1 _16614_ (.B1(_11713_),
    .Y(_11714_),
    .A1(net2578),
    .A2(net5062));
 sg13g2_o21ai_1 _16615_ (.B1(_11706_),
    .Y(_00902_),
    .A1(net4722),
    .A2(_11714_));
 sg13g2_nand2_1 _16616_ (.Y(_11715_),
    .A(net6374),
    .B(net3159));
 sg13g2_o21ai_1 _16617_ (.B1(_11458_),
    .Y(_11716_),
    .A1(\soc_inst.core_instr_data[9] ),
    .A2(_11560_));
 sg13g2_o21ai_1 _16618_ (.B1(_11607_),
    .Y(_11717_),
    .A1(net5997),
    .A2(_11571_));
 sg13g2_nand2_1 _16619_ (.Y(_11718_),
    .A(_11486_),
    .B(_11689_));
 sg13g2_a21oi_1 _16620_ (.A1(\soc_inst.core_instr_data[9] ),
    .A2(_11436_),
    .Y(_11719_),
    .B1(_11718_));
 sg13g2_a21o_1 _16621_ (.A2(_11719_),
    .A1(_11717_),
    .B1(_11686_),
    .X(_11720_));
 sg13g2_nand3_1 _16622_ (.B(_11716_),
    .C(_11720_),
    .A(net5062),
    .Y(_11721_));
 sg13g2_o21ai_1 _16623_ (.B1(_11721_),
    .Y(_11722_),
    .A1(net2576),
    .A2(net5062));
 sg13g2_o21ai_1 _16624_ (.B1(_11715_),
    .Y(_00903_),
    .A1(net4719),
    .A2(_11722_));
 sg13g2_nand2_1 _16625_ (.Y(_11723_),
    .A(net6373),
    .B(net2729));
 sg13g2_o21ai_1 _16626_ (.B1(_11458_),
    .Y(_11724_),
    .A1(net6520),
    .A2(_11560_));
 sg13g2_nor2_1 _16627_ (.A(_11606_),
    .B(_11718_),
    .Y(_11725_));
 sg13g2_nand2_1 _16628_ (.Y(_11726_),
    .A(net6520),
    .B(_11436_));
 sg13g2_a21o_1 _16629_ (.A2(_11726_),
    .A1(_11725_),
    .B1(_11686_),
    .X(_11727_));
 sg13g2_nand3_1 _16630_ (.B(_11724_),
    .C(_11727_),
    .A(net5062),
    .Y(_11728_));
 sg13g2_o21ai_1 _16631_ (.B1(_11728_),
    .Y(_11729_),
    .A1(net2503),
    .A2(net5062));
 sg13g2_o21ai_1 _16632_ (.B1(_11723_),
    .Y(_00904_),
    .A1(net4722),
    .A2(_11729_));
 sg13g2_nand2_1 _16633_ (.Y(_11730_),
    .A(net6362),
    .B(net2743));
 sg13g2_a21oi_1 _16634_ (.A1(net6518),
    .A2(_09959_),
    .Y(_11731_),
    .B1(_09977_));
 sg13g2_a21oi_1 _16635_ (.A1(net6523),
    .A2(_11436_),
    .Y(_11732_),
    .B1(_11731_));
 sg13g2_a21oi_1 _16636_ (.A1(_11725_),
    .A2(_11732_),
    .Y(_11733_),
    .B1(_11686_));
 sg13g2_nand2b_1 _16637_ (.Y(_11734_),
    .B(net5130),
    .A_N(net1848));
 sg13g2_o21ai_1 _16638_ (.B1(_11734_),
    .Y(_11735_),
    .A1(net5130),
    .A2(_11733_));
 sg13g2_o21ai_1 _16639_ (.B1(_11730_),
    .Y(_00905_),
    .A1(net4722),
    .A2(_11735_));
 sg13g2_nand2_1 _16640_ (.Y(_11736_),
    .A(net6330),
    .B(net3325));
 sg13g2_nand2b_1 _16641_ (.Y(_11737_),
    .B(net5130),
    .A_N(net1446));
 sg13g2_a21oi_1 _16642_ (.A1(_11549_),
    .A2(_11725_),
    .Y(_11738_),
    .B1(_11686_));
 sg13g2_o21ai_1 _16643_ (.B1(_11737_),
    .Y(_11739_),
    .A1(net5130),
    .A2(_11738_));
 sg13g2_o21ai_1 _16644_ (.B1(_11736_),
    .Y(_00906_),
    .A1(net4722),
    .A2(_11739_));
 sg13g2_a22oi_1 _16645_ (.Y(_00907_),
    .B1(net4754),
    .B2(_07818_),
    .A2(_07910_),
    .A1(net6362));
 sg13g2_a22oi_1 _16646_ (.Y(_00908_),
    .B1(net4753),
    .B2(_07820_),
    .A2(_07909_),
    .A1(net6375));
 sg13g2_a22oi_1 _16647_ (.Y(_00909_),
    .B1(net4753),
    .B2(_07822_),
    .A2(_07912_),
    .A1(net6376));
 sg13g2_a22oi_1 _16648_ (.Y(_00910_),
    .B1(net4754),
    .B2(_07824_),
    .A2(_07911_),
    .A1(net6371));
 sg13g2_a22oi_1 _16649_ (.Y(_00911_),
    .B1(net4754),
    .B2(_07826_),
    .A2(_07913_),
    .A1(net6361));
 sg13g2_a22oi_1 _16650_ (.Y(_00912_),
    .B1(net4753),
    .B2(_07828_),
    .A2(_07914_),
    .A1(net6407));
 sg13g2_a22oi_1 _16651_ (.Y(_00913_),
    .B1(net4753),
    .B2(_07830_),
    .A2(_07915_),
    .A1(net6406));
 sg13g2_a22oi_1 _16652_ (.Y(_00914_),
    .B1(net4753),
    .B2(_07832_),
    .A2(_07916_),
    .A1(net6370));
 sg13g2_a22oi_1 _16653_ (.Y(_00915_),
    .B1(net4751),
    .B2(_07834_),
    .A2(_07917_),
    .A1(net6368));
 sg13g2_a22oi_1 _16654_ (.Y(_00916_),
    .B1(net4753),
    .B2(_07836_),
    .A2(_07918_),
    .A1(net6368));
 sg13g2_a22oi_1 _16655_ (.Y(_00917_),
    .B1(net4751),
    .B2(_07838_),
    .A2(_07919_),
    .A1(net6391));
 sg13g2_a22oi_1 _16656_ (.Y(_00918_),
    .B1(net4751),
    .B2(_07840_),
    .A2(_07920_),
    .A1(net6404));
 sg13g2_a22oi_1 _16657_ (.Y(_00919_),
    .B1(net4752),
    .B2(_07842_),
    .A2(_07921_),
    .A1(net6351));
 sg13g2_a22oi_1 _16658_ (.Y(_00920_),
    .B1(net4751),
    .B2(_07844_),
    .A2(_07922_),
    .A1(net6350));
 sg13g2_a22oi_1 _16659_ (.Y(_00921_),
    .B1(net4751),
    .B2(_07846_),
    .A2(_07923_),
    .A1(net6350));
 sg13g2_a22oi_1 _16660_ (.Y(_00922_),
    .B1(net4750),
    .B2(_07848_),
    .A2(_07924_),
    .A1(net6350));
 sg13g2_a22oi_1 _16661_ (.Y(_00923_),
    .B1(net4750),
    .B2(_07850_),
    .A2(_07925_),
    .A1(net6337));
 sg13g2_a22oi_1 _16662_ (.Y(_00924_),
    .B1(net4750),
    .B2(_07852_),
    .A2(_07926_),
    .A1(net6337));
 sg13g2_a22oi_1 _16663_ (.Y(_00925_),
    .B1(net4750),
    .B2(_07854_),
    .A2(_07927_),
    .A1(net6338));
 sg13g2_a22oi_1 _16664_ (.Y(_00926_),
    .B1(net4750),
    .B2(_07856_),
    .A2(_07928_),
    .A1(net6338));
 sg13g2_a22oi_1 _16665_ (.Y(_00927_),
    .B1(net4750),
    .B2(_07858_),
    .A2(_07929_),
    .A1(net6344));
 sg13g2_a22oi_1 _16666_ (.Y(_00928_),
    .B1(net4750),
    .B2(_07860_),
    .A2(_07930_),
    .A1(net6345));
 sg13g2_a22oi_1 _16667_ (.Y(_00929_),
    .B1(net4750),
    .B2(_07862_),
    .A2(_07931_),
    .A1(net6344));
 sg13g2_a22oi_1 _16668_ (.Y(_00930_),
    .B1(net4752),
    .B2(_07864_),
    .A2(_07932_),
    .A1(net6333));
 sg13g2_nor2_1 _16669_ (.A(net2451),
    .B(net4753),
    .Y(_11740_));
 sg13g2_a21oi_1 _16670_ (.A1(net5132),
    .A2(net4753),
    .Y(_00931_),
    .B1(_11740_));
 sg13g2_mux2_1 _16671_ (.A0(net644),
    .A1(net1936),
    .S(net6365),
    .X(_00932_));
 sg13g2_mux2_1 _16672_ (.A0(net394),
    .A1(net1893),
    .S(net6365),
    .X(_00933_));
 sg13g2_mux2_1 _16673_ (.A0(\soc_inst.cpu_core.ex_rs1_data[2] ),
    .A1(net1738),
    .S(net6359),
    .X(_00934_));
 sg13g2_mux2_1 _16674_ (.A0(net316),
    .A1(net1598),
    .S(net6374),
    .X(_00935_));
 sg13g2_mux2_1 _16675_ (.A0(net257),
    .A1(net1786),
    .S(net6365),
    .X(_00936_));
 sg13g2_mux2_1 _16676_ (.A0(net519),
    .A1(net1664),
    .S(net6379),
    .X(_00937_));
 sg13g2_mux2_1 _16677_ (.A0(net455),
    .A1(net2113),
    .S(net6330),
    .X(_00938_));
 sg13g2_mux2_1 _16678_ (.A0(net1197),
    .A1(net2390),
    .S(net6335),
    .X(_00939_));
 sg13g2_mux2_1 _16679_ (.A0(net260),
    .A1(net1413),
    .S(net6335),
    .X(_00940_));
 sg13g2_mux2_1 _16680_ (.A0(net206),
    .A1(net1456),
    .S(net6362),
    .X(_00941_));
 sg13g2_mux2_1 _16681_ (.A0(net243),
    .A1(net1479),
    .S(net6334),
    .X(_00942_));
 sg13g2_mux2_1 _16682_ (.A0(net326),
    .A1(net1582),
    .S(net6335),
    .X(_00943_));
 sg13g2_mux2_1 _16683_ (.A0(net231),
    .A1(net1299),
    .S(net6324),
    .X(_00944_));
 sg13g2_mux2_1 _16684_ (.A0(net288),
    .A1(net1452),
    .S(net6325),
    .X(_00945_));
 sg13g2_mux2_1 _16685_ (.A0(net367),
    .A1(net1378),
    .S(net6336),
    .X(_00946_));
 sg13g2_mux2_1 _16686_ (.A0(net729),
    .A1(net2221),
    .S(net6336),
    .X(_00947_));
 sg13g2_mux2_1 _16687_ (.A0(net275),
    .A1(net1787),
    .S(net6337),
    .X(_00948_));
 sg13g2_mux2_1 _16688_ (.A0(net217),
    .A1(net1716),
    .S(net6336),
    .X(_00949_));
 sg13g2_mux2_1 _16689_ (.A0(net1033),
    .A1(net2700),
    .S(net6338),
    .X(_00950_));
 sg13g2_mux2_1 _16690_ (.A0(net524),
    .A1(net1772),
    .S(net6337),
    .X(_00951_));
 sg13g2_mux2_1 _16691_ (.A0(net891),
    .A1(net2260),
    .S(net6343),
    .X(_00952_));
 sg13g2_mux2_1 _16692_ (.A0(net2223),
    .A1(net2445),
    .S(net6343),
    .X(_00953_));
 sg13g2_mux2_1 _16693_ (.A0(net885),
    .A1(net2337),
    .S(net6337),
    .X(_00954_));
 sg13g2_mux2_1 _16694_ (.A0(net1368),
    .A1(net2599),
    .S(net6336),
    .X(_00955_));
 sg13g2_mux2_1 _16695_ (.A0(net1279),
    .A1(net2674),
    .S(net6337),
    .X(_00956_));
 sg13g2_mux2_1 _16696_ (.A0(net732),
    .A1(net2145),
    .S(net6336),
    .X(_00957_));
 sg13g2_mux2_1 _16697_ (.A0(net214),
    .A1(net1504),
    .S(net6397),
    .X(_00958_));
 sg13g2_mux2_1 _16698_ (.A0(net320),
    .A1(net1591),
    .S(net6339),
    .X(_00959_));
 sg13g2_mux2_1 _16699_ (.A0(net328),
    .A1(net1627),
    .S(net6341),
    .X(_00960_));
 sg13g2_mux2_1 _16700_ (.A0(\soc_inst.cpu_core.ex_rs1_data[29] ),
    .A1(net2672),
    .S(net6317),
    .X(_00961_));
 sg13g2_mux2_1 _16701_ (.A0(net374),
    .A1(net1348),
    .S(net6336),
    .X(_00962_));
 sg13g2_mux2_1 _16702_ (.A0(net381),
    .A1(net1398),
    .S(net6353),
    .X(_00963_));
 sg13g2_a22oi_1 _16703_ (.Y(_11741_),
    .B1(net5307),
    .B2(net1886),
    .A2(net6375),
    .A1(net2480));
 sg13g2_inv_1 _16704_ (.Y(_00964_),
    .A(_11741_));
 sg13g2_a22oi_1 _16705_ (.Y(_11742_),
    .B1(net5307),
    .B2(net2013),
    .A2(net6375),
    .A1(net2833));
 sg13g2_inv_1 _16706_ (.Y(_00965_),
    .A(_11742_));
 sg13g2_a22oi_1 _16707_ (.Y(_11743_),
    .B1(net2936),
    .B2(net5311),
    .A2(net3016),
    .A1(net6373));
 sg13g2_inv_1 _16708_ (.Y(_00966_),
    .A(_11743_));
 sg13g2_a22oi_1 _16709_ (.Y(_11744_),
    .B1(net3065),
    .B2(net5305),
    .A2(net3051),
    .A1(net6375));
 sg13g2_inv_1 _16710_ (.Y(_00967_),
    .A(_11744_));
 sg13g2_a22oi_1 _16711_ (.Y(_11745_),
    .B1(net5305),
    .B2(net2877),
    .A2(net6413),
    .A1(net3050));
 sg13g2_inv_1 _16712_ (.Y(_00968_),
    .A(_11745_));
 sg13g2_a22oi_1 _16713_ (.Y(_11746_),
    .B1(net3174),
    .B2(net5309),
    .A2(net3182),
    .A1(net6414));
 sg13g2_inv_1 _16714_ (.Y(_00969_),
    .A(_11746_));
 sg13g2_a22oi_1 _16715_ (.Y(_11747_),
    .B1(net6452),
    .B2(net5308),
    .A2(net6306),
    .A1(net6413));
 sg13g2_inv_1 _16716_ (.Y(_00970_),
    .A(_11747_));
 sg13g2_a22oi_1 _16717_ (.Y(_11748_),
    .B1(net5305),
    .B2(net1906),
    .A2(net2416),
    .A1(net6378));
 sg13g2_inv_1 _16718_ (.Y(_00971_),
    .A(_11748_));
 sg13g2_a22oi_1 _16719_ (.Y(_11749_),
    .B1(net5306),
    .B2(net1270),
    .A2(net2345),
    .A1(net6378));
 sg13g2_inv_1 _16720_ (.Y(_00972_),
    .A(_11749_));
 sg13g2_a22oi_1 _16721_ (.Y(_11750_),
    .B1(net5306),
    .B2(net1265),
    .A2(net2153),
    .A1(net6377));
 sg13g2_inv_1 _16722_ (.Y(_00973_),
    .A(_11750_));
 sg13g2_a22oi_1 _16723_ (.Y(_11751_),
    .B1(net5306),
    .B2(net873),
    .A2(net1652),
    .A1(net6378));
 sg13g2_inv_1 _16724_ (.Y(_00974_),
    .A(_11751_));
 sg13g2_a22oi_1 _16725_ (.Y(_11752_),
    .B1(net5306),
    .B2(net1248),
    .A2(net1835),
    .A1(net6377));
 sg13g2_inv_1 _16726_ (.Y(_00975_),
    .A(_11752_));
 sg13g2_a22oi_1 _16727_ (.Y(_11753_),
    .B1(net3014),
    .B2(net5310),
    .A2(net3155),
    .A1(net6410));
 sg13g2_inv_1 _16728_ (.Y(_00976_),
    .A(_11753_));
 sg13g2_a22oi_1 _16729_ (.Y(_11754_),
    .B1(net2924),
    .B2(net5303),
    .A2(net3119),
    .A1(net6409));
 sg13g2_inv_1 _16730_ (.Y(_00977_),
    .A(_11754_));
 sg13g2_a22oi_1 _16731_ (.Y(_11755_),
    .B1(net2945),
    .B2(net5308),
    .A2(net2234),
    .A1(net6404));
 sg13g2_inv_1 _16732_ (.Y(_00978_),
    .A(_11755_));
 sg13g2_a22oi_1 _16733_ (.Y(_11756_),
    .B1(net5303),
    .B2(net6450),
    .A2(net360),
    .A1(net6395));
 sg13g2_inv_1 _16734_ (.Y(_00979_),
    .A(_11756_));
 sg13g2_a22oi_1 _16735_ (.Y(_11757_),
    .B1(net5307),
    .B2(net6448),
    .A2(net1350),
    .A1(net6360));
 sg13g2_inv_1 _16736_ (.Y(_00980_),
    .A(_11757_));
 sg13g2_a22oi_1 _16737_ (.Y(_11758_),
    .B1(net5300),
    .B2(net6445),
    .A2(net1545),
    .A1(net6391));
 sg13g2_inv_1 _16738_ (.Y(_00981_),
    .A(_11758_));
 sg13g2_a22oi_1 _16739_ (.Y(_11759_),
    .B1(net5307),
    .B2(net6444),
    .A2(net1363),
    .A1(net6367));
 sg13g2_inv_1 _16740_ (.Y(_00982_),
    .A(_11759_));
 sg13g2_a22oi_1 _16741_ (.Y(_11760_),
    .B1(net5307),
    .B2(net6443),
    .A2(net1864),
    .A1(net6369));
 sg13g2_inv_1 _16742_ (.Y(_00983_),
    .A(_11760_));
 sg13g2_and2_1 _16743_ (.A(net6438),
    .B(net5309),
    .X(_11761_));
 sg13g2_a21o_1 _16744_ (.A2(net630),
    .A1(net6388),
    .B1(net5102),
    .X(_00984_));
 sg13g2_a22oi_1 _16745_ (.Y(_11762_),
    .B1(net6436),
    .B2(net5304),
    .A2(net2501),
    .A1(net6353));
 sg13g2_inv_1 _16746_ (.Y(_00985_),
    .A(_11762_));
 sg13g2_a22oi_1 _16747_ (.Y(_11763_),
    .B1(net6435),
    .B2(net5300),
    .A2(net2556),
    .A1(net6355));
 sg13g2_inv_1 _16748_ (.Y(_00986_),
    .A(_11763_));
 sg13g2_a22oi_1 _16749_ (.Y(_11764_),
    .B1(net6433),
    .B2(net5303),
    .A2(net2885),
    .A1(net6392));
 sg13g2_inv_1 _16750_ (.Y(_00987_),
    .A(_11764_));
 sg13g2_a22oi_1 _16751_ (.Y(_11765_),
    .B1(net6431),
    .B2(net5304),
    .A2(net2286),
    .A1(net6354));
 sg13g2_inv_1 _16752_ (.Y(_00988_),
    .A(_11765_));
 sg13g2_a22oi_1 _16753_ (.Y(_11766_),
    .B1(net2838),
    .B2(net5300),
    .A2(net1121),
    .A1(net6352));
 sg13g2_inv_1 _16754_ (.Y(_00989_),
    .A(_11766_));
 sg13g2_a22oi_1 _16755_ (.Y(_11767_),
    .B1(\soc_inst.cpu_core.if_funct7[1] ),
    .B2(net5300),
    .A2(net2698),
    .A1(net6352));
 sg13g2_inv_1 _16756_ (.Y(_00990_),
    .A(net2699));
 sg13g2_a22oi_1 _16757_ (.Y(_11768_),
    .B1(net2649),
    .B2(net5300),
    .A2(net2613),
    .A1(net6352));
 sg13g2_inv_1 _16758_ (.Y(_00991_),
    .A(_11768_));
 sg13g2_a22oi_1 _16759_ (.Y(_11769_),
    .B1(\soc_inst.cpu_core.if_funct7[3] ),
    .B2(net5303),
    .A2(net2893),
    .A1(net6391));
 sg13g2_inv_1 _16760_ (.Y(_00992_),
    .A(net2894));
 sg13g2_a22oi_1 _16761_ (.Y(_11770_),
    .B1(net2729),
    .B2(net5300),
    .A2(net2609),
    .A1(net6356));
 sg13g2_inv_1 _16762_ (.Y(_00993_),
    .A(_11770_));
 sg13g2_nand2_1 _16763_ (.Y(_11771_),
    .A(net2743),
    .B(net5309));
 sg13g2_a22oi_1 _16764_ (.Y(_02607_),
    .B1(net2743),
    .B2(net5300),
    .A2(net2566),
    .A1(net6354));
 sg13g2_inv_1 _16765_ (.Y(_00994_),
    .A(_02607_));
 sg13g2_nand2_1 _16766_ (.Y(_02608_),
    .A(\soc_inst.cpu_core.if_funct7[6] ),
    .B(net5308));
 sg13g2_a22oi_1 _16767_ (.Y(_02609_),
    .B1(\soc_inst.cpu_core.if_funct7[6] ),
    .B2(net5300),
    .A2(net2726),
    .A1(net6367));
 sg13g2_inv_1 _16768_ (.Y(_00995_),
    .A(net2727));
 sg13g2_nand2b_2 _16769_ (.Y(_02610_),
    .B(net6445),
    .A_N(net6444));
 sg13g2_nand2_2 _16770_ (.Y(_02611_),
    .A(net6449),
    .B(net6446));
 sg13g2_nor3_1 _16771_ (.A(net6987),
    .B(_02610_),
    .C(_02611_),
    .Y(_02612_));
 sg13g2_nand2_1 _16772_ (.Y(_02613_),
    .A(\soc_inst.cpu_core.register_file.registers[23][0] ),
    .B(net5993));
 sg13g2_nor4_1 _16773_ (.A(net6449),
    .B(net6446),
    .C(_08135_),
    .D(_02610_),
    .Y(_02614_));
 sg13g2_nor2_1 _16774_ (.A(net6445),
    .B(net6444),
    .Y(_02615_));
 sg13g2_nand2b_2 _16775_ (.Y(_02616_),
    .B(net6446),
    .A_N(net6450));
 sg13g2_nor4_1 _16776_ (.A(net6445),
    .B(net6444),
    .C(net6442),
    .D(_02616_),
    .Y(_02617_));
 sg13g2_nand2b_2 _16777_ (.Y(_02618_),
    .B(net6444),
    .A_N(net6445));
 sg13g2_nand2b_2 _16778_ (.Y(_02619_),
    .B(net6450),
    .A_N(net6447));
 sg13g2_nor3_1 _16779_ (.A(net6441),
    .B(_02618_),
    .C(_02619_),
    .Y(_02620_));
 sg13g2_nand2_2 _16780_ (.Y(_02621_),
    .A(net6445),
    .B(net6444));
 sg13g2_nor3_1 _16781_ (.A(net6987),
    .B(_02611_),
    .C(_02621_),
    .Y(_02622_));
 sg13g2_nor3_1 _16782_ (.A(net6440),
    .B(_02610_),
    .C(_02616_),
    .Y(_02623_));
 sg13g2_nor3_1 _16783_ (.A(net6440),
    .B(_02616_),
    .C(_02621_),
    .Y(_02624_));
 sg13g2_nor3_1 _16784_ (.A(net6987),
    .B(_02616_),
    .C(_02618_),
    .Y(_02625_));
 sg13g2_nor3_1 _16785_ (.A(net6440),
    .B(_02611_),
    .C(_02618_),
    .Y(_02626_));
 sg13g2_nand2_2 _16786_ (.Y(_02627_),
    .A(net6442),
    .B(_02615_));
 sg13g2_nor2_1 _16787_ (.A(_02611_),
    .B(_02627_),
    .Y(_02628_));
 sg13g2_nor3_1 _16788_ (.A(net6440),
    .B(_02611_),
    .C(_02621_),
    .Y(_02629_));
 sg13g2_nor3_1 _16789_ (.A(net6987),
    .B(_02610_),
    .C(_02616_),
    .Y(_02630_));
 sg13g2_nor4_1 _16790_ (.A(\soc_inst.cpu_core.if_instr[17] ),
    .B(\soc_inst.cpu_core.if_instr[18] ),
    .C(net6442),
    .D(_02611_),
    .Y(_02631_));
 sg13g2_a22oi_1 _16791_ (.Y(_02632_),
    .B1(net5938),
    .B2(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][0] ));
 sg13g2_nor3_1 _16792_ (.A(_08135_),
    .B(_02616_),
    .C(_02621_),
    .Y(_02633_));
 sg13g2_nor2_1 _16793_ (.A(_02616_),
    .B(_02627_),
    .Y(_02634_));
 sg13g2_or2_1 _16794_ (.X(_02635_),
    .B(_02619_),
    .A(_08135_));
 sg13g2_nor2_1 _16795_ (.A(_02619_),
    .B(_02627_),
    .Y(_02636_));
 sg13g2_nor4_1 _16796_ (.A(net6449),
    .B(net6446),
    .C(net6440),
    .D(_02610_),
    .Y(_02637_));
 sg13g2_nor3_1 _16797_ (.A(net6449),
    .B(net6446),
    .C(_02627_),
    .Y(_02638_));
 sg13g2_nor2_1 _16798_ (.A(_02618_),
    .B(_02635_),
    .Y(_02639_));
 sg13g2_nor4_1 _16799_ (.A(net6448),
    .B(\soc_inst.cpu_core.if_instr[17] ),
    .C(\soc_inst.cpu_core.if_instr[18] ),
    .D(net6443),
    .Y(_02640_));
 sg13g2_nand3b_1 _16800_ (.B(net6987),
    .C(_02615_),
    .Y(_02641_),
    .A_N(net6447));
 sg13g2_nor2_1 _16801_ (.A(_02610_),
    .B(_02635_),
    .Y(_02642_));
 sg13g2_nor3_1 _16802_ (.A(net6441),
    .B(_02619_),
    .C(_02621_),
    .Y(_02643_));
 sg13g2_nor3_1 _16803_ (.A(net6987),
    .B(_02611_),
    .C(_02618_),
    .Y(_02644_));
 sg13g2_nor4_1 _16804_ (.A(net6449),
    .B(net6446),
    .C(net6987),
    .D(_02618_),
    .Y(_02645_));
 sg13g2_nor4_1 _16805_ (.A(net6449),
    .B(net6446),
    .C(net6440),
    .D(_02618_),
    .Y(_02646_));
 sg13g2_nor3_1 _16806_ (.A(net6441),
    .B(_02610_),
    .C(_02611_),
    .Y(_02647_));
 sg13g2_nor4_1 _16807_ (.A(net6449),
    .B(net6446),
    .C(net6440),
    .D(_02621_),
    .Y(_02648_));
 sg13g2_nor3_1 _16808_ (.A(net6440),
    .B(_02616_),
    .C(_02618_),
    .Y(_02649_));
 sg13g2_nor3_1 _16809_ (.A(net6441),
    .B(_02610_),
    .C(_02619_),
    .Y(_02650_));
 sg13g2_nor2_1 _16810_ (.A(_02621_),
    .B(_02635_),
    .Y(_02651_));
 sg13g2_nor4_1 _16811_ (.A(net6449),
    .B(net6447),
    .C(net6987),
    .D(_02621_),
    .Y(_02652_));
 sg13g2_a22oi_1 _16812_ (.Y(_02653_),
    .B1(net5907),
    .B2(\soc_inst.cpu_core.register_file.registers[24][0] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][0] ));
 sg13g2_a22oi_1 _16813_ (.Y(_02654_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][0] ));
 sg13g2_a22oi_1 _16814_ (.Y(_02655_),
    .B1(net5953),
    .B2(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][0] ));
 sg13g2_a22oi_1 _16815_ (.Y(_02656_),
    .B1(net5917),
    .B2(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][0] ));
 sg13g2_a22oi_1 _16816_ (.Y(_02657_),
    .B1(net5483),
    .B2(\soc_inst.cpu_core.register_file.registers[29][0] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][0] ));
 sg13g2_nand4_1 _16817_ (.B(_02653_),
    .C(_02656_),
    .A(_02632_),
    .Y(_02658_),
    .D(_02657_));
 sg13g2_a22oi_1 _16818_ (.Y(_02659_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][0] ));
 sg13g2_a22oi_1 _16819_ (.Y(_02660_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .A2(net5498),
    .A1(\soc_inst.cpu_core.register_file.registers[16][0] ));
 sg13g2_nand4_1 _16820_ (.B(_02655_),
    .C(_02659_),
    .A(_02613_),
    .Y(_02661_),
    .D(_02660_));
 sg13g2_a21oi_1 _16821_ (.A1(\soc_inst.cpu_core.register_file.registers[25][0] ),
    .A2(net5493),
    .Y(_02662_),
    .B1(net6082));
 sg13g2_a22oi_1 _16822_ (.Y(_02663_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][0] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][0] ));
 sg13g2_a22oi_1 _16823_ (.Y(_02664_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][0] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][0] ));
 sg13g2_nand4_1 _16824_ (.B(_02662_),
    .C(_02663_),
    .A(_02654_),
    .Y(_02665_),
    .D(_02664_));
 sg13g2_a22oi_1 _16825_ (.Y(_02666_),
    .B1(net5508),
    .B2(\soc_inst.cpu_core.register_file.registers[18][0] ),
    .A2(net5978),
    .A1(\soc_inst.cpu_core.register_file.registers[9][0] ));
 sg13g2_a22oi_1 _16826_ (.Y(_02667_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][0] ),
    .A2(net5968),
    .A1(\soc_inst.cpu_core.register_file.registers[6][0] ));
 sg13g2_a22oi_1 _16827_ (.Y(_02668_),
    .B1(net5948),
    .B2(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .A2(net5963),
    .A1(\soc_inst.cpu_core.register_file.registers[14][0] ));
 sg13g2_a22oi_1 _16828_ (.Y(_02669_),
    .B1(net5912),
    .B2(\soc_inst.cpu_core.register_file.registers[27][0] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][0] ));
 sg13g2_nand4_1 _16829_ (.B(_02667_),
    .C(_02668_),
    .A(_02666_),
    .Y(_02670_),
    .D(_02669_));
 sg13g2_or2_1 _16830_ (.X(_02671_),
    .B(_02670_),
    .A(_02665_));
 sg13g2_nor3_1 _16831_ (.A(_02658_),
    .B(_02661_),
    .C(_02671_),
    .Y(_02672_));
 sg13g2_nor2_1 _16832_ (.A(net6450),
    .B(net5921),
    .Y(_02673_));
 sg13g2_nor3_1 _16833_ (.A(net6395),
    .B(_11390_),
    .C(_02673_),
    .Y(_02674_));
 sg13g2_nand2b_2 _16834_ (.Y(_02675_),
    .B(net5303),
    .A_N(_02673_));
 sg13g2_o21ai_1 _16835_ (.B1(net5297),
    .Y(_02676_),
    .A1(net1209),
    .A2(net5924));
 sg13g2_or2_1 _16836_ (.X(_02677_),
    .B(_02676_),
    .A(_02672_));
 sg13g2_o21ai_1 _16837_ (.B1(_02677_),
    .Y(_00996_),
    .A1(net6152),
    .A2(_08029_));
 sg13g2_nand2_1 _16838_ (.Y(_02678_),
    .A(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .B(net5978));
 sg13g2_a22oi_1 _16839_ (.Y(_02679_),
    .B1(net5958),
    .B2(\soc_inst.cpu_core.register_file.registers[26][1] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][1] ));
 sg13g2_a22oi_1 _16840_ (.Y(_02680_),
    .B1(net5907),
    .B2(\soc_inst.cpu_core.register_file.registers[24][1] ),
    .A2(net5917),
    .A1(\soc_inst.cpu_core.register_file.registers[13][1] ));
 sg13g2_a22oi_1 _16841_ (.Y(_02681_),
    .B1(net5508),
    .B2(\soc_inst.cpu_core.register_file.registers[18][1] ),
    .A2(net5963),
    .A1(\soc_inst.cpu_core.register_file.registers[14][1] ));
 sg13g2_a22oi_1 _16842_ (.Y(_02682_),
    .B1(net5493),
    .B2(\soc_inst.cpu_core.register_file.registers[25][1] ),
    .A2(net5948),
    .A1(\soc_inst.cpu_core.register_file.registers[15][1] ));
 sg13g2_a22oi_1 _16843_ (.Y(_02683_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][1] ),
    .A2(net5938),
    .A1(\soc_inst.cpu_core.register_file.registers[3][1] ));
 sg13g2_a22oi_1 _16844_ (.Y(_02684_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][1] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][1] ));
 sg13g2_nand4_1 _16845_ (.B(_02682_),
    .C(_02683_),
    .A(_02679_),
    .Y(_02685_),
    .D(_02684_));
 sg13g2_a22oi_1 _16846_ (.Y(_02686_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][1] ));
 sg13g2_nand4_1 _16847_ (.B(_02680_),
    .C(_02681_),
    .A(_02678_),
    .Y(_02687_),
    .D(_02686_));
 sg13g2_nor2_1 _16848_ (.A(_02685_),
    .B(_02687_),
    .Y(_02688_));
 sg13g2_a21oi_1 _16849_ (.A1(\soc_inst.cpu_core.register_file.registers[20][1] ),
    .A2(net5988),
    .Y(_02689_),
    .B1(net6082));
 sg13g2_a22oi_1 _16850_ (.Y(_02690_),
    .B1(net5498),
    .B2(\soc_inst.cpu_core.register_file.registers[16][1] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][1] ));
 sg13g2_a22oi_1 _16851_ (.Y(_02691_),
    .B1(net5483),
    .B2(\soc_inst.cpu_core.register_file.registers[29][1] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][1] ));
 sg13g2_a22oi_1 _16852_ (.Y(_02692_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][1] ));
 sg13g2_nand4_1 _16853_ (.B(_02690_),
    .C(_02691_),
    .A(_02689_),
    .Y(_02693_),
    .D(_02692_));
 sg13g2_a22oi_1 _16854_ (.Y(_02694_),
    .B1(net5912),
    .B2(\soc_inst.cpu_core.register_file.registers[27][1] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][1] ));
 sg13g2_a22oi_1 _16855_ (.Y(_02695_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .A2(net5953),
    .A1(\soc_inst.cpu_core.register_file.registers[11][1] ));
 sg13g2_a22oi_1 _16856_ (.Y(_02696_),
    .B1(net5968),
    .B2(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][1] ));
 sg13g2_a22oi_1 _16857_ (.Y(_02697_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][1] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][1] ));
 sg13g2_nand4_1 _16858_ (.B(_02695_),
    .C(_02696_),
    .A(_02694_),
    .Y(_02698_),
    .D(_02697_));
 sg13g2_nor2_1 _16859_ (.A(_02693_),
    .B(_02698_),
    .Y(_02699_));
 sg13g2_o21ai_1 _16860_ (.B1(net5299),
    .Y(_02700_),
    .A1(net1139),
    .A2(net5924));
 sg13g2_a21oi_2 _16861_ (.B1(_02700_),
    .Y(_02701_),
    .A2(_02699_),
    .A1(_02688_));
 sg13g2_a21o_1 _16862_ (.A2(net3189),
    .A1(net6422),
    .B1(_02701_),
    .X(_00997_));
 sg13g2_a22oi_1 _16863_ (.Y(_02702_),
    .B1(net5948),
    .B2(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][2] ));
 sg13g2_nand2_1 _16864_ (.Y(_02703_),
    .A(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .B(net5978));
 sg13g2_a22oi_1 _16865_ (.Y(_02704_),
    .B1(net5508),
    .B2(\soc_inst.cpu_core.register_file.registers[18][2] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][2] ));
 sg13g2_a22oi_1 _16866_ (.Y(_02705_),
    .B1(net5917),
    .B2(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][2] ));
 sg13g2_a22oi_1 _16867_ (.Y(_02706_),
    .B1(net5493),
    .B2(\soc_inst.cpu_core.register_file.registers[25][2] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][2] ));
 sg13g2_a22oi_1 _16868_ (.Y(_02707_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .A2(net5498),
    .A1(\soc_inst.cpu_core.register_file.registers[16][2] ));
 sg13g2_a22oi_1 _16869_ (.Y(_02708_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][2] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][2] ));
 sg13g2_a22oi_1 _16870_ (.Y(_02709_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][2] ));
 sg13g2_a22oi_1 _16871_ (.Y(_02710_),
    .B1(net5953),
    .B2(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][2] ));
 sg13g2_a22oi_1 _16872_ (.Y(_02711_),
    .B1(net5912),
    .B2(\soc_inst.cpu_core.register_file.registers[27][2] ),
    .A2(net5968),
    .A1(\soc_inst.cpu_core.register_file.registers[6][2] ));
 sg13g2_nand4_1 _16873_ (.B(_02709_),
    .C(_02710_),
    .A(_02706_),
    .Y(_02712_),
    .D(_02711_));
 sg13g2_a22oi_1 _16874_ (.Y(_02713_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][2] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][2] ));
 sg13g2_nand4_1 _16875_ (.B(_02707_),
    .C(_02708_),
    .A(_02703_),
    .Y(_02714_),
    .D(_02713_));
 sg13g2_nor2_1 _16876_ (.A(_02712_),
    .B(_02714_),
    .Y(_02715_));
 sg13g2_a21oi_1 _16877_ (.A1(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .A2(net5938),
    .Y(_02716_),
    .B1(net6082));
 sg13g2_a22oi_1 _16878_ (.Y(_02717_),
    .B1(net5963),
    .B2(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][2] ));
 sg13g2_a22oi_1 _16879_ (.Y(_02718_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][2] ),
    .A2(net5483),
    .A1(\soc_inst.cpu_core.register_file.registers[29][2] ));
 sg13g2_nand4_1 _16880_ (.B(_02716_),
    .C(_02717_),
    .A(_02704_),
    .Y(_02719_),
    .D(_02718_));
 sg13g2_a22oi_1 _16881_ (.Y(_02720_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .A2(net5907),
    .A1(\soc_inst.cpu_core.register_file.registers[24][2] ));
 sg13g2_a22oi_1 _16882_ (.Y(_02721_),
    .B1(net5503),
    .B2(\soc_inst.cpu_core.register_file.registers[17][2] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][2] ));
 sg13g2_nand4_1 _16883_ (.B(_02705_),
    .C(_02720_),
    .A(_02702_),
    .Y(_02722_),
    .D(_02721_));
 sg13g2_nor2_1 _16884_ (.A(_02719_),
    .B(_02722_),
    .Y(_02723_));
 sg13g2_o21ai_1 _16885_ (.B1(net5297),
    .Y(_02724_),
    .A1(net507),
    .A2(net5923));
 sg13g2_a21oi_2 _16886_ (.B1(_02724_),
    .Y(_02725_),
    .A2(_02723_),
    .A1(_02715_));
 sg13g2_a21o_1 _16887_ (.A2(net3283),
    .A1(net6424),
    .B1(_02725_),
    .X(_00998_));
 sg13g2_a22oi_1 _16888_ (.Y(_02726_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][3] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][3] ));
 sg13g2_a22oi_1 _16889_ (.Y(_02727_),
    .B1(net5972),
    .B2(\soc_inst.cpu_core.register_file.registers[31][3] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][3] ));
 sg13g2_nand2_1 _16890_ (.Y(_02728_),
    .A(\soc_inst.cpu_core.register_file.registers[27][3] ),
    .B(net5911));
 sg13g2_a22oi_1 _16891_ (.Y(_02729_),
    .B1(net5901),
    .B2(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .A2(net5927),
    .A1(\soc_inst.cpu_core.register_file.registers[4][3] ));
 sg13g2_a22oi_1 _16892_ (.Y(_02730_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][3] ));
 sg13g2_a22oi_1 _16893_ (.Y(_02731_),
    .B1(net5957),
    .B2(\soc_inst.cpu_core.register_file.registers[26][3] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][3] ));
 sg13g2_a22oi_1 _16894_ (.Y(_02732_),
    .B1(net5906),
    .B2(\soc_inst.cpu_core.register_file.registers[24][3] ),
    .A2(net5502),
    .A1(\soc_inst.cpu_core.register_file.registers[17][3] ));
 sg13g2_a22oi_1 _16895_ (.Y(_02733_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][3] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][3] ));
 sg13g2_nand4_1 _16896_ (.B(_02731_),
    .C(_02732_),
    .A(_02727_),
    .Y(_02734_),
    .D(_02733_));
 sg13g2_a22oi_1 _16897_ (.Y(_02735_),
    .B1(net5891),
    .B2(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][3] ));
 sg13g2_a22oi_1 _16898_ (.Y(_02736_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][3] ),
    .A2(net5916),
    .A1(\soc_inst.cpu_core.register_file.registers[13][3] ));
 sg13g2_nand4_1 _16899_ (.B(_02729_),
    .C(_02735_),
    .A(_02728_),
    .Y(_02737_),
    .D(_02736_));
 sg13g2_a21oi_1 _16900_ (.A1(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .A2(net5967),
    .Y(_02738_),
    .B1(net6081));
 sg13g2_a22oi_1 _16901_ (.Y(_02739_),
    .B1(net5487),
    .B2(\soc_inst.cpu_core.register_file.registers[21][3] ),
    .A2(net5942),
    .A1(\soc_inst.cpu_core.register_file.registers[22][3] ));
 sg13g2_nand4_1 _16902_ (.B(_02730_),
    .C(_02738_),
    .A(_02726_),
    .Y(_02740_),
    .D(_02739_));
 sg13g2_a22oi_1 _16903_ (.Y(_02741_),
    .B1(net5492),
    .B2(\soc_inst.cpu_core.register_file.registers[25][3] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][3] ));
 sg13g2_a22oi_1 _16904_ (.Y(_02742_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .A2(net5932),
    .A1(\soc_inst.cpu_core.register_file.registers[30][3] ));
 sg13g2_a22oi_1 _16905_ (.Y(_02743_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][3] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][3] ));
 sg13g2_a22oi_1 _16906_ (.Y(_02744_),
    .B1(net5507),
    .B2(\soc_inst.cpu_core.register_file.registers[18][3] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][3] ));
 sg13g2_nand4_1 _16907_ (.B(_02742_),
    .C(_02743_),
    .A(_02741_),
    .Y(_02745_),
    .D(_02744_));
 sg13g2_or2_1 _16908_ (.X(_02746_),
    .B(_02745_),
    .A(_02740_));
 sg13g2_nor3_2 _16909_ (.A(_02734_),
    .B(_02737_),
    .C(_02746_),
    .Y(_02747_));
 sg13g2_o21ai_1 _16910_ (.B1(net5297),
    .Y(_02748_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .A2(net5922));
 sg13g2_or2_1 _16911_ (.X(_02749_),
    .B(_02748_),
    .A(_02747_));
 sg13g2_o21ai_1 _16912_ (.B1(_02749_),
    .Y(_00999_),
    .A1(net6145),
    .A2(_08031_));
 sg13g2_a22oi_1 _16913_ (.Y(_02750_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][4] ));
 sg13g2_nand2_1 _16914_ (.Y(_02751_),
    .A(\soc_inst.cpu_core.register_file.registers[23][4] ),
    .B(net5994));
 sg13g2_a22oi_1 _16915_ (.Y(_02752_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .A2(net5929),
    .A1(\soc_inst.cpu_core.register_file.registers[4][4] ));
 sg13g2_a22oi_1 _16916_ (.Y(_02753_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][4] ),
    .A2(net5504),
    .A1(\soc_inst.cpu_core.register_file.registers[17][4] ));
 sg13g2_a22oi_1 _16917_ (.Y(_02754_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .A2(net5494),
    .A1(\soc_inst.cpu_core.register_file.registers[25][4] ));
 sg13g2_a22oi_1 _16918_ (.Y(_02755_),
    .B1(net5939),
    .B2(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][4] ));
 sg13g2_a22oi_1 _16919_ (.Y(_02756_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][4] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][4] ));
 sg13g2_nand4_1 _16920_ (.B(_02753_),
    .C(_02755_),
    .A(_02752_),
    .Y(_02757_),
    .D(_02756_));
 sg13g2_a22oi_1 _16921_ (.Y(_02758_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .A2(net5903),
    .A1(\soc_inst.cpu_core.register_file.registers[8][4] ));
 sg13g2_a22oi_1 _16922_ (.Y(_02759_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][4] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][4] ));
 sg13g2_nand4_1 _16923_ (.B(_02751_),
    .C(_02758_),
    .A(_02750_),
    .Y(_02760_),
    .D(_02759_));
 sg13g2_a21oi_1 _16924_ (.A1(\soc_inst.cpu_core.register_file.registers[20][4] ),
    .A2(net5989),
    .Y(_02761_),
    .B1(net6083));
 sg13g2_a22oi_1 _16925_ (.Y(_02762_),
    .B1(net5969),
    .B2(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][4] ));
 sg13g2_a22oi_1 _16926_ (.Y(_02763_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][4] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][4] ));
 sg13g2_nand4_1 _16927_ (.B(_02761_),
    .C(_02762_),
    .A(_02754_),
    .Y(_02764_),
    .D(_02763_));
 sg13g2_a22oi_1 _16928_ (.Y(_02765_),
    .B1(net5509),
    .B2(\soc_inst.cpu_core.register_file.registers[18][4] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][4] ));
 sg13g2_a22oi_1 _16929_ (.Y(_02766_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .A2(net5489),
    .A1(\soc_inst.cpu_core.register_file.registers[21][4] ));
 sg13g2_a22oi_1 _16930_ (.Y(_02767_),
    .B1(net5949),
    .B2(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][4] ));
 sg13g2_a22oi_1 _16931_ (.Y(_02768_),
    .B1(net5913),
    .B2(\soc_inst.cpu_core.register_file.registers[27][4] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][4] ));
 sg13g2_nand4_1 _16932_ (.B(_02766_),
    .C(_02767_),
    .A(_02765_),
    .Y(_02769_),
    .D(_02768_));
 sg13g2_or2_1 _16933_ (.X(_02770_),
    .B(_02769_),
    .A(_02764_));
 sg13g2_nor3_2 _16934_ (.A(_02757_),
    .B(_02760_),
    .C(_02770_),
    .Y(_02771_));
 sg13g2_o21ai_1 _16935_ (.B1(net5299),
    .Y(_02772_),
    .A1(net444),
    .A2(net5926));
 sg13g2_or2_1 _16936_ (.X(_02773_),
    .B(_02772_),
    .A(_02771_));
 sg13g2_o21ai_1 _16937_ (.B1(_02773_),
    .Y(_01000_),
    .A1(net6152),
    .A2(_08039_));
 sg13g2_nand2_1 _16938_ (.Y(_02774_),
    .A(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .B(net5885));
 sg13g2_a22oi_1 _16939_ (.Y(_02775_),
    .B1(net5971),
    .B2(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .A2(net5981),
    .A1(\soc_inst.cpu_core.register_file.registers[9][5] ));
 sg13g2_a22oi_1 _16940_ (.Y(_02776_),
    .B1(net5511),
    .B2(\soc_inst.cpu_core.register_file.registers[18][5] ),
    .A2(net5991),
    .A1(\soc_inst.cpu_core.register_file.registers[20][5] ));
 sg13g2_a22oi_1 _16941_ (.Y(_02777_),
    .B1(net5931),
    .B2(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .A2(net5951),
    .A1(\soc_inst.cpu_core.register_file.registers[15][5] ));
 sg13g2_a22oi_1 _16942_ (.Y(_02778_),
    .B1(net5900),
    .B2(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .A2(net5961),
    .A1(\soc_inst.cpu_core.register_file.registers[26][5] ));
 sg13g2_a22oi_1 _16943_ (.Y(_02779_),
    .B1(net5491),
    .B2(\soc_inst.cpu_core.register_file.registers[21][5] ),
    .A2(net5941),
    .A1(\soc_inst.cpu_core.register_file.registers[3][5] ));
 sg13g2_a22oi_1 _16944_ (.Y(_02780_),
    .B1(net5915),
    .B2(\soc_inst.cpu_core.register_file.registers[27][5] ),
    .A2(net5516),
    .A1(\soc_inst.cpu_core.register_file.registers[19][5] ));
 sg13g2_nand4_1 _16945_ (.B(_02778_),
    .C(_02779_),
    .A(_02775_),
    .Y(_02781_),
    .D(_02780_));
 sg13g2_a22oi_1 _16946_ (.Y(_02782_),
    .B1(net5895),
    .B2(\soc_inst.cpu_core.register_file.registers[12][5] ),
    .A2(net5501),
    .A1(\soc_inst.cpu_core.register_file.registers[16][5] ));
 sg13g2_a22oi_1 _16947_ (.Y(_02783_),
    .B1(net5880),
    .B2(\soc_inst.cpu_core.register_file.registers[28][5] ),
    .A2(net5486),
    .A1(\soc_inst.cpu_core.register_file.registers[29][5] ));
 sg13g2_nand4_1 _16948_ (.B(_02777_),
    .C(_02782_),
    .A(_02774_),
    .Y(_02784_),
    .D(_02783_));
 sg13g2_nor2_1 _16949_ (.A(_02781_),
    .B(_02784_),
    .Y(_02785_));
 sg13g2_a21oi_1 _16950_ (.A1(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .A2(net5890),
    .Y(_02786_),
    .B1(net6085));
 sg13g2_a22oi_1 _16951_ (.Y(_02787_),
    .B1(net5496),
    .B2(\soc_inst.cpu_core.register_file.registers[25][5] ),
    .A2(net5936),
    .A1(\soc_inst.cpu_core.register_file.registers[30][5] ));
 sg13g2_a22oi_1 _16952_ (.Y(_02788_),
    .B1(net5946),
    .B2(\soc_inst.cpu_core.register_file.registers[22][5] ),
    .A2(net5976),
    .A1(\soc_inst.cpu_core.register_file.registers[31][5] ));
 sg13g2_nand4_1 _16953_ (.B(_02786_),
    .C(_02787_),
    .A(_02776_),
    .Y(_02789_),
    .D(_02788_));
 sg13g2_a22oi_1 _16954_ (.Y(_02790_),
    .B1(net5986),
    .B2(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .A2(net5996),
    .A1(\soc_inst.cpu_core.register_file.registers[23][5] ));
 sg13g2_a22oi_1 _16955_ (.Y(_02791_),
    .B1(net5910),
    .B2(\soc_inst.cpu_core.register_file.registers[24][5] ),
    .A2(net5956),
    .A1(\soc_inst.cpu_core.register_file.registers[11][5] ));
 sg13g2_a22oi_1 _16956_ (.Y(_02792_),
    .B1(net5920),
    .B2(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .A2(net5506),
    .A1(\soc_inst.cpu_core.register_file.registers[17][5] ));
 sg13g2_a22oi_1 _16957_ (.Y(_02793_),
    .B1(net5905),
    .B2(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][5] ));
 sg13g2_nand4_1 _16958_ (.B(_02791_),
    .C(_02792_),
    .A(_02790_),
    .Y(_02794_),
    .D(_02793_));
 sg13g2_nor2_1 _16959_ (.A(_02789_),
    .B(_02794_),
    .Y(_02795_));
 sg13g2_a21oi_2 _16960_ (.B1(_02675_),
    .Y(_02796_),
    .A2(_02795_),
    .A1(_02785_));
 sg13g2_o21ai_1 _16961_ (.B1(_02796_),
    .Y(_02797_),
    .A1(net1044),
    .A2(net5924));
 sg13g2_o21ai_1 _16962_ (.B1(_02797_),
    .Y(_01001_),
    .A1(net6153),
    .A2(_08037_));
 sg13g2_a22oi_1 _16963_ (.Y(_02798_),
    .B1(net5483),
    .B2(\soc_inst.cpu_core.register_file.registers[29][6] ),
    .A2(net5917),
    .A1(\soc_inst.cpu_core.register_file.registers[13][6] ));
 sg13g2_nand2_1 _16964_ (.Y(_02799_),
    .A(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .B(net5978));
 sg13g2_a22oi_1 _16965_ (.Y(_02800_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .A2(net5498),
    .A1(\soc_inst.cpu_core.register_file.registers[16][6] ));
 sg13g2_a22oi_1 _16966_ (.Y(_02801_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][6] ),
    .A2(net5953),
    .A1(\soc_inst.cpu_core.register_file.registers[11][6] ));
 sg13g2_a22oi_1 _16967_ (.Y(_02802_),
    .B1(net5907),
    .B2(\soc_inst.cpu_core.register_file.registers[24][6] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][6] ));
 sg13g2_a22oi_1 _16968_ (.Y(_02803_),
    .B1(net5948),
    .B2(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][6] ));
 sg13g2_a22oi_1 _16969_ (.Y(_02804_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .A2(net5963),
    .A1(\soc_inst.cpu_core.register_file.registers[14][6] ));
 sg13g2_a22oi_1 _16970_ (.Y(_02805_),
    .B1(net5513),
    .B2(\soc_inst.cpu_core.register_file.registers[19][6] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][6] ));
 sg13g2_a22oi_1 _16971_ (.Y(_02806_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][6] ));
 sg13g2_a22oi_1 _16972_ (.Y(_02807_),
    .B1(net5968),
    .B2(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][6] ));
 sg13g2_a22oi_1 _16973_ (.Y(_02808_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][6] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][6] ));
 sg13g2_nand4_1 _16974_ (.B(_02806_),
    .C(_02807_),
    .A(_02802_),
    .Y(_02809_),
    .D(_02808_));
 sg13g2_a22oi_1 _16975_ (.Y(_02810_),
    .B1(net5493),
    .B2(\soc_inst.cpu_core.register_file.registers[25][6] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][6] ));
 sg13g2_nand4_1 _16976_ (.B(_02803_),
    .C(_02804_),
    .A(_02799_),
    .Y(_02811_),
    .D(_02810_));
 sg13g2_nor2_1 _16977_ (.A(_02809_),
    .B(_02811_),
    .Y(_02812_));
 sg13g2_a21oi_1 _16978_ (.A1(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .A2(net5938),
    .Y(_02813_),
    .B1(net6082));
 sg13g2_a22oi_1 _16979_ (.Y(_02814_),
    .B1(net5928),
    .B2(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .A2(net5508),
    .A1(\soc_inst.cpu_core.register_file.registers[18][6] ));
 sg13g2_nand4_1 _16980_ (.B(_02805_),
    .C(_02813_),
    .A(_02798_),
    .Y(_02815_),
    .D(_02814_));
 sg13g2_a22oi_1 _16981_ (.Y(_02816_),
    .B1(net5912),
    .B2(\soc_inst.cpu_core.register_file.registers[27][6] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][6] ));
 sg13g2_a22oi_1 _16982_ (.Y(_02817_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][6] ));
 sg13g2_nand4_1 _16983_ (.B(_02801_),
    .C(_02816_),
    .A(_02800_),
    .Y(_02818_),
    .D(_02817_));
 sg13g2_nor2_1 _16984_ (.A(_02815_),
    .B(_02818_),
    .Y(_02819_));
 sg13g2_a21oi_2 _16985_ (.B1(_02675_),
    .Y(_02820_),
    .A2(_02819_),
    .A1(_02812_));
 sg13g2_o21ai_1 _16986_ (.B1(_02820_),
    .Y(_02821_),
    .A1(net1094),
    .A2(net5924));
 sg13g2_o21ai_1 _16987_ (.B1(_02821_),
    .Y(_01002_),
    .A1(net6152),
    .A2(_08035_));
 sg13g2_nand2_1 _16988_ (.Y(_02822_),
    .A(\soc_inst.cpu_core.register_file.registers[9][7] ),
    .B(net5979));
 sg13g2_a22oi_1 _16989_ (.Y(_02823_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][7] ),
    .A2(net5494),
    .A1(\soc_inst.cpu_core.register_file.registers[25][7] ));
 sg13g2_a22oi_1 _16990_ (.Y(_02824_),
    .B1(net5934),
    .B2(\soc_inst.cpu_core.register_file.registers[30][7] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][7] ));
 sg13g2_a22oi_1 _16991_ (.Y(_02825_),
    .B1(net5949),
    .B2(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][7] ));
 sg13g2_a22oi_1 _16992_ (.Y(_02826_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][7] ));
 sg13g2_a22oi_1 _16993_ (.Y(_02827_),
    .B1(net5969),
    .B2(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][7] ));
 sg13g2_a22oi_1 _16994_ (.Y(_02828_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][7] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][7] ));
 sg13g2_nand4_1 _16995_ (.B(_02826_),
    .C(_02827_),
    .A(_02823_),
    .Y(_02829_),
    .D(_02828_));
 sg13g2_a22oi_1 _16996_ (.Y(_02830_),
    .B1(net5489),
    .B2(\soc_inst.cpu_core.register_file.registers[21][7] ),
    .A2(net5509),
    .A1(\soc_inst.cpu_core.register_file.registers[18][7] ));
 sg13g2_a22oi_1 _16997_ (.Y(_02831_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .A2(net5965),
    .A1(\soc_inst.cpu_core.register_file.registers[14][7] ));
 sg13g2_nand4_1 _16998_ (.B(_02825_),
    .C(_02830_),
    .A(_02822_),
    .Y(_02832_),
    .D(_02831_));
 sg13g2_nor2_1 _16999_ (.A(_02829_),
    .B(_02832_),
    .Y(_02833_));
 sg13g2_a21oi_1 _17000_ (.A1(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .A2(net5939),
    .Y(_02834_),
    .B1(net6083));
 sg13g2_a22oi_1 _17001_ (.Y(_02835_),
    .B1(net5929),
    .B2(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][7] ));
 sg13g2_a22oi_1 _17002_ (.Y(_02836_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .A2(net5504),
    .A1(\soc_inst.cpu_core.register_file.registers[17][7] ));
 sg13g2_nand4_1 _17003_ (.B(_02834_),
    .C(_02835_),
    .A(_02824_),
    .Y(_02837_),
    .D(_02836_));
 sg13g2_a22oi_1 _17004_ (.Y(_02838_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][7] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][7] ));
 sg13g2_a22oi_1 _17005_ (.Y(_02839_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .A2(net5903),
    .A1(\soc_inst.cpu_core.register_file.registers[8][7] ));
 sg13g2_a22oi_1 _17006_ (.Y(_02840_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .A2(net5913),
    .A1(\soc_inst.cpu_core.register_file.registers[27][7] ));
 sg13g2_a22oi_1 _17007_ (.Y(_02841_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][7] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][7] ));
 sg13g2_nand4_1 _17008_ (.B(_02839_),
    .C(_02840_),
    .A(_02838_),
    .Y(_02842_),
    .D(_02841_));
 sg13g2_nor2_1 _17009_ (.A(_02837_),
    .B(_02842_),
    .Y(_02843_));
 sg13g2_a21oi_2 _17010_ (.B1(_02675_),
    .Y(_02844_),
    .A2(_02843_),
    .A1(_02833_));
 sg13g2_o21ai_1 _17011_ (.B1(_02844_),
    .Y(_02845_),
    .A1(net798),
    .A2(net5923));
 sg13g2_o21ai_1 _17012_ (.B1(_02845_),
    .Y(_01003_),
    .A1(net6152),
    .A2(_08033_));
 sg13g2_nand2_1 _17013_ (.Y(_02846_),
    .A(\soc_inst.cpu_core.register_file.registers[27][8] ),
    .B(net5912));
 sg13g2_a22oi_1 _17014_ (.Y(_02847_),
    .B1(net5963),
    .B2(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][8] ));
 sg13g2_a22oi_1 _17015_ (.Y(_02848_),
    .B1(net5907),
    .B2(\soc_inst.cpu_core.register_file.registers[24][8] ),
    .A2(net5948),
    .A1(\soc_inst.cpu_core.register_file.registers[15][8] ));
 sg13g2_a22oi_1 _17016_ (.Y(_02849_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][8] ));
 sg13g2_a22oi_1 _17017_ (.Y(_02850_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][8] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][8] ));
 sg13g2_a22oi_1 _17018_ (.Y(_02851_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][8] ));
 sg13g2_a22oi_1 _17019_ (.Y(_02852_),
    .B1(net5917),
    .B2(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .A2(net5938),
    .A1(\soc_inst.cpu_core.register_file.registers[3][8] ));
 sg13g2_a22oi_1 _17020_ (.Y(_02853_),
    .B1(net5493),
    .B2(\soc_inst.cpu_core.register_file.registers[25][8] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][8] ));
 sg13g2_nand4_1 _17021_ (.B(_02850_),
    .C(_02852_),
    .A(_02849_),
    .Y(_02854_),
    .D(_02853_));
 sg13g2_a22oi_1 _17022_ (.Y(_02855_),
    .B1(net5508),
    .B2(\soc_inst.cpu_core.register_file.registers[18][8] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][8] ));
 sg13g2_a22oi_1 _17023_ (.Y(_02856_),
    .B1(net5498),
    .B2(\soc_inst.cpu_core.register_file.registers[16][8] ),
    .A2(net5953),
    .A1(\soc_inst.cpu_core.register_file.registers[11][8] ));
 sg13g2_nand4_1 _17024_ (.B(_02851_),
    .C(_02855_),
    .A(_02846_),
    .Y(_02857_),
    .D(_02856_));
 sg13g2_a21oi_1 _17025_ (.A1(\soc_inst.cpu_core.register_file.registers[29][8] ),
    .A2(net5483),
    .Y(_02858_),
    .B1(net6082));
 sg13g2_a22oi_1 _17026_ (.Y(_02859_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][8] ));
 sg13g2_a22oi_1 _17027_ (.Y(_02860_),
    .B1(net5968),
    .B2(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][8] ));
 sg13g2_a22oi_1 _17028_ (.Y(_02861_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][8] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][8] ));
 sg13g2_nand4_1 _17029_ (.B(_02859_),
    .C(_02860_),
    .A(_02858_),
    .Y(_02862_),
    .D(_02861_));
 sg13g2_a22oi_1 _17030_ (.Y(_02863_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][8] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][8] ));
 sg13g2_a22oi_1 _17031_ (.Y(_02864_),
    .B1(net5943),
    .B2(\soc_inst.cpu_core.register_file.registers[22][8] ),
    .A2(net5978),
    .A1(\soc_inst.cpu_core.register_file.registers[9][8] ));
 sg13g2_nand4_1 _17032_ (.B(_02848_),
    .C(_02863_),
    .A(_02847_),
    .Y(_02865_),
    .D(_02864_));
 sg13g2_or2_1 _17033_ (.X(_02866_),
    .B(_02865_),
    .A(_02862_));
 sg13g2_nor3_2 _17034_ (.A(_02854_),
    .B(_02857_),
    .C(_02866_),
    .Y(_02867_));
 sg13g2_o21ai_1 _17035_ (.B1(net5297),
    .Y(_02868_),
    .A1(net488),
    .A2(net5923));
 sg13g2_or2_1 _17036_ (.X(_02869_),
    .B(_02868_),
    .A(_02867_));
 sg13g2_o21ai_1 _17037_ (.B1(_02869_),
    .Y(_01004_),
    .A1(net6148),
    .A2(_08054_));
 sg13g2_a22oi_1 _17038_ (.Y(_02870_),
    .B1(net5889),
    .B2(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .A2(net5510),
    .A1(\soc_inst.cpu_core.register_file.registers[18][9] ));
 sg13g2_a22oi_1 _17039_ (.Y(_02871_),
    .B1(net5930),
    .B2(\soc_inst.cpu_core.register_file.registers[4][9] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][9] ));
 sg13g2_nand2_1 _17040_ (.Y(_02872_),
    .A(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .B(net5904));
 sg13g2_a22oi_1 _17041_ (.Y(_02873_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .A2(net5960),
    .A1(\soc_inst.cpu_core.register_file.registers[26][9] ));
 sg13g2_a22oi_1 _17042_ (.Y(_02874_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][9] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][9] ));
 sg13g2_a22oi_1 _17043_ (.Y(_02875_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][9] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][9] ));
 sg13g2_a22oi_1 _17044_ (.Y(_02876_),
    .B1(net5964),
    .B2(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][9] ));
 sg13g2_nand4_1 _17045_ (.B(_02871_),
    .C(_02873_),
    .A(_02870_),
    .Y(_02877_),
    .D(_02876_));
 sg13g2_a22oi_1 _17046_ (.Y(_02878_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][9] ),
    .A2(net5950),
    .A1(\soc_inst.cpu_core.register_file.registers[15][9] ));
 sg13g2_a22oi_1 _17047_ (.Y(_02879_),
    .B1(net5495),
    .B2(\soc_inst.cpu_core.register_file.registers[25][9] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][9] ));
 sg13g2_nand4_1 _17048_ (.B(_02875_),
    .C(_02878_),
    .A(_02872_),
    .Y(_02880_),
    .D(_02879_));
 sg13g2_a21oi_1 _17049_ (.A1(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .A2(net5894),
    .Y(_02881_),
    .B1(net6084));
 sg13g2_a22oi_1 _17050_ (.Y(_02882_),
    .B1(net5485),
    .B2(\soc_inst.cpu_core.register_file.registers[29][9] ),
    .A2(net5935),
    .A1(\soc_inst.cpu_core.register_file.registers[30][9] ));
 sg13g2_a22oi_1 _17051_ (.Y(_02883_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][9] ));
 sg13g2_nand4_1 _17052_ (.B(_02881_),
    .C(_02882_),
    .A(_02874_),
    .Y(_02884_),
    .D(_02883_));
 sg13g2_a22oi_1 _17053_ (.Y(_02885_),
    .B1(net5505),
    .B2(\soc_inst.cpu_core.register_file.registers[17][9] ),
    .A2(net5945),
    .A1(\soc_inst.cpu_core.register_file.registers[22][9] ));
 sg13g2_a22oi_1 _17054_ (.Y(_02886_),
    .B1(net5940),
    .B2(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .A2(net5515),
    .A1(\soc_inst.cpu_core.register_file.registers[19][9] ));
 sg13g2_a22oi_1 _17055_ (.Y(_02887_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][9] ),
    .A2(net5970),
    .A1(\soc_inst.cpu_core.register_file.registers[6][9] ));
 sg13g2_a22oi_1 _17056_ (.Y(_02888_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .A2(net5914),
    .A1(\soc_inst.cpu_core.register_file.registers[27][9] ));
 sg13g2_nand4_1 _17057_ (.B(_02886_),
    .C(_02887_),
    .A(_02885_),
    .Y(_02889_),
    .D(_02888_));
 sg13g2_or2_1 _17058_ (.X(_02890_),
    .B(_02889_),
    .A(_02884_));
 sg13g2_nor3_2 _17059_ (.A(_02877_),
    .B(_02880_),
    .C(_02890_),
    .Y(_02891_));
 sg13g2_o21ai_1 _17060_ (.B1(net5297),
    .Y(_02892_),
    .A1(net673),
    .A2(net5923));
 sg13g2_or2_1 _17061_ (.X(_02893_),
    .B(_02892_),
    .A(_02891_));
 sg13g2_o21ai_1 _17062_ (.B1(_02893_),
    .Y(_01005_),
    .A1(net6155),
    .A2(_08052_));
 sg13g2_nand2_1 _17063_ (.Y(_02894_),
    .A(\soc_inst.cpu_core.register_file.registers[25][10] ),
    .B(net5495));
 sg13g2_a22oi_1 _17064_ (.Y(_02895_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .A2(net5515),
    .A1(\soc_inst.cpu_core.register_file.registers[19][10] ));
 sg13g2_a22oi_1 _17065_ (.Y(_02896_),
    .B1(net5980),
    .B2(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][10] ));
 sg13g2_a22oi_1 _17066_ (.Y(_02897_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][10] ),
    .A2(net5505),
    .A1(\soc_inst.cpu_core.register_file.registers[17][10] ));
 sg13g2_a22oi_1 _17067_ (.Y(_02898_),
    .B1(net5940),
    .B2(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .A2(net5945),
    .A1(\soc_inst.cpu_core.register_file.registers[22][10] ));
 sg13g2_a22oi_1 _17068_ (.Y(_02899_),
    .B1(net5485),
    .B2(\soc_inst.cpu_core.register_file.registers[29][10] ),
    .A2(net5889),
    .A1(\soc_inst.cpu_core.register_file.registers[10][10] ));
 sg13g2_a22oi_1 _17069_ (.Y(_02900_),
    .B1(net5935),
    .B2(\soc_inst.cpu_core.register_file.registers[30][10] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][10] ));
 sg13g2_nand4_1 _17070_ (.B(_02898_),
    .C(_02899_),
    .A(_02897_),
    .Y(_02901_),
    .D(_02900_));
 sg13g2_a22oi_1 _17071_ (.Y(_02902_),
    .B1(net5894),
    .B2(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .A2(net5510),
    .A1(\soc_inst.cpu_core.register_file.registers[18][10] ));
 sg13g2_a22oi_1 _17072_ (.Y(_02903_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][10] ));
 sg13g2_a22oi_1 _17073_ (.Y(_02904_),
    .B1(net5960),
    .B2(\soc_inst.cpu_core.register_file.registers[26][10] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][10] ));
 sg13g2_a22oi_1 _17074_ (.Y(_02905_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][10] ),
    .A2(net5970),
    .A1(\soc_inst.cpu_core.register_file.registers[6][10] ));
 sg13g2_nand4_1 _17075_ (.B(_02903_),
    .C(_02904_),
    .A(_02896_),
    .Y(_02906_),
    .D(_02905_));
 sg13g2_a22oi_1 _17076_ (.Y(_02907_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][10] ),
    .A2(net5914),
    .A1(\soc_inst.cpu_core.register_file.registers[27][10] ));
 sg13g2_a22oi_1 _17077_ (.Y(_02908_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][10] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][10] ));
 sg13g2_nand4_1 _17078_ (.B(_02902_),
    .C(_02907_),
    .A(_02894_),
    .Y(_02909_),
    .D(_02908_));
 sg13g2_or2_1 _17079_ (.X(_02910_),
    .B(_02909_),
    .A(_02906_));
 sg13g2_a21oi_1 _17080_ (.A1(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .A2(net5904),
    .Y(_02911_),
    .B1(net6084));
 sg13g2_a22oi_1 _17081_ (.Y(_02912_),
    .B1(net5950),
    .B2(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][10] ));
 sg13g2_a22oi_1 _17082_ (.Y(_02913_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .A2(net5930),
    .A1(\soc_inst.cpu_core.register_file.registers[4][10] ));
 sg13g2_nand4_1 _17083_ (.B(_02911_),
    .C(_02912_),
    .A(_02895_),
    .Y(_02914_),
    .D(_02913_));
 sg13g2_nor3_2 _17084_ (.A(_02901_),
    .B(_02910_),
    .C(_02914_),
    .Y(_02915_));
 sg13g2_o21ai_1 _17085_ (.B1(net5299),
    .Y(_02916_),
    .A1(net684),
    .A2(net5923));
 sg13g2_or2_1 _17086_ (.X(_02917_),
    .B(_02916_),
    .A(_02915_));
 sg13g2_o21ai_1 _17087_ (.B1(_02917_),
    .Y(_01006_),
    .A1(net6155),
    .A2(_08050_));
 sg13g2_nand2_1 _17088_ (.Y(_02918_),
    .A(\soc_inst.cpu_core.register_file.registers[24][11] ),
    .B(net5907));
 sg13g2_a22oi_1 _17089_ (.Y(_02919_),
    .B1(net5978),
    .B2(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][11] ));
 sg13g2_a22oi_1 _17090_ (.Y(_02920_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .A2(net5933),
    .A1(\soc_inst.cpu_core.register_file.registers[30][11] ));
 sg13g2_a22oi_1 _17091_ (.Y(_02921_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][11] ));
 sg13g2_a22oi_1 _17092_ (.Y(_02922_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .A2(net5983),
    .A1(\soc_inst.cpu_core.register_file.registers[2][11] ));
 sg13g2_a22oi_1 _17093_ (.Y(_02923_),
    .B1(net5968),
    .B2(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][11] ));
 sg13g2_a22oi_1 _17094_ (.Y(_02924_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][11] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][11] ));
 sg13g2_nand4_1 _17095_ (.B(_02922_),
    .C(_02923_),
    .A(_02919_),
    .Y(_02925_),
    .D(_02924_));
 sg13g2_a22oi_1 _17096_ (.Y(_02926_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .A2(net5902),
    .A1(\soc_inst.cpu_core.register_file.registers[8][11] ));
 sg13g2_a22oi_1 _17097_ (.Y(_02927_),
    .B1(net5498),
    .B2(\soc_inst.cpu_core.register_file.registers[16][11] ),
    .A2(net5953),
    .A1(\soc_inst.cpu_core.register_file.registers[11][11] ));
 sg13g2_nand4_1 _17098_ (.B(_02921_),
    .C(_02926_),
    .A(_02918_),
    .Y(_02928_),
    .D(_02927_));
 sg13g2_a21oi_1 _17099_ (.A1(\soc_inst.cpu_core.register_file.registers[29][11] ),
    .A2(net5483),
    .Y(_02929_),
    .B1(net6082));
 sg13g2_a22oi_1 _17100_ (.Y(_02930_),
    .B1(net5948),
    .B2(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .A2(net5963),
    .A1(\soc_inst.cpu_core.register_file.registers[14][11] ));
 sg13g2_a22oi_1 _17101_ (.Y(_02931_),
    .B1(net5917),
    .B2(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][11] ));
 sg13g2_nand4_1 _17102_ (.B(_02929_),
    .C(_02930_),
    .A(_02920_),
    .Y(_02932_),
    .D(_02931_));
 sg13g2_a22oi_1 _17103_ (.Y(_02933_),
    .B1(net5938),
    .B2(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][11] ));
 sg13g2_a22oi_1 _17104_ (.Y(_02934_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][11] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][11] ));
 sg13g2_a22oi_1 _17105_ (.Y(_02935_),
    .B1(net5508),
    .B2(\soc_inst.cpu_core.register_file.registers[18][11] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][11] ));
 sg13g2_a22oi_1 _17106_ (.Y(_02936_),
    .B1(net5912),
    .B2(\soc_inst.cpu_core.register_file.registers[27][11] ),
    .A2(net5493),
    .A1(\soc_inst.cpu_core.register_file.registers[25][11] ));
 sg13g2_nand4_1 _17107_ (.B(_02934_),
    .C(_02935_),
    .A(_02933_),
    .Y(_02937_),
    .D(_02936_));
 sg13g2_or2_1 _17108_ (.X(_02938_),
    .B(_02937_),
    .A(_02932_));
 sg13g2_nor3_2 _17109_ (.A(_02925_),
    .B(_02928_),
    .C(_02938_),
    .Y(_02939_));
 sg13g2_o21ai_1 _17110_ (.B1(net5299),
    .Y(_02940_),
    .A1(net991),
    .A2(net5923));
 sg13g2_or2_1 _17111_ (.X(_02941_),
    .B(_02940_),
    .A(_02939_));
 sg13g2_o21ai_1 _17112_ (.B1(_02941_),
    .Y(_01007_),
    .A1(net6145),
    .A2(_08049_));
 sg13g2_nand2_1 _17113_ (.Y(_02942_),
    .A(\soc_inst.cpu_core.register_file.registers[24][12] ),
    .B(net5908));
 sg13g2_a22oi_1 _17114_ (.Y(_02943_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][12] ),
    .A2(net5965),
    .A1(\soc_inst.cpu_core.register_file.registers[14][12] ));
 sg13g2_a22oi_1 _17115_ (.Y(_02944_),
    .B1(net5949),
    .B2(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .A2(net5969),
    .A1(\soc_inst.cpu_core.register_file.registers[6][12] ));
 sg13g2_a22oi_1 _17116_ (.Y(_02945_),
    .B1(net5903),
    .B2(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][12] ));
 sg13g2_a22oi_1 _17117_ (.Y(_02946_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][12] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][12] ));
 sg13g2_a22oi_1 _17118_ (.Y(_02947_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][12] ));
 sg13g2_a22oi_1 _17119_ (.Y(_02948_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][12] ),
    .A2(net5504),
    .A1(\soc_inst.cpu_core.register_file.registers[17][12] ));
 sg13g2_nand4_1 _17120_ (.B(_02946_),
    .C(_02947_),
    .A(_02943_),
    .Y(_02949_),
    .D(_02948_));
 sg13g2_a22oi_1 _17121_ (.Y(_02950_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][12] ));
 sg13g2_a22oi_1 _17122_ (.Y(_02951_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .A2(net5939),
    .A1(\soc_inst.cpu_core.register_file.registers[3][12] ));
 sg13g2_nand4_1 _17123_ (.B(_02945_),
    .C(_02950_),
    .A(_02942_),
    .Y(_02952_),
    .D(_02951_));
 sg13g2_a21oi_1 _17124_ (.A1(\soc_inst.cpu_core.register_file.registers[16][12] ),
    .A2(net5499),
    .Y(_02953_),
    .B1(net6083));
 sg13g2_a22oi_1 _17125_ (.Y(_02954_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][12] ));
 sg13g2_a22oi_1 _17126_ (.Y(_02955_),
    .B1(net5929),
    .B2(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][12] ));
 sg13g2_nand4_1 _17127_ (.B(_02953_),
    .C(_02954_),
    .A(_02944_),
    .Y(_02956_),
    .D(_02955_));
 sg13g2_a22oi_1 _17128_ (.Y(_02957_),
    .B1(net5489),
    .B2(\soc_inst.cpu_core.register_file.registers[21][12] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][12] ));
 sg13g2_a22oi_1 _17129_ (.Y(_02958_),
    .B1(net5959),
    .B2(\soc_inst.cpu_core.register_file.registers[26][12] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][12] ));
 sg13g2_a22oi_1 _17130_ (.Y(_02959_),
    .B1(net5509),
    .B2(\soc_inst.cpu_core.register_file.registers[18][12] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][12] ));
 sg13g2_a22oi_1 _17131_ (.Y(_02960_),
    .B1(net5913),
    .B2(\soc_inst.cpu_core.register_file.registers[27][12] ),
    .A2(net5494),
    .A1(\soc_inst.cpu_core.register_file.registers[25][12] ));
 sg13g2_nand4_1 _17132_ (.B(_02958_),
    .C(_02959_),
    .A(_02957_),
    .Y(_02961_),
    .D(_02960_));
 sg13g2_or2_1 _17133_ (.X(_02962_),
    .B(_02961_),
    .A(_02956_));
 sg13g2_nor3_2 _17134_ (.A(_02949_),
    .B(_02952_),
    .C(_02962_),
    .Y(_02963_));
 sg13g2_o21ai_1 _17135_ (.B1(net5296),
    .Y(_02964_),
    .A1(net479),
    .A2(net5922));
 sg13g2_or2_1 _17136_ (.X(_02965_),
    .B(_02964_),
    .A(_02963_));
 sg13g2_o21ai_1 _17137_ (.B1(_02965_),
    .Y(_01008_),
    .A1(net6148),
    .A2(_08047_));
 sg13g2_nand2_1 _17138_ (.Y(_02966_),
    .A(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .B(net5903));
 sg13g2_a22oi_1 _17139_ (.Y(_02967_),
    .B1(net5914),
    .B2(\soc_inst.cpu_core.register_file.registers[27][13] ),
    .A2(net5970),
    .A1(\soc_inst.cpu_core.register_file.registers[6][13] ));
 sg13g2_a22oi_1 _17140_ (.Y(_02968_),
    .B1(net5894),
    .B2(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .A2(net5908),
    .A1(\soc_inst.cpu_core.register_file.registers[24][13] ));
 sg13g2_a22oi_1 _17141_ (.Y(_02969_),
    .B1(net5505),
    .B2(\soc_inst.cpu_core.register_file.registers[17][13] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][13] ));
 sg13g2_a22oi_1 _17142_ (.Y(_02970_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][13] ));
 sg13g2_a22oi_1 _17143_ (.Y(_02971_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][13] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][13] ));
 sg13g2_a22oi_1 _17144_ (.Y(_02972_),
    .B1(net5939),
    .B2(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][13] ));
 sg13g2_a22oi_1 _17145_ (.Y(_02973_),
    .B1(net5965),
    .B2(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][13] ));
 sg13g2_a22oi_1 _17146_ (.Y(_02974_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .A2(net5509),
    .A1(\soc_inst.cpu_core.register_file.registers[18][13] ));
 sg13g2_nand4_1 _17147_ (.B(_02972_),
    .C(_02973_),
    .A(_02970_),
    .Y(_02975_),
    .D(_02974_));
 sg13g2_a22oi_1 _17148_ (.Y(_02976_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][13] ),
    .A2(net5949),
    .A1(\soc_inst.cpu_core.register_file.registers[15][13] ));
 sg13g2_a22oi_1 _17149_ (.Y(_02977_),
    .B1(net5494),
    .B2(\soc_inst.cpu_core.register_file.registers[25][13] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][13] ));
 sg13g2_nand4_1 _17150_ (.B(_02971_),
    .C(_02976_),
    .A(_02966_),
    .Y(_02978_),
    .D(_02977_));
 sg13g2_or2_1 _17151_ (.X(_02979_),
    .B(_02978_),
    .A(_02975_));
 sg13g2_a21oi_1 _17152_ (.A1(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .A2(net5899),
    .Y(_02980_),
    .B1(net6084));
 sg13g2_a22oi_1 _17153_ (.Y(_02981_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][13] ),
    .A2(net5935),
    .A1(\soc_inst.cpu_core.register_file.registers[30][13] ));
 sg13g2_a22oi_1 _17154_ (.Y(_02982_),
    .B1(net5485),
    .B2(\soc_inst.cpu_core.register_file.registers[29][13] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][13] ));
 sg13g2_nand4_1 _17155_ (.B(_02980_),
    .C(_02981_),
    .A(_02967_),
    .Y(_02983_),
    .D(_02982_));
 sg13g2_a22oi_1 _17156_ (.Y(_02984_),
    .B1(net5945),
    .B2(\soc_inst.cpu_core.register_file.registers[22][13] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][13] ));
 sg13g2_a22oi_1 _17157_ (.Y(_02985_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .A2(net5930),
    .A1(\soc_inst.cpu_core.register_file.registers[4][13] ));
 sg13g2_nand4_1 _17158_ (.B(_02969_),
    .C(_02984_),
    .A(_02968_),
    .Y(_02986_),
    .D(_02985_));
 sg13g2_nor3_2 _17159_ (.A(_02979_),
    .B(_02983_),
    .C(_02986_),
    .Y(_02987_));
 sg13g2_o21ai_1 _17160_ (.B1(net5296),
    .Y(_02988_),
    .A1(net808),
    .A2(net5921));
 sg13g2_or2_1 _17161_ (.X(_02989_),
    .B(_02988_),
    .A(_02987_));
 sg13g2_o21ai_1 _17162_ (.B1(_02989_),
    .Y(_01009_),
    .A1(net6143),
    .A2(_08045_));
 sg13g2_a22oi_1 _17163_ (.Y(_02990_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][14] ),
    .A2(net5497),
    .A1(\soc_inst.cpu_core.register_file.registers[16][14] ));
 sg13g2_nand2_1 _17164_ (.Y(_02991_),
    .A(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .B(net5977));
 sg13g2_a22oi_1 _17165_ (.Y(_02992_),
    .B1(net5492),
    .B2(\soc_inst.cpu_core.register_file.registers[25][14] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][14] ));
 sg13g2_a22oi_1 _17166_ (.Y(_02993_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][14] ));
 sg13g2_a22oi_1 _17167_ (.Y(_02994_),
    .B1(net5901),
    .B2(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][14] ));
 sg13g2_a22oi_1 _17168_ (.Y(_02995_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .A2(net5927),
    .A1(\soc_inst.cpu_core.register_file.registers[4][14] ));
 sg13g2_a22oi_1 _17169_ (.Y(_02996_),
    .B1(net5947),
    .B2(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .A2(net5967),
    .A1(\soc_inst.cpu_core.register_file.registers[6][14] ));
 sg13g2_a22oi_1 _17170_ (.Y(_02997_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][14] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][14] ));
 sg13g2_a22oi_1 _17171_ (.Y(_02998_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][14] ),
    .A2(net5942),
    .A1(\soc_inst.cpu_core.register_file.registers[22][14] ));
 sg13g2_a22oi_1 _17172_ (.Y(_02999_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .A2(net5502),
    .A1(\soc_inst.cpu_core.register_file.registers[17][14] ));
 sg13g2_nand4_1 _17173_ (.B(_02997_),
    .C(_02998_),
    .A(_02993_),
    .Y(_03000_),
    .D(_02999_));
 sg13g2_a22oi_1 _17174_ (.Y(_03001_),
    .B1(net5891),
    .B2(\soc_inst.cpu_core.register_file.registers[12][14] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][14] ));
 sg13g2_nand4_1 _17175_ (.B(_02994_),
    .C(_02995_),
    .A(_02991_),
    .Y(_03002_),
    .D(_03001_));
 sg13g2_nor2_1 _17176_ (.A(_03000_),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_a21oi_1 _17177_ (.A1(\soc_inst.cpu_core.register_file.registers[21][14] ),
    .A2(net5487),
    .Y(_03004_),
    .B1(net6081));
 sg13g2_a22oi_1 _17178_ (.Y(_03005_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][14] ));
 sg13g2_a22oi_1 _17179_ (.Y(_03006_),
    .B1(net5932),
    .B2(\soc_inst.cpu_core.register_file.registers[30][14] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][14] ));
 sg13g2_nand4_1 _17180_ (.B(_03004_),
    .C(_03005_),
    .A(_02992_),
    .Y(_03007_),
    .D(_03006_));
 sg13g2_a22oi_1 _17181_ (.Y(_03008_),
    .B1(net5906),
    .B2(\soc_inst.cpu_core.register_file.registers[24][14] ),
    .A2(net5507),
    .A1(\soc_inst.cpu_core.register_file.registers[18][14] ));
 sg13g2_a22oi_1 _17182_ (.Y(_03009_),
    .B1(net5957),
    .B2(\soc_inst.cpu_core.register_file.registers[26][14] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][14] ));
 sg13g2_nand4_1 _17183_ (.B(_02996_),
    .C(_03008_),
    .A(_02990_),
    .Y(_03010_),
    .D(_03009_));
 sg13g2_nor2_1 _17184_ (.A(_03007_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_o21ai_1 _17185_ (.B1(net5296),
    .Y(_03012_),
    .A1(net839),
    .A2(net5921));
 sg13g2_a21o_2 _17186_ (.A2(_03011_),
    .A1(_03003_),
    .B1(_03012_),
    .X(_03013_));
 sg13g2_o21ai_1 _17187_ (.B1(_03013_),
    .Y(_01010_),
    .A1(net6146),
    .A2(_08043_));
 sg13g2_nand2_1 _17188_ (.Y(_03014_),
    .A(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .B(net5903));
 sg13g2_a22oi_1 _17189_ (.Y(_03015_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][15] ));
 sg13g2_a22oi_1 _17190_ (.Y(_03016_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .A2(net5929),
    .A1(\soc_inst.cpu_core.register_file.registers[4][15] ));
 sg13g2_a22oi_1 _17191_ (.Y(_03017_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][15] ));
 sg13g2_a22oi_1 _17192_ (.Y(_03018_),
    .B1(net5913),
    .B2(\soc_inst.cpu_core.register_file.registers[27][15] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][15] ));
 sg13g2_a22oi_1 _17193_ (.Y(_03019_),
    .B1(net5494),
    .B2(\soc_inst.cpu_core.register_file.registers[25][15] ),
    .A2(net5939),
    .A1(\soc_inst.cpu_core.register_file.registers[3][15] ));
 sg13g2_a22oi_1 _17194_ (.Y(_03020_),
    .B1(net5489),
    .B2(\soc_inst.cpu_core.register_file.registers[21][15] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][15] ));
 sg13g2_a22oi_1 _17195_ (.Y(_03021_),
    .B1(net5965),
    .B2(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][15] ));
 sg13g2_a22oi_1 _17196_ (.Y(_03022_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][15] ));
 sg13g2_nand4_1 _17197_ (.B(_03020_),
    .C(_03021_),
    .A(_03016_),
    .Y(_03023_),
    .D(_03022_));
 sg13g2_a22oi_1 _17198_ (.Y(_03024_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][15] ),
    .A2(net5949),
    .A1(\soc_inst.cpu_core.register_file.registers[15][15] ));
 sg13g2_a22oi_1 _17199_ (.Y(_03025_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][15] ));
 sg13g2_nand4_1 _17200_ (.B(_03019_),
    .C(_03024_),
    .A(_03014_),
    .Y(_03026_),
    .D(_03025_));
 sg13g2_or2_1 _17201_ (.X(_03027_),
    .B(_03026_),
    .A(_03023_));
 sg13g2_a21oi_1 _17202_ (.A1(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .A2(net5969),
    .Y(_03028_),
    .B1(net6083));
 sg13g2_a22oi_1 _17203_ (.Y(_03029_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][15] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][15] ));
 sg13g2_a22oi_1 _17204_ (.Y(_03030_),
    .B1(net5504),
    .B2(\soc_inst.cpu_core.register_file.registers[17][15] ),
    .A2(net5509),
    .A1(\soc_inst.cpu_core.register_file.registers[18][15] ));
 sg13g2_nand4_1 _17205_ (.B(_03028_),
    .C(_03029_),
    .A(_03015_),
    .Y(_03031_),
    .D(_03030_));
 sg13g2_a22oi_1 _17206_ (.Y(_03032_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][15] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][15] ));
 sg13g2_a22oi_1 _17207_ (.Y(_03033_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][15] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][15] ));
 sg13g2_nand4_1 _17208_ (.B(_03018_),
    .C(_03032_),
    .A(_03017_),
    .Y(_03034_),
    .D(_03033_));
 sg13g2_nor3_2 _17209_ (.A(_03027_),
    .B(_03031_),
    .C(_03034_),
    .Y(_03035_));
 sg13g2_o21ai_1 _17210_ (.B1(net5296),
    .Y(_03036_),
    .A1(net641),
    .A2(net5921));
 sg13g2_or2_1 _17211_ (.X(_03037_),
    .B(_03036_),
    .A(_03035_));
 sg13g2_o21ai_1 _17212_ (.B1(_03037_),
    .Y(_01011_),
    .A1(net6144),
    .A2(_08041_));
 sg13g2_nand2_1 _17213_ (.Y(_03038_),
    .A(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .B(net5903));
 sg13g2_a22oi_1 _17214_ (.Y(_03039_),
    .B1(net5929),
    .B2(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][16] ));
 sg13g2_a22oi_1 _17215_ (.Y(_03040_),
    .B1(net5514),
    .B2(\soc_inst.cpu_core.register_file.registers[19][16] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][16] ));
 sg13g2_a22oi_1 _17216_ (.Y(_03041_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][16] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][16] ));
 sg13g2_a22oi_1 _17217_ (.Y(_03042_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][16] ),
    .A2(net5504),
    .A1(\soc_inst.cpu_core.register_file.registers[17][16] ));
 sg13g2_a22oi_1 _17218_ (.Y(_03043_),
    .B1(net5939),
    .B2(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][16] ));
 sg13g2_nand4_1 _17219_ (.B(_03041_),
    .C(_03042_),
    .A(_03040_),
    .Y(_03044_),
    .D(_03043_));
 sg13g2_a22oi_1 _17220_ (.Y(_03045_),
    .B1(net5509),
    .B2(\soc_inst.cpu_core.register_file.registers[18][16] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][16] ));
 sg13g2_a22oi_1 _17221_ (.Y(_03046_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .A2(net5494),
    .A1(\soc_inst.cpu_core.register_file.registers[25][16] ));
 sg13g2_a22oi_1 _17222_ (.Y(_03047_),
    .B1(net5965),
    .B2(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][16] ));
 sg13g2_a22oi_1 _17223_ (.Y(_03048_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .A2(net5489),
    .A1(\soc_inst.cpu_core.register_file.registers[21][16] ));
 sg13g2_nand4_1 _17224_ (.B(_03046_),
    .C(_03047_),
    .A(_03039_),
    .Y(_03049_),
    .D(_03048_));
 sg13g2_a22oi_1 _17225_ (.Y(_03050_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][16] ),
    .A2(net5949),
    .A1(\soc_inst.cpu_core.register_file.registers[15][16] ));
 sg13g2_a22oi_1 _17226_ (.Y(_03051_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][16] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][16] ));
 sg13g2_nand4_1 _17227_ (.B(_03045_),
    .C(_03050_),
    .A(_03038_),
    .Y(_03052_),
    .D(_03051_));
 sg13g2_or2_1 _17228_ (.X(_03053_),
    .B(_03052_),
    .A(_03049_));
 sg13g2_a21oi_1 _17229_ (.A1(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .A2(net5969),
    .Y(_03054_),
    .B1(net6083));
 sg13g2_a22oi_1 _17230_ (.Y(_03055_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .A2(net5913),
    .A1(\soc_inst.cpu_core.register_file.registers[27][16] ));
 sg13g2_a22oi_1 _17231_ (.Y(_03056_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][16] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][16] ));
 sg13g2_a22oi_1 _17232_ (.Y(_03057_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][16] ));
 sg13g2_nand4_1 _17233_ (.B(_03055_),
    .C(_03056_),
    .A(_03054_),
    .Y(_03058_),
    .D(_03057_));
 sg13g2_nor3_2 _17234_ (.A(_03044_),
    .B(_03053_),
    .C(_03058_),
    .Y(_03059_));
 sg13g2_o21ai_1 _17235_ (.B1(net5296),
    .Y(_03060_),
    .A1(net1734),
    .A2(net5921));
 sg13g2_or2_1 _17236_ (.X(_03061_),
    .B(_03060_),
    .A(_03059_));
 sg13g2_o21ai_1 _17237_ (.B1(_03061_),
    .Y(_01012_),
    .A1(net6143),
    .A2(_08080_));
 sg13g2_a22oi_1 _17238_ (.Y(_03062_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][17] ));
 sg13g2_a22oi_1 _17239_ (.Y(_03063_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][17] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][17] ));
 sg13g2_nand2_1 _17240_ (.Y(_03064_),
    .A(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .B(net5901));
 sg13g2_a22oi_1 _17241_ (.Y(_03065_),
    .B1(net5952),
    .B2(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][17] ));
 sg13g2_a22oi_1 _17242_ (.Y(_03066_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .A2(net5492),
    .A1(\soc_inst.cpu_core.register_file.registers[25][17] ));
 sg13g2_a22oi_1 _17243_ (.Y(_03067_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][17] ),
    .A2(net5507),
    .A1(\soc_inst.cpu_core.register_file.registers[18][17] ));
 sg13g2_a22oi_1 _17244_ (.Y(_03068_),
    .B1(net5957),
    .B2(\soc_inst.cpu_core.register_file.registers[26][17] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][17] ));
 sg13g2_a22oi_1 _17245_ (.Y(_03069_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][17] ),
    .A2(net5967),
    .A1(\soc_inst.cpu_core.register_file.registers[6][17] ));
 sg13g2_a22oi_1 _17246_ (.Y(_03070_),
    .B1(net5927),
    .B2(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][17] ));
 sg13g2_a22oi_1 _17247_ (.Y(_03071_),
    .B1(net5962),
    .B2(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][17] ));
 sg13g2_a22oi_1 _17248_ (.Y(_03072_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .A2(net5487),
    .A1(\soc_inst.cpu_core.register_file.registers[21][17] ));
 sg13g2_nand4_1 _17249_ (.B(_03070_),
    .C(_03071_),
    .A(_03066_),
    .Y(_03073_),
    .D(_03072_));
 sg13g2_nand4_1 _17250_ (.B(_03064_),
    .C(_03067_),
    .A(_03063_),
    .Y(_03074_),
    .D(_03068_));
 sg13g2_nor2_1 _17251_ (.A(_03073_),
    .B(_03074_),
    .Y(_03075_));
 sg13g2_a21oi_1 _17252_ (.A1(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .A2(net5891),
    .Y(_03076_),
    .B1(net6081));
 sg13g2_a22oi_1 _17253_ (.Y(_03077_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][17] ),
    .A2(net5932),
    .A1(\soc_inst.cpu_core.register_file.registers[30][17] ));
 sg13g2_a22oi_1 _17254_ (.Y(_03078_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][17] ));
 sg13g2_nand4_1 _17255_ (.B(_03076_),
    .C(_03077_),
    .A(_03065_),
    .Y(_03079_),
    .D(_03078_));
 sg13g2_a22oi_1 _17256_ (.Y(_03080_),
    .B1(net5937),
    .B2(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .A2(net5942),
    .A1(\soc_inst.cpu_core.register_file.registers[22][17] ));
 sg13g2_a22oi_1 _17257_ (.Y(_03081_),
    .B1(net5906),
    .B2(\soc_inst.cpu_core.register_file.registers[24][17] ),
    .A2(net5502),
    .A1(\soc_inst.cpu_core.register_file.registers[17][17] ));
 sg13g2_nand4_1 _17258_ (.B(_03069_),
    .C(_03080_),
    .A(_03062_),
    .Y(_03082_),
    .D(_03081_));
 sg13g2_nor2_1 _17259_ (.A(_03079_),
    .B(_03082_),
    .Y(_03083_));
 sg13g2_o21ai_1 _17260_ (.B1(net5298),
    .Y(_03084_),
    .A1(net1196),
    .A2(net5925));
 sg13g2_a21o_2 _17261_ (.A2(_03083_),
    .A1(_03075_),
    .B1(_03084_),
    .X(_03085_));
 sg13g2_o21ai_1 _17262_ (.B1(_03085_),
    .Y(_01013_),
    .A1(net6146),
    .A2(_08078_));
 sg13g2_nand2_1 _17263_ (.Y(_03086_),
    .A(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .B(net5904));
 sg13g2_a22oi_1 _17264_ (.Y(_03087_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][18] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][18] ));
 sg13g2_a22oi_1 _17265_ (.Y(_03088_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][18] ),
    .A2(net5940),
    .A1(\soc_inst.cpu_core.register_file.registers[3][18] ));
 sg13g2_a22oi_1 _17266_ (.Y(_03089_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][18] ));
 sg13g2_a22oi_1 _17267_ (.Y(_03090_),
    .B1(net5913),
    .B2(\soc_inst.cpu_core.register_file.registers[27][18] ),
    .A2(net5969),
    .A1(\soc_inst.cpu_core.register_file.registers[6][18] ));
 sg13g2_a22oi_1 _17268_ (.Y(_03091_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][18] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][18] ));
 sg13g2_a22oi_1 _17269_ (.Y(_03092_),
    .B1(net5960),
    .B2(\soc_inst.cpu_core.register_file.registers[26][18] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][18] ));
 sg13g2_nand4_1 _17270_ (.B(_03090_),
    .C(_03091_),
    .A(_03089_),
    .Y(_03093_),
    .D(_03092_));
 sg13g2_a22oi_1 _17271_ (.Y(_03094_),
    .B1(net5495),
    .B2(\soc_inst.cpu_core.register_file.registers[25][18] ),
    .A2(net5929),
    .A1(\soc_inst.cpu_core.register_file.registers[4][18] ));
 sg13g2_a22oi_1 _17272_ (.Y(_03095_),
    .B1(net5489),
    .B2(\soc_inst.cpu_core.register_file.registers[21][18] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][18] ));
 sg13g2_a22oi_1 _17273_ (.Y(_03096_),
    .B1(net5965),
    .B2(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][18] ));
 sg13g2_a22oi_1 _17274_ (.Y(_03097_),
    .B1(net5889),
    .B2(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][18] ));
 sg13g2_nand4_1 _17275_ (.B(_03095_),
    .C(_03096_),
    .A(_03088_),
    .Y(_03098_),
    .D(_03097_));
 sg13g2_a22oi_1 _17276_ (.Y(_03099_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][18] ),
    .A2(net5950),
    .A1(\soc_inst.cpu_core.register_file.registers[15][18] ));
 sg13g2_a22oi_1 _17277_ (.Y(_03100_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][18] ),
    .A2(net5918),
    .A1(\soc_inst.cpu_core.register_file.registers[13][18] ));
 sg13g2_nand4_1 _17278_ (.B(_03094_),
    .C(_03099_),
    .A(_03086_),
    .Y(_03101_),
    .D(_03100_));
 sg13g2_or2_1 _17279_ (.X(_03102_),
    .B(_03101_),
    .A(_03098_));
 sg13g2_a21oi_1 _17280_ (.A1(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .A2(net5893),
    .Y(_03103_),
    .B1(net6083));
 sg13g2_a22oi_1 _17281_ (.Y(_03104_),
    .B1(net5510),
    .B2(\soc_inst.cpu_core.register_file.registers[18][18] ),
    .A2(net5515),
    .A1(\soc_inst.cpu_core.register_file.registers[19][18] ));
 sg13g2_a22oi_1 _17282_ (.Y(_03105_),
    .B1(net5504),
    .B2(\soc_inst.cpu_core.register_file.registers[17][18] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][18] ));
 sg13g2_nand4_1 _17283_ (.B(_03103_),
    .C(_03104_),
    .A(_03087_),
    .Y(_03106_),
    .D(_03105_));
 sg13g2_nor3_2 _17284_ (.A(_03093_),
    .B(_03102_),
    .C(_03106_),
    .Y(_03107_));
 sg13g2_o21ai_1 _17285_ (.B1(net5296),
    .Y(_03108_),
    .A1(net1036),
    .A2(net5921));
 sg13g2_or2_1 _17286_ (.X(_03109_),
    .B(_03108_),
    .A(_03107_));
 sg13g2_o21ai_1 _17287_ (.B1(_03109_),
    .Y(_01014_),
    .A1(net6150),
    .A2(_08076_));
 sg13g2_nand2_1 _17288_ (.Y(_03110_),
    .A(\soc_inst.cpu_core.register_file.registers[29][19] ),
    .B(net5484));
 sg13g2_a22oi_1 _17289_ (.Y(_03111_),
    .B1(net5878),
    .B2(\soc_inst.cpu_core.register_file.registers[28][19] ),
    .A2(net5903),
    .A1(\soc_inst.cpu_core.register_file.registers[8][19] ));
 sg13g2_a22oi_1 _17290_ (.Y(_03112_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .A2(net5913),
    .A1(\soc_inst.cpu_core.register_file.registers[27][19] ));
 sg13g2_a22oi_1 _17291_ (.Y(_03113_),
    .B1(net5504),
    .B2(\soc_inst.cpu_core.register_file.registers[17][19] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][19] ));
 sg13g2_a22oi_1 _17292_ (.Y(_03114_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .A2(net5494),
    .A1(\soc_inst.cpu_core.register_file.registers[25][19] ));
 sg13g2_a22oi_1 _17293_ (.Y(_03115_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][19] ),
    .A2(net5954),
    .A1(\soc_inst.cpu_core.register_file.registers[11][19] ));
 sg13g2_a22oi_1 _17294_ (.Y(_03116_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][19] ));
 sg13g2_a22oi_1 _17295_ (.Y(_03117_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][19] ),
    .A2(net5489),
    .A1(\soc_inst.cpu_core.register_file.registers[21][19] ));
 sg13g2_a22oi_1 _17296_ (.Y(_03118_),
    .B1(net5934),
    .B2(\soc_inst.cpu_core.register_file.registers[30][19] ),
    .A2(net5969),
    .A1(\soc_inst.cpu_core.register_file.registers[6][19] ));
 sg13g2_nand4_1 _17297_ (.B(_03116_),
    .C(_03117_),
    .A(_03113_),
    .Y(_03119_),
    .D(_03118_));
 sg13g2_a22oi_1 _17298_ (.Y(_03120_),
    .B1(net5509),
    .B2(\soc_inst.cpu_core.register_file.registers[18][19] ),
    .A2(net5514),
    .A1(\soc_inst.cpu_core.register_file.registers[19][19] ));
 sg13g2_nand4_1 _17299_ (.B(_03114_),
    .C(_03115_),
    .A(_03110_),
    .Y(_03121_),
    .D(_03120_));
 sg13g2_nor2_1 _17300_ (.A(_03119_),
    .B(_03121_),
    .Y(_03122_));
 sg13g2_a21oi_1 _17301_ (.A1(\soc_inst.cpu_core.register_file.registers[23][19] ),
    .A2(net5994),
    .Y(_03123_),
    .B1(net6083));
 sg13g2_a22oi_1 _17302_ (.Y(_03124_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][19] ));
 sg13g2_a22oi_1 _17303_ (.Y(_03125_),
    .B1(net5949),
    .B2(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .A2(net5965),
    .A1(\soc_inst.cpu_core.register_file.registers[14][19] ));
 sg13g2_a22oi_1 _17304_ (.Y(_03126_),
    .B1(net5929),
    .B2(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .A2(net5939),
    .A1(\soc_inst.cpu_core.register_file.registers[3][19] ));
 sg13g2_nand4_1 _17305_ (.B(_03124_),
    .C(_03125_),
    .A(_03123_),
    .Y(_03127_),
    .D(_03126_));
 sg13g2_a22oi_1 _17306_ (.Y(_03128_),
    .B1(net5959),
    .B2(\soc_inst.cpu_core.register_file.registers[26][19] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][19] ));
 sg13g2_a22oi_1 _17307_ (.Y(_03129_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][19] ));
 sg13g2_nand4_1 _17308_ (.B(_03112_),
    .C(_03128_),
    .A(_03111_),
    .Y(_03130_),
    .D(_03129_));
 sg13g2_nor2_1 _17309_ (.A(_03127_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_o21ai_1 _17310_ (.B1(net5298),
    .Y(_03132_),
    .A1(net392),
    .A2(net5925));
 sg13g2_a21o_2 _17311_ (.A2(_03131_),
    .A1(_03122_),
    .B1(_03132_),
    .X(_03133_));
 sg13g2_o21ai_1 _17312_ (.B1(_03133_),
    .Y(_01015_),
    .A1(net6150),
    .A2(_08074_));
 sg13g2_nand2_1 _17313_ (.Y(_03134_),
    .A(\soc_inst.cpu_core.register_file.registers[29][20] ),
    .B(net5485));
 sg13g2_a22oi_1 _17314_ (.Y(_03135_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][20] ),
    .A2(net5945),
    .A1(\soc_inst.cpu_core.register_file.registers[22][20] ));
 sg13g2_a22oi_1 _17315_ (.Y(_03136_),
    .B1(net5889),
    .B2(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .A2(net5505),
    .A1(\soc_inst.cpu_core.register_file.registers[17][20] ));
 sg13g2_a22oi_1 _17316_ (.Y(_03137_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][20] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][20] ));
 sg13g2_a22oi_1 _17317_ (.Y(_03138_),
    .B1(net5894),
    .B2(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .A2(net5495),
    .A1(\soc_inst.cpu_core.register_file.registers[25][20] ));
 sg13g2_a22oi_1 _17318_ (.Y(_03139_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][20] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][20] ));
 sg13g2_a22oi_1 _17319_ (.Y(_03140_),
    .B1(net5960),
    .B2(\soc_inst.cpu_core.register_file.registers[26][20] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][20] ));
 sg13g2_a22oi_1 _17320_ (.Y(_03141_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][20] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][20] ));
 sg13g2_a22oi_1 _17321_ (.Y(_03142_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .A2(net5904),
    .A1(\soc_inst.cpu_core.register_file.registers[8][20] ));
 sg13g2_a22oi_1 _17322_ (.Y(_03143_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][20] ),
    .A2(net5914),
    .A1(\soc_inst.cpu_core.register_file.registers[27][20] ));
 sg13g2_nand4_1 _17323_ (.B(_03141_),
    .C(_03142_),
    .A(_03140_),
    .Y(_03144_),
    .D(_03143_));
 sg13g2_a22oi_1 _17324_ (.Y(_03145_),
    .B1(net5970),
    .B2(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][20] ));
 sg13g2_a22oi_1 _17325_ (.Y(_03146_),
    .B1(net5515),
    .B2(\soc_inst.cpu_core.register_file.registers[19][20] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][20] ));
 sg13g2_a22oi_1 _17326_ (.Y(_03147_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][20] ),
    .A2(net5935),
    .A1(\soc_inst.cpu_core.register_file.registers[30][20] ));
 sg13g2_nand4_1 _17327_ (.B(_03145_),
    .C(_03146_),
    .A(_03137_),
    .Y(_03148_),
    .D(_03147_));
 sg13g2_nand4_1 _17328_ (.B(_03135_),
    .C(_03138_),
    .A(_03134_),
    .Y(_03149_),
    .D(_03139_));
 sg13g2_a21oi_1 _17329_ (.A1(\soc_inst.cpu_core.register_file.registers[18][20] ),
    .A2(net5510),
    .Y(_03150_),
    .B1(net6084));
 sg13g2_a22oi_1 _17330_ (.Y(_03151_),
    .B1(net5950),
    .B2(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][20] ));
 sg13g2_a22oi_1 _17331_ (.Y(_03152_),
    .B1(net5930),
    .B2(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .A2(net5940),
    .A1(\soc_inst.cpu_core.register_file.registers[3][20] ));
 sg13g2_nand4_1 _17332_ (.B(_03150_),
    .C(_03151_),
    .A(_03136_),
    .Y(_03153_),
    .D(_03152_));
 sg13g2_nor4_2 _17333_ (.A(_03144_),
    .B(_03148_),
    .C(_03149_),
    .Y(_03154_),
    .D(_03153_));
 sg13g2_nor2_1 _17334_ (.A(_02675_),
    .B(_03154_),
    .Y(_03155_));
 sg13g2_o21ai_1 _17335_ (.B1(_03155_),
    .Y(_03156_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .A2(net5926));
 sg13g2_o21ai_1 _17336_ (.B1(_03156_),
    .Y(_01016_),
    .A1(net6146),
    .A2(_08073_));
 sg13g2_a22oi_1 _17337_ (.Y(_03157_),
    .B1(net5910),
    .B2(\soc_inst.cpu_core.register_file.registers[24][21] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][21] ));
 sg13g2_nand2_1 _17338_ (.Y(_03158_),
    .A(\soc_inst.cpu_core.register_file.registers[27][21] ),
    .B(net5914));
 sg13g2_a22oi_1 _17339_ (.Y(_03159_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][21] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][21] ));
 sg13g2_a22oi_1 _17340_ (.Y(_03160_),
    .B1(net5904),
    .B2(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .A2(net5981),
    .A1(\soc_inst.cpu_core.register_file.registers[9][21] ));
 sg13g2_a22oi_1 _17341_ (.Y(_03161_),
    .B1(net5940),
    .B2(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .A2(net5991),
    .A1(\soc_inst.cpu_core.register_file.registers[20][21] ));
 sg13g2_a22oi_1 _17342_ (.Y(_03162_),
    .B1(net5495),
    .B2(\soc_inst.cpu_core.register_file.registers[25][21] ),
    .A2(net5936),
    .A1(\soc_inst.cpu_core.register_file.registers[30][21] ));
 sg13g2_a22oi_1 _17343_ (.Y(_03163_),
    .B1(net5895),
    .B2(\soc_inst.cpu_core.register_file.registers[12][21] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][21] ));
 sg13g2_nand4_1 _17344_ (.B(_03161_),
    .C(_03162_),
    .A(_03159_),
    .Y(_03164_),
    .D(_03163_));
 sg13g2_a22oi_1 _17345_ (.Y(_03165_),
    .B1(net5510),
    .B2(\soc_inst.cpu_core.register_file.registers[18][21] ),
    .A2(net5515),
    .A1(\soc_inst.cpu_core.register_file.registers[19][21] ));
 sg13g2_a22oi_1 _17346_ (.Y(_03166_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .A2(net5930),
    .A1(\soc_inst.cpu_core.register_file.registers[4][21] ));
 sg13g2_nand4_1 _17347_ (.B(_03160_),
    .C(_03165_),
    .A(_03158_),
    .Y(_03167_),
    .D(_03166_));
 sg13g2_nor2_1 _17348_ (.A(_03164_),
    .B(_03167_),
    .Y(_03168_));
 sg13g2_a21oi_1 _17349_ (.A1(\soc_inst.cpu_core.register_file.registers[16][21] ),
    .A2(net5501),
    .Y(_03169_),
    .B1(net6084));
 sg13g2_a22oi_1 _17350_ (.Y(_03170_),
    .B1(net5951),
    .B2(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .A2(net5970),
    .A1(\soc_inst.cpu_core.register_file.registers[6][21] ));
 sg13g2_a22oi_1 _17351_ (.Y(_03171_),
    .B1(net5890),
    .B2(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .A2(net5961),
    .A1(\soc_inst.cpu_core.register_file.registers[26][21] ));
 sg13g2_a22oi_1 _17352_ (.Y(_03172_),
    .B1(net5486),
    .B2(\soc_inst.cpu_core.register_file.registers[29][21] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][21] ));
 sg13g2_nand4_1 _17353_ (.B(_03170_),
    .C(_03171_),
    .A(_03169_),
    .Y(_03173_),
    .D(_03172_));
 sg13g2_a22oi_1 _17354_ (.Y(_03174_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .A2(net5946),
    .A1(\soc_inst.cpu_core.register_file.registers[22][21] ));
 sg13g2_a22oi_1 _17355_ (.Y(_03175_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][21] ),
    .A2(net5506),
    .A1(\soc_inst.cpu_core.register_file.registers[17][21] ));
 sg13g2_a22oi_1 _17356_ (.Y(_03176_),
    .B1(net5920),
    .B2(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .A2(net5986),
    .A1(\soc_inst.cpu_core.register_file.registers[2][21] ));
 sg13g2_nand4_1 _17357_ (.B(_03174_),
    .C(_03175_),
    .A(_03157_),
    .Y(_03177_),
    .D(_03176_));
 sg13g2_nor2_1 _17358_ (.A(_03173_),
    .B(_03177_),
    .Y(_03178_));
 sg13g2_o21ai_1 _17359_ (.B1(net5298),
    .Y(_03179_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][21] ),
    .A2(net5925));
 sg13g2_a21oi_2 _17360_ (.B1(_03179_),
    .Y(_03180_),
    .A2(_03178_),
    .A1(_03168_));
 sg13g2_a21o_1 _17361_ (.A2(net3276),
    .A1(net6384),
    .B1(_03180_),
    .X(_01017_));
 sg13g2_a22oi_1 _17362_ (.Y(_03181_),
    .B1(net5492),
    .B2(\soc_inst.cpu_core.register_file.registers[25][22] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][22] ));
 sg13g2_nand2_1 _17363_ (.Y(_03182_),
    .A(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .B(net5901));
 sg13g2_a22oi_1 _17364_ (.Y(_03183_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .A2(net5967),
    .A1(\soc_inst.cpu_core.register_file.registers[6][22] ));
 sg13g2_a22oi_1 _17365_ (.Y(_03184_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][22] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][22] ));
 sg13g2_a22oi_1 _17366_ (.Y(_03185_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][22] ),
    .A2(net5881),
    .A1(\soc_inst.cpu_core.register_file.registers[5][22] ));
 sg13g2_a22oi_1 _17367_ (.Y(_03186_),
    .B1(net5507),
    .B2(\soc_inst.cpu_core.register_file.registers[18][22] ),
    .A2(net5932),
    .A1(\soc_inst.cpu_core.register_file.registers[30][22] ));
 sg13g2_a22oi_1 _17368_ (.Y(_03187_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][22] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][22] ));
 sg13g2_a22oi_1 _17369_ (.Y(_03188_),
    .B1(net5512),
    .B2(\soc_inst.cpu_core.register_file.registers[19][22] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][22] ));
 sg13g2_a22oi_1 _17370_ (.Y(_03189_),
    .B1(net5927),
    .B2(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][22] ));
 sg13g2_a22oi_1 _17371_ (.Y(_03190_),
    .B1(net5962),
    .B2(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][22] ));
 sg13g2_a22oi_1 _17372_ (.Y(_03191_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .A2(net5487),
    .A1(\soc_inst.cpu_core.register_file.registers[21][22] ));
 sg13g2_nand4_1 _17373_ (.B(_03189_),
    .C(_03190_),
    .A(_03185_),
    .Y(_03192_),
    .D(_03191_));
 sg13g2_a22oi_1 _17374_ (.Y(_03193_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][22] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][22] ));
 sg13g2_nand4_1 _17375_ (.B(_03186_),
    .C(_03187_),
    .A(_03182_),
    .Y(_03194_),
    .D(_03193_));
 sg13g2_nor2_1 _17376_ (.A(_03192_),
    .B(_03194_),
    .Y(_03195_));
 sg13g2_a21oi_1 _17377_ (.A1(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .A2(net5891),
    .Y(_03196_),
    .B1(net6081));
 sg13g2_a22oi_1 _17378_ (.Y(_03197_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][22] ));
 sg13g2_nand4_1 _17379_ (.B(_03188_),
    .C(_03196_),
    .A(_03181_),
    .Y(_03198_),
    .D(_03197_));
 sg13g2_a22oi_1 _17380_ (.Y(_03199_),
    .B1(net5906),
    .B2(\soc_inst.cpu_core.register_file.registers[24][22] ),
    .A2(net5502),
    .A1(\soc_inst.cpu_core.register_file.registers[17][22] ));
 sg13g2_a22oi_1 _17381_ (.Y(_03200_),
    .B1(net5942),
    .B2(\soc_inst.cpu_core.register_file.registers[22][22] ),
    .A2(net5957),
    .A1(\soc_inst.cpu_core.register_file.registers[26][22] ));
 sg13g2_nand4_1 _17382_ (.B(_03184_),
    .C(_03199_),
    .A(_03183_),
    .Y(_03201_),
    .D(_03200_));
 sg13g2_nor2_1 _17383_ (.A(_03198_),
    .B(_03201_),
    .Y(_03202_));
 sg13g2_o21ai_1 _17384_ (.B1(net5296),
    .Y(_03203_),
    .A1(net635),
    .A2(net5921));
 sg13g2_a21o_2 _17385_ (.A2(_03202_),
    .A1(_03195_),
    .B1(_03203_),
    .X(_03204_));
 sg13g2_o21ai_1 _17386_ (.B1(_03204_),
    .Y(_01018_),
    .A1(net6146),
    .A2(_08070_));
 sg13g2_a22oi_1 _17387_ (.Y(_03205_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][23] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][23] ));
 sg13g2_a22oi_1 _17388_ (.Y(_03206_),
    .B1(net5495),
    .B2(\soc_inst.cpu_core.register_file.registers[25][23] ),
    .A2(net5930),
    .A1(\soc_inst.cpu_core.register_file.registers[4][23] ));
 sg13g2_nand2_1 _17389_ (.Y(_03207_),
    .A(\soc_inst.cpu_core.register_file.registers[26][23] ),
    .B(net5960));
 sg13g2_a22oi_1 _17390_ (.Y(_03208_),
    .B1(net5485),
    .B2(\soc_inst.cpu_core.register_file.registers[29][23] ),
    .A2(net5889),
    .A1(\soc_inst.cpu_core.register_file.registers[10][23] ));
 sg13g2_a22oi_1 _17391_ (.Y(_03209_),
    .B1(net5505),
    .B2(\soc_inst.cpu_core.register_file.registers[17][23] ),
    .A2(net5510),
    .A1(\soc_inst.cpu_core.register_file.registers[18][23] ));
 sg13g2_a22oi_1 _17392_ (.Y(_03210_),
    .B1(net5894),
    .B2(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][23] ));
 sg13g2_a22oi_1 _17393_ (.Y(_03211_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .A2(net5940),
    .A1(\soc_inst.cpu_core.register_file.registers[3][23] ));
 sg13g2_a22oi_1 _17394_ (.Y(_03212_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .A2(net5904),
    .A1(\soc_inst.cpu_core.register_file.registers[8][23] ));
 sg13g2_nand4_1 _17395_ (.B(_03209_),
    .C(_03211_),
    .A(_03206_),
    .Y(_03213_),
    .D(_03212_));
 sg13g2_a22oi_1 _17396_ (.Y(_03214_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][23] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][23] ));
 sg13g2_a22oi_1 _17397_ (.Y(_03215_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][23] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][23] ));
 sg13g2_nand4_1 _17398_ (.B(_03210_),
    .C(_03214_),
    .A(_03207_),
    .Y(_03216_),
    .D(_03215_));
 sg13g2_a21oi_1 _17399_ (.A1(\soc_inst.cpu_core.register_file.registers[30][23] ),
    .A2(net5935),
    .Y(_03217_),
    .B1(net6084));
 sg13g2_a22oi_1 _17400_ (.Y(_03218_),
    .B1(net5970),
    .B2(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][23] ));
 sg13g2_a22oi_1 _17401_ (.Y(_03219_),
    .B1(net5884),
    .B2(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .A2(net5914),
    .A1(\soc_inst.cpu_core.register_file.registers[27][23] ));
 sg13g2_nand4_1 _17402_ (.B(_03217_),
    .C(_03218_),
    .A(_03208_),
    .Y(_03220_),
    .D(_03219_));
 sg13g2_a22oi_1 _17403_ (.Y(_03221_),
    .B1(net5515),
    .B2(\soc_inst.cpu_core.register_file.registers[19][23] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][23] ));
 sg13g2_a22oi_1 _17404_ (.Y(_03222_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][23] ),
    .A2(net5945),
    .A1(\soc_inst.cpu_core.register_file.registers[22][23] ));
 sg13g2_a22oi_1 _17405_ (.Y(_03223_),
    .B1(net5950),
    .B2(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][23] ));
 sg13g2_nand4_1 _17406_ (.B(_03221_),
    .C(_03222_),
    .A(_03205_),
    .Y(_03224_),
    .D(_03223_));
 sg13g2_or2_1 _17407_ (.X(_03225_),
    .B(_03224_),
    .A(_03220_));
 sg13g2_nor3_2 _17408_ (.A(_03213_),
    .B(_03216_),
    .C(_03225_),
    .Y(_03226_));
 sg13g2_o21ai_1 _17409_ (.B1(net5298),
    .Y(_03227_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][23] ),
    .A2(net5925));
 sg13g2_or2_1 _17410_ (.X(_03228_),
    .B(_03227_),
    .A(_03226_));
 sg13g2_o21ai_1 _17411_ (.B1(_03228_),
    .Y(_01019_),
    .A1(net6143),
    .A2(_08068_));
 sg13g2_a22oi_1 _17412_ (.Y(_03229_),
    .B1(net5967),
    .B2(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][24] ));
 sg13g2_nand2_1 _17413_ (.Y(_03230_),
    .A(\soc_inst.cpu_core.register_file.registers[28][24] ),
    .B(net5876));
 sg13g2_a22oi_1 _17414_ (.Y(_03231_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][24] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][24] ));
 sg13g2_a22oi_1 _17415_ (.Y(_03232_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][24] ));
 sg13g2_a22oi_1 _17416_ (.Y(_03233_),
    .B1(net5901),
    .B2(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .A2(net5487),
    .A1(\soc_inst.cpu_core.register_file.registers[21][24] ));
 sg13g2_a22oi_1 _17417_ (.Y(_03234_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .A2(net5911),
    .A1(\soc_inst.cpu_core.register_file.registers[27][24] ));
 sg13g2_a22oi_1 _17418_ (.Y(_03235_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][24] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][24] ));
 sg13g2_a22oi_1 _17419_ (.Y(_03236_),
    .B1(net5927),
    .B2(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][24] ));
 sg13g2_a22oi_1 _17420_ (.Y(_03237_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][24] ));
 sg13g2_nand4_1 _17421_ (.B(_03235_),
    .C(_03236_),
    .A(_03232_),
    .Y(_03238_),
    .D(_03237_));
 sg13g2_nand4_1 _17422_ (.B(_03230_),
    .C(_03233_),
    .A(_03229_),
    .Y(_03239_),
    .D(_03234_));
 sg13g2_nor2_1 _17423_ (.A(_03238_),
    .B(_03239_),
    .Y(_03240_));
 sg13g2_a21oi_1 _17424_ (.A1(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .A2(net5891),
    .Y(_03241_),
    .B1(net6081));
 sg13g2_a22oi_1 _17425_ (.Y(_03242_),
    .B1(net5492),
    .B2(\soc_inst.cpu_core.register_file.registers[25][24] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][24] ));
 sg13g2_a22oi_1 _17426_ (.Y(_03243_),
    .B1(net5942),
    .B2(\soc_inst.cpu_core.register_file.registers[22][24] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][24] ));
 sg13g2_nand4_1 _17427_ (.B(_03241_),
    .C(_03242_),
    .A(_03231_),
    .Y(_03244_),
    .D(_03243_));
 sg13g2_a22oi_1 _17428_ (.Y(_03245_),
    .B1(net5507),
    .B2(\soc_inst.cpu_core.register_file.registers[18][24] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][24] ));
 sg13g2_a22oi_1 _17429_ (.Y(_03246_),
    .B1(net5932),
    .B2(\soc_inst.cpu_core.register_file.registers[30][24] ),
    .A2(net5957),
    .A1(\soc_inst.cpu_core.register_file.registers[26][24] ));
 sg13g2_a22oi_1 _17430_ (.Y(_03247_),
    .B1(net5502),
    .B2(\soc_inst.cpu_core.register_file.registers[17][24] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][24] ));
 sg13g2_a22oi_1 _17431_ (.Y(_03248_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .A2(net5906),
    .A1(\soc_inst.cpu_core.register_file.registers[24][24] ));
 sg13g2_nand4_1 _17432_ (.B(_03246_),
    .C(_03247_),
    .A(_03245_),
    .Y(_03249_),
    .D(_03248_));
 sg13g2_nor2_1 _17433_ (.A(_03244_),
    .B(_03249_),
    .Y(_03250_));
 sg13g2_o21ai_1 _17434_ (.B1(net5298),
    .Y(_03251_),
    .A1(net1304),
    .A2(net5925));
 sg13g2_a21o_2 _17435_ (.A2(_03250_),
    .A1(_03240_),
    .B1(_03251_),
    .X(_03252_));
 sg13g2_o21ai_1 _17436_ (.B1(_03252_),
    .Y(_01020_),
    .A1(net6146),
    .A2(_08066_));
 sg13g2_nand2_1 _17437_ (.Y(_03253_),
    .A(\soc_inst.cpu_core.register_file.registers[21][25] ),
    .B(net5487));
 sg13g2_a22oi_1 _17438_ (.Y(_03254_),
    .B1(net5502),
    .B2(\soc_inst.cpu_core.register_file.registers[17][25] ),
    .A2(net5942),
    .A1(\soc_inst.cpu_core.register_file.registers[22][25] ));
 sg13g2_a22oi_1 _17439_ (.Y(_03255_),
    .B1(net5932),
    .B2(\soc_inst.cpu_core.register_file.registers[30][25] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][25] ));
 sg13g2_a22oi_1 _17440_ (.Y(_03256_),
    .B1(net5947),
    .B2(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][25] ));
 sg13g2_a22oi_1 _17441_ (.Y(_03257_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][25] ),
    .A2(net5901),
    .A1(\soc_inst.cpu_core.register_file.registers[8][25] ));
 sg13g2_a22oi_1 _17442_ (.Y(_03258_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .A2(net5906),
    .A1(\soc_inst.cpu_core.register_file.registers[24][25] ));
 sg13g2_a22oi_1 _17443_ (.Y(_03259_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][25] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][25] ));
 sg13g2_a22oi_1 _17444_ (.Y(_03260_),
    .B1(net5507),
    .B2(\soc_inst.cpu_core.register_file.registers[18][25] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][25] ));
 sg13g2_a22oi_1 _17445_ (.Y(_03261_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][25] ));
 sg13g2_a22oi_1 _17446_ (.Y(_03262_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .A2(net5927),
    .A1(\soc_inst.cpu_core.register_file.registers[4][25] ));
 sg13g2_nand4_1 _17447_ (.B(_03260_),
    .C(_03261_),
    .A(_03256_),
    .Y(_03263_),
    .D(_03262_));
 sg13g2_a22oi_1 _17448_ (.Y(_03264_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][25] ));
 sg13g2_nand4_1 _17449_ (.B(_03257_),
    .C(_03258_),
    .A(_03253_),
    .Y(_03265_),
    .D(_03264_));
 sg13g2_nor2_1 _17450_ (.A(_03263_),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_a21oi_1 _17451_ (.A1(\soc_inst.cpu_core.register_file.registers[28][25] ),
    .A2(net5876),
    .Y(_03267_),
    .B1(net6081));
 sg13g2_a22oi_1 _17452_ (.Y(_03268_),
    .B1(net5957),
    .B2(\soc_inst.cpu_core.register_file.registers[26][25] ),
    .A2(net5967),
    .A1(\soc_inst.cpu_core.register_file.registers[6][25] ));
 sg13g2_a22oi_1 _17453_ (.Y(_03269_),
    .B1(net5977),
    .B2(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][25] ));
 sg13g2_nand4_1 _17454_ (.B(_03267_),
    .C(_03268_),
    .A(_03259_),
    .Y(_03270_),
    .D(_03269_));
 sg13g2_a22oi_1 _17455_ (.Y(_03271_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][25] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][25] ));
 sg13g2_a22oi_1 _17456_ (.Y(_03272_),
    .B1(net5891),
    .B2(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .A2(net5492),
    .A1(\soc_inst.cpu_core.register_file.registers[25][25] ));
 sg13g2_nand4_1 _17457_ (.B(_03255_),
    .C(_03271_),
    .A(_03254_),
    .Y(_03273_),
    .D(_03272_));
 sg13g2_nor2_1 _17458_ (.A(_03270_),
    .B(_03273_),
    .Y(_03274_));
 sg13g2_o21ai_1 _17459_ (.B1(net5296),
    .Y(_03275_),
    .A1(net1097),
    .A2(net5921));
 sg13g2_a21o_2 _17460_ (.A2(_03274_),
    .A1(_03266_),
    .B1(_03275_),
    .X(_03276_));
 sg13g2_o21ai_1 _17461_ (.B1(_03276_),
    .Y(_01021_),
    .A1(net6150),
    .A2(_08065_));
 sg13g2_a22oi_1 _17462_ (.Y(_03277_),
    .B1(net5898),
    .B2(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .A2(net5969),
    .A1(\soc_inst.cpu_core.register_file.registers[6][26] ));
 sg13g2_a22oi_1 _17463_ (.Y(_03278_),
    .B1(net5913),
    .B2(\soc_inst.cpu_core.register_file.registers[27][26] ),
    .A2(net5489),
    .A1(\soc_inst.cpu_core.register_file.registers[21][26] ));
 sg13g2_nand2_1 _17464_ (.Y(_03279_),
    .A(\soc_inst.cpu_core.register_file.registers[19][26] ),
    .B(net5514));
 sg13g2_a22oi_1 _17465_ (.Y(_03280_),
    .B1(net5908),
    .B2(\soc_inst.cpu_core.register_file.registers[24][26] ),
    .A2(net5934),
    .A1(\soc_inst.cpu_core.register_file.registers[30][26] ));
 sg13g2_a22oi_1 _17466_ (.Y(_03281_),
    .B1(net5949),
    .B2(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .A2(net5965),
    .A1(\soc_inst.cpu_core.register_file.registers[14][26] ));
 sg13g2_a22oi_1 _17467_ (.Y(_03282_),
    .B1(net5499),
    .B2(\soc_inst.cpu_core.register_file.registers[16][26] ),
    .A2(net5509),
    .A1(\soc_inst.cpu_core.register_file.registers[18][26] ));
 sg13g2_a22oi_1 _17468_ (.Y(_03283_),
    .B1(net5888),
    .B2(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .A2(net5959),
    .A1(\soc_inst.cpu_core.register_file.registers[26][26] ));
 sg13g2_a22oi_1 _17469_ (.Y(_03284_),
    .B1(net5883),
    .B2(\soc_inst.cpu_core.register_file.registers[5][26] ),
    .A2(net5979),
    .A1(\soc_inst.cpu_core.register_file.registers[9][26] ));
 sg13g2_nand4_1 _17470_ (.B(_03282_),
    .C(_03283_),
    .A(_03281_),
    .Y(_03285_),
    .D(_03284_));
 sg13g2_a22oi_1 _17471_ (.Y(_03286_),
    .B1(net5893),
    .B2(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .A2(net5903),
    .A1(\soc_inst.cpu_core.register_file.registers[8][26] ));
 sg13g2_a22oi_1 _17472_ (.Y(_03287_),
    .B1(net5504),
    .B2(\soc_inst.cpu_core.register_file.registers[17][26] ),
    .A2(net5944),
    .A1(\soc_inst.cpu_core.register_file.registers[22][26] ));
 sg13g2_a22oi_1 _17473_ (.Y(_03288_),
    .B1(net5484),
    .B2(\soc_inst.cpu_core.register_file.registers[29][26] ),
    .A2(net5989),
    .A1(\soc_inst.cpu_core.register_file.registers[20][26] ));
 sg13g2_a22oi_1 _17474_ (.Y(_03289_),
    .B1(net5918),
    .B2(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .A2(net5929),
    .A1(\soc_inst.cpu_core.register_file.registers[4][26] ));
 sg13g2_nand4_1 _17475_ (.B(_03287_),
    .C(_03288_),
    .A(_03280_),
    .Y(_03290_),
    .D(_03289_));
 sg13g2_a22oi_1 _17476_ (.Y(_03291_),
    .B1(net5939),
    .B2(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .A2(net5984),
    .A1(\soc_inst.cpu_core.register_file.registers[2][26] ));
 sg13g2_a22oi_1 _17477_ (.Y(_03292_),
    .B1(net5954),
    .B2(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .A2(net5994),
    .A1(\soc_inst.cpu_core.register_file.registers[23][26] ));
 sg13g2_nand4_1 _17478_ (.B(_03286_),
    .C(_03291_),
    .A(_03279_),
    .Y(_03293_),
    .D(_03292_));
 sg13g2_or2_1 _17479_ (.X(_03294_),
    .B(_03293_),
    .A(_03290_));
 sg13g2_a21oi_1 _17480_ (.A1(\soc_inst.cpu_core.register_file.registers[28][26] ),
    .A2(net5878),
    .Y(_03295_),
    .B1(net6083));
 sg13g2_a22oi_1 _17481_ (.Y(_03296_),
    .B1(net5494),
    .B2(\soc_inst.cpu_core.register_file.registers[25][26] ),
    .A2(net5974),
    .A1(\soc_inst.cpu_core.register_file.registers[31][26] ));
 sg13g2_nand4_1 _17482_ (.B(_03278_),
    .C(_03295_),
    .A(_03277_),
    .Y(_03297_),
    .D(_03296_));
 sg13g2_nor3_1 _17483_ (.A(_03285_),
    .B(_03294_),
    .C(_03297_),
    .Y(_03298_));
 sg13g2_o21ai_1 _17484_ (.B1(net5298),
    .Y(_03299_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][26] ),
    .A2(net5925));
 sg13g2_or2_1 _17485_ (.X(_03300_),
    .B(_03299_),
    .A(_03298_));
 sg13g2_o21ai_1 _17486_ (.B1(_03300_),
    .Y(_01022_),
    .A1(net6150),
    .A2(_08063_));
 sg13g2_a22oi_1 _17487_ (.Y(_03301_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][27] ));
 sg13g2_a22oi_1 _17488_ (.Y(_03302_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][27] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][27] ));
 sg13g2_a21oi_1 _17489_ (.A1(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .A2(net5891),
    .Y(_03303_),
    .B1(net6081));
 sg13g2_nand2_1 _17490_ (.Y(_03304_),
    .A(\soc_inst.cpu_core.register_file.registers[25][27] ),
    .B(net5492));
 sg13g2_a22oi_1 _17491_ (.Y(_03305_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][27] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][27] ));
 sg13g2_a22oi_1 _17492_ (.Y(_03306_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][27] ),
    .A2(net5507),
    .A1(\soc_inst.cpu_core.register_file.registers[18][27] ));
 sg13g2_a22oi_1 _17493_ (.Y(_03307_),
    .B1(net5512),
    .B2(\soc_inst.cpu_core.register_file.registers[19][27] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][27] ));
 sg13g2_a22oi_1 _17494_ (.Y(_03308_),
    .B1(net5502),
    .B2(\soc_inst.cpu_core.register_file.registers[17][27] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][27] ));
 sg13g2_a22oi_1 _17495_ (.Y(_03309_),
    .B1(net5967),
    .B2(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][27] ));
 sg13g2_a22oi_1 _17496_ (.Y(_03310_),
    .B1(net5906),
    .B2(\soc_inst.cpu_core.register_file.registers[24][27] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][27] ));
 sg13g2_a22oi_1 _17497_ (.Y(_03311_),
    .B1(net5927),
    .B2(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .A2(net5937),
    .A1(\soc_inst.cpu_core.register_file.registers[3][27] ));
 sg13g2_a22oi_1 _17498_ (.Y(_03312_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][27] ),
    .A2(net5886),
    .A1(\soc_inst.cpu_core.register_file.registers[10][27] ));
 sg13g2_nand4_1 _17499_ (.B(_03310_),
    .C(_03311_),
    .A(_03301_),
    .Y(_03313_),
    .D(_03312_));
 sg13g2_nand4_1 _17500_ (.B(_03304_),
    .C(_03306_),
    .A(_03302_),
    .Y(_03314_),
    .D(_03307_));
 sg13g2_nor2_1 _17501_ (.A(_03313_),
    .B(_03314_),
    .Y(_03315_));
 sg13g2_a22oi_1 _17502_ (.Y(_03316_),
    .B1(net5487),
    .B2(\soc_inst.cpu_core.register_file.registers[21][27] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][27] ));
 sg13g2_a22oi_1 _17503_ (.Y(_03317_),
    .B1(net5932),
    .B2(\soc_inst.cpu_core.register_file.registers[30][27] ),
    .A2(net5957),
    .A1(\soc_inst.cpu_core.register_file.registers[26][27] ));
 sg13g2_nand4_1 _17504_ (.B(_03305_),
    .C(_03316_),
    .A(_03303_),
    .Y(_03318_),
    .D(_03317_));
 sg13g2_a22oi_1 _17505_ (.Y(_03319_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .A2(net5901),
    .A1(\soc_inst.cpu_core.register_file.registers[8][27] ));
 sg13g2_a22oi_1 _17506_ (.Y(_03320_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][27] ),
    .A2(net5942),
    .A1(\soc_inst.cpu_core.register_file.registers[22][27] ));
 sg13g2_nand4_1 _17507_ (.B(_03309_),
    .C(_03319_),
    .A(_03308_),
    .Y(_03321_),
    .D(_03320_));
 sg13g2_nor2_1 _17508_ (.A(_03318_),
    .B(_03321_),
    .Y(_03322_));
 sg13g2_o21ai_1 _17509_ (.B1(net5297),
    .Y(_03323_),
    .A1(net829),
    .A2(net5922));
 sg13g2_a21o_2 _17510_ (.A2(_03322_),
    .A1(_03315_),
    .B1(_03323_),
    .X(_03324_));
 sg13g2_o21ai_1 _17511_ (.B1(_03324_),
    .Y(_01023_),
    .A1(net6146),
    .A2(_08061_));
 sg13g2_nand2_1 _17512_ (.Y(_03325_),
    .A(\soc_inst.cpu_core.register_file.registers[17][28] ),
    .B(net5502));
 sg13g2_a22oi_1 _17513_ (.Y(_03326_),
    .B1(net5937),
    .B2(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .A2(net5962),
    .A1(\soc_inst.cpu_core.register_file.registers[14][28] ));
 sg13g2_a22oi_1 _17514_ (.Y(_03327_),
    .B1(net5901),
    .B2(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .A2(net5972),
    .A1(\soc_inst.cpu_core.register_file.registers[31][28] ));
 sg13g2_a22oi_1 _17515_ (.Y(_03328_),
    .B1(net5896),
    .B2(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .A2(net5487),
    .A1(\soc_inst.cpu_core.register_file.registers[21][28] ));
 sg13g2_a22oi_1 _17516_ (.Y(_03329_),
    .B1(net5497),
    .B2(\soc_inst.cpu_core.register_file.registers[16][28] ),
    .A2(net5952),
    .A1(\soc_inst.cpu_core.register_file.registers[11][28] ));
 sg13g2_a22oi_1 _17517_ (.Y(_03330_),
    .B1(net5911),
    .B2(\soc_inst.cpu_core.register_file.registers[27][28] ),
    .A2(net5947),
    .A1(\soc_inst.cpu_core.register_file.registers[15][28] ));
 sg13g2_a22oi_1 _17518_ (.Y(_03331_),
    .B1(net5916),
    .B2(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .A2(net5927),
    .A1(\soc_inst.cpu_core.register_file.registers[4][28] ));
 sg13g2_a22oi_1 _17519_ (.Y(_03332_),
    .B1(net5886),
    .B2(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .A2(net5492),
    .A1(\soc_inst.cpu_core.register_file.registers[25][28] ));
 sg13g2_nand4_1 _17520_ (.B(_03330_),
    .C(_03331_),
    .A(_03326_),
    .Y(_03333_),
    .D(_03332_));
 sg13g2_a22oi_1 _17521_ (.Y(_03334_),
    .B1(net5881),
    .B2(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .A2(net5982),
    .A1(\soc_inst.cpu_core.register_file.registers[2][28] ));
 sg13g2_nand4_1 _17522_ (.B(_03327_),
    .C(_03328_),
    .A(_03325_),
    .Y(_03335_),
    .D(_03334_));
 sg13g2_nor2_1 _17523_ (.A(_03333_),
    .B(_03335_),
    .Y(_03336_));
 sg13g2_a21oi_1 _17524_ (.A1(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .A2(net5891),
    .Y(_03337_),
    .B1(net6081));
 sg13g2_a22oi_1 _17525_ (.Y(_03338_),
    .B1(net5942),
    .B2(\soc_inst.cpu_core.register_file.registers[22][28] ),
    .A2(net5512),
    .A1(\soc_inst.cpu_core.register_file.registers[19][28] ));
 sg13g2_a22oi_1 _17526_ (.Y(_03339_),
    .B1(net5482),
    .B2(\soc_inst.cpu_core.register_file.registers[29][28] ),
    .A2(net5906),
    .A1(\soc_inst.cpu_core.register_file.registers[24][28] ));
 sg13g2_nand4_1 _17527_ (.B(_03337_),
    .C(_03338_),
    .A(_03329_),
    .Y(_03340_),
    .D(_03339_));
 sg13g2_a22oi_1 _17528_ (.Y(_03341_),
    .B1(net5932),
    .B2(\soc_inst.cpu_core.register_file.registers[30][28] ),
    .A2(net5987),
    .A1(\soc_inst.cpu_core.register_file.registers[20][28] ));
 sg13g2_a22oi_1 _17529_ (.Y(_03342_),
    .B1(net5507),
    .B2(\soc_inst.cpu_core.register_file.registers[18][28] ),
    .A2(net5992),
    .A1(\soc_inst.cpu_core.register_file.registers[23][28] ));
 sg13g2_a22oi_1 _17530_ (.Y(_03343_),
    .B1(net5876),
    .B2(\soc_inst.cpu_core.register_file.registers[28][28] ),
    .A2(net5967),
    .A1(\soc_inst.cpu_core.register_file.registers[6][28] ));
 sg13g2_a22oi_1 _17531_ (.Y(_03344_),
    .B1(net5957),
    .B2(\soc_inst.cpu_core.register_file.registers[26][28] ),
    .A2(net5977),
    .A1(\soc_inst.cpu_core.register_file.registers[9][28] ));
 sg13g2_nand4_1 _17532_ (.B(_03342_),
    .C(_03343_),
    .A(_03341_),
    .Y(_03345_),
    .D(_03344_));
 sg13g2_nor2_1 _17533_ (.A(_03340_),
    .B(_03345_),
    .Y(_03346_));
 sg13g2_o21ai_1 _17534_ (.B1(net5298),
    .Y(_03347_),
    .A1(net484),
    .A2(net5925));
 sg13g2_a21o_2 _17535_ (.A2(_03346_),
    .A1(_03336_),
    .B1(_03347_),
    .X(_03348_));
 sg13g2_o21ai_1 _17536_ (.B1(_03348_),
    .Y(_01024_),
    .A1(net6146),
    .A2(_08060_));
 sg13g2_nand2_1 _17537_ (.Y(_03349_),
    .A(\soc_inst.cpu_core.register_file.registers[27][29] ),
    .B(net5912));
 sg13g2_a22oi_1 _17538_ (.Y(_03350_),
    .B1(net5917),
    .B2(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .A2(net5498),
    .A1(\soc_inst.cpu_core.register_file.registers[16][29] ));
 sg13g2_a22oi_1 _17539_ (.Y(_03351_),
    .B1(net5897),
    .B2(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .A2(net5928),
    .A1(\soc_inst.cpu_core.register_file.registers[4][29] ));
 sg13g2_a22oi_1 _17540_ (.Y(_03352_),
    .B1(net5907),
    .B2(\soc_inst.cpu_core.register_file.registers[24][29] ),
    .A2(net5513),
    .A1(\soc_inst.cpu_core.register_file.registers[19][29] ));
 sg13g2_a22oi_1 _17541_ (.Y(_03353_),
    .B1(net5948),
    .B2(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .A2(net5968),
    .A1(\soc_inst.cpu_core.register_file.registers[6][29] ));
 sg13g2_a22oi_1 _17542_ (.Y(_03354_),
    .B1(net5983),
    .B2(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .A2(net5988),
    .A1(\soc_inst.cpu_core.register_file.registers[20][29] ));
 sg13g2_a22oi_1 _17543_ (.Y(_03355_),
    .B1(net5933),
    .B2(\soc_inst.cpu_core.register_file.registers[30][29] ),
    .A2(net5938),
    .A1(\soc_inst.cpu_core.register_file.registers[3][29] ));
 sg13g2_nand4_1 _17544_ (.B(_03353_),
    .C(_03354_),
    .A(_03350_),
    .Y(_03356_),
    .D(_03355_));
 sg13g2_a22oi_1 _17545_ (.Y(_03357_),
    .B1(net5483),
    .B2(\soc_inst.cpu_core.register_file.registers[29][29] ),
    .A2(net5973),
    .A1(\soc_inst.cpu_core.register_file.registers[31][29] ));
 sg13g2_a22oi_1 _17546_ (.Y(_03358_),
    .B1(net5493),
    .B2(\soc_inst.cpu_core.register_file.registers[25][29] ),
    .A2(net5508),
    .A1(\soc_inst.cpu_core.register_file.registers[18][29] ));
 sg13g2_nand4_1 _17547_ (.B(_03352_),
    .C(_03357_),
    .A(_03349_),
    .Y(_03359_),
    .D(_03358_));
 sg13g2_nor2_1 _17548_ (.A(_03356_),
    .B(_03359_),
    .Y(_03360_));
 sg13g2_a21oi_1 _17549_ (.A1(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .A2(net5902),
    .Y(_03361_),
    .B1(net6082));
 sg13g2_a22oi_1 _17550_ (.Y(_03362_),
    .B1(net5877),
    .B2(\soc_inst.cpu_core.register_file.registers[28][29] ),
    .A2(net5958),
    .A1(\soc_inst.cpu_core.register_file.registers[26][29] ));
 sg13g2_a22oi_1 _17551_ (.Y(_03363_),
    .B1(net5488),
    .B2(\soc_inst.cpu_core.register_file.registers[21][29] ),
    .A2(net5993),
    .A1(\soc_inst.cpu_core.register_file.registers[23][29] ));
 sg13g2_nand4_1 _17552_ (.B(_03361_),
    .C(_03362_),
    .A(_03351_),
    .Y(_03364_),
    .D(_03363_));
 sg13g2_a22oi_1 _17553_ (.Y(_03365_),
    .B1(net5887),
    .B2(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .A2(net5953),
    .A1(\soc_inst.cpu_core.register_file.registers[11][29] ));
 sg13g2_a22oi_1 _17554_ (.Y(_03366_),
    .B1(net5892),
    .B2(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .A2(net5943),
    .A1(\soc_inst.cpu_core.register_file.registers[22][29] ));
 sg13g2_a22oi_1 _17555_ (.Y(_03367_),
    .B1(net5963),
    .B2(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .A2(net5978),
    .A1(\soc_inst.cpu_core.register_file.registers[9][29] ));
 sg13g2_a22oi_1 _17556_ (.Y(_03368_),
    .B1(net5882),
    .B2(\soc_inst.cpu_core.register_file.registers[5][29] ),
    .A2(net5503),
    .A1(\soc_inst.cpu_core.register_file.registers[17][29] ));
 sg13g2_nand4_1 _17557_ (.B(_03366_),
    .C(_03367_),
    .A(_03365_),
    .Y(_03369_),
    .D(_03368_));
 sg13g2_nor2_1 _17558_ (.A(_03364_),
    .B(_03369_),
    .Y(_03370_));
 sg13g2_o21ai_1 _17559_ (.B1(net5297),
    .Y(_03371_),
    .A1(net741),
    .A2(net5923));
 sg13g2_a21oi_2 _17560_ (.B1(_03371_),
    .Y(_03372_),
    .A2(_03370_),
    .A1(_03360_));
 sg13g2_a21o_1 _17561_ (.A2(net3163),
    .A1(net6400),
    .B1(_03372_),
    .X(_01025_));
 sg13g2_nand2_1 _17562_ (.Y(_03373_),
    .A(\soc_inst.cpu_core.register_file.registers[17][30] ),
    .B(net5505));
 sg13g2_a22oi_1 _17563_ (.Y(_03374_),
    .B1(net5495),
    .B2(\soc_inst.cpu_core.register_file.registers[25][30] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][30] ));
 sg13g2_a22oi_1 _17564_ (.Y(_03375_),
    .B1(net5894),
    .B2(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .A2(net5900),
    .A1(\soc_inst.cpu_core.register_file.registers[7][30] ));
 sg13g2_a22oi_1 _17565_ (.Y(_03376_),
    .B1(net5515),
    .B2(\soc_inst.cpu_core.register_file.registers[19][30] ),
    .A2(net5970),
    .A1(\soc_inst.cpu_core.register_file.registers[6][30] ));
 sg13g2_a22oi_1 _17566_ (.Y(_03377_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][30] ),
    .A2(net5945),
    .A1(\soc_inst.cpu_core.register_file.registers[22][30] ));
 sg13g2_a22oi_1 _17567_ (.Y(_03378_),
    .B1(net5904),
    .B2(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .A2(net5950),
    .A1(\soc_inst.cpu_core.register_file.registers[15][30] ));
 sg13g2_a22oi_1 _17568_ (.Y(_03379_),
    .B1(net5510),
    .B2(\soc_inst.cpu_core.register_file.registers[18][30] ),
    .A2(net5995),
    .A1(\soc_inst.cpu_core.register_file.registers[23][30] ));
 sg13g2_a22oi_1 _17569_ (.Y(_03380_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .A2(net5960),
    .A1(\soc_inst.cpu_core.register_file.registers[26][30] ));
 sg13g2_a22oi_1 _17570_ (.Y(_03381_),
    .B1(net5485),
    .B2(\soc_inst.cpu_core.register_file.registers[29][30] ),
    .A2(net5940),
    .A1(\soc_inst.cpu_core.register_file.registers[3][30] ));
 sg13g2_nand4_1 _17571_ (.B(_03379_),
    .C(_03380_),
    .A(_03374_),
    .Y(_03382_),
    .D(_03381_));
 sg13g2_a22oi_1 _17572_ (.Y(_03383_),
    .B1(net5930),
    .B2(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][30] ));
 sg13g2_a22oi_1 _17573_ (.Y(_03384_),
    .B1(net5490),
    .B2(\soc_inst.cpu_core.register_file.registers[21][30] ),
    .A2(net5955),
    .A1(\soc_inst.cpu_core.register_file.registers[11][30] ));
 sg13g2_nand4_1 _17574_ (.B(_03375_),
    .C(_03383_),
    .A(_03373_),
    .Y(_03385_),
    .D(_03384_));
 sg13g2_or2_1 _17575_ (.X(_03386_),
    .B(_03385_),
    .A(_03382_));
 sg13g2_a21oi_1 _17576_ (.A1(\soc_inst.cpu_core.register_file.registers[16][30] ),
    .A2(net5500),
    .Y(_03387_),
    .B1(net6085));
 sg13g2_a22oi_1 _17577_ (.Y(_03388_),
    .B1(net5889),
    .B2(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .A2(net5966),
    .A1(\soc_inst.cpu_core.register_file.registers[14][30] ));
 sg13g2_a22oi_1 _17578_ (.Y(_03389_),
    .B1(net5880),
    .B2(\soc_inst.cpu_core.register_file.registers[28][30] ),
    .A2(net5884),
    .A1(\soc_inst.cpu_core.register_file.registers[5][30] ));
 sg13g2_nand4_1 _17579_ (.B(_03387_),
    .C(_03388_),
    .A(_03378_),
    .Y(_03390_),
    .D(_03389_));
 sg13g2_a22oi_1 _17580_ (.Y(_03391_),
    .B1(net5914),
    .B2(\soc_inst.cpu_core.register_file.registers[27][30] ),
    .A2(net5975),
    .A1(\soc_inst.cpu_core.register_file.registers[31][30] ));
 sg13g2_a22oi_1 _17581_ (.Y(_03392_),
    .B1(net5935),
    .B2(\soc_inst.cpu_core.register_file.registers[30][30] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][30] ));
 sg13g2_nand4_1 _17582_ (.B(_03377_),
    .C(_03391_),
    .A(_03376_),
    .Y(_03393_),
    .D(_03392_));
 sg13g2_nor3_2 _17583_ (.A(_03386_),
    .B(_03390_),
    .C(_03393_),
    .Y(_03394_));
 sg13g2_o21ai_1 _17584_ (.B1(net5298),
    .Y(_03395_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][30] ),
    .A2(net5925));
 sg13g2_or2_1 _17585_ (.X(_03396_),
    .B(_03395_),
    .A(_03394_));
 sg13g2_o21ai_1 _17586_ (.B1(_03396_),
    .Y(_01026_),
    .A1(net6148),
    .A2(_08058_));
 sg13g2_nand2_1 _17587_ (.Y(_03397_),
    .A(\soc_inst.cpu_core.register_file.registers[27][31] ),
    .B(net5915));
 sg13g2_a22oi_1 _17588_ (.Y(_03398_),
    .B1(net5500),
    .B2(\soc_inst.cpu_core.register_file.registers[16][31] ),
    .A2(net5956),
    .A1(\soc_inst.cpu_core.register_file.registers[11][31] ));
 sg13g2_a22oi_1 _17589_ (.Y(_03399_),
    .B1(net5505),
    .B2(\soc_inst.cpu_core.register_file.registers[17][31] ),
    .A2(net5950),
    .A1(\soc_inst.cpu_core.register_file.registers[15][31] ));
 sg13g2_a22oi_1 _17590_ (.Y(_03400_),
    .B1(net5905),
    .B2(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .A2(net5516),
    .A1(\soc_inst.cpu_core.register_file.registers[19][31] ));
 sg13g2_a22oi_1 _17591_ (.Y(_03401_),
    .B1(net5899),
    .B2(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .A2(net5971),
    .A1(\soc_inst.cpu_core.register_file.registers[6][31] ));
 sg13g2_a22oi_1 _17592_ (.Y(_03402_),
    .B1(net5945),
    .B2(\soc_inst.cpu_core.register_file.registers[22][31] ),
    .A2(net5980),
    .A1(\soc_inst.cpu_core.register_file.registers[9][31] ));
 sg13g2_a22oi_1 _17593_ (.Y(_03403_),
    .B1(net5976),
    .B2(\soc_inst.cpu_core.register_file.registers[31][31] ),
    .A2(net5990),
    .A1(\soc_inst.cpu_core.register_file.registers[20][31] ));
 sg13g2_nand4_1 _17594_ (.B(_03401_),
    .C(_03402_),
    .A(_03400_),
    .Y(_03404_),
    .D(_03403_));
 sg13g2_a22oi_1 _17595_ (.Y(_03405_),
    .B1(net5909),
    .B2(\soc_inst.cpu_core.register_file.registers[24][31] ),
    .A2(net5491),
    .A1(\soc_inst.cpu_core.register_file.registers[21][31] ));
 sg13g2_a22oi_1 _17596_ (.Y(_03406_),
    .B1(net5511),
    .B2(\soc_inst.cpu_core.register_file.registers[18][31] ),
    .A2(net5960),
    .A1(\soc_inst.cpu_core.register_file.registers[26][31] ));
 sg13g2_a22oi_1 _17597_ (.Y(_03407_),
    .B1(net5919),
    .B2(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .A2(net5964),
    .A1(\soc_inst.cpu_core.register_file.registers[14][31] ));
 sg13g2_a22oi_1 _17598_ (.Y(_03408_),
    .B1(net5931),
    .B2(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .A2(net5941),
    .A1(\soc_inst.cpu_core.register_file.registers[3][31] ));
 sg13g2_nand4_1 _17599_ (.B(_03406_),
    .C(_03407_),
    .A(_03399_),
    .Y(_03409_),
    .D(_03408_));
 sg13g2_a22oi_1 _17600_ (.Y(_03410_),
    .B1(net5885),
    .B2(\soc_inst.cpu_core.register_file.registers[5][31] ),
    .A2(net5985),
    .A1(\soc_inst.cpu_core.register_file.registers[2][31] ));
 sg13g2_a22oi_1 _17601_ (.Y(_03411_),
    .B1(net5496),
    .B2(\soc_inst.cpu_core.register_file.registers[25][31] ),
    .A2(net5996),
    .A1(\soc_inst.cpu_core.register_file.registers[23][31] ));
 sg13g2_nand4_1 _17602_ (.B(_03405_),
    .C(_03410_),
    .A(_03397_),
    .Y(_03412_),
    .D(_03411_));
 sg13g2_a21oi_1 _17603_ (.A1(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .A2(net5894),
    .Y(_03413_),
    .B1(net6084));
 sg13g2_a22oi_1 _17604_ (.Y(_03414_),
    .B1(net5889),
    .B2(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .A2(net5935),
    .A1(\soc_inst.cpu_core.register_file.registers[30][31] ));
 sg13g2_a22oi_1 _17605_ (.Y(_03415_),
    .B1(net5879),
    .B2(\soc_inst.cpu_core.register_file.registers[28][31] ),
    .A2(net5485),
    .A1(\soc_inst.cpu_core.register_file.registers[29][31] ));
 sg13g2_nand4_1 _17606_ (.B(_03413_),
    .C(_03414_),
    .A(_03398_),
    .Y(_03416_),
    .D(_03415_));
 sg13g2_nor4_2 _17607_ (.A(_03404_),
    .B(_03409_),
    .C(_03412_),
    .Y(_03417_),
    .D(_03416_));
 sg13g2_nor2_1 _17608_ (.A(_02675_),
    .B(_03417_),
    .Y(_03418_));
 sg13g2_o21ai_1 _17609_ (.B1(_03418_),
    .Y(_03419_),
    .A1(\soc_inst.cpu_core.register_file.registers[1][31] ),
    .A2(net5923));
 sg13g2_o21ai_1 _17610_ (.B1(_03419_),
    .Y(_01027_),
    .A1(net6143),
    .A2(_08057_));
 sg13g2_mux2_1 _17611_ (.A0(_00261_),
    .A1(net2301),
    .S(net6327),
    .X(_01028_));
 sg13g2_mux2_1 _17612_ (.A0(_00262_),
    .A1(net2582),
    .S(net6328),
    .X(_01029_));
 sg13g2_mux2_1 _17613_ (.A0(\soc_inst.cpu_core.ex_instr[2] ),
    .A1(net1982),
    .S(net6328),
    .X(_01030_));
 sg13g2_mux2_1 _17614_ (.A0(\soc_inst.cpu_core.ex_instr[3] ),
    .A1(net2275),
    .S(net6328),
    .X(_01031_));
 sg13g2_nand2_1 _17615_ (.Y(_03420_),
    .A(net1831),
    .B(net6364));
 sg13g2_o21ai_1 _17616_ (.B1(_03420_),
    .Y(_01032_),
    .A1(_07791_),
    .A2(net6364));
 sg13g2_mux2_1 _17617_ (.A0(net2774),
    .A1(\soc_inst.cpu_core.mem_instr[5] ),
    .S(net6369),
    .X(_01033_));
 sg13g2_mux2_1 _17618_ (.A0(\soc_inst.cpu_core.ex_instr[6] ),
    .A1(net3023),
    .S(net6364),
    .X(_01034_));
 sg13g2_mux2_1 _17619_ (.A0(net2130),
    .A1(net3231),
    .S(net6417),
    .X(_01035_));
 sg13g2_mux2_1 _17620_ (.A0(net2978),
    .A1(net6305),
    .S(net6366),
    .X(_01036_));
 sg13g2_nor2_1 _17621_ (.A(net3028),
    .B(net6360),
    .Y(_03421_));
 sg13g2_a21oi_1 _17622_ (.A1(net6173),
    .A2(net6359),
    .Y(_01037_),
    .B1(_03421_));
 sg13g2_nor2_1 _17623_ (.A(net1756),
    .B(net6359),
    .Y(_03422_));
 sg13g2_a21oi_1 _17624_ (.A1(net6169),
    .A2(net6359),
    .Y(_01038_),
    .B1(_03422_));
 sg13g2_nand2_1 _17625_ (.Y(_03423_),
    .A(net6351),
    .B(net1083));
 sg13g2_o21ai_1 _17626_ (.B1(_03423_),
    .Y(_01039_),
    .A1(net6333),
    .A2(_08173_));
 sg13g2_mux2_1 _17627_ (.A0(\soc_inst.cpu_core.ex_instr[16] ),
    .A1(net2384),
    .S(net6360),
    .X(_01040_));
 sg13g2_nand2_1 _17628_ (.Y(_03424_),
    .A(net6351),
    .B(\soc_inst.cpu_core.mem_instr[17] ));
 sg13g2_o21ai_1 _17629_ (.B1(_03424_),
    .Y(_01041_),
    .A1(net6351),
    .A2(_08175_));
 sg13g2_mux2_1 _17630_ (.A0(\soc_inst.cpu_core.ex_instr[18] ),
    .A1(net2282),
    .S(net6366),
    .X(_01042_));
 sg13g2_mux2_1 _17631_ (.A0(\soc_inst.cpu_core.ex_instr[19] ),
    .A1(net1404),
    .S(net6364),
    .X(_01043_));
 sg13g2_nand2_1 _17632_ (.Y(_03425_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .B(net6348));
 sg13g2_o21ai_1 _17633_ (.B1(_03425_),
    .Y(_01044_),
    .A1(net6340),
    .A2(_08176_));
 sg13g2_mux2_1 _17634_ (.A0(net2487),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .S(net6390),
    .X(_01045_));
 sg13g2_nor2_1 _17635_ (.A(net6333),
    .B(net1281),
    .Y(_03426_));
 sg13g2_a21oi_1 _17636_ (.A1(_07805_),
    .A2(net6333),
    .Y(_01046_),
    .B1(_03426_));
 sg13g2_mux2_1 _17637_ (.A0(net2715),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .S(net6388),
    .X(_01047_));
 sg13g2_mux2_1 _17638_ (.A0(net2661),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .S(net6351),
    .X(_01048_));
 sg13g2_nand2_1 _17639_ (.Y(_03427_),
    .A(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .B(net6333));
 sg13g2_o21ai_1 _17640_ (.B1(_03427_),
    .Y(_01049_),
    .A1(net6333),
    .A2(_08179_));
 sg13g2_mux2_1 _17641_ (.A0(net2338),
    .A1(net2444),
    .S(net6348),
    .X(_01050_));
 sg13g2_mux2_1 _17642_ (.A0(net2393),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .S(net6349),
    .X(_01051_));
 sg13g2_nor2_1 _17643_ (.A(net6333),
    .B(\soc_inst.cpu_core.ex_funct7[3] ),
    .Y(_03428_));
 sg13g2_a21oi_1 _17644_ (.A1(_07807_),
    .A2(net6325),
    .Y(_01052_),
    .B1(_03428_));
 sg13g2_mux2_1 _17645_ (.A0(net2371),
    .A1(net2572),
    .S(net6352),
    .X(_01053_));
 sg13g2_mux2_1 _17646_ (.A0(net2098),
    .A1(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .S(net6350),
    .X(_01054_));
 sg13g2_mux2_1 _17647_ (.A0(net2785),
    .A1(net2808),
    .S(net6389),
    .X(_01055_));
 sg13g2_nor4_2 _17648_ (.A(net6431),
    .B(net6436),
    .C(net6435),
    .Y(_03429_),
    .D(net6433));
 sg13g2_nor3_2 _17649_ (.A(net6401),
    .B(_11390_),
    .C(net6076),
    .Y(_03430_));
 sg13g2_a21oi_1 _17650_ (.A1(net1209),
    .A2(net5103),
    .Y(_03431_),
    .B1(net5293));
 sg13g2_nand2b_2 _17651_ (.Y(_03432_),
    .B(net6434),
    .A_N(net6432));
 sg13g2_nor4_1 _17652_ (.A(net6430),
    .B(net6436),
    .C(net6438),
    .D(_03432_),
    .Y(_03433_));
 sg13g2_nor2_1 _17653_ (.A(net6141),
    .B(net6436),
    .Y(_03434_));
 sg13g2_nand2_2 _17654_ (.Y(_03435_),
    .A(net6438),
    .B(_03434_));
 sg13g2_nand2b_2 _17655_ (.Y(_03436_),
    .B(net6432),
    .A_N(net6434));
 sg13g2_nor2_1 _17656_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 sg13g2_nand2_2 _17657_ (.Y(_03438_),
    .A(net6437),
    .B(net6438));
 sg13g2_nand2_2 _17658_ (.Y(_03439_),
    .A(net6435),
    .B(net6432));
 sg13g2_nor3_1 _17659_ (.A(net6141),
    .B(_03438_),
    .C(_03439_),
    .Y(_03440_));
 sg13g2_nor3_1 _17660_ (.A(net6141),
    .B(_03432_),
    .C(_03438_),
    .Y(_03441_));
 sg13g2_nor4_1 _17661_ (.A(net6141),
    .B(net6434),
    .C(net6432),
    .D(_03438_),
    .Y(_03442_));
 sg13g2_nand2b_2 _17662_ (.Y(_03443_),
    .B(_03434_),
    .A_N(net6439));
 sg13g2_nor3_1 _17663_ (.A(net6434),
    .B(net6432),
    .C(_03443_),
    .Y(_03444_));
 sg13g2_nor4_1 _17664_ (.A(net6430),
    .B(net6437),
    .C(net6439),
    .D(_03439_),
    .Y(_03445_));
 sg13g2_nand3_1 _17665_ (.B(_08132_),
    .C(net6439),
    .A(_08131_),
    .Y(_03446_));
 sg13g2_nor2_1 _17666_ (.A(_03432_),
    .B(_03446_),
    .Y(_03447_));
 sg13g2_nand2b_2 _17667_ (.Y(_03448_),
    .B(net6437),
    .A_N(net6439));
 sg13g2_nor4_1 _17668_ (.A(net6429),
    .B(net6434),
    .C(net6432),
    .D(_03448_),
    .Y(_03449_));
 sg13g2_nor2_1 _17669_ (.A(_03432_),
    .B(_03443_),
    .Y(_03450_));
 sg13g2_nor3_1 _17670_ (.A(net6141),
    .B(_03436_),
    .C(_03448_),
    .Y(_03451_));
 sg13g2_nor3_1 _17671_ (.A(net6429),
    .B(_03436_),
    .C(_03448_),
    .Y(_03452_));
 sg13g2_nor3_1 _17672_ (.A(net6429),
    .B(_03439_),
    .C(_03448_),
    .Y(_03453_));
 sg13g2_nor3_1 _17673_ (.A(net6141),
    .B(_03439_),
    .C(_03448_),
    .Y(_03454_));
 sg13g2_nor4_1 _17674_ (.A(net6141),
    .B(net6434),
    .C(net6432),
    .D(_03448_),
    .Y(_03455_));
 sg13g2_nor3_1 _17675_ (.A(net6434),
    .B(net6433),
    .C(_03435_),
    .Y(_03456_));
 sg13g2_nor4_1 _17676_ (.A(net6430),
    .B(net6437),
    .C(net6439),
    .D(_03436_),
    .Y(_03457_));
 sg13g2_nor3_1 _17677_ (.A(net6429),
    .B(_03436_),
    .C(_03438_),
    .Y(_03458_));
 sg13g2_nor2_1 _17678_ (.A(_03436_),
    .B(_03446_),
    .Y(_03459_));
 sg13g2_nor3_1 _17679_ (.A(_08131_),
    .B(_03436_),
    .C(_03438_),
    .Y(_03460_));
 sg13g2_nor2_1 _17680_ (.A(_03432_),
    .B(_03435_),
    .Y(_03461_));
 sg13g2_nand2_1 _17681_ (.Y(_03462_),
    .A(\soc_inst.cpu_core.register_file.registers[21][0] ),
    .B(net5267));
 sg13g2_nor3_1 _17682_ (.A(net6429),
    .B(_03438_),
    .C(_03439_),
    .Y(_03463_));
 sg13g2_nor2_1 _17683_ (.A(_03439_),
    .B(_03446_),
    .Y(_03464_));
 sg13g2_nor2_1 _17684_ (.A(_03435_),
    .B(_03439_),
    .Y(_03465_));
 sg13g2_nor3_1 _17685_ (.A(net6141),
    .B(_03432_),
    .C(_03448_),
    .Y(_03466_));
 sg13g2_nor3_1 _17686_ (.A(net6429),
    .B(_03432_),
    .C(_03448_),
    .Y(_03467_));
 sg13g2_nor2_1 _17687_ (.A(_03439_),
    .B(_03443_),
    .Y(_03468_));
 sg13g2_nor2_1 _17688_ (.A(_03436_),
    .B(_03443_),
    .Y(_03469_));
 sg13g2_a22oi_1 _17689_ (.Y(_03470_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][0] ),
    .A2(net5257),
    .A1(\soc_inst.cpu_core.register_file.registers[28][0] ));
 sg13g2_nor4_1 _17690_ (.A(net6429),
    .B(net6434),
    .C(net6432),
    .D(_03438_),
    .Y(_03471_));
 sg13g2_nor3_1 _17691_ (.A(net6429),
    .B(_03432_),
    .C(_03438_),
    .Y(_03472_));
 sg13g2_a22oi_1 _17692_ (.Y(_03473_),
    .B1(net5832),
    .B2(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][0] ));
 sg13g2_a22oi_1 _17693_ (.Y(_03474_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .A2(net5807),
    .A1(\soc_inst.cpu_core.register_file.registers[27][0] ));
 sg13g2_a22oi_1 _17694_ (.Y(_03475_),
    .B1(net5797),
    .B2(\soc_inst.cpu_core.register_file.registers[22][0] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][0] ));
 sg13g2_a22oi_1 _17695_ (.Y(_03476_),
    .B1(net5852),
    .B2(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][0] ));
 sg13g2_a22oi_1 _17696_ (.Y(_03477_),
    .B1(net5812),
    .B2(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .A2(net5867),
    .A1(\soc_inst.cpu_core.register_file.registers[31][0] ));
 sg13g2_a22oi_1 _17697_ (.Y(_03478_),
    .B1(net5837),
    .B2(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .A2(net5842),
    .A1(\soc_inst.cpu_core.register_file.registers[26][0] ));
 sg13g2_a22oi_1 _17698_ (.Y(_03479_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .A2(net5872),
    .A1(\soc_inst.cpu_core.register_file.registers[4][0] ));
 sg13g2_a22oi_1 _17699_ (.Y(_03480_),
    .B1(net5827),
    .B2(\soc_inst.cpu_core.register_file.registers[30][0] ),
    .A2(net5277),
    .A1(\soc_inst.cpu_core.register_file.registers[20][0] ));
 sg13g2_a22oi_1 _17700_ (.Y(_03481_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .A2(net5272),
    .A1(\soc_inst.cpu_core.register_file.registers[17][0] ));
 sg13g2_nand4_1 _17701_ (.B(_03479_),
    .C(_03480_),
    .A(_03475_),
    .Y(_03482_),
    .D(_03481_));
 sg13g2_a22oi_1 _17702_ (.Y(_03483_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .A2(net5817),
    .A1(\soc_inst.cpu_core.register_file.registers[8][0] ));
 sg13g2_nand4_1 _17703_ (.B(_03476_),
    .C(_03477_),
    .A(_03462_),
    .Y(_03484_),
    .D(_03483_));
 sg13g2_nor2_1 _17704_ (.A(_03482_),
    .B(_03484_),
    .Y(_03485_));
 sg13g2_a21oi_1 _17705_ (.A1(\soc_inst.cpu_core.register_file.registers[29][0] ),
    .A2(net5262),
    .Y(_03486_),
    .B1(net6077));
 sg13g2_a22oi_1 _17706_ (.Y(_03487_),
    .B1(net5792),
    .B2(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .A2(net5847),
    .A1(\soc_inst.cpu_core.register_file.registers[2][0] ));
 sg13g2_nand4_1 _17707_ (.B(_03478_),
    .C(_03486_),
    .A(_03470_),
    .Y(_03488_),
    .D(_03487_));
 sg13g2_a22oi_1 _17708_ (.Y(_03489_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][0] ),
    .A2(net5478),
    .A1(\soc_inst.cpu_core.register_file.registers[5][0] ));
 sg13g2_a22oi_1 _17709_ (.Y(_03490_),
    .B1(net5473),
    .B2(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][0] ));
 sg13g2_nand4_1 _17710_ (.B(_03474_),
    .C(_03489_),
    .A(_03473_),
    .Y(_03491_),
    .D(_03490_));
 sg13g2_nor2_1 _17711_ (.A(_03488_),
    .B(_03491_),
    .Y(_03492_));
 sg13g2_a21oi_2 _17712_ (.B1(_03431_),
    .Y(_03493_),
    .A2(_03492_),
    .A1(_03485_));
 sg13g2_a21o_1 _17713_ (.A2(net1491),
    .A1(net6423),
    .B1(_03493_),
    .X(_01056_));
 sg13g2_a21oi_1 _17714_ (.A1(net1139),
    .A2(net5103),
    .Y(_03494_),
    .B1(net5293));
 sg13g2_nand2_1 _17715_ (.Y(_03495_),
    .A(\soc_inst.cpu_core.register_file.registers[28][1] ),
    .B(net5257));
 sg13g2_a22oi_1 _17716_ (.Y(_03496_),
    .B1(net5812),
    .B2(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][1] ));
 sg13g2_a22oi_1 _17717_ (.Y(_03497_),
    .B1(net5262),
    .B2(\soc_inst.cpu_core.register_file.registers[29][1] ),
    .A2(net5852),
    .A1(\soc_inst.cpu_core.register_file.registers[12][1] ));
 sg13g2_a22oi_1 _17718_ (.Y(_03498_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][1] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][1] ));
 sg13g2_a22oi_1 _17719_ (.Y(_03499_),
    .B1(net5797),
    .B2(\soc_inst.cpu_core.register_file.registers[22][1] ),
    .A2(net5837),
    .A1(\soc_inst.cpu_core.register_file.registers[10][1] ));
 sg13g2_a22oi_1 _17720_ (.Y(_03500_),
    .B1(net5277),
    .B2(\soc_inst.cpu_core.register_file.registers[20][1] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][1] ));
 sg13g2_a22oi_1 _17721_ (.Y(_03501_),
    .B1(net5473),
    .B2(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .A2(net5842),
    .A1(\soc_inst.cpu_core.register_file.registers[26][1] ));
 sg13g2_a22oi_1 _17722_ (.Y(_03502_),
    .B1(net5792),
    .B2(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .A2(net5827),
    .A1(\soc_inst.cpu_core.register_file.registers[30][1] ));
 sg13g2_a22oi_1 _17723_ (.Y(_03503_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][1] ),
    .A2(net5267),
    .A1(\soc_inst.cpu_core.register_file.registers[21][1] ));
 sg13g2_a22oi_1 _17724_ (.Y(_03504_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .A2(net5832),
    .A1(\soc_inst.cpu_core.register_file.registers[14][1] ));
 sg13g2_nand4_1 _17725_ (.B(_03502_),
    .C(_03503_),
    .A(_03501_),
    .Y(_03505_),
    .D(_03504_));
 sg13g2_a22oi_1 _17726_ (.Y(_03506_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .A2(net5872),
    .A1(\soc_inst.cpu_core.register_file.registers[4][1] ));
 sg13g2_a22oi_1 _17727_ (.Y(_03507_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][1] ),
    .A2(net5867),
    .A1(\soc_inst.cpu_core.register_file.registers[31][1] ));
 sg13g2_nand4_1 _17728_ (.B(_03500_),
    .C(_03506_),
    .A(_03498_),
    .Y(_03508_),
    .D(_03507_));
 sg13g2_a22oi_1 _17729_ (.Y(_03509_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .A2(net5817),
    .A1(\soc_inst.cpu_core.register_file.registers[8][1] ));
 sg13g2_nand4_1 _17730_ (.B(_03496_),
    .C(_03497_),
    .A(_03495_),
    .Y(_03510_),
    .D(_03509_));
 sg13g2_a21oi_1 _17731_ (.A1(\soc_inst.cpu_core.register_file.registers[23][1] ),
    .A2(net5862),
    .Y(_03511_),
    .B1(net6077));
 sg13g2_a22oi_1 _17732_ (.Y(_03512_),
    .B1(net5847),
    .B2(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .A2(net5478),
    .A1(\soc_inst.cpu_core.register_file.registers[5][1] ));
 sg13g2_a22oi_1 _17733_ (.Y(_03513_),
    .B1(net5807),
    .B2(\soc_inst.cpu_core.register_file.registers[27][1] ),
    .A2(net5272),
    .A1(\soc_inst.cpu_core.register_file.registers[17][1] ));
 sg13g2_nand4_1 _17734_ (.B(_03511_),
    .C(_03512_),
    .A(_03499_),
    .Y(_03514_),
    .D(_03513_));
 sg13g2_nor4_1 _17735_ (.A(_03505_),
    .B(_03508_),
    .C(_03510_),
    .D(_03514_),
    .Y(_03515_));
 sg13g2_nor2_2 _17736_ (.A(_03494_),
    .B(_03515_),
    .Y(_03516_));
 sg13g2_a21o_1 _17737_ (.A2(net1466),
    .A1(net6423),
    .B1(_03516_),
    .X(_01057_));
 sg13g2_a21oi_1 _17738_ (.A1(net507),
    .A2(net5103),
    .Y(_03517_),
    .B1(net5292));
 sg13g2_nand2_1 _17739_ (.Y(_03518_),
    .A(\soc_inst.cpu_core.register_file.registers[25][2] ),
    .B(net5287));
 sg13g2_a22oi_1 _17740_ (.Y(_03519_),
    .B1(net5827),
    .B2(\soc_inst.cpu_core.register_file.registers[30][2] ),
    .A2(net5837),
    .A1(\soc_inst.cpu_core.register_file.registers[10][2] ));
 sg13g2_a22oi_1 _17741_ (.Y(_03520_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][2] ),
    .A2(net5842),
    .A1(\soc_inst.cpu_core.register_file.registers[26][2] ));
 sg13g2_a22oi_1 _17742_ (.Y(_03521_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][2] ),
    .A2(net5812),
    .A1(\soc_inst.cpu_core.register_file.registers[11][2] ));
 sg13g2_a22oi_1 _17743_ (.Y(_03522_),
    .B1(net5852),
    .B2(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][2] ));
 sg13g2_a22oi_1 _17744_ (.Y(_03523_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .A2(net5872),
    .A1(\soc_inst.cpu_core.register_file.registers[4][2] ));
 sg13g2_a22oi_1 _17745_ (.Y(_03524_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .A2(net5272),
    .A1(\soc_inst.cpu_core.register_file.registers[17][2] ));
 sg13g2_a22oi_1 _17746_ (.Y(_03525_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .A2(net5817),
    .A1(\soc_inst.cpu_core.register_file.registers[8][2] ));
 sg13g2_nand4_1 _17747_ (.B(_03523_),
    .C(_03524_),
    .A(_03520_),
    .Y(_03526_),
    .D(_03525_));
 sg13g2_a22oi_1 _17748_ (.Y(_03527_),
    .B1(net5267),
    .B2(\soc_inst.cpu_core.register_file.registers[21][2] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][2] ));
 sg13g2_nand4_1 _17749_ (.B(_03521_),
    .C(_03522_),
    .A(_03518_),
    .Y(_03528_),
    .D(_03527_));
 sg13g2_nor2_1 _17750_ (.A(_03526_),
    .B(_03528_),
    .Y(_03529_));
 sg13g2_a21oi_1 _17751_ (.A1(\soc_inst.cpu_core.register_file.registers[29][2] ),
    .A2(net5262),
    .Y(_03530_),
    .B1(net6077));
 sg13g2_a22oi_1 _17752_ (.Y(_03531_),
    .B1(net5847),
    .B2(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .A2(net5478),
    .A1(\soc_inst.cpu_core.register_file.registers[5][2] ));
 sg13g2_a22oi_1 _17753_ (.Y(_03532_),
    .B1(net5792),
    .B2(\soc_inst.cpu_core.register_file.registers[6][2] ),
    .A2(net5807),
    .A1(\soc_inst.cpu_core.register_file.registers[27][2] ));
 sg13g2_nand4_1 _17754_ (.B(_03530_),
    .C(_03531_),
    .A(_03519_),
    .Y(_03533_),
    .D(_03532_));
 sg13g2_a22oi_1 _17755_ (.Y(_03534_),
    .B1(net5473),
    .B2(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][2] ));
 sg13g2_a22oi_1 _17756_ (.Y(_03535_),
    .B1(net5257),
    .B2(\soc_inst.cpu_core.register_file.registers[28][2] ),
    .A2(net5797),
    .A1(\soc_inst.cpu_core.register_file.registers[22][2] ));
 sg13g2_a22oi_1 _17757_ (.Y(_03536_),
    .B1(net5277),
    .B2(\soc_inst.cpu_core.register_file.registers[20][2] ),
    .A2(net5867),
    .A1(\soc_inst.cpu_core.register_file.registers[31][2] ));
 sg13g2_a22oi_1 _17758_ (.Y(_03537_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .A2(net5832),
    .A1(\soc_inst.cpu_core.register_file.registers[14][2] ));
 sg13g2_nand4_1 _17759_ (.B(_03535_),
    .C(_03536_),
    .A(_03534_),
    .Y(_03538_),
    .D(_03537_));
 sg13g2_nor2_1 _17760_ (.A(_03533_),
    .B(_03538_),
    .Y(_03539_));
 sg13g2_a21oi_2 _17761_ (.B1(_03517_),
    .Y(_03540_),
    .A2(_03539_),
    .A1(_03529_));
 sg13g2_a21o_1 _17762_ (.A2(net1291),
    .A1(net6418),
    .B1(_03540_),
    .X(_01058_));
 sg13g2_a22oi_1 _17763_ (.Y(_03541_),
    .B1(net5786),
    .B2(\soc_inst.cpu_core.register_file.registers[3][3] ),
    .A2(net5261),
    .A1(\soc_inst.cpu_core.register_file.registers[29][3] ));
 sg13g2_and2_1 _17764_ (.A(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .B(net5831),
    .X(_03542_));
 sg13g2_a22oi_1 _17765_ (.Y(_03543_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .A2(net5816),
    .A1(\soc_inst.cpu_core.register_file.registers[8][3] ));
 sg13g2_a22oi_1 _17766_ (.Y(_03544_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][3] ),
    .A2(net5276),
    .A1(\soc_inst.cpu_core.register_file.registers[20][3] ));
 sg13g2_nand3_1 _17767_ (.B(_03543_),
    .C(_03544_),
    .A(_03541_),
    .Y(_03545_));
 sg13g2_a221oi_1 _17768_ (.B2(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .C1(_03545_),
    .B1(net5801),
    .A1(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .Y(_03546_),
    .A2(net5836));
 sg13g2_a22oi_1 _17769_ (.Y(_03547_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][3] ),
    .A2(net5266),
    .A1(\soc_inst.cpu_core.register_file.registers[21][3] ));
 sg13g2_a22oi_1 _17770_ (.Y(_03548_),
    .B1(net5467),
    .B2(\soc_inst.cpu_core.register_file.registers[13][3] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][3] ));
 sg13g2_a221oi_1 _17771_ (.B2(\soc_inst.cpu_core.register_file.registers[27][3] ),
    .C1(_03542_),
    .B1(net5806),
    .A1(\soc_inst.cpu_core.register_file.registers[25][3] ),
    .Y(_03549_),
    .A2(net5286));
 sg13g2_nand4_1 _17772_ (.B(_03547_),
    .C(_03548_),
    .A(_03546_),
    .Y(_03550_),
    .D(_03549_));
 sg13g2_a21oi_1 _17773_ (.A1(\soc_inst.cpu_core.register_file.registers[23][3] ),
    .A2(net5861),
    .Y(_03551_),
    .B1(net6076));
 sg13g2_a22oi_1 _17774_ (.Y(_03552_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][3] ));
 sg13g2_a22oi_1 _17775_ (.Y(_03553_),
    .B1(net5841),
    .B2(\soc_inst.cpu_core.register_file.registers[26][3] ),
    .A2(net5846),
    .A1(\soc_inst.cpu_core.register_file.registers[2][3] ));
 sg13g2_a22oi_1 _17776_ (.Y(_03554_),
    .B1(net5821),
    .B2(\soc_inst.cpu_core.register_file.registers[18][3] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][3] ));
 sg13g2_nand4_1 _17777_ (.B(_03552_),
    .C(_03553_),
    .A(_03551_),
    .Y(_03555_),
    .D(_03554_));
 sg13g2_a22oi_1 _17778_ (.Y(_03556_),
    .B1(net5271),
    .B2(\soc_inst.cpu_core.register_file.registers[17][3] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][3] ));
 sg13g2_a22oi_1 _17779_ (.Y(_03557_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .A2(net5851),
    .A1(\soc_inst.cpu_core.register_file.registers[12][3] ));
 sg13g2_a22oi_1 _17780_ (.Y(_03558_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][3] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][3] ));
 sg13g2_a22oi_1 _17781_ (.Y(_03559_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .A2(net5871),
    .A1(\soc_inst.cpu_core.register_file.registers[4][3] ));
 sg13g2_nand4_1 _17782_ (.B(_03557_),
    .C(_03558_),
    .A(_03556_),
    .Y(_03560_),
    .D(_03559_));
 sg13g2_nor3_2 _17783_ (.A(_03550_),
    .B(_03555_),
    .C(_03560_),
    .Y(_03561_));
 sg13g2_a21oi_1 _17784_ (.A1(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .A2(net5104),
    .Y(_03562_),
    .B1(net5294));
 sg13g2_or2_1 _17785_ (.X(_03563_),
    .B(_03562_),
    .A(_03561_));
 sg13g2_o21ai_1 _17786_ (.B1(_03563_),
    .Y(_01059_),
    .A1(net6145),
    .A2(_08032_));
 sg13g2_a22oi_1 _17787_ (.Y(_03564_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .A2(net5808),
    .A1(\soc_inst.cpu_core.register_file.registers[27][4] ));
 sg13g2_and2_1 _17788_ (.A(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .B(net5788),
    .X(_03565_));
 sg13g2_a22oi_1 _17789_ (.Y(_03566_),
    .B1(net5803),
    .B2(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .A2(net5278),
    .A1(\soc_inst.cpu_core.register_file.registers[20][4] ));
 sg13g2_a22oi_1 _17790_ (.Y(_03567_),
    .B1(net5273),
    .B2(\soc_inst.cpu_core.register_file.registers[17][4] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][4] ));
 sg13g2_a22oi_1 _17791_ (.Y(_03568_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][4] ),
    .A2(net5813),
    .A1(\soc_inst.cpu_core.register_file.registers[11][4] ));
 sg13g2_a22oi_1 _17792_ (.Y(_03569_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .A2(net5479),
    .A1(\soc_inst.cpu_core.register_file.registers[5][4] ));
 sg13g2_a22oi_1 _17793_ (.Y(_03570_),
    .B1(net5838),
    .B2(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][4] ));
 sg13g2_nand3_1 _17794_ (.B(_03569_),
    .C(_03570_),
    .A(_03568_),
    .Y(_03571_));
 sg13g2_a221oi_1 _17795_ (.B2(\soc_inst.cpu_core.register_file.registers[30][4] ),
    .C1(_03571_),
    .B1(net5828),
    .A1(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .Y(_03572_),
    .A2(net5848));
 sg13g2_a22oi_1 _17796_ (.Y(_03573_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][4] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][4] ));
 sg13g2_a22oi_1 _17797_ (.Y(_03574_),
    .B1(net5474),
    .B2(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][4] ));
 sg13g2_a221oi_1 _17798_ (.B2(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .C1(_03565_),
    .B1(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[25][4] ),
    .Y(_03575_),
    .A2(net5288));
 sg13g2_nand4_1 _17799_ (.B(_03573_),
    .C(_03574_),
    .A(_03572_),
    .Y(_03576_),
    .D(_03575_));
 sg13g2_a21oi_1 _17800_ (.A1(\soc_inst.cpu_core.register_file.registers[24][4] ),
    .A2(net5253),
    .Y(_03577_),
    .B1(net6078));
 sg13g2_a22oi_1 _17801_ (.Y(_03578_),
    .B1(net5258),
    .B2(\soc_inst.cpu_core.register_file.registers[28][4] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][4] ));
 sg13g2_a22oi_1 _17802_ (.Y(_03579_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][4] ));
 sg13g2_nand4_1 _17803_ (.B(_03577_),
    .C(_03578_),
    .A(_03566_),
    .Y(_03580_),
    .D(_03579_));
 sg13g2_a22oi_1 _17804_ (.Y(_03581_),
    .B1(net5467),
    .B2(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .A2(net5863),
    .A1(\soc_inst.cpu_core.register_file.registers[23][4] ));
 sg13g2_a22oi_1 _17805_ (.Y(_03582_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][4] ),
    .A2(net5843),
    .A1(\soc_inst.cpu_core.register_file.registers[26][4] ));
 sg13g2_nand4_1 _17806_ (.B(_03567_),
    .C(_03581_),
    .A(_03564_),
    .Y(_03583_),
    .D(_03582_));
 sg13g2_nor3_2 _17807_ (.A(_03576_),
    .B(_03580_),
    .C(_03583_),
    .Y(_03584_));
 sg13g2_a21oi_1 _17808_ (.A1(net444),
    .A2(net5106),
    .Y(_03585_),
    .B1(_03430_));
 sg13g2_or2_1 _17809_ (.X(_03586_),
    .B(_03585_),
    .A(_03584_));
 sg13g2_o21ai_1 _17810_ (.B1(_03586_),
    .Y(_01060_),
    .A1(net6153),
    .A2(_08040_));
 sg13g2_a22oi_1 _17811_ (.Y(_03587_),
    .B1(net5260),
    .B2(\soc_inst.cpu_core.register_file.registers[28][5] ),
    .A2(net5794),
    .A1(\soc_inst.cpu_core.register_file.registers[6][5] ));
 sg13g2_and2_1 _17812_ (.A(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .B(net5481),
    .X(_03588_));
 sg13g2_a22oi_1 _17813_ (.Y(_03589_),
    .B1(net5805),
    .B2(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .A2(net5273),
    .A1(\soc_inst.cpu_core.register_file.registers[17][5] ));
 sg13g2_a22oi_1 _17814_ (.Y(_03590_),
    .B1(net5790),
    .B2(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .A2(net5810),
    .A1(\soc_inst.cpu_core.register_file.registers[27][5] ));
 sg13g2_a22oi_1 _17815_ (.Y(_03591_),
    .B1(net5820),
    .B2(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .A2(net5865),
    .A1(\soc_inst.cpu_core.register_file.registers[23][5] ));
 sg13g2_a22oi_1 _17816_ (.Y(_03592_),
    .B1(net5800),
    .B2(\soc_inst.cpu_core.register_file.registers[22][5] ),
    .A2(net5825),
    .A1(\soc_inst.cpu_core.register_file.registers[18][5] ));
 sg13g2_a22oi_1 _17817_ (.Y(_03593_),
    .B1(net5270),
    .B2(\soc_inst.cpu_core.register_file.registers[21][5] ),
    .A2(net5850),
    .A1(\soc_inst.cpu_core.register_file.registers[2][5] ));
 sg13g2_nand3_1 _17818_ (.B(_03592_),
    .C(_03593_),
    .A(_03591_),
    .Y(_03594_));
 sg13g2_a221oi_1 _17819_ (.B2(\soc_inst.cpu_core.register_file.registers[29][5] ),
    .C1(_03594_),
    .B1(net5265),
    .A1(\soc_inst.cpu_core.register_file.registers[31][5] ),
    .Y(_03595_),
    .A2(net5870));
 sg13g2_a221oi_1 _17820_ (.B2(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .C1(_03588_),
    .B1(net5815),
    .A1(\soc_inst.cpu_core.register_file.registers[16][5] ),
    .Y(_03596_),
    .A2(net5285));
 sg13g2_nand4_1 _17821_ (.B(_03590_),
    .C(_03595_),
    .A(_03589_),
    .Y(_03597_),
    .D(_03596_));
 sg13g2_a21oi_1 _17822_ (.A1(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .A2(net5833),
    .Y(_03598_),
    .B1(net6079));
 sg13g2_a22oi_1 _17823_ (.Y(_03599_),
    .B1(net5785),
    .B2(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .A2(net5860),
    .A1(\soc_inst.cpu_core.register_file.registers[19][5] ));
 sg13g2_a22oi_1 _17824_ (.Y(_03600_),
    .B1(net5476),
    .B2(\soc_inst.cpu_core.register_file.registers[9][5] ),
    .A2(net5280),
    .A1(\soc_inst.cpu_core.register_file.registers[20][5] ));
 sg13g2_nand4_1 _17825_ (.B(_03598_),
    .C(_03599_),
    .A(_03587_),
    .Y(_03601_),
    .D(_03600_));
 sg13g2_a22oi_1 _17826_ (.Y(_03602_),
    .B1(net5840),
    .B2(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .A2(net5855),
    .A1(\soc_inst.cpu_core.register_file.registers[12][5] ));
 sg13g2_a22oi_1 _17827_ (.Y(_03603_),
    .B1(net5255),
    .B2(\soc_inst.cpu_core.register_file.registers[24][5] ),
    .A2(net5844),
    .A1(\soc_inst.cpu_core.register_file.registers[26][5] ));
 sg13g2_a22oi_1 _17828_ (.Y(_03604_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .A2(net5874),
    .A1(\soc_inst.cpu_core.register_file.registers[4][5] ));
 sg13g2_a22oi_1 _17829_ (.Y(_03605_),
    .B1(net5830),
    .B2(\soc_inst.cpu_core.register_file.registers[30][5] ),
    .A2(net5290),
    .A1(\soc_inst.cpu_core.register_file.registers[25][5] ));
 sg13g2_nand4_1 _17830_ (.B(_03603_),
    .C(_03604_),
    .A(_03602_),
    .Y(_03606_),
    .D(_03605_));
 sg13g2_nor3_2 _17831_ (.A(_03597_),
    .B(_03601_),
    .C(_03606_),
    .Y(_03607_));
 sg13g2_a21oi_1 _17832_ (.A1(net1044),
    .A2(net5106),
    .Y(_03608_),
    .B1(net5293));
 sg13g2_or2_1 _17833_ (.X(_03609_),
    .B(_03608_),
    .A(_03607_));
 sg13g2_o21ai_1 _17834_ (.B1(_03609_),
    .Y(_01061_),
    .A1(net6154),
    .A2(_08038_));
 sg13g2_and2_1 _17835_ (.A(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .B(net5832),
    .X(_03610_));
 sg13g2_a22oi_1 _17836_ (.Y(_03611_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .A2(net5827),
    .A1(\soc_inst.cpu_core.register_file.registers[30][6] ));
 sg13g2_a22oi_1 _17837_ (.Y(_03612_),
    .B1(net5257),
    .B2(\soc_inst.cpu_core.register_file.registers[28][6] ),
    .A2(net5473),
    .A1(\soc_inst.cpu_core.register_file.registers[9][6] ));
 sg13g2_a22oi_1 _17838_ (.Y(_03613_),
    .B1(net5478),
    .B2(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][6] ));
 sg13g2_a22oi_1 _17839_ (.Y(_03614_),
    .B1(net5807),
    .B2(\soc_inst.cpu_core.register_file.registers[27][6] ),
    .A2(net5847),
    .A1(\soc_inst.cpu_core.register_file.registers[2][6] ));
 sg13g2_nand3_1 _17840_ (.B(_03613_),
    .C(_03614_),
    .A(_03612_),
    .Y(_03615_));
 sg13g2_a221oi_1 _17841_ (.B2(\soc_inst.cpu_core.register_file.registers[29][6] ),
    .C1(_03615_),
    .B1(net5262),
    .A1(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .Y(_03616_),
    .A2(net5468));
 sg13g2_a22oi_1 _17842_ (.Y(_03617_),
    .B1(net5267),
    .B2(\soc_inst.cpu_core.register_file.registers[21][6] ),
    .A2(net5812),
    .A1(\soc_inst.cpu_core.register_file.registers[11][6] ));
 sg13g2_a22oi_1 _17843_ (.Y(_03618_),
    .B1(net5272),
    .B2(\soc_inst.cpu_core.register_file.registers[17][6] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][6] ));
 sg13g2_a221oi_1 _17844_ (.B2(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .C1(_03610_),
    .B1(net5782),
    .A1(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .Y(_03619_),
    .A2(net5787));
 sg13g2_nand4_1 _17845_ (.B(_03617_),
    .C(_03618_),
    .A(_03616_),
    .Y(_03620_),
    .D(_03619_));
 sg13g2_a21oi_1 _17846_ (.A1(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .A2(net5792),
    .Y(_03621_),
    .B1(net6079));
 sg13g2_a22oi_1 _17847_ (.Y(_03622_),
    .B1(net5797),
    .B2(\soc_inst.cpu_core.register_file.registers[22][6] ),
    .A2(net5277),
    .A1(\soc_inst.cpu_core.register_file.registers[20][6] ));
 sg13g2_a22oi_1 _17848_ (.Y(_03623_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][6] ),
    .A2(net5872),
    .A1(\soc_inst.cpu_core.register_file.registers[4][6] ));
 sg13g2_nand4_1 _17849_ (.B(_03621_),
    .C(_03622_),
    .A(_03611_),
    .Y(_03624_),
    .D(_03623_));
 sg13g2_a22oi_1 _17850_ (.Y(_03625_),
    .B1(net5817),
    .B2(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .A2(net5837),
    .A1(\soc_inst.cpu_core.register_file.registers[10][6] ));
 sg13g2_a22oi_1 _17851_ (.Y(_03626_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][6] ),
    .A2(net5842),
    .A1(\soc_inst.cpu_core.register_file.registers[26][6] ));
 sg13g2_a22oi_1 _17852_ (.Y(_03627_),
    .B1(net5852),
    .B2(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][6] ));
 sg13g2_a22oi_1 _17853_ (.Y(_03628_),
    .B1(net5867),
    .B2(\soc_inst.cpu_core.register_file.registers[31][6] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][6] ));
 sg13g2_nand4_1 _17854_ (.B(_03626_),
    .C(_03627_),
    .A(_03625_),
    .Y(_03629_),
    .D(_03628_));
 sg13g2_nor3_2 _17855_ (.A(_03620_),
    .B(_03624_),
    .C(_03629_),
    .Y(_03630_));
 sg13g2_a21oi_1 _17856_ (.A1(net1094),
    .A2(net5103),
    .Y(_03631_),
    .B1(net5293));
 sg13g2_or2_1 _17857_ (.X(_03632_),
    .B(_03631_),
    .A(_03630_));
 sg13g2_o21ai_1 _17858_ (.B1(_03632_),
    .Y(_01062_),
    .A1(net6152),
    .A2(_08036_));
 sg13g2_and2_1 _17859_ (.A(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .B(net5479),
    .X(_03633_));
 sg13g2_a22oi_1 _17860_ (.Y(_03634_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][7] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][7] ));
 sg13g2_a22oi_1 _17861_ (.Y(_03635_),
    .B1(net5788),
    .B2(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][7] ));
 sg13g2_a22oi_1 _17862_ (.Y(_03636_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .A2(net5474),
    .A1(\soc_inst.cpu_core.register_file.registers[9][7] ));
 sg13g2_a22oi_1 _17863_ (.Y(_03637_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][7] ));
 sg13g2_a22oi_1 _17864_ (.Y(_03638_),
    .B1(net5469),
    .B2(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .A2(net5274),
    .A1(\soc_inst.cpu_core.register_file.registers[17][7] ));
 sg13g2_a22oi_1 _17865_ (.Y(_03639_),
    .B1(net5793),
    .B2(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][7] ));
 sg13g2_a22oi_1 _17866_ (.Y(_03640_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][7] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][7] ));
 sg13g2_a22oi_1 _17867_ (.Y(_03641_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][7] ),
    .A2(net5838),
    .A1(\soc_inst.cpu_core.register_file.registers[10][7] ));
 sg13g2_nand3_1 _17868_ (.B(_03640_),
    .C(_03641_),
    .A(_03639_),
    .Y(_03642_));
 sg13g2_a221oi_1 _17869_ (.B2(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .C1(_03642_),
    .B1(net5803),
    .A1(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .Y(_03643_),
    .A2(net5834));
 sg13g2_a221oi_1 _17870_ (.B2(\soc_inst.cpu_core.register_file.registers[28][7] ),
    .C1(_03633_),
    .B1(net5258),
    .A1(\soc_inst.cpu_core.register_file.registers[19][7] ),
    .Y(_03644_),
    .A2(net5858));
 sg13g2_a22oi_1 _17871_ (.Y(_03645_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][7] ),
    .A2(net5848),
    .A1(\soc_inst.cpu_core.register_file.registers[2][7] ));
 sg13g2_nand4_1 _17872_ (.B(_03643_),
    .C(_03644_),
    .A(_03638_),
    .Y(_03646_),
    .D(_03645_));
 sg13g2_a21oi_1 _17873_ (.A1(\soc_inst.cpu_core.register_file.registers[30][7] ),
    .A2(net5828),
    .Y(_03647_),
    .B1(net6078));
 sg13g2_a22oi_1 _17874_ (.Y(_03648_),
    .B1(net5813),
    .B2(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .A2(net5278),
    .A1(\soc_inst.cpu_core.register_file.registers[20][7] ));
 sg13g2_nand4_1 _17875_ (.B(_03635_),
    .C(_03647_),
    .A(_03634_),
    .Y(_03649_),
    .D(_03648_));
 sg13g2_a22oi_1 _17876_ (.Y(_03650_),
    .B1(net5843),
    .B2(\soc_inst.cpu_core.register_file.registers[26][7] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][7] ));
 sg13g2_a22oi_1 _17877_ (.Y(_03651_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][7] ),
    .A2(net5863),
    .A1(\soc_inst.cpu_core.register_file.registers[23][7] ));
 sg13g2_nand4_1 _17878_ (.B(_03637_),
    .C(_03650_),
    .A(_03636_),
    .Y(_03652_),
    .D(_03651_));
 sg13g2_nor3_2 _17879_ (.A(_03646_),
    .B(_03649_),
    .C(_03652_),
    .Y(_03653_));
 sg13g2_a21oi_1 _17880_ (.A1(net798),
    .A2(net5103),
    .Y(_03654_),
    .B1(net5292));
 sg13g2_or2_1 _17881_ (.X(_03655_),
    .B(_03654_),
    .A(_03653_));
 sg13g2_o21ai_1 _17882_ (.B1(_03655_),
    .Y(_01063_),
    .A1(net6152),
    .A2(_08034_));
 sg13g2_and2_1 _17883_ (.A(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .B(net5817),
    .X(_03656_));
 sg13g2_a22oi_1 _17884_ (.Y(_03657_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .A2(net5478),
    .A1(\soc_inst.cpu_core.register_file.registers[5][8] ));
 sg13g2_a22oi_1 _17885_ (.Y(_03658_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][8] ),
    .A2(net5827),
    .A1(\soc_inst.cpu_core.register_file.registers[30][8] ));
 sg13g2_a22oi_1 _17886_ (.Y(_03659_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][8] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][8] ));
 sg13g2_a22oi_1 _17887_ (.Y(_03660_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .A2(net5837),
    .A1(\soc_inst.cpu_core.register_file.registers[10][8] ));
 sg13g2_nand3_1 _17888_ (.B(_03659_),
    .C(_03660_),
    .A(_03658_),
    .Y(_03661_));
 sg13g2_a221oi_1 _17889_ (.B2(\soc_inst.cpu_core.register_file.registers[24][8] ),
    .C1(_03661_),
    .B1(net5252),
    .A1(\soc_inst.cpu_core.register_file.registers[27][8] ),
    .Y(_03662_),
    .A2(net5807));
 sg13g2_a22oi_1 _17890_ (.Y(_03663_),
    .B1(net5847),
    .B2(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][8] ));
 sg13g2_a22oi_1 _17891_ (.Y(_03664_),
    .B1(net5812),
    .B2(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][8] ));
 sg13g2_a221oi_1 _17892_ (.B2(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .C1(_03656_),
    .B1(net5473),
    .A1(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .Y(_03665_),
    .A2(net5832));
 sg13g2_nand4_1 _17893_ (.B(_03663_),
    .C(_03664_),
    .A(_03662_),
    .Y(_03666_),
    .D(_03665_));
 sg13g2_a21oi_1 _17894_ (.A1(\soc_inst.cpu_core.register_file.registers[31][8] ),
    .A2(net5867),
    .Y(_03667_),
    .B1(net6077));
 sg13g2_a22oi_1 _17895_ (.Y(_03668_),
    .B1(net5792),
    .B2(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .A2(net5267),
    .A1(\soc_inst.cpu_core.register_file.registers[21][8] ));
 sg13g2_a22oi_1 _17896_ (.Y(_03669_),
    .B1(net5262),
    .B2(\soc_inst.cpu_core.register_file.registers[29][8] ),
    .A2(net5842),
    .A1(\soc_inst.cpu_core.register_file.registers[26][8] ));
 sg13g2_nand4_1 _17897_ (.B(_03667_),
    .C(_03668_),
    .A(_03657_),
    .Y(_03670_),
    .D(_03669_));
 sg13g2_a22oi_1 _17898_ (.Y(_03671_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .A2(net5852),
    .A1(\soc_inst.cpu_core.register_file.registers[12][8] ));
 sg13g2_a22oi_1 _17899_ (.Y(_03672_),
    .B1(net5797),
    .B2(\soc_inst.cpu_core.register_file.registers[22][8] ),
    .A2(net5277),
    .A1(\soc_inst.cpu_core.register_file.registers[20][8] ));
 sg13g2_a22oi_1 _17900_ (.Y(_03673_),
    .B1(net5282),
    .B2(\soc_inst.cpu_core.register_file.registers[16][8] ),
    .A2(net5872),
    .A1(\soc_inst.cpu_core.register_file.registers[4][8] ));
 sg13g2_a22oi_1 _17901_ (.Y(_03674_),
    .B1(net5257),
    .B2(\soc_inst.cpu_core.register_file.registers[28][8] ),
    .A2(net5272),
    .A1(\soc_inst.cpu_core.register_file.registers[17][8] ));
 sg13g2_nand4_1 _17902_ (.B(_03672_),
    .C(_03673_),
    .A(_03671_),
    .Y(_03675_),
    .D(_03674_));
 sg13g2_nor3_2 _17903_ (.A(_03666_),
    .B(_03670_),
    .C(_03675_),
    .Y(_03676_));
 sg13g2_a21oi_1 _17904_ (.A1(net488),
    .A2(net5103),
    .Y(_03677_),
    .B1(net5292));
 sg13g2_or2_1 _17905_ (.X(_03678_),
    .B(_03677_),
    .A(_03676_));
 sg13g2_o21ai_1 _17906_ (.B1(_03678_),
    .Y(_01064_),
    .A1(net6144),
    .A2(_08055_));
 sg13g2_and2_1 _17907_ (.A(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .B(net5839),
    .X(_03679_));
 sg13g2_a22oi_1 _17908_ (.Y(_03680_),
    .B1(net5476),
    .B2(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .A2(net5854),
    .A1(\soc_inst.cpu_core.register_file.registers[12][9] ));
 sg13g2_a22oi_1 _17909_ (.Y(_03681_),
    .B1(net5280),
    .B2(\soc_inst.cpu_core.register_file.registers[20][9] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][9] ));
 sg13g2_a22oi_1 _17910_ (.Y(_03682_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][9] ),
    .A2(net5480),
    .A1(\soc_inst.cpu_core.register_file.registers[5][9] ));
 sg13g2_a22oi_1 _17911_ (.Y(_03683_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .A2(net5819),
    .A1(\soc_inst.cpu_core.register_file.registers[8][9] ));
 sg13g2_a22oi_1 _17912_ (.Y(_03684_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][9] ));
 sg13g2_a22oi_1 _17913_ (.Y(_03685_),
    .B1(net5265),
    .B2(\soc_inst.cpu_core.register_file.registers[29][9] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][9] ));
 sg13g2_nand3_1 _17914_ (.B(_03684_),
    .C(_03685_),
    .A(_03683_),
    .Y(_03686_));
 sg13g2_a221oi_1 _17915_ (.B2(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .C1(_03686_),
    .B1(net5794),
    .A1(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .Y(_03687_),
    .A2(net5850));
 sg13g2_a22oi_1 _17916_ (.Y(_03688_),
    .B1(net5830),
    .B2(\soc_inst.cpu_core.register_file.registers[30][9] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][9] ));
 sg13g2_a22oi_1 _17917_ (.Y(_03689_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .A2(net5845),
    .A1(\soc_inst.cpu_core.register_file.registers[26][9] ));
 sg13g2_a221oi_1 _17918_ (.B2(\soc_inst.cpu_core.register_file.registers[24][9] ),
    .C1(_03679_),
    .B1(net5254),
    .A1(\soc_inst.cpu_core.register_file.registers[27][9] ),
    .Y(_03690_),
    .A2(net5810));
 sg13g2_nand4_1 _17919_ (.B(_03688_),
    .C(_03689_),
    .A(_03687_),
    .Y(_03691_),
    .D(_03690_));
 sg13g2_a21oi_1 _17920_ (.A1(\soc_inst.cpu_core.register_file.registers[23][9] ),
    .A2(net5864),
    .Y(_03692_),
    .B1(net6079));
 sg13g2_a22oi_1 _17921_ (.Y(_03693_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][9] ),
    .A2(net5290),
    .A1(\soc_inst.cpu_core.register_file.registers[25][9] ));
 sg13g2_a22oi_1 _17922_ (.Y(_03694_),
    .B1(net5273),
    .B2(\soc_inst.cpu_core.register_file.registers[17][9] ),
    .A2(net5824),
    .A1(\soc_inst.cpu_core.register_file.registers[18][9] ));
 sg13g2_nand4_1 _17923_ (.B(_03692_),
    .C(_03693_),
    .A(_03680_),
    .Y(_03695_),
    .D(_03694_));
 sg13g2_a22oi_1 _17924_ (.Y(_03696_),
    .B1(net5814),
    .B2(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .A2(net5875),
    .A1(\soc_inst.cpu_core.register_file.registers[4][9] ));
 sg13g2_a22oi_1 _17925_ (.Y(_03697_),
    .B1(net5799),
    .B2(\soc_inst.cpu_core.register_file.registers[22][9] ),
    .A2(net5804),
    .A1(\soc_inst.cpu_core.register_file.registers[15][9] ));
 sg13g2_nand4_1 _17926_ (.B(_03682_),
    .C(_03696_),
    .A(_03681_),
    .Y(_03698_),
    .D(_03697_));
 sg13g2_nor3_2 _17927_ (.A(_03691_),
    .B(_03695_),
    .C(_03698_),
    .Y(_03699_));
 sg13g2_a21oi_1 _17928_ (.A1(net673),
    .A2(net5103),
    .Y(_03700_),
    .B1(net5292));
 sg13g2_or2_1 _17929_ (.X(_03701_),
    .B(_03700_),
    .A(_03699_));
 sg13g2_o21ai_1 _17930_ (.B1(_03701_),
    .Y(_01065_),
    .A1(net6148),
    .A2(_08053_));
 sg13g2_and2_1 _17931_ (.A(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .B(net5854),
    .X(_03702_));
 sg13g2_a22oi_1 _17932_ (.Y(_03703_),
    .B1(net5849),
    .B2(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][10] ));
 sg13g2_a22oi_1 _17933_ (.Y(_03704_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .A2(net5804),
    .A1(\soc_inst.cpu_core.register_file.registers[15][10] ));
 sg13g2_a22oi_1 _17934_ (.Y(_03705_),
    .B1(net5819),
    .B2(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .A2(net5844),
    .A1(\soc_inst.cpu_core.register_file.registers[26][10] ));
 sg13g2_a22oi_1 _17935_ (.Y(_03706_),
    .B1(net5809),
    .B2(\soc_inst.cpu_core.register_file.registers[27][10] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][10] ));
 sg13g2_nand3_1 _17936_ (.B(_03705_),
    .C(_03706_),
    .A(_03704_),
    .Y(_03707_));
 sg13g2_a221oi_1 _17937_ (.B2(\soc_inst.cpu_core.register_file.registers[22][10] ),
    .C1(_03707_),
    .B1(net5799),
    .A1(\soc_inst.cpu_core.register_file.registers[23][10] ),
    .Y(_03708_),
    .A2(net5864));
 sg13g2_a22oi_1 _17938_ (.Y(_03709_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .A2(net5839),
    .A1(\soc_inst.cpu_core.register_file.registers[10][10] ));
 sg13g2_a22oi_1 _17939_ (.Y(_03710_),
    .B1(net5264),
    .B2(\soc_inst.cpu_core.register_file.registers[29][10] ),
    .A2(net5480),
    .A1(\soc_inst.cpu_core.register_file.registers[5][10] ));
 sg13g2_a221oi_1 _17940_ (.B2(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .C1(_03702_),
    .B1(net5794),
    .A1(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .Y(_03711_),
    .A2(net5475));
 sg13g2_nand4_1 _17941_ (.B(_03709_),
    .C(_03710_),
    .A(_03708_),
    .Y(_03712_),
    .D(_03711_));
 sg13g2_a21oi_1 _17942_ (.A1(\soc_inst.cpu_core.register_file.registers[17][10] ),
    .A2(net5273),
    .Y(_03713_),
    .B1(net6079));
 sg13g2_a22oi_1 _17943_ (.Y(_03714_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][10] ),
    .A2(net5289),
    .A1(\soc_inst.cpu_core.register_file.registers[25][10] ));
 sg13g2_a22oi_1 _17944_ (.Y(_03715_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][10] ),
    .A2(net5829),
    .A1(\soc_inst.cpu_core.register_file.registers[30][10] ));
 sg13g2_nand4_1 _17945_ (.B(_03713_),
    .C(_03714_),
    .A(_03703_),
    .Y(_03716_),
    .D(_03715_));
 sg13g2_a22oi_1 _17946_ (.Y(_03717_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][10] ),
    .A2(net5279),
    .A1(\soc_inst.cpu_core.register_file.registers[20][10] ));
 sg13g2_a22oi_1 _17947_ (.Y(_03718_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][10] ));
 sg13g2_a22oi_1 _17948_ (.Y(_03719_),
    .B1(net5814),
    .B2(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .A2(net5874),
    .A1(\soc_inst.cpu_core.register_file.registers[4][10] ));
 sg13g2_a22oi_1 _17949_ (.Y(_03720_),
    .B1(net5824),
    .B2(\soc_inst.cpu_core.register_file.registers[18][10] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][10] ));
 sg13g2_nand4_1 _17950_ (.B(_03718_),
    .C(_03719_),
    .A(_03717_),
    .Y(_03721_),
    .D(_03720_));
 sg13g2_nor3_2 _17951_ (.A(_03712_),
    .B(_03716_),
    .C(_03721_),
    .Y(_03722_));
 sg13g2_a21oi_1 _17952_ (.A1(net684),
    .A2(net5103),
    .Y(_03723_),
    .B1(net5292));
 sg13g2_or2_1 _17953_ (.X(_03724_),
    .B(_03723_),
    .A(_03722_));
 sg13g2_o21ai_1 _17954_ (.B1(_03724_),
    .Y(_01066_),
    .A1(net6148),
    .A2(_08051_));
 sg13g2_a21oi_1 _17955_ (.A1(net991),
    .A2(net5105),
    .Y(_03725_),
    .B1(net5292));
 sg13g2_nand2_1 _17956_ (.Y(_03726_),
    .A(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .B(net5872));
 sg13g2_a22oi_1 _17957_ (.Y(_03727_),
    .B1(net5842),
    .B2(\soc_inst.cpu_core.register_file.registers[26][11] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][11] ));
 sg13g2_a22oi_1 _17958_ (.Y(_03728_),
    .B1(net5262),
    .B2(\soc_inst.cpu_core.register_file.registers[29][11] ),
    .A2(net5473),
    .A1(\soc_inst.cpu_core.register_file.registers[9][11] ));
 sg13g2_a22oi_1 _17959_ (.Y(_03729_),
    .B1(net5478),
    .B2(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][11] ));
 sg13g2_a22oi_1 _17960_ (.Y(_03730_),
    .B1(net5257),
    .B2(\soc_inst.cpu_core.register_file.registers[28][11] ),
    .A2(net5817),
    .A1(\soc_inst.cpu_core.register_file.registers[8][11] ));
 sg13g2_a22oi_1 _17961_ (.Y(_03731_),
    .B1(net5837),
    .B2(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][11] ));
 sg13g2_a22oi_1 _17962_ (.Y(_03732_),
    .B1(net5277),
    .B2(\soc_inst.cpu_core.register_file.registers[20][11] ),
    .A2(net5852),
    .A1(\soc_inst.cpu_core.register_file.registers[12][11] ));
 sg13g2_nand4_1 _17963_ (.B(_03730_),
    .C(_03731_),
    .A(_03728_),
    .Y(_03733_),
    .D(_03732_));
 sg13g2_a22oi_1 _17964_ (.Y(_03734_),
    .B1(net5797),
    .B2(\soc_inst.cpu_core.register_file.registers[22][11] ),
    .A2(net5267),
    .A1(\soc_inst.cpu_core.register_file.registers[21][11] ));
 sg13g2_a22oi_1 _17965_ (.Y(_03735_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .A2(net5822),
    .A1(\soc_inst.cpu_core.register_file.registers[18][11] ));
 sg13g2_nand4_1 _17966_ (.B(_03727_),
    .C(_03734_),
    .A(_03726_),
    .Y(_03736_),
    .D(_03735_));
 sg13g2_nor2_1 _17967_ (.A(_03733_),
    .B(_03736_),
    .Y(_03737_));
 sg13g2_a21oi_1 _17968_ (.A1(\soc_inst.cpu_core.register_file.registers[19][11] ),
    .A2(net5857),
    .Y(_03738_),
    .B1(net6077));
 sg13g2_a22oi_1 _17969_ (.Y(_03739_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .A2(net5272),
    .A1(\soc_inst.cpu_core.register_file.registers[17][11] ));
 sg13g2_a22oi_1 _17970_ (.Y(_03740_),
    .B1(net5807),
    .B2(\soc_inst.cpu_core.register_file.registers[27][11] ),
    .A2(net5867),
    .A1(\soc_inst.cpu_core.register_file.registers[31][11] ));
 sg13g2_nand4_1 _17971_ (.B(_03738_),
    .C(_03739_),
    .A(_03729_),
    .Y(_03741_),
    .D(_03740_));
 sg13g2_a22oi_1 _17972_ (.Y(_03742_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .A2(net5812),
    .A1(\soc_inst.cpu_core.register_file.registers[11][11] ));
 sg13g2_a22oi_1 _17973_ (.Y(_03743_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .A2(net5847),
    .A1(\soc_inst.cpu_core.register_file.registers[2][11] ));
 sg13g2_a22oi_1 _17974_ (.Y(_03744_),
    .B1(net5827),
    .B2(\soc_inst.cpu_core.register_file.registers[30][11] ),
    .A2(net5832),
    .A1(\soc_inst.cpu_core.register_file.registers[14][11] ));
 sg13g2_a22oi_1 _17975_ (.Y(_03745_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][11] ),
    .A2(net5792),
    .A1(\soc_inst.cpu_core.register_file.registers[6][11] ));
 sg13g2_nand4_1 _17976_ (.B(_03743_),
    .C(_03744_),
    .A(_03742_),
    .Y(_03746_),
    .D(_03745_));
 sg13g2_nor2_1 _17977_ (.A(_03741_),
    .B(_03746_),
    .Y(_03747_));
 sg13g2_a21oi_2 _17978_ (.B1(_03725_),
    .Y(_03748_),
    .A2(_03747_),
    .A1(_03737_));
 sg13g2_a21o_1 _17979_ (.A2(net1726),
    .A1(net6419),
    .B1(_03748_),
    .X(_01067_));
 sg13g2_and2_1 _17980_ (.A(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .B(net5848),
    .X(_03749_));
 sg13g2_a22oi_1 _17981_ (.Y(_03750_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][12] ));
 sg13g2_a22oi_1 _17982_ (.Y(_03751_),
    .B1(net5793),
    .B2(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .A2(net5479),
    .A1(\soc_inst.cpu_core.register_file.registers[5][12] ));
 sg13g2_a22oi_1 _17983_ (.Y(_03752_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][12] ),
    .A2(net5274),
    .A1(\soc_inst.cpu_core.register_file.registers[17][12] ));
 sg13g2_a22oi_1 _17984_ (.Y(_03753_),
    .B1(net5278),
    .B2(\soc_inst.cpu_core.register_file.registers[20][12] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][12] ));
 sg13g2_a22oi_1 _17985_ (.Y(_03754_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][12] ));
 sg13g2_nand3_1 _17986_ (.B(_03753_),
    .C(_03754_),
    .A(_03752_),
    .Y(_03755_));
 sg13g2_a221oi_1 _17987_ (.B2(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .C1(_03755_),
    .B1(net5803),
    .A1(\soc_inst.cpu_core.register_file.registers[16][12] ),
    .Y(_03756_),
    .A2(net5283));
 sg13g2_a22oi_1 _17988_ (.Y(_03757_),
    .B1(net5813),
    .B2(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .A2(net5874),
    .A1(\soc_inst.cpu_core.register_file.registers[4][12] ));
 sg13g2_a22oi_1 _17989_ (.Y(_03758_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][12] ),
    .A2(net5828),
    .A1(\soc_inst.cpu_core.register_file.registers[30][12] ));
 sg13g2_a221oi_1 _17990_ (.B2(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .C1(_03749_),
    .B1(net5788),
    .A1(\soc_inst.cpu_core.register_file.registers[26][12] ),
    .Y(_03759_),
    .A2(net5844));
 sg13g2_nand4_1 _17991_ (.B(_03757_),
    .C(_03758_),
    .A(_03756_),
    .Y(_03760_),
    .D(_03759_));
 sg13g2_a21oi_1 _17992_ (.A1(\soc_inst.cpu_core.register_file.registers[23][12] ),
    .A2(net5863),
    .Y(_03761_),
    .B1(net6078));
 sg13g2_a22oi_1 _17993_ (.Y(_03762_),
    .B1(net5469),
    .B2(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][12] ));
 sg13g2_nand4_1 _17994_ (.B(_03751_),
    .C(_03761_),
    .A(_03750_),
    .Y(_03763_),
    .D(_03762_));
 sg13g2_a22oi_1 _17995_ (.Y(_03764_),
    .B1(net5474),
    .B2(\soc_inst.cpu_core.register_file.registers[9][12] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][12] ));
 sg13g2_a22oi_1 _17996_ (.Y(_03765_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][12] ),
    .A2(net5268),
    .A1(\soc_inst.cpu_core.register_file.registers[21][12] ));
 sg13g2_a22oi_1 _17997_ (.Y(_03766_),
    .B1(net5823),
    .B2(\soc_inst.cpu_core.register_file.registers[18][12] ),
    .A2(net5838),
    .A1(\soc_inst.cpu_core.register_file.registers[10][12] ));
 sg13g2_a22oi_1 _17998_ (.Y(_03767_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][12] ),
    .A2(net5258),
    .A1(\soc_inst.cpu_core.register_file.registers[28][12] ));
 sg13g2_nand4_1 _17999_ (.B(_03765_),
    .C(_03766_),
    .A(_03764_),
    .Y(_03768_),
    .D(_03767_));
 sg13g2_nor3_2 _18000_ (.A(_03760_),
    .B(_03763_),
    .C(_03768_),
    .Y(_03769_));
 sg13g2_a21oi_1 _18001_ (.A1(net479),
    .A2(net5104),
    .Y(_03770_),
    .B1(net5291));
 sg13g2_or2_1 _18002_ (.X(_03771_),
    .B(_03770_),
    .A(_03769_));
 sg13g2_o21ai_1 _18003_ (.B1(_03771_),
    .Y(_01068_),
    .A1(net6143),
    .A2(_08048_));
 sg13g2_a22oi_1 _18004_ (.Y(_03772_),
    .B1(net5480),
    .B2(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][13] ));
 sg13g2_and2_1 _18005_ (.A(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .B(net5474),
    .X(_03773_));
 sg13g2_a22oi_1 _18006_ (.Y(_03774_),
    .B1(net5799),
    .B2(\soc_inst.cpu_core.register_file.registers[22][13] ),
    .A2(net5824),
    .A1(\soc_inst.cpu_core.register_file.registers[18][13] ));
 sg13g2_a22oi_1 _18007_ (.Y(_03775_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .A2(net5863),
    .A1(\soc_inst.cpu_core.register_file.registers[23][13] ));
 sg13g2_a22oi_1 _18008_ (.Y(_03776_),
    .B1(net5803),
    .B2(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][13] ));
 sg13g2_a22oi_1 _18009_ (.Y(_03777_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][13] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][13] ));
 sg13g2_nand3_1 _18010_ (.B(_03776_),
    .C(_03777_),
    .A(_03775_),
    .Y(_03778_));
 sg13g2_a221oi_1 _18011_ (.B2(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .C1(_03778_),
    .B1(net5838),
    .A1(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .Y(_03779_),
    .A2(net5848));
 sg13g2_a22oi_1 _18012_ (.Y(_03780_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][13] ));
 sg13g2_a221oi_1 _18013_ (.B2(\soc_inst.cpu_core.register_file.registers[29][13] ),
    .C1(_03773_),
    .B1(net5264),
    .A1(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .Y(_03781_),
    .A2(net5469));
 sg13g2_nand4_1 _18014_ (.B(_03779_),
    .C(_03780_),
    .A(_03772_),
    .Y(_03782_),
    .D(_03781_));
 sg13g2_a21oi_1 _18015_ (.A1(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .A2(net5814),
    .Y(_03783_),
    .B1(net6078));
 sg13g2_a22oi_1 _18016_ (.Y(_03784_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .A2(net5274),
    .A1(\soc_inst.cpu_core.register_file.registers[17][13] ));
 sg13g2_a22oi_1 _18017_ (.Y(_03785_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][13] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][13] ));
 sg13g2_nand4_1 _18018_ (.B(_03783_),
    .C(_03784_),
    .A(_03774_),
    .Y(_03786_),
    .D(_03785_));
 sg13g2_a22oi_1 _18019_ (.Y(_03787_),
    .B1(net5258),
    .B2(\soc_inst.cpu_core.register_file.registers[28][13] ),
    .A2(net5793),
    .A1(\soc_inst.cpu_core.register_file.registers[6][13] ));
 sg13g2_a22oi_1 _18020_ (.Y(_03788_),
    .B1(net5279),
    .B2(\soc_inst.cpu_core.register_file.registers[20][13] ),
    .A2(net5854),
    .A1(\soc_inst.cpu_core.register_file.registers[12][13] ));
 sg13g2_a22oi_1 _18021_ (.Y(_03789_),
    .B1(net5809),
    .B2(\soc_inst.cpu_core.register_file.registers[27][13] ),
    .A2(net5843),
    .A1(\soc_inst.cpu_core.register_file.registers[26][13] ));
 sg13g2_a22oi_1 _18022_ (.Y(_03790_),
    .B1(net5829),
    .B2(\soc_inst.cpu_core.register_file.registers[30][13] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][13] ));
 sg13g2_nand4_1 _18023_ (.B(_03788_),
    .C(_03789_),
    .A(_03787_),
    .Y(_03791_),
    .D(_03790_));
 sg13g2_nor3_2 _18024_ (.A(_03782_),
    .B(_03786_),
    .C(_03791_),
    .Y(_03792_));
 sg13g2_a21oi_1 _18025_ (.A1(net808),
    .A2(net5102),
    .Y(_03793_),
    .B1(net5291));
 sg13g2_or2_1 _18026_ (.X(_03794_),
    .B(_03793_),
    .A(_03792_));
 sg13g2_o21ai_1 _18027_ (.B1(_03794_),
    .Y(_01069_),
    .A1(net6144),
    .A2(_08046_));
 sg13g2_a22oi_1 _18028_ (.Y(_03795_),
    .B1(net5786),
    .B2(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][14] ));
 sg13g2_and2_1 _18029_ (.A(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .B(net5467),
    .X(_03796_));
 sg13g2_a22oi_1 _18030_ (.Y(_03797_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .A2(net5276),
    .A1(\soc_inst.cpu_core.register_file.registers[20][14] ));
 sg13g2_a22oi_1 _18031_ (.Y(_03798_),
    .B1(net5846),
    .B2(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][14] ));
 sg13g2_a22oi_1 _18032_ (.Y(_03799_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][14] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][14] ));
 sg13g2_a22oi_1 _18033_ (.Y(_03800_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .A2(net5831),
    .A1(\soc_inst.cpu_core.register_file.registers[14][14] ));
 sg13g2_nand3_1 _18034_ (.B(_03799_),
    .C(_03800_),
    .A(_03798_),
    .Y(_03801_));
 sg13g2_a221oi_1 _18035_ (.B2(\soc_inst.cpu_core.register_file.registers[27][14] ),
    .C1(_03801_),
    .B1(net5806),
    .A1(\soc_inst.cpu_core.register_file.registers[23][14] ),
    .Y(_03802_),
    .A2(net5861));
 sg13g2_a22oi_1 _18036_ (.Y(_03803_),
    .B1(net5816),
    .B2(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .A2(net5841),
    .A1(\soc_inst.cpu_core.register_file.registers[26][14] ));
 sg13g2_a22oi_1 _18037_ (.Y(_03804_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][14] ));
 sg13g2_a221oi_1 _18038_ (.B2(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .C1(_03796_),
    .B1(net5801),
    .A1(\soc_inst.cpu_core.register_file.registers[25][14] ),
    .Y(_03805_),
    .A2(net5286));
 sg13g2_nand4_1 _18039_ (.B(_03803_),
    .C(_03804_),
    .A(_03802_),
    .Y(_03806_),
    .D(_03805_));
 sg13g2_a21oi_1 _18040_ (.A1(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .A2(net5871),
    .Y(_03807_),
    .B1(net6076));
 sg13g2_a22oi_1 _18041_ (.Y(_03808_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][14] ),
    .A2(net5851),
    .A1(\soc_inst.cpu_core.register_file.registers[12][14] ));
 sg13g2_a22oi_1 _18042_ (.Y(_03809_),
    .B1(net5271),
    .B2(\soc_inst.cpu_core.register_file.registers[17][14] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][14] ));
 sg13g2_nand4_1 _18043_ (.B(_03807_),
    .C(_03808_),
    .A(_03797_),
    .Y(_03810_),
    .D(_03809_));
 sg13g2_a22oi_1 _18044_ (.Y(_03811_),
    .B1(net5821),
    .B2(\soc_inst.cpu_core.register_file.registers[18][14] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][14] ));
 sg13g2_a22oi_1 _18045_ (.Y(_03812_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .A2(net5261),
    .A1(\soc_inst.cpu_core.register_file.registers[29][14] ));
 sg13g2_a22oi_1 _18046_ (.Y(_03813_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][14] ),
    .A2(net5266),
    .A1(\soc_inst.cpu_core.register_file.registers[21][14] ));
 sg13g2_nand4_1 _18047_ (.B(_03811_),
    .C(_03812_),
    .A(_03795_),
    .Y(_03814_),
    .D(_03813_));
 sg13g2_nor3_1 _18048_ (.A(_03806_),
    .B(_03810_),
    .C(_03814_),
    .Y(_03815_));
 sg13g2_a21oi_1 _18049_ (.A1(net839),
    .A2(net5102),
    .Y(_03816_),
    .B1(net5291));
 sg13g2_or2_1 _18050_ (.X(_03817_),
    .B(_03816_),
    .A(_03815_));
 sg13g2_o21ai_1 _18051_ (.B1(_03817_),
    .Y(_01070_),
    .A1(net6143),
    .A2(_08044_));
 sg13g2_and2_1 _18052_ (.A(\soc_inst.cpu_core.register_file.registers[31][15] ),
    .B(net5868),
    .X(_03818_));
 sg13g2_a22oi_1 _18053_ (.Y(_03819_),
    .B1(net5813),
    .B2(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][15] ));
 sg13g2_a22oi_1 _18054_ (.Y(_03820_),
    .B1(net5828),
    .B2(\soc_inst.cpu_core.register_file.registers[30][15] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][15] ));
 sg13g2_a22oi_1 _18055_ (.Y(_03821_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][15] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][15] ));
 sg13g2_a22oi_1 _18056_ (.Y(_03822_),
    .B1(net5474),
    .B2(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .A2(net5863),
    .A1(\soc_inst.cpu_core.register_file.registers[23][15] ));
 sg13g2_nand3_1 _18057_ (.B(_03821_),
    .C(_03822_),
    .A(_03820_),
    .Y(_03823_));
 sg13g2_a221oi_1 _18058_ (.B2(\soc_inst.cpu_core.register_file.registers[29][15] ),
    .C1(_03823_),
    .B1(net5263),
    .A1(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .Y(_03824_),
    .A2(net5848));
 sg13g2_a22oi_1 _18059_ (.Y(_03825_),
    .B1(net5803),
    .B2(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .A2(net5818),
    .A1(\soc_inst.cpu_core.register_file.registers[8][15] ));
 sg13g2_a22oi_1 _18060_ (.Y(_03826_),
    .B1(net5788),
    .B2(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .A2(net5258),
    .A1(\soc_inst.cpu_core.register_file.registers[28][15] ));
 sg13g2_a221oi_1 _18061_ (.B2(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .C1(_03818_),
    .B1(net5793),
    .A1(\soc_inst.cpu_core.register_file.registers[17][15] ),
    .Y(_03827_),
    .A2(net5274));
 sg13g2_nand4_1 _18062_ (.B(_03825_),
    .C(_03826_),
    .A(_03824_),
    .Y(_03828_),
    .D(_03827_));
 sg13g2_a21oi_1 _18063_ (.A1(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .A2(net5873),
    .Y(_03829_),
    .B1(net6078));
 sg13g2_a22oi_1 _18064_ (.Y(_03830_),
    .B1(net5838),
    .B2(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][15] ));
 sg13g2_a22oi_1 _18065_ (.Y(_03831_),
    .B1(net5469),
    .B2(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .A2(net5843),
    .A1(\soc_inst.cpu_core.register_file.registers[26][15] ));
 sg13g2_nand4_1 _18066_ (.B(_03829_),
    .C(_03830_),
    .A(_03819_),
    .Y(_03832_),
    .D(_03831_));
 sg13g2_a22oi_1 _18067_ (.Y(_03833_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][15] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][15] ));
 sg13g2_a22oi_1 _18068_ (.Y(_03834_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][15] ),
    .A2(net5479),
    .A1(\soc_inst.cpu_core.register_file.registers[5][15] ));
 sg13g2_a22oi_1 _18069_ (.Y(_03835_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .A2(net5808),
    .A1(\soc_inst.cpu_core.register_file.registers[27][15] ));
 sg13g2_a22oi_1 _18070_ (.Y(_03836_),
    .B1(net5278),
    .B2(\soc_inst.cpu_core.register_file.registers[20][15] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][15] ));
 sg13g2_nand4_1 _18071_ (.B(_03834_),
    .C(_03835_),
    .A(_03833_),
    .Y(_03837_),
    .D(_03836_));
 sg13g2_nor3_2 _18072_ (.A(_03828_),
    .B(_03832_),
    .C(_03837_),
    .Y(_03838_));
 sg13g2_a21oi_1 _18073_ (.A1(net641),
    .A2(net5102),
    .Y(_03839_),
    .B1(net5291));
 sg13g2_or2_1 _18074_ (.X(_03840_),
    .B(_03839_),
    .A(_03838_));
 sg13g2_o21ai_1 _18075_ (.B1(_03840_),
    .Y(_01071_),
    .A1(net6144),
    .A2(_08042_));
 sg13g2_and2_1 _18076_ (.A(\soc_inst.cpu_core.register_file.registers[23][16] ),
    .B(net5863),
    .X(_03841_));
 sg13g2_a22oi_1 _18077_ (.Y(_03842_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][16] ),
    .A2(net5839),
    .A1(\soc_inst.cpu_core.register_file.registers[10][16] ));
 sg13g2_a22oi_1 _18078_ (.Y(_03843_),
    .B1(net5828),
    .B2(\soc_inst.cpu_core.register_file.registers[30][16] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][16] ));
 sg13g2_a22oi_1 _18079_ (.Y(_03844_),
    .B1(net5474),
    .B2(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .A2(net5274),
    .A1(\soc_inst.cpu_core.register_file.registers[17][16] ));
 sg13g2_a22oi_1 _18080_ (.Y(_03845_),
    .B1(net5793),
    .B2(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .A2(net5278),
    .A1(\soc_inst.cpu_core.register_file.registers[20][16] ));
 sg13g2_nand3_1 _18081_ (.B(_03844_),
    .C(_03845_),
    .A(_03843_),
    .Y(_03846_));
 sg13g2_a221oi_1 _18082_ (.B2(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .C1(_03846_),
    .B1(net5469),
    .A1(\soc_inst.cpu_core.register_file.registers[31][16] ),
    .Y(_03847_),
    .A2(net5868));
 sg13g2_a22oi_1 _18083_ (.Y(_03848_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][16] ));
 sg13g2_a22oi_1 _18084_ (.Y(_03849_),
    .B1(net5258),
    .B2(\soc_inst.cpu_core.register_file.registers[28][16] ),
    .A2(net5263),
    .A1(\soc_inst.cpu_core.register_file.registers[29][16] ));
 sg13g2_a221oi_1 _18085_ (.B2(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .C1(_03841_),
    .B1(net5784),
    .A1(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .Y(_03850_),
    .A2(net5479));
 sg13g2_nand4_1 _18086_ (.B(_03848_),
    .C(_03849_),
    .A(_03847_),
    .Y(_03851_),
    .D(_03850_));
 sg13g2_a21oi_1 _18087_ (.A1(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .A2(net5788),
    .Y(_03852_),
    .B1(net6080));
 sg13g2_a22oi_1 _18088_ (.Y(_03853_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][16] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][16] ));
 sg13g2_a22oi_1 _18089_ (.Y(_03854_),
    .B1(net5834),
    .B2(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .A2(net5848),
    .A1(\soc_inst.cpu_core.register_file.registers[2][16] ));
 sg13g2_nand4_1 _18090_ (.B(_03852_),
    .C(_03853_),
    .A(_03842_),
    .Y(_03855_),
    .D(_03854_));
 sg13g2_a22oi_1 _18091_ (.Y(_03856_),
    .B1(net5843),
    .B2(\soc_inst.cpu_core.register_file.registers[26][16] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][16] ));
 sg13g2_a22oi_1 _18092_ (.Y(_03857_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][16] ),
    .A2(net5803),
    .A1(\soc_inst.cpu_core.register_file.registers[15][16] ));
 sg13g2_a22oi_1 _18093_ (.Y(_03858_),
    .B1(net5813),
    .B2(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][16] ));
 sg13g2_a22oi_1 _18094_ (.Y(_03859_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][16] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][16] ));
 sg13g2_nand4_1 _18095_ (.B(_03857_),
    .C(_03858_),
    .A(_03856_),
    .Y(_03860_),
    .D(_03859_));
 sg13g2_nor3_2 _18096_ (.A(_03851_),
    .B(_03855_),
    .C(_03860_),
    .Y(_03861_));
 sg13g2_a21oi_1 _18097_ (.A1(net1734),
    .A2(net5102),
    .Y(_03862_),
    .B1(net5291));
 sg13g2_or2_1 _18098_ (.X(_03863_),
    .B(_03862_),
    .A(_03861_));
 sg13g2_o21ai_1 _18099_ (.B1(_03863_),
    .Y(_01072_),
    .A1(net6150),
    .A2(_08081_));
 sg13g2_and2_1 _18100_ (.A(\soc_inst.cpu_core.register_file.registers[22][17] ),
    .B(net5796),
    .X(_03864_));
 sg13g2_a22oi_1 _18101_ (.Y(_03865_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][17] ));
 sg13g2_a22oi_1 _18102_ (.Y(_03866_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][17] ),
    .A2(net5831),
    .A1(\soc_inst.cpu_core.register_file.registers[14][17] ));
 sg13g2_a22oi_1 _18103_ (.Y(_03867_),
    .B1(net5786),
    .B2(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][17] ));
 sg13g2_a22oi_1 _18104_ (.Y(_03868_),
    .B1(net5276),
    .B2(\soc_inst.cpu_core.register_file.registers[20][17] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][17] ));
 sg13g2_a22oi_1 _18105_ (.Y(_03869_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][17] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][17] ));
 sg13g2_a22oi_1 _18106_ (.Y(_03870_),
    .B1(net5806),
    .B2(\soc_inst.cpu_core.register_file.registers[27][17] ),
    .A2(net5841),
    .A1(\soc_inst.cpu_core.register_file.registers[26][17] ));
 sg13g2_nand3_1 _18107_ (.B(_03869_),
    .C(_03870_),
    .A(_03868_),
    .Y(_03871_));
 sg13g2_a221oi_1 _18108_ (.B2(\soc_inst.cpu_core.register_file.registers[17][17] ),
    .C1(_03871_),
    .B1(net5271),
    .A1(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .Y(_03872_),
    .A2(net5871));
 sg13g2_a22oi_1 _18109_ (.Y(_03873_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .A2(net5811),
    .A1(\soc_inst.cpu_core.register_file.registers[11][17] ));
 sg13g2_a22oi_1 _18110_ (.Y(_03874_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .A2(net5846),
    .A1(\soc_inst.cpu_core.register_file.registers[2][17] ));
 sg13g2_a221oi_1 _18111_ (.B2(\soc_inst.cpu_core.register_file.registers[21][17] ),
    .C1(_03864_),
    .B1(net5266),
    .A1(\soc_inst.cpu_core.register_file.registers[18][17] ),
    .Y(_03875_),
    .A2(net5821));
 sg13g2_nand4_1 _18112_ (.B(_03873_),
    .C(_03874_),
    .A(_03872_),
    .Y(_03876_),
    .D(_03875_));
 sg13g2_a21oi_1 _18113_ (.A1(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .A2(net5467),
    .Y(_03877_),
    .B1(net6076));
 sg13g2_a22oi_1 _18114_ (.Y(_03878_),
    .B1(net5856),
    .B2(\soc_inst.cpu_core.register_file.registers[19][17] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][17] ));
 sg13g2_a22oi_1 _18115_ (.Y(_03879_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .A2(net5816),
    .A1(\soc_inst.cpu_core.register_file.registers[8][17] ));
 sg13g2_nand4_1 _18116_ (.B(_03877_),
    .C(_03878_),
    .A(_03865_),
    .Y(_03880_),
    .D(_03879_));
 sg13g2_a22oi_1 _18117_ (.Y(_03881_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][17] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][17] ));
 sg13g2_a22oi_1 _18118_ (.Y(_03882_),
    .B1(net5851),
    .B2(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][17] ));
 sg13g2_nand4_1 _18119_ (.B(_03867_),
    .C(_03881_),
    .A(_03866_),
    .Y(_03883_),
    .D(_03882_));
 sg13g2_nor3_2 _18120_ (.A(_03876_),
    .B(_03880_),
    .C(_03883_),
    .Y(_03884_));
 sg13g2_a21oi_1 _18121_ (.A1(net1196),
    .A2(net5105),
    .Y(_03885_),
    .B1(net5294));
 sg13g2_or2_1 _18122_ (.X(_03886_),
    .B(_03885_),
    .A(_03884_));
 sg13g2_o21ai_1 _18123_ (.B1(_03886_),
    .Y(_01073_),
    .A1(net6146),
    .A2(_08079_));
 sg13g2_a22oi_1 _18124_ (.Y(_03887_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][18] ),
    .A2(net5813),
    .A1(\soc_inst.cpu_core.register_file.registers[11][18] ));
 sg13g2_and2_1 _18125_ (.A(\soc_inst.cpu_core.register_file.registers[19][18] ),
    .B(net5859),
    .X(_03888_));
 sg13g2_a22oi_1 _18126_ (.Y(_03889_),
    .B1(net5804),
    .B2(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][18] ));
 sg13g2_a22oi_1 _18127_ (.Y(_03890_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][18] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][18] ));
 sg13g2_a22oi_1 _18128_ (.Y(_03891_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][18] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][18] ));
 sg13g2_a22oi_1 _18129_ (.Y(_03892_),
    .B1(net5819),
    .B2(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][18] ));
 sg13g2_a22oi_1 _18130_ (.Y(_03893_),
    .B1(net5274),
    .B2(\soc_inst.cpu_core.register_file.registers[17][18] ),
    .A2(net5479),
    .A1(\soc_inst.cpu_core.register_file.registers[5][18] ));
 sg13g2_nand3_1 _18131_ (.B(_03892_),
    .C(_03893_),
    .A(_03891_),
    .Y(_03894_));
 sg13g2_a221oi_1 _18132_ (.B2(\soc_inst.cpu_core.register_file.registers[30][18] ),
    .C1(_03894_),
    .B1(net5828),
    .A1(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .Y(_03895_),
    .A2(net5849));
 sg13g2_a22oi_1 _18133_ (.Y(_03896_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][18] ),
    .A2(net5469),
    .A1(\soc_inst.cpu_core.register_file.registers[13][18] ));
 sg13g2_a22oi_1 _18134_ (.Y(_03897_),
    .B1(net5793),
    .B2(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .A2(net5798),
    .A1(\soc_inst.cpu_core.register_file.registers[22][18] ));
 sg13g2_a221oi_1 _18135_ (.B2(\soc_inst.cpu_core.register_file.registers[20][18] ),
    .C1(_03888_),
    .B1(net5278),
    .A1(\soc_inst.cpu_core.register_file.registers[25][18] ),
    .Y(_03898_),
    .A2(net5289));
 sg13g2_nand4_1 _18136_ (.B(_03896_),
    .C(_03897_),
    .A(_03895_),
    .Y(_03899_),
    .D(_03898_));
 sg13g2_a21oi_1 _18137_ (.A1(\soc_inst.cpu_core.register_file.registers[26][18] ),
    .A2(net5843),
    .Y(_03900_),
    .B1(net6078));
 sg13g2_a22oi_1 _18138_ (.Y(_03901_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .A2(net5864),
    .A1(\soc_inst.cpu_core.register_file.registers[23][18] ));
 sg13g2_nand4_1 _18139_ (.B(_03890_),
    .C(_03900_),
    .A(_03889_),
    .Y(_03902_),
    .D(_03901_));
 sg13g2_a22oi_1 _18140_ (.Y(_03903_),
    .B1(net5853),
    .B2(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][18] ));
 sg13g2_a22oi_1 _18141_ (.Y(_03904_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][18] ),
    .A2(net5475),
    .A1(\soc_inst.cpu_core.register_file.registers[9][18] ));
 sg13g2_a22oi_1 _18142_ (.Y(_03905_),
    .B1(net5788),
    .B2(\soc_inst.cpu_core.register_file.registers[3][18] ),
    .A2(net5838),
    .A1(\soc_inst.cpu_core.register_file.registers[10][18] ));
 sg13g2_nand4_1 _18143_ (.B(_03903_),
    .C(_03904_),
    .A(_03887_),
    .Y(_03906_),
    .D(_03905_));
 sg13g2_nor3_2 _18144_ (.A(_03899_),
    .B(_03902_),
    .C(_03906_),
    .Y(_03907_));
 sg13g2_a21oi_1 _18145_ (.A1(net1036),
    .A2(net5102),
    .Y(_03908_),
    .B1(net5291));
 sg13g2_or2_1 _18146_ (.X(_03909_),
    .B(_03908_),
    .A(_03907_));
 sg13g2_o21ai_1 _18147_ (.B1(_03909_),
    .Y(_01074_),
    .A1(net6147),
    .A2(_08077_));
 sg13g2_and2_1 _18148_ (.A(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .B(net5813),
    .X(_03910_));
 sg13g2_a22oi_1 _18149_ (.Y(_03911_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][19] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][19] ));
 sg13g2_a22oi_1 _18150_ (.Y(_03912_),
    .B1(net5469),
    .B2(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][19] ));
 sg13g2_a22oi_1 _18151_ (.Y(_03913_),
    .B1(net5803),
    .B2(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .A2(net5474),
    .A1(\soc_inst.cpu_core.register_file.registers[9][19] ));
 sg13g2_a22oi_1 _18152_ (.Y(_03914_),
    .B1(net5838),
    .B2(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][19] ));
 sg13g2_a22oi_1 _18153_ (.Y(_03915_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][19] ),
    .A2(net5843),
    .A1(\soc_inst.cpu_core.register_file.registers[26][19] ));
 sg13g2_a22oi_1 _18154_ (.Y(_03916_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][19] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][19] ));
 sg13g2_a22oi_1 _18155_ (.Y(_03917_),
    .B1(net5258),
    .B2(\soc_inst.cpu_core.register_file.registers[28][19] ),
    .A2(net5848),
    .A1(\soc_inst.cpu_core.register_file.registers[2][19] ));
 sg13g2_nand3_1 _18156_ (.B(_03916_),
    .C(_03917_),
    .A(_03915_),
    .Y(_03918_));
 sg13g2_a221oi_1 _18157_ (.B2(\soc_inst.cpu_core.register_file.registers[24][19] ),
    .C1(_03918_),
    .B1(net5253),
    .A1(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .Y(_03919_),
    .A2(net5873));
 sg13g2_a22oi_1 _18158_ (.Y(_03920_),
    .B1(net5818),
    .B2(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][19] ));
 sg13g2_a22oi_1 _18159_ (.Y(_03921_),
    .B1(net5788),
    .B2(\soc_inst.cpu_core.register_file.registers[3][19] ),
    .A2(net5288),
    .A1(\soc_inst.cpu_core.register_file.registers[25][19] ));
 sg13g2_a221oi_1 _18160_ (.B2(\soc_inst.cpu_core.register_file.registers[30][19] ),
    .C1(_03910_),
    .B1(net5828),
    .A1(\soc_inst.cpu_core.register_file.registers[20][19] ),
    .Y(_03922_),
    .A2(net5278));
 sg13g2_nand4_1 _18161_ (.B(_03920_),
    .C(_03921_),
    .A(_03919_),
    .Y(_03923_),
    .D(_03922_));
 sg13g2_a21oi_1 _18162_ (.A1(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .A2(net5479),
    .Y(_03924_),
    .B1(net6078));
 sg13g2_a22oi_1 _18163_ (.Y(_03925_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][19] ),
    .A2(net5823),
    .A1(\soc_inst.cpu_core.register_file.registers[18][19] ));
 sg13g2_nand4_1 _18164_ (.B(_03912_),
    .C(_03924_),
    .A(_03911_),
    .Y(_03926_),
    .D(_03925_));
 sg13g2_a22oi_1 _18165_ (.Y(_03927_),
    .B1(net5274),
    .B2(\soc_inst.cpu_core.register_file.registers[17][19] ),
    .A2(net5863),
    .A1(\soc_inst.cpu_core.register_file.registers[23][19] ));
 sg13g2_a22oi_1 _18166_ (.Y(_03928_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .A2(net5793),
    .A1(\soc_inst.cpu_core.register_file.registers[6][19] ));
 sg13g2_nand4_1 _18167_ (.B(_03914_),
    .C(_03927_),
    .A(_03913_),
    .Y(_03929_),
    .D(_03928_));
 sg13g2_nor3_1 _18168_ (.A(_03923_),
    .B(_03926_),
    .C(_03929_),
    .Y(_03930_));
 sg13g2_a21oi_1 _18169_ (.A1(net392),
    .A2(net5105),
    .Y(_03931_),
    .B1(net5295));
 sg13g2_or2_1 _18170_ (.X(_03932_),
    .B(_03931_),
    .A(_03930_));
 sg13g2_o21ai_1 _18171_ (.B1(_03932_),
    .Y(_01075_),
    .A1(net6147),
    .A2(_08075_));
 sg13g2_a21oi_1 _18172_ (.A1(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .A2(net5105),
    .Y(_03933_),
    .B1(net5295));
 sg13g2_a22oi_1 _18173_ (.Y(_03934_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][20] ),
    .A2(net5289),
    .A1(\soc_inst.cpu_core.register_file.registers[25][20] ));
 sg13g2_a22oi_1 _18174_ (.Y(_03935_),
    .B1(net5854),
    .B2(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][20] ));
 sg13g2_a22oi_1 _18175_ (.Y(_03936_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][20] ),
    .A2(net5470),
    .A1(\soc_inst.cpu_core.register_file.registers[13][20] ));
 sg13g2_nand2_1 _18176_ (.Y(_03937_),
    .A(\soc_inst.cpu_core.register_file.registers[23][20] ),
    .B(net5864));
 sg13g2_a22oi_1 _18177_ (.Y(_03938_),
    .B1(net5804),
    .B2(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .A2(net5839),
    .A1(\soc_inst.cpu_core.register_file.registers[10][20] ));
 sg13g2_a22oi_1 _18178_ (.Y(_03939_),
    .B1(net5829),
    .B2(\soc_inst.cpu_core.register_file.registers[30][20] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][20] ));
 sg13g2_a22oi_1 _18179_ (.Y(_03940_),
    .B1(net5475),
    .B2(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .A2(net5279),
    .A1(\soc_inst.cpu_core.register_file.registers[20][20] ));
 sg13g2_a22oi_1 _18180_ (.Y(_03941_),
    .B1(net5273),
    .B2(\soc_inst.cpu_core.register_file.registers[17][20] ),
    .A2(net5844),
    .A1(\soc_inst.cpu_core.register_file.registers[26][20] ));
 sg13g2_a22oi_1 _18181_ (.Y(_03942_),
    .B1(net5814),
    .B2(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][20] ));
 sg13g2_a22oi_1 _18182_ (.Y(_03943_),
    .B1(net5849),
    .B2(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .A2(net5480),
    .A1(\soc_inst.cpu_core.register_file.registers[5][20] ));
 sg13g2_nand4_1 _18183_ (.B(_03936_),
    .C(_03942_),
    .A(_03935_),
    .Y(_03944_),
    .D(_03943_));
 sg13g2_a22oi_1 _18184_ (.Y(_03945_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][20] ),
    .A2(net5264),
    .A1(\soc_inst.cpu_core.register_file.registers[29][20] ));
 sg13g2_nand4_1 _18185_ (.B(_03940_),
    .C(_03941_),
    .A(_03937_),
    .Y(_03946_),
    .D(_03945_));
 sg13g2_nor2_2 _18186_ (.A(_03944_),
    .B(_03946_),
    .Y(_03947_));
 sg13g2_a21oi_1 _18187_ (.A1(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .A2(net5874),
    .Y(_03948_),
    .B1(net6079));
 sg13g2_a22oi_1 _18188_ (.Y(_03949_),
    .B1(net5794),
    .B2(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .A2(net5824),
    .A1(\soc_inst.cpu_core.register_file.registers[18][20] ));
 sg13g2_a22oi_1 _18189_ (.Y(_03950_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][20] ),
    .A2(net5809),
    .A1(\soc_inst.cpu_core.register_file.registers[27][20] ));
 sg13g2_nand4_1 _18190_ (.B(_03948_),
    .C(_03949_),
    .A(_03934_),
    .Y(_03951_),
    .D(_03950_));
 sg13g2_a22oi_1 _18191_ (.Y(_03952_),
    .B1(net5819),
    .B2(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][20] ));
 sg13g2_a22oi_1 _18192_ (.Y(_03953_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .A2(net5799),
    .A1(\soc_inst.cpu_core.register_file.registers[22][20] ));
 sg13g2_nand4_1 _18193_ (.B(_03939_),
    .C(_03952_),
    .A(_03938_),
    .Y(_03954_),
    .D(_03953_));
 sg13g2_nor2_2 _18194_ (.A(_03951_),
    .B(_03954_),
    .Y(_03955_));
 sg13g2_a21oi_2 _18195_ (.B1(_03933_),
    .Y(_03956_),
    .A2(_03955_),
    .A1(_03947_));
 sg13g2_a21o_1 _18196_ (.A2(net3359),
    .A1(net6386),
    .B1(_03956_),
    .X(_01076_));
 sg13g2_a21oi_1 _18197_ (.A1(net878),
    .A2(net5106),
    .Y(_03957_),
    .B1(net5295));
 sg13g2_a22oi_1 _18198_ (.Y(_03958_),
    .B1(net5260),
    .B2(\soc_inst.cpu_core.register_file.registers[28][21] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][21] ));
 sg13g2_a22oi_1 _18199_ (.Y(_03959_),
    .B1(net5800),
    .B2(\soc_inst.cpu_core.register_file.registers[22][21] ),
    .A2(net5825),
    .A1(\soc_inst.cpu_core.register_file.registers[18][21] ));
 sg13g2_nand2_1 _18200_ (.Y(_03960_),
    .A(\soc_inst.cpu_core.register_file.registers[17][21] ),
    .B(net5273));
 sg13g2_a22oi_1 _18201_ (.Y(_03961_),
    .B1(net5264),
    .B2(\soc_inst.cpu_core.register_file.registers[29][21] ),
    .A2(net5279),
    .A1(\soc_inst.cpu_core.register_file.registers[20][21] ));
 sg13g2_a22oi_1 _18202_ (.Y(_03962_),
    .B1(net5255),
    .B2(\soc_inst.cpu_core.register_file.registers[24][21] ),
    .A2(net5854),
    .A1(\soc_inst.cpu_core.register_file.registers[12][21] ));
 sg13g2_a22oi_1 _18203_ (.Y(_03963_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][21] ),
    .A2(net5814),
    .A1(\soc_inst.cpu_core.register_file.registers[11][21] ));
 sg13g2_a22oi_1 _18204_ (.Y(_03964_),
    .B1(net5480),
    .B2(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .A2(net5289),
    .A1(\soc_inst.cpu_core.register_file.registers[25][21] ));
 sg13g2_a22oi_1 _18205_ (.Y(_03965_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .A2(net5809),
    .A1(\soc_inst.cpu_core.register_file.registers[27][21] ));
 sg13g2_a22oi_1 _18206_ (.Y(_03966_),
    .B1(net5833),
    .B2(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .A2(net5840),
    .A1(\soc_inst.cpu_core.register_file.registers[10][21] ));
 sg13g2_a22oi_1 _18207_ (.Y(_03967_),
    .B1(net5849),
    .B2(\soc_inst.cpu_core.register_file.registers[2][21] ),
    .A2(net5875),
    .A1(\soc_inst.cpu_core.register_file.registers[4][21] ));
 sg13g2_nand4_1 _18208_ (.B(_03965_),
    .C(_03966_),
    .A(_03959_),
    .Y(_03968_),
    .D(_03967_));
 sg13g2_a22oi_1 _18209_ (.Y(_03969_),
    .B1(net5794),
    .B2(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][21] ));
 sg13g2_a22oi_1 _18210_ (.Y(_03970_),
    .B1(net5475),
    .B2(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .A2(net5865),
    .A1(\soc_inst.cpu_core.register_file.registers[23][21] ));
 sg13g2_nand4_1 _18211_ (.B(_03964_),
    .C(_03969_),
    .A(_03960_),
    .Y(_03971_),
    .D(_03970_));
 sg13g2_nor2_1 _18212_ (.A(_03968_),
    .B(_03971_),
    .Y(_03972_));
 sg13g2_a21oi_1 _18213_ (.A1(\soc_inst.cpu_core.register_file.registers[30][21] ),
    .A2(net5829),
    .Y(_03973_),
    .B1(net6079));
 sg13g2_a22oi_1 _18214_ (.Y(_03974_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .A2(net5845),
    .A1(\soc_inst.cpu_core.register_file.registers[26][21] ));
 sg13g2_nand4_1 _18215_ (.B(_03961_),
    .C(_03973_),
    .A(_03958_),
    .Y(_03975_),
    .D(_03974_));
 sg13g2_a22oi_1 _18216_ (.Y(_03976_),
    .B1(net5805),
    .B2(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .A2(net5819),
    .A1(\soc_inst.cpu_core.register_file.registers[8][21] ));
 sg13g2_a22oi_1 _18217_ (.Y(_03977_),
    .B1(net5790),
    .B2(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .A2(net5285),
    .A1(\soc_inst.cpu_core.register_file.registers[16][21] ));
 sg13g2_nand4_1 _18218_ (.B(_03963_),
    .C(_03976_),
    .A(_03962_),
    .Y(_03978_),
    .D(_03977_));
 sg13g2_nor2_1 _18219_ (.A(_03975_),
    .B(_03978_),
    .Y(_03979_));
 sg13g2_a21oi_2 _18220_ (.B1(_03957_),
    .Y(_03980_),
    .A2(_03979_),
    .A1(_03972_));
 sg13g2_a21o_1 _18221_ (.A2(net3112),
    .A1(net6397),
    .B1(_03980_),
    .X(_01077_));
 sg13g2_a21oi_1 _18222_ (.A1(net635),
    .A2(net5104),
    .Y(_03981_),
    .B1(net5291));
 sg13g2_a22oi_1 _18223_ (.Y(_03982_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][22] ),
    .A2(net5821),
    .A1(\soc_inst.cpu_core.register_file.registers[18][22] ));
 sg13g2_nand2_1 _18224_ (.Y(_03983_),
    .A(\soc_inst.cpu_core.register_file.registers[24][22] ),
    .B(net5251));
 sg13g2_a22oi_1 _18225_ (.Y(_03984_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][22] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][22] ));
 sg13g2_a22oi_1 _18226_ (.Y(_03985_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .A2(net5851),
    .A1(\soc_inst.cpu_core.register_file.registers[12][22] ));
 sg13g2_a22oi_1 _18227_ (.Y(_03986_),
    .B1(net5266),
    .B2(\soc_inst.cpu_core.register_file.registers[21][22] ),
    .A2(net5271),
    .A1(\soc_inst.cpu_core.register_file.registers[17][22] ));
 sg13g2_a22oi_1 _18228_ (.Y(_03987_),
    .B1(net5806),
    .B2(\soc_inst.cpu_core.register_file.registers[27][22] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][22] ));
 sg13g2_a22oi_1 _18229_ (.Y(_03988_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .A2(net5276),
    .A1(\soc_inst.cpu_core.register_file.registers[20][22] ));
 sg13g2_a22oi_1 _18230_ (.Y(_03989_),
    .B1(net5831),
    .B2(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][22] ));
 sg13g2_a22oi_1 _18231_ (.Y(_03990_),
    .B1(net5846),
    .B2(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .A2(net5871),
    .A1(\soc_inst.cpu_core.register_file.registers[4][22] ));
 sg13g2_nand4_1 _18232_ (.B(_03988_),
    .C(_03989_),
    .A(_03982_),
    .Y(_03991_),
    .D(_03990_));
 sg13g2_a22oi_1 _18233_ (.Y(_03992_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][22] ));
 sg13g2_a22oi_1 _18234_ (.Y(_03993_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][22] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][22] ));
 sg13g2_nand4_1 _18235_ (.B(_03984_),
    .C(_03992_),
    .A(_03983_),
    .Y(_03994_),
    .D(_03993_));
 sg13g2_nor2_1 _18236_ (.A(_03991_),
    .B(_03994_),
    .Y(_03995_));
 sg13g2_a21oi_1 _18237_ (.A1(\soc_inst.cpu_core.register_file.registers[26][22] ),
    .A2(net5841),
    .Y(_03996_),
    .B1(net6076));
 sg13g2_a22oi_1 _18238_ (.Y(_03997_),
    .B1(net5826),
    .B2(\soc_inst.cpu_core.register_file.registers[30][22] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][22] ));
 sg13g2_a22oi_1 _18239_ (.Y(_03998_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][22] ),
    .A2(net5467),
    .A1(\soc_inst.cpu_core.register_file.registers[13][22] ));
 sg13g2_nand4_1 _18240_ (.B(_03996_),
    .C(_03997_),
    .A(_03987_),
    .Y(_03999_),
    .D(_03998_));
 sg13g2_a22oi_1 _18241_ (.Y(_04000_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .A2(net5816),
    .A1(\soc_inst.cpu_core.register_file.registers[8][22] ));
 sg13g2_a22oi_1 _18242_ (.Y(_04001_),
    .B1(net5786),
    .B2(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][22] ));
 sg13g2_nand4_1 _18243_ (.B(_03986_),
    .C(_04000_),
    .A(_03985_),
    .Y(_04002_),
    .D(_04001_));
 sg13g2_nor2_1 _18244_ (.A(_03999_),
    .B(_04002_),
    .Y(_04003_));
 sg13g2_a21oi_2 _18245_ (.B1(_03981_),
    .Y(_04004_),
    .A2(_04003_),
    .A1(_03995_));
 sg13g2_a21o_1 _18246_ (.A2(net3100),
    .A1(net6398),
    .B1(_04004_),
    .X(_01078_));
 sg13g2_a21oi_1 _18247_ (.A1(net390),
    .A2(net5106),
    .Y(_04005_),
    .B1(net5295));
 sg13g2_a22oi_1 _18248_ (.Y(_04006_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][23] ),
    .A2(net5269),
    .A1(\soc_inst.cpu_core.register_file.registers[21][23] ));
 sg13g2_nand2_1 _18249_ (.Y(_04007_),
    .A(\soc_inst.cpu_core.register_file.registers[17][23] ),
    .B(net5273));
 sg13g2_a22oi_1 _18250_ (.Y(_04008_),
    .B1(net5264),
    .B2(\soc_inst.cpu_core.register_file.registers[29][23] ),
    .A2(net5470),
    .A1(\soc_inst.cpu_core.register_file.registers[13][23] ));
 sg13g2_a22oi_1 _18251_ (.Y(_04009_),
    .B1(net5809),
    .B2(\soc_inst.cpu_core.register_file.registers[27][23] ),
    .A2(net5829),
    .A1(\soc_inst.cpu_core.register_file.registers[30][23] ));
 sg13g2_a22oi_1 _18252_ (.Y(_04010_),
    .B1(net5824),
    .B2(\soc_inst.cpu_core.register_file.registers[18][23] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][23] ));
 sg13g2_a22oi_1 _18253_ (.Y(_04011_),
    .B1(net5814),
    .B2(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .A2(net5854),
    .A1(\soc_inst.cpu_core.register_file.registers[12][23] ));
 sg13g2_a22oi_1 _18254_ (.Y(_04012_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][23] ),
    .A2(net5480),
    .A1(\soc_inst.cpu_core.register_file.registers[5][23] ));
 sg13g2_a22oi_1 _18255_ (.Y(_04013_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .A2(net5279),
    .A1(\soc_inst.cpu_core.register_file.registers[20][23] ));
 sg13g2_a22oi_1 _18256_ (.Y(_04014_),
    .B1(net5839),
    .B2(\soc_inst.cpu_core.register_file.registers[10][23] ),
    .A2(net5864),
    .A1(\soc_inst.cpu_core.register_file.registers[23][23] ));
 sg13g2_a22oi_1 _18257_ (.Y(_04015_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][23] ),
    .A2(net5849),
    .A1(\soc_inst.cpu_core.register_file.registers[2][23] ));
 sg13g2_nand4_1 _18258_ (.B(_04013_),
    .C(_04014_),
    .A(_04010_),
    .Y(_04016_),
    .D(_04015_));
 sg13g2_a22oi_1 _18259_ (.Y(_04017_),
    .B1(net5794),
    .B2(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][23] ));
 sg13g2_a22oi_1 _18260_ (.Y(_04018_),
    .B1(net5799),
    .B2(\soc_inst.cpu_core.register_file.registers[22][23] ),
    .A2(net5819),
    .A1(\soc_inst.cpu_core.register_file.registers[8][23] ));
 sg13g2_nand4_1 _18261_ (.B(_04012_),
    .C(_04017_),
    .A(_04007_),
    .Y(_04019_),
    .D(_04018_));
 sg13g2_nor2_2 _18262_ (.A(_04016_),
    .B(_04019_),
    .Y(_04020_));
 sg13g2_a21oi_1 _18263_ (.A1(\soc_inst.cpu_core.register_file.registers[4][23] ),
    .A2(net5874),
    .Y(_04021_),
    .B1(net6079));
 sg13g2_a22oi_1 _18264_ (.Y(_04022_),
    .B1(net5869),
    .B2(\soc_inst.cpu_core.register_file.registers[31][23] ),
    .A2(net5289),
    .A1(\soc_inst.cpu_core.register_file.registers[25][23] ));
 sg13g2_nand4_1 _18265_ (.B(_04009_),
    .C(_04021_),
    .A(_04008_),
    .Y(_04023_),
    .D(_04022_));
 sg13g2_a22oi_1 _18266_ (.Y(_04024_),
    .B1(net5804),
    .B2(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .A2(net5475),
    .A1(\soc_inst.cpu_core.register_file.registers[9][23] ));
 sg13g2_a22oi_1 _18267_ (.Y(_04025_),
    .B1(net5844),
    .B2(\soc_inst.cpu_core.register_file.registers[26][23] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][23] ));
 sg13g2_nand4_1 _18268_ (.B(_04011_),
    .C(_04024_),
    .A(_04006_),
    .Y(_04026_),
    .D(_04025_));
 sg13g2_nor2_2 _18269_ (.A(_04023_),
    .B(_04026_),
    .Y(_04027_));
 sg13g2_a21oi_2 _18270_ (.B1(_04005_),
    .Y(_04028_),
    .A2(_04027_),
    .A1(_04020_));
 sg13g2_a21o_1 _18271_ (.A2(net3237),
    .A1(net6398),
    .B1(_04028_),
    .X(_01079_));
 sg13g2_a21oi_1 _18272_ (.A1(net1304),
    .A2(net5105),
    .Y(_04029_),
    .B1(net5295));
 sg13g2_a22oi_1 _18273_ (.Y(_04030_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .A2(net5841),
    .A1(\soc_inst.cpu_core.register_file.registers[26][24] ));
 sg13g2_nand2_1 _18274_ (.Y(_04031_),
    .A(\soc_inst.cpu_core.register_file.registers[27][24] ),
    .B(net5806));
 sg13g2_a22oi_1 _18275_ (.Y(_04032_),
    .B1(net5276),
    .B2(\soc_inst.cpu_core.register_file.registers[20][24] ),
    .A2(net5846),
    .A1(\soc_inst.cpu_core.register_file.registers[2][24] ));
 sg13g2_a22oi_1 _18276_ (.Y(_04033_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][24] ),
    .A2(net5472),
    .A1(\soc_inst.cpu_core.register_file.registers[9][24] ));
 sg13g2_a22oi_1 _18277_ (.Y(_04034_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][24] ));
 sg13g2_a22oi_1 _18278_ (.Y(_04035_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][24] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][24] ));
 sg13g2_a22oi_1 _18279_ (.Y(_04036_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][24] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][24] ));
 sg13g2_a22oi_1 _18280_ (.Y(_04037_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][24] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][24] ));
 sg13g2_a22oi_1 _18281_ (.Y(_04038_),
    .B1(net5831),
    .B2(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][24] ));
 sg13g2_nand4_1 _18282_ (.B(_04036_),
    .C(_04037_),
    .A(_04035_),
    .Y(_04039_),
    .D(_04038_));
 sg13g2_a22oi_1 _18283_ (.Y(_04040_),
    .B1(net5266),
    .B2(\soc_inst.cpu_core.register_file.registers[21][24] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][24] ));
 sg13g2_a22oi_1 _18284_ (.Y(_04041_),
    .B1(net5821),
    .B2(\soc_inst.cpu_core.register_file.registers[18][24] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][24] ));
 sg13g2_nand4_1 _18285_ (.B(_04033_),
    .C(_04040_),
    .A(_04031_),
    .Y(_04042_),
    .D(_04041_));
 sg13g2_nor2_1 _18286_ (.A(_04039_),
    .B(_04042_),
    .Y(_04043_));
 sg13g2_a21oi_1 _18287_ (.A1(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .A2(net5467),
    .Y(_04044_),
    .B1(net6077));
 sg13g2_a22oi_1 _18288_ (.Y(_04045_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .A2(net5786),
    .A1(\soc_inst.cpu_core.register_file.registers[3][24] ));
 sg13g2_a22oi_1 _18289_ (.Y(_04046_),
    .B1(net5816),
    .B2(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][24] ));
 sg13g2_nand4_1 _18290_ (.B(_04044_),
    .C(_04045_),
    .A(_04032_),
    .Y(_04047_),
    .D(_04046_));
 sg13g2_a22oi_1 _18291_ (.Y(_04048_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .A2(net5271),
    .A1(\soc_inst.cpu_core.register_file.registers[17][24] ));
 sg13g2_a22oi_1 _18292_ (.Y(_04049_),
    .B1(net5851),
    .B2(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .A2(net5871),
    .A1(\soc_inst.cpu_core.register_file.registers[4][24] ));
 sg13g2_nand4_1 _18293_ (.B(_04034_),
    .C(_04048_),
    .A(_04030_),
    .Y(_04050_),
    .D(_04049_));
 sg13g2_nor2_1 _18294_ (.A(_04047_),
    .B(_04050_),
    .Y(_04051_));
 sg13g2_a21oi_2 _18295_ (.B1(_04029_),
    .Y(_04052_),
    .A2(_04051_),
    .A1(_04043_));
 sg13g2_a21o_1 _18296_ (.A2(net3115),
    .A1(net6400),
    .B1(_04052_),
    .X(_01080_));
 sg13g2_a21oi_1 _18297_ (.A1(net1097),
    .A2(net5102),
    .Y(_04053_),
    .B1(net5291));
 sg13g2_a22oi_1 _18298_ (.Y(_04054_),
    .B1(net5271),
    .B2(\soc_inst.cpu_core.register_file.registers[17][25] ),
    .A2(net5831),
    .A1(\soc_inst.cpu_core.register_file.registers[14][25] ));
 sg13g2_nand2_1 _18299_ (.Y(_04055_),
    .A(\soc_inst.cpu_core.register_file.registers[20][25] ),
    .B(net5276));
 sg13g2_a22oi_1 _18300_ (.Y(_04056_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .A2(net5786),
    .A1(\soc_inst.cpu_core.register_file.registers[3][25] ));
 sg13g2_a22oi_1 _18301_ (.Y(_04057_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][25] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][25] ));
 sg13g2_a22oi_1 _18302_ (.Y(_04058_),
    .B1(net5266),
    .B2(\soc_inst.cpu_core.register_file.registers[21][25] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][25] ));
 sg13g2_a22oi_1 _18303_ (.Y(_04059_),
    .B1(net5791),
    .B2(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .A2(net5806),
    .A1(\soc_inst.cpu_core.register_file.registers[27][25] ));
 sg13g2_a22oi_1 _18304_ (.Y(_04060_),
    .B1(net5821),
    .B2(\soc_inst.cpu_core.register_file.registers[18][25] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][25] ));
 sg13g2_a22oi_1 _18305_ (.Y(_04061_),
    .B1(net5841),
    .B2(\soc_inst.cpu_core.register_file.registers[26][25] ),
    .A2(net5851),
    .A1(\soc_inst.cpu_core.register_file.registers[12][25] ));
 sg13g2_a22oi_1 _18306_ (.Y(_04062_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .A2(net5811),
    .A1(\soc_inst.cpu_core.register_file.registers[11][25] ));
 sg13g2_nand4_1 _18307_ (.B(_04060_),
    .C(_04061_),
    .A(_04058_),
    .Y(_04063_),
    .D(_04062_));
 sg13g2_a22oi_1 _18308_ (.Y(_04064_),
    .B1(net5467),
    .B2(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .A2(net5846),
    .A1(\soc_inst.cpu_core.register_file.registers[2][25] ));
 sg13g2_a22oi_1 _18309_ (.Y(_04065_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][25] ));
 sg13g2_nand4_1 _18310_ (.B(_04059_),
    .C(_04064_),
    .A(_04055_),
    .Y(_04066_),
    .D(_04065_));
 sg13g2_nor2_1 _18311_ (.A(_04063_),
    .B(_04066_),
    .Y(_04067_));
 sg13g2_a21oi_1 _18312_ (.A1(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .A2(net5816),
    .Y(_04068_),
    .B1(net6076));
 sg13g2_a22oi_1 _18313_ (.Y(_04069_),
    .B1(net5826),
    .B2(\soc_inst.cpu_core.register_file.registers[30][25] ),
    .A2(net5871),
    .A1(\soc_inst.cpu_core.register_file.registers[4][25] ));
 sg13g2_a22oi_1 _18314_ (.Y(_04070_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][25] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][25] ));
 sg13g2_nand4_1 _18315_ (.B(_04068_),
    .C(_04069_),
    .A(_04056_),
    .Y(_04071_),
    .D(_04070_));
 sg13g2_a22oi_1 _18316_ (.Y(_04072_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][25] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][25] ));
 sg13g2_a22oi_1 _18317_ (.Y(_04073_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][25] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][25] ));
 sg13g2_nand4_1 _18318_ (.B(_04057_),
    .C(_04072_),
    .A(_04054_),
    .Y(_04074_),
    .D(_04073_));
 sg13g2_nor2_1 _18319_ (.A(_04071_),
    .B(_04074_),
    .Y(_04075_));
 sg13g2_a21oi_1 _18320_ (.A1(_04067_),
    .A2(_04075_),
    .Y(_04076_),
    .B1(_04053_));
 sg13g2_a21o_1 _18321_ (.A2(net3362),
    .A1(net6399),
    .B1(_04076_),
    .X(_01081_));
 sg13g2_a21oi_1 _18322_ (.A1(net912),
    .A2(net5105),
    .Y(_04077_),
    .B1(net5295));
 sg13g2_a22oi_1 _18323_ (.Y(_04078_),
    .B1(net5258),
    .B2(\soc_inst.cpu_core.register_file.registers[28][26] ),
    .A2(net5479),
    .A1(\soc_inst.cpu_core.register_file.registers[5][26] ));
 sg13g2_nand2_1 _18324_ (.Y(_04079_),
    .A(\soc_inst.cpu_core.register_file.registers[23][26] ),
    .B(net5863));
 sg13g2_a22oi_1 _18325_ (.Y(_04080_),
    .B1(net5469),
    .B2(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .A2(net5873),
    .A1(\soc_inst.cpu_core.register_file.registers[4][26] ));
 sg13g2_a22oi_1 _18326_ (.Y(_04081_),
    .B1(net5268),
    .B2(\soc_inst.cpu_core.register_file.registers[21][26] ),
    .A2(net5834),
    .A1(\soc_inst.cpu_core.register_file.registers[14][26] ));
 sg13g2_a22oi_1 _18327_ (.Y(_04082_),
    .B1(net5793),
    .B2(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .A2(net5818),
    .A1(\soc_inst.cpu_core.register_file.registers[8][26] ));
 sg13g2_a22oi_1 _18328_ (.Y(_04083_),
    .B1(net5783),
    .B2(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .A2(net5278),
    .A1(\soc_inst.cpu_core.register_file.registers[20][26] ));
 sg13g2_a22oi_1 _18329_ (.Y(_04084_),
    .B1(net5808),
    .B2(\soc_inst.cpu_core.register_file.registers[27][26] ),
    .A2(net5828),
    .A1(\soc_inst.cpu_core.register_file.registers[30][26] ));
 sg13g2_a22oi_1 _18330_ (.Y(_04085_),
    .B1(net5788),
    .B2(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .A2(net5848),
    .A1(\soc_inst.cpu_core.register_file.registers[2][26] ));
 sg13g2_nand4_1 _18331_ (.B(_04080_),
    .C(_04084_),
    .A(_04078_),
    .Y(_04086_),
    .D(_04085_));
 sg13g2_a22oi_1 _18332_ (.Y(_04087_),
    .B1(net5813),
    .B2(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .A2(net5853),
    .A1(\soc_inst.cpu_core.register_file.registers[12][26] ));
 sg13g2_nand4_1 _18333_ (.B(_04082_),
    .C(_04083_),
    .A(_04079_),
    .Y(_04088_),
    .D(_04087_));
 sg13g2_nor2_1 _18334_ (.A(_04086_),
    .B(_04088_),
    .Y(_04089_));
 sg13g2_a21oi_1 _18335_ (.A1(\soc_inst.cpu_core.register_file.registers[25][26] ),
    .A2(net5288),
    .Y(_04090_),
    .B1(net6078));
 sg13g2_a22oi_1 _18336_ (.Y(_04091_),
    .B1(net5823),
    .B2(\soc_inst.cpu_core.register_file.registers[18][26] ),
    .A2(net5838),
    .A1(\soc_inst.cpu_core.register_file.registers[10][26] ));
 sg13g2_a22oi_1 _18337_ (.Y(_04092_),
    .B1(net5803),
    .B2(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .A2(net5283),
    .A1(\soc_inst.cpu_core.register_file.registers[16][26] ));
 sg13g2_nand4_1 _18338_ (.B(_04090_),
    .C(_04091_),
    .A(_04081_),
    .Y(_04093_),
    .D(_04092_));
 sg13g2_a22oi_1 _18339_ (.Y(_04094_),
    .B1(net5253),
    .B2(\soc_inst.cpu_core.register_file.registers[24][26] ),
    .A2(net5274),
    .A1(\soc_inst.cpu_core.register_file.registers[17][26] ));
 sg13g2_a22oi_1 _18340_ (.Y(_04095_),
    .B1(net5474),
    .B2(\soc_inst.cpu_core.register_file.registers[9][26] ),
    .A2(net5858),
    .A1(\soc_inst.cpu_core.register_file.registers[19][26] ));
 sg13g2_a22oi_1 _18341_ (.Y(_04096_),
    .B1(net5798),
    .B2(\soc_inst.cpu_core.register_file.registers[22][26] ),
    .A2(net5843),
    .A1(\soc_inst.cpu_core.register_file.registers[26][26] ));
 sg13g2_a22oi_1 _18342_ (.Y(_04097_),
    .B1(net5263),
    .B2(\soc_inst.cpu_core.register_file.registers[29][26] ),
    .A2(net5868),
    .A1(\soc_inst.cpu_core.register_file.registers[31][26] ));
 sg13g2_nand4_1 _18343_ (.B(_04095_),
    .C(_04096_),
    .A(_04094_),
    .Y(_04098_),
    .D(_04097_));
 sg13g2_nor2_1 _18344_ (.A(_04093_),
    .B(_04098_),
    .Y(_04099_));
 sg13g2_a21oi_2 _18345_ (.B1(_04077_),
    .Y(_04100_),
    .A2(_04099_),
    .A1(_04089_));
 sg13g2_a21o_1 _18346_ (.A2(net3134),
    .A1(net6400),
    .B1(_04100_),
    .X(_01082_));
 sg13g2_a21oi_1 _18347_ (.A1(net829),
    .A2(net5102),
    .Y(_04101_),
    .B1(net5294));
 sg13g2_nand2_1 _18348_ (.Y(_04102_),
    .A(\soc_inst.cpu_core.register_file.registers[3][27] ),
    .B(net5786));
 sg13g2_a22oi_1 _18349_ (.Y(_04103_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][27] ));
 sg13g2_a22oi_1 _18350_ (.Y(_04104_),
    .B1(net5841),
    .B2(\soc_inst.cpu_core.register_file.registers[26][27] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][27] ));
 sg13g2_a22oi_1 _18351_ (.Y(_04105_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][27] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][27] ));
 sg13g2_a22oi_1 _18352_ (.Y(_04106_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][27] ));
 sg13g2_a22oi_1 _18353_ (.Y(_04107_),
    .B1(net5266),
    .B2(\soc_inst.cpu_core.register_file.registers[21][27] ),
    .A2(net5271),
    .A1(\soc_inst.cpu_core.register_file.registers[17][27] ));
 sg13g2_a22oi_1 _18354_ (.Y(_04108_),
    .B1(net5856),
    .B2(\soc_inst.cpu_core.register_file.registers[19][27] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][27] ));
 sg13g2_a22oi_1 _18355_ (.Y(_04109_),
    .B1(net5806),
    .B2(\soc_inst.cpu_core.register_file.registers[27][27] ),
    .A2(net5276),
    .A1(\soc_inst.cpu_core.register_file.registers[20][27] ));
 sg13g2_a22oi_1 _18356_ (.Y(_04110_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .A2(net5816),
    .A1(\soc_inst.cpu_core.register_file.registers[8][27] ));
 sg13g2_nand4_1 _18357_ (.B(_04108_),
    .C(_04109_),
    .A(_04105_),
    .Y(_04111_),
    .D(_04110_));
 sg13g2_a22oi_1 _18358_ (.Y(_04112_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .A2(net5831),
    .A1(\soc_inst.cpu_core.register_file.registers[14][27] ));
 sg13g2_a22oi_1 _18359_ (.Y(_04113_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][27] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][27] ));
 sg13g2_nand4_1 _18360_ (.B(_04107_),
    .C(_04112_),
    .A(_04102_),
    .Y(_04114_),
    .D(_04113_));
 sg13g2_nor2_1 _18361_ (.A(_04111_),
    .B(_04114_),
    .Y(_04115_));
 sg13g2_a21oi_1 _18362_ (.A1(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .A2(net5851),
    .Y(_04116_),
    .B1(net6076));
 sg13g2_a22oi_1 _18363_ (.Y(_04117_),
    .B1(net5467),
    .B2(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .A2(net5871),
    .A1(\soc_inst.cpu_core.register_file.registers[4][27] ));
 sg13g2_a22oi_1 _18364_ (.Y(_04118_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][27] ),
    .A2(net5821),
    .A1(\soc_inst.cpu_core.register_file.registers[18][27] ));
 sg13g2_nand4_1 _18365_ (.B(_04116_),
    .C(_04117_),
    .A(_04106_),
    .Y(_04119_),
    .D(_04118_));
 sg13g2_a22oi_1 _18366_ (.Y(_04120_),
    .B1(net5846),
    .B2(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .A2(net5477),
    .A1(\soc_inst.cpu_core.register_file.registers[5][27] ));
 sg13g2_a22oi_1 _18367_ (.Y(_04121_),
    .B1(net5256),
    .B2(\soc_inst.cpu_core.register_file.registers[28][27] ),
    .A2(net5791),
    .A1(\soc_inst.cpu_core.register_file.registers[6][27] ));
 sg13g2_nand4_1 _18368_ (.B(_04104_),
    .C(_04120_),
    .A(_04103_),
    .Y(_04122_),
    .D(_04121_));
 sg13g2_nor2_1 _18369_ (.A(_04119_),
    .B(_04122_),
    .Y(_04123_));
 sg13g2_a21oi_2 _18370_ (.B1(_04101_),
    .Y(_04124_),
    .A2(_04123_),
    .A1(_04115_));
 sg13g2_a21o_1 _18371_ (.A2(net3132),
    .A1(net6401),
    .B1(_04124_),
    .X(_01083_));
 sg13g2_a21oi_1 _18372_ (.A1(net484),
    .A2(net5105),
    .Y(_04125_),
    .B1(net5295));
 sg13g2_nand2_1 _18373_ (.Y(_04126_),
    .A(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .B(net5871));
 sg13g2_a22oi_1 _18374_ (.Y(_04127_),
    .B1(net5841),
    .B2(\soc_inst.cpu_core.register_file.registers[26][28] ),
    .A2(net5866),
    .A1(\soc_inst.cpu_core.register_file.registers[31][28] ));
 sg13g2_a22oi_1 _18375_ (.Y(_04128_),
    .B1(net5271),
    .B2(\soc_inst.cpu_core.register_file.registers[17][28] ),
    .A2(net5281),
    .A1(\soc_inst.cpu_core.register_file.registers[16][28] ));
 sg13g2_a22oi_1 _18376_ (.Y(_04129_),
    .B1(net5251),
    .B2(\soc_inst.cpu_core.register_file.registers[24][28] ),
    .A2(net5266),
    .A1(\soc_inst.cpu_core.register_file.registers[21][28] ));
 sg13g2_a22oi_1 _18377_ (.Y(_04130_),
    .B1(net5792),
    .B2(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .A2(net5806),
    .A1(\soc_inst.cpu_core.register_file.registers[27][28] ));
 sg13g2_a22oi_1 _18378_ (.Y(_04131_),
    .B1(net5781),
    .B2(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .A2(net5856),
    .A1(\soc_inst.cpu_core.register_file.registers[19][28] ));
 sg13g2_a22oi_1 _18379_ (.Y(_04132_),
    .B1(net5801),
    .B2(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .A2(net5816),
    .A1(\soc_inst.cpu_core.register_file.registers[8][28] ));
 sg13g2_a22oi_1 _18380_ (.Y(_04133_),
    .B1(net5811),
    .B2(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .A2(net5851),
    .A1(\soc_inst.cpu_core.register_file.registers[12][28] ));
 sg13g2_nand4_1 _18381_ (.B(_04131_),
    .C(_04132_),
    .A(_04128_),
    .Y(_04134_),
    .D(_04133_));
 sg13g2_a22oi_1 _18382_ (.Y(_04135_),
    .B1(net5261),
    .B2(\soc_inst.cpu_core.register_file.registers[29][28] ),
    .A2(net5826),
    .A1(\soc_inst.cpu_core.register_file.registers[30][28] ));
 sg13g2_nand4_1 _18383_ (.B(_04129_),
    .C(_04130_),
    .A(_04126_),
    .Y(_04136_),
    .D(_04135_));
 sg13g2_nor2_1 _18384_ (.A(_04134_),
    .B(_04136_),
    .Y(_04137_));
 sg13g2_a21oi_1 _18385_ (.A1(\soc_inst.cpu_core.register_file.registers[28][28] ),
    .A2(net5256),
    .Y(_04138_),
    .B1(net6076));
 sg13g2_a22oi_1 _18386_ (.Y(_04139_),
    .B1(net5468),
    .B2(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .A2(net5276),
    .A1(\soc_inst.cpu_core.register_file.registers[20][28] ));
 sg13g2_a22oi_1 _18387_ (.Y(_04140_),
    .B1(net5796),
    .B2(\soc_inst.cpu_core.register_file.registers[22][28] ),
    .A2(net5821),
    .A1(\soc_inst.cpu_core.register_file.registers[18][28] ));
 sg13g2_nand4_1 _18388_ (.B(_04138_),
    .C(_04139_),
    .A(_04127_),
    .Y(_04141_),
    .D(_04140_));
 sg13g2_a22oi_1 _18389_ (.Y(_04142_),
    .B1(net5786),
    .B2(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .A2(net5846),
    .A1(\soc_inst.cpu_core.register_file.registers[2][28] ));
 sg13g2_a22oi_1 _18390_ (.Y(_04143_),
    .B1(net5831),
    .B2(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .A2(net5836),
    .A1(\soc_inst.cpu_core.register_file.registers[10][28] ));
 sg13g2_a22oi_1 _18391_ (.Y(_04144_),
    .B1(net5472),
    .B2(\soc_inst.cpu_core.register_file.registers[9][28] ),
    .A2(net5861),
    .A1(\soc_inst.cpu_core.register_file.registers[23][28] ));
 sg13g2_a22oi_1 _18392_ (.Y(_04145_),
    .B1(net5477),
    .B2(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .A2(net5286),
    .A1(\soc_inst.cpu_core.register_file.registers[25][28] ));
 sg13g2_nand4_1 _18393_ (.B(_04143_),
    .C(_04144_),
    .A(_04142_),
    .Y(_04146_),
    .D(_04145_));
 sg13g2_nor2_1 _18394_ (.A(_04141_),
    .B(_04146_),
    .Y(_04147_));
 sg13g2_a21oi_2 _18395_ (.B1(_04125_),
    .Y(_04148_),
    .A2(_04147_),
    .A1(_04137_));
 sg13g2_a21o_1 _18396_ (.A2(net1318),
    .A1(net6401),
    .B1(_04148_),
    .X(_01084_));
 sg13g2_a21oi_1 _18397_ (.A1(net741),
    .A2(net5105),
    .Y(_04149_),
    .B1(net5292));
 sg13g2_nand2_1 _18398_ (.Y(_04150_),
    .A(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .B(net5872));
 sg13g2_a22oi_1 _18399_ (.Y(_04151_),
    .B1(net5257),
    .B2(\soc_inst.cpu_core.register_file.registers[28][29] ),
    .A2(net5797),
    .A1(\soc_inst.cpu_core.register_file.registers[22][29] ));
 sg13g2_a22oi_1 _18400_ (.Y(_04152_),
    .B1(net5473),
    .B2(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .A2(net5478),
    .A1(\soc_inst.cpu_core.register_file.registers[5][29] ));
 sg13g2_a22oi_1 _18401_ (.Y(_04153_),
    .B1(net5272),
    .B2(\soc_inst.cpu_core.register_file.registers[17][29] ),
    .A2(net5282),
    .A1(\soc_inst.cpu_core.register_file.registers[16][29] ));
 sg13g2_a22oi_1 _18402_ (.Y(_04154_),
    .B1(net5252),
    .B2(\soc_inst.cpu_core.register_file.registers[24][29] ),
    .A2(net5267),
    .A1(\soc_inst.cpu_core.register_file.registers[21][29] ));
 sg13g2_a22oi_1 _18403_ (.Y(_04155_),
    .B1(net5782),
    .B2(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .A2(net5262),
    .A1(\soc_inst.cpu_core.register_file.registers[29][29] ));
 sg13g2_a22oi_1 _18404_ (.Y(_04156_),
    .B1(net5807),
    .B2(\soc_inst.cpu_core.register_file.registers[27][29] ),
    .A2(net5827),
    .A1(\soc_inst.cpu_core.register_file.registers[30][29] ));
 sg13g2_a22oi_1 _18405_ (.Y(_04157_),
    .B1(net5795),
    .B2(\soc_inst.cpu_core.register_file.registers[6][29] ),
    .A2(net5857),
    .A1(\soc_inst.cpu_core.register_file.registers[19][29] ));
 sg13g2_a22oi_1 _18406_ (.Y(_04158_),
    .B1(net5802),
    .B2(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .A2(net5817),
    .A1(\soc_inst.cpu_core.register_file.registers[8][29] ));
 sg13g2_a22oi_1 _18407_ (.Y(_04159_),
    .B1(net5812),
    .B2(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .A2(net5852),
    .A1(\soc_inst.cpu_core.register_file.registers[12][29] ));
 sg13g2_nand4_1 _18408_ (.B(_04157_),
    .C(_04158_),
    .A(_04153_),
    .Y(_04160_),
    .D(_04159_));
 sg13g2_a22oi_1 _18409_ (.Y(_04161_),
    .B1(net5842),
    .B2(\soc_inst.cpu_core.register_file.registers[26][29] ),
    .A2(net5277),
    .A1(\soc_inst.cpu_core.register_file.registers[20][29] ));
 sg13g2_nand4_1 _18410_ (.B(_04154_),
    .C(_04155_),
    .A(_04150_),
    .Y(_04162_),
    .D(_04161_));
 sg13g2_nor2_1 _18411_ (.A(_04160_),
    .B(_04162_),
    .Y(_04163_));
 sg13g2_a21oi_1 _18412_ (.A1(\soc_inst.cpu_core.register_file.registers[31][29] ),
    .A2(net5867),
    .Y(_04164_),
    .B1(net6077));
 sg13g2_a22oi_1 _18413_ (.Y(_04165_),
    .B1(net5822),
    .B2(\soc_inst.cpu_core.register_file.registers[18][29] ),
    .A2(net5862),
    .A1(\soc_inst.cpu_core.register_file.registers[23][29] ));
 sg13g2_a22oi_1 _18414_ (.Y(_04166_),
    .B1(net5471),
    .B2(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .A2(net5287),
    .A1(\soc_inst.cpu_core.register_file.registers[25][29] ));
 sg13g2_nand4_1 _18415_ (.B(_04164_),
    .C(_04165_),
    .A(_04156_),
    .Y(_04167_),
    .D(_04166_));
 sg13g2_a22oi_1 _18416_ (.Y(_04168_),
    .B1(net5787),
    .B2(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .A2(net5847),
    .A1(\soc_inst.cpu_core.register_file.registers[2][29] ));
 sg13g2_a22oi_1 _18417_ (.Y(_04169_),
    .B1(net5832),
    .B2(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .A2(net5837),
    .A1(\soc_inst.cpu_core.register_file.registers[10][29] ));
 sg13g2_nand4_1 _18418_ (.B(_04152_),
    .C(_04168_),
    .A(_04151_),
    .Y(_04170_),
    .D(_04169_));
 sg13g2_nor2_1 _18419_ (.A(_04167_),
    .B(_04170_),
    .Y(_04171_));
 sg13g2_a21oi_2 _18420_ (.B1(_04149_),
    .Y(_04172_),
    .A2(_04171_),
    .A1(_04163_));
 sg13g2_a21o_1 _18421_ (.A2(net1343),
    .A1(net6401),
    .B1(_04172_),
    .X(_01085_));
 sg13g2_a21oi_2 _18422_ (.B1(net5295),
    .Y(_04173_),
    .A2(net5106),
    .A1(\soc_inst.cpu_core.register_file.registers[1][30] ));
 sg13g2_nand2_1 _18423_ (.Y(_04174_),
    .A(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .B(net5874));
 sg13g2_a22oi_1 _18424_ (.Y(_04175_),
    .B1(net5814),
    .B2(\soc_inst.cpu_core.register_file.registers[11][30] ),
    .A2(net5854),
    .A1(\soc_inst.cpu_core.register_file.registers[12][30] ));
 sg13g2_a22oi_1 _18425_ (.Y(_04176_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][30] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][30] ));
 sg13g2_a22oi_1 _18426_ (.Y(_04177_),
    .B1(net5799),
    .B2(\soc_inst.cpu_core.register_file.registers[22][30] ),
    .A2(net5859),
    .A1(\soc_inst.cpu_core.register_file.registers[19][30] ));
 sg13g2_a22oi_1 _18427_ (.Y(_04178_),
    .B1(net5784),
    .B2(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .A2(net5864),
    .A1(\soc_inst.cpu_core.register_file.registers[23][30] ));
 sg13g2_a22oi_1 _18428_ (.Y(_04179_),
    .B1(net5804),
    .B2(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .A2(net5820),
    .A1(\soc_inst.cpu_core.register_file.registers[8][30] ));
 sg13g2_nand4_1 _18429_ (.B(_04176_),
    .C(_04178_),
    .A(_04175_),
    .Y(_04180_),
    .D(_04179_));
 sg13g2_a22oi_1 _18430_ (.Y(_04181_),
    .B1(net5279),
    .B2(\soc_inst.cpu_core.register_file.registers[20][30] ),
    .A2(net5289),
    .A1(\soc_inst.cpu_core.register_file.registers[25][30] ));
 sg13g2_a22oi_1 _18431_ (.Y(_04182_),
    .B1(net5794),
    .B2(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .A2(net5264),
    .A1(\soc_inst.cpu_core.register_file.registers[29][30] ));
 sg13g2_nand4_1 _18432_ (.B(_04177_),
    .C(_04181_),
    .A(_04174_),
    .Y(_04183_),
    .D(_04182_));
 sg13g2_nor2_1 _18433_ (.A(_04180_),
    .B(_04183_),
    .Y(_04184_));
 sg13g2_a21oi_1 _18434_ (.A1(\soc_inst.cpu_core.register_file.registers[30][30] ),
    .A2(net5829),
    .Y(_04185_),
    .B1(net6080));
 sg13g2_a22oi_1 _18435_ (.Y(_04186_),
    .B1(net5809),
    .B2(\soc_inst.cpu_core.register_file.registers[27][30] ),
    .A2(net5869),
    .A1(\soc_inst.cpu_core.register_file.registers[31][30] ));
 sg13g2_a22oi_1 _18436_ (.Y(_04187_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .A2(net5844),
    .A1(\soc_inst.cpu_core.register_file.registers[26][30] ));
 sg13g2_a22oi_1 _18437_ (.Y(_04188_),
    .B1(net5269),
    .B2(\soc_inst.cpu_core.register_file.registers[21][30] ),
    .A2(net5824),
    .A1(\soc_inst.cpu_core.register_file.registers[18][30] ));
 sg13g2_nand4_1 _18438_ (.B(_04186_),
    .C(_04187_),
    .A(_04185_),
    .Y(_04189_),
    .D(_04188_));
 sg13g2_a22oi_1 _18439_ (.Y(_04190_),
    .B1(net5835),
    .B2(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .A2(net5839),
    .A1(\soc_inst.cpu_core.register_file.registers[10][30] ));
 sg13g2_a22oi_1 _18440_ (.Y(_04191_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .A2(net5849),
    .A1(\soc_inst.cpu_core.register_file.registers[2][30] ));
 sg13g2_a22oi_1 _18441_ (.Y(_04192_),
    .B1(net5475),
    .B2(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .A2(net5275),
    .A1(\soc_inst.cpu_core.register_file.registers[17][30] ));
 sg13g2_a22oi_1 _18442_ (.Y(_04193_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][30] ),
    .A2(net5481),
    .A1(\soc_inst.cpu_core.register_file.registers[5][30] ));
 sg13g2_nand4_1 _18443_ (.B(_04191_),
    .C(_04192_),
    .A(_04190_),
    .Y(_04194_),
    .D(_04193_));
 sg13g2_nor2_1 _18444_ (.A(_04189_),
    .B(_04194_),
    .Y(_04195_));
 sg13g2_a21oi_2 _18445_ (.B1(_04173_),
    .Y(_04196_),
    .A2(_04195_),
    .A1(_04184_));
 sg13g2_a21o_1 _18446_ (.A2(net3360),
    .A1(net6400),
    .B1(_04196_),
    .X(_01086_));
 sg13g2_and2_1 _18447_ (.A(\soc_inst.cpu_core.register_file.registers[30][31] ),
    .B(net5829),
    .X(_04197_));
 sg13g2_a22oi_1 _18448_ (.Y(_04198_),
    .B1(net5264),
    .B2(\soc_inst.cpu_core.register_file.registers[29][31] ),
    .A2(net5475),
    .A1(\soc_inst.cpu_core.register_file.registers[9][31] ));
 sg13g2_a22oi_1 _18449_ (.Y(_04199_),
    .B1(net5824),
    .B2(\soc_inst.cpu_core.register_file.registers[18][31] ),
    .A2(net5480),
    .A1(\soc_inst.cpu_core.register_file.registers[5][31] ));
 sg13g2_a22oi_1 _18450_ (.Y(_04200_),
    .B1(net5254),
    .B2(\soc_inst.cpu_core.register_file.registers[24][31] ),
    .A2(net5855),
    .A1(\soc_inst.cpu_core.register_file.registers[12][31] ));
 sg13g2_a22oi_1 _18451_ (.Y(_04201_),
    .B1(net5794),
    .B2(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .A2(net5799),
    .A1(\soc_inst.cpu_core.register_file.registers[22][31] ));
 sg13g2_a22oi_1 _18452_ (.Y(_04202_),
    .B1(net5259),
    .B2(\soc_inst.cpu_core.register_file.registers[28][31] ),
    .A2(net5860),
    .A1(\soc_inst.cpu_core.register_file.registers[19][31] ));
 sg13g2_a22oi_1 _18453_ (.Y(_04203_),
    .B1(net5470),
    .B2(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .A2(net5870),
    .A1(\soc_inst.cpu_core.register_file.registers[31][31] ));
 sg13g2_a22oi_1 _18454_ (.Y(_04204_),
    .B1(net5864),
    .B2(\soc_inst.cpu_core.register_file.registers[23][31] ),
    .A2(net5874),
    .A1(\soc_inst.cpu_core.register_file.registers[4][31] ));
 sg13g2_nand3_1 _18455_ (.B(_04203_),
    .C(_04204_),
    .A(_04202_),
    .Y(_04205_));
 sg13g2_a221oi_1 _18456_ (.B2(\soc_inst.cpu_core.register_file.registers[27][31] ),
    .C1(_04205_),
    .B1(net5809),
    .A1(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .Y(_04206_),
    .A2(net5849));
 sg13g2_a22oi_1 _18457_ (.Y(_04207_),
    .B1(net5804),
    .B2(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .A2(net5833),
    .A1(\soc_inst.cpu_core.register_file.registers[14][31] ));
 sg13g2_a221oi_1 _18458_ (.B2(\soc_inst.cpu_core.register_file.registers[21][31] ),
    .C1(_04197_),
    .B1(net5270),
    .A1(\soc_inst.cpu_core.register_file.registers[25][31] ),
    .Y(_04208_),
    .A2(net5289));
 sg13g2_nand4_1 _18459_ (.B(_04206_),
    .C(_04207_),
    .A(_04198_),
    .Y(_04209_),
    .D(_04208_));
 sg13g2_a21oi_1 _18460_ (.A1(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .A2(net5785),
    .Y(_04210_),
    .B1(net6079));
 sg13g2_a22oi_1 _18461_ (.Y(_04211_),
    .B1(net5815),
    .B2(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .A2(net5844),
    .A1(\soc_inst.cpu_core.register_file.registers[26][31] ));
 sg13g2_a22oi_1 _18462_ (.Y(_04212_),
    .B1(net5839),
    .B2(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .A2(net5284),
    .A1(\soc_inst.cpu_core.register_file.registers[16][31] ));
 sg13g2_nand4_1 _18463_ (.B(_04210_),
    .C(_04211_),
    .A(_04201_),
    .Y(_04213_),
    .D(_04212_));
 sg13g2_a22oi_1 _18464_ (.Y(_04214_),
    .B1(net5819),
    .B2(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .A2(net5273),
    .A1(\soc_inst.cpu_core.register_file.registers[17][31] ));
 sg13g2_a22oi_1 _18465_ (.Y(_04215_),
    .B1(net5789),
    .B2(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .A2(net5279),
    .A1(\soc_inst.cpu_core.register_file.registers[20][31] ));
 sg13g2_nand4_1 _18466_ (.B(_04200_),
    .C(_04214_),
    .A(_04199_),
    .Y(_04216_),
    .D(_04215_));
 sg13g2_nor3_2 _18467_ (.A(_04209_),
    .B(_04213_),
    .C(_04216_),
    .Y(_04217_));
 sg13g2_a21oi_1 _18468_ (.A1(net555),
    .A2(net5104),
    .Y(_04218_),
    .B1(net5292));
 sg13g2_or2_1 _18469_ (.X(_04219_),
    .B(_04218_),
    .A(_04217_));
 sg13g2_o21ai_1 _18470_ (.B1(_04219_),
    .Y(_01087_),
    .A1(net6150),
    .A2(_08056_));
 sg13g2_and2_1 _18471_ (.A(_00254_),
    .B(\soc_inst.cpu_core.if_instr[5] ),
    .X(_04220_));
 sg13g2_nor2_1 _18472_ (.A(_00253_),
    .B(_00252_),
    .Y(_04221_));
 sg13g2_nor4_2 _18473_ (.A(net2013),
    .B(net1886),
    .C(net3065),
    .Y(_04222_),
    .D(net2936));
 sg13g2_and2_1 _18474_ (.A(net6140),
    .B(_04222_),
    .X(_04223_));
 sg13g2_nand2_2 _18475_ (.Y(_04224_),
    .A(net6140),
    .B(_04222_));
 sg13g2_and2_1 _18476_ (.A(_04220_),
    .B(_04222_),
    .X(_04225_));
 sg13g2_and2_1 _18477_ (.A(net6140),
    .B(net5775),
    .X(_04226_));
 sg13g2_and4_1 _18478_ (.A(\soc_inst.cpu_core.if_instr[2] ),
    .B(net6451),
    .C(_04220_),
    .D(_04221_),
    .X(_04227_));
 sg13g2_nand4_1 _18479_ (.B(net6451),
    .C(_04220_),
    .A(\soc_inst.cpu_core.if_instr[2] ),
    .Y(_04228_),
    .D(_04221_));
 sg13g2_o21ai_1 _18480_ (.B1(_04228_),
    .Y(_04229_),
    .A1(\soc_inst.cpu_core.if_instr[5] ),
    .A2(net5779));
 sg13g2_nor2b_2 _18481_ (.A(\soc_inst.cpu_core.if_instr[3] ),
    .B_N(_04229_),
    .Y(_04230_));
 sg13g2_inv_1 _18482_ (.Y(_04231_),
    .A(_04230_));
 sg13g2_a22oi_1 _18483_ (.Y(_04232_),
    .B1(_04230_),
    .B2(net6438),
    .A2(_04226_),
    .A1(net1906));
 sg13g2_inv_1 _18484_ (.Y(_04233_),
    .A(_04232_));
 sg13g2_a22oi_1 _18485_ (.Y(_04234_),
    .B1(net5305),
    .B2(_04233_),
    .A2(net3047),
    .A1(net6377));
 sg13g2_inv_1 _18486_ (.Y(_01088_),
    .A(_04234_));
 sg13g2_a22oi_1 _18487_ (.Y(_04235_),
    .B1(_04229_),
    .B2(net6436),
    .A2(net5775),
    .A1(net1270));
 sg13g2_inv_1 _18488_ (.Y(_04236_),
    .A(_04235_));
 sg13g2_a22oi_1 _18489_ (.Y(_04237_),
    .B1(net5305),
    .B2(_04236_),
    .A2(net3098),
    .A1(net6377));
 sg13g2_inv_1 _18490_ (.Y(_01089_),
    .A(_04237_));
 sg13g2_a22oi_1 _18491_ (.Y(_04238_),
    .B1(_04229_),
    .B2(net6435),
    .A2(_04225_),
    .A1(net1265));
 sg13g2_inv_1 _18492_ (.Y(_04239_),
    .A(_04238_));
 sg13g2_a22oi_1 _18493_ (.Y(_04240_),
    .B1(net5305),
    .B2(_04239_),
    .A2(net3099),
    .A1(net6377));
 sg13g2_inv_1 _18494_ (.Y(_01090_),
    .A(_04240_));
 sg13g2_nand3_1 _18495_ (.B(net5309),
    .C(_04229_),
    .A(net6433),
    .Y(_04241_));
 sg13g2_nand3_1 _18496_ (.B(net5306),
    .C(net5775),
    .A(net873),
    .Y(_04242_));
 sg13g2_and2_1 _18497_ (.A(_04241_),
    .B(_04242_),
    .X(_04243_));
 sg13g2_o21ai_1 _18498_ (.B1(_04243_),
    .Y(_01091_),
    .A1(net6152),
    .A2(_08086_));
 sg13g2_nand3_1 _18499_ (.B(net5305),
    .C(_04229_),
    .A(net6431),
    .Y(_04244_));
 sg13g2_nand3_1 _18500_ (.B(net5306),
    .C(net5775),
    .A(net1248),
    .Y(_04245_));
 sg13g2_and2_1 _18501_ (.A(_04244_),
    .B(_04245_),
    .X(_04246_));
 sg13g2_o21ai_1 _18502_ (.B1(_04246_),
    .Y(_01092_),
    .A1(net6153),
    .A2(_08088_));
 sg13g2_or2_1 _18503_ (.X(_04247_),
    .B(_04229_),
    .A(net5775));
 sg13g2_inv_1 _18504_ (.Y(_04248_),
    .A(_04247_));
 sg13g2_nand3_1 _18505_ (.B(net5309),
    .C(_04247_),
    .A(net2838),
    .Y(_04249_));
 sg13g2_o21ai_1 _18506_ (.B1(_04249_),
    .Y(_01093_),
    .A1(net6153),
    .A2(_08090_));
 sg13g2_nand3_1 _18507_ (.B(net5309),
    .C(_04247_),
    .A(\soc_inst.cpu_core.if_funct7[1] ),
    .Y(_04250_));
 sg13g2_o21ai_1 _18508_ (.B1(_04250_),
    .Y(_01094_),
    .A1(net6152),
    .A2(_08092_));
 sg13g2_nand3_1 _18509_ (.B(net5308),
    .C(_04247_),
    .A(net2649),
    .Y(_04251_));
 sg13g2_o21ai_1 _18510_ (.B1(_04251_),
    .Y(_01095_),
    .A1(net6154),
    .A2(_08094_));
 sg13g2_nand3_1 _18511_ (.B(net5308),
    .C(_04247_),
    .A(net3159),
    .Y(_04252_));
 sg13g2_o21ai_1 _18512_ (.B1(_04252_),
    .Y(_01096_),
    .A1(net6155),
    .A2(_08096_));
 sg13g2_nand3_1 _18513_ (.B(net5308),
    .C(_04247_),
    .A(net2729),
    .Y(_04253_));
 sg13g2_o21ai_1 _18514_ (.B1(_04253_),
    .Y(_01097_),
    .A1(net6155),
    .A2(_08098_));
 sg13g2_nand3_1 _18515_ (.B(net5308),
    .C(_04247_),
    .A(net2743),
    .Y(_04254_));
 sg13g2_o21ai_1 _18516_ (.B1(_04254_),
    .Y(_01098_),
    .A1(net6155),
    .A2(_08100_));
 sg13g2_nor2_1 _18517_ (.A(_04226_),
    .B(_04230_),
    .Y(_04255_));
 sg13g2_nor2_1 _18518_ (.A(\soc_inst.cpu_core.if_funct7[6] ),
    .B(_04255_),
    .Y(_04256_));
 sg13g2_and2_1 _18519_ (.A(\soc_inst.cpu_core.if_instr[3] ),
    .B(_04227_),
    .X(_04257_));
 sg13g2_nand2_2 _18520_ (.Y(_04258_),
    .A(\soc_inst.cpu_core.if_instr[3] ),
    .B(_04227_));
 sg13g2_and2_1 _18521_ (.A(net6451),
    .B(net5775),
    .X(_04259_));
 sg13g2_a22oi_1 _18522_ (.Y(_04260_),
    .B1(_04259_),
    .B2(net1906),
    .A2(net5466),
    .A1(net6438));
 sg13g2_a21oi_1 _18523_ (.A1(_04255_),
    .A2(_04260_),
    .Y(_04261_),
    .B1(_04256_));
 sg13g2_inv_1 _18524_ (.Y(_04262_),
    .A(_04261_));
 sg13g2_a22oi_1 _18525_ (.Y(_04263_),
    .B1(net5305),
    .B2(_04261_),
    .A2(net3274),
    .A1(net6413));
 sg13g2_inv_1 _18526_ (.Y(_01099_),
    .A(net3275));
 sg13g2_nor3_1 _18527_ (.A(_00254_),
    .B(\soc_inst.cpu_core.if_instr[3] ),
    .C(net6451),
    .Y(_04264_));
 sg13g2_nand3_1 _18528_ (.B(_04221_),
    .C(_04264_),
    .A(\soc_inst.cpu_core.if_instr[2] ),
    .Y(_04265_));
 sg13g2_nand2_1 _18529_ (.Y(_04266_),
    .A(_04258_),
    .B(_04265_));
 sg13g2_nand2_1 _18530_ (.Y(_04267_),
    .A(net3014),
    .B(net5250));
 sg13g2_a21oi_2 _18531_ (.B1(_04230_),
    .Y(_04268_),
    .A2(net5775),
    .A1(\soc_inst.cpu_core.if_funct7[6] ));
 sg13g2_o21ai_1 _18532_ (.B1(net5308),
    .Y(_04269_),
    .A1(\soc_inst.cpu_core.if_funct7[6] ),
    .A2(_04231_));
 sg13g2_a21oi_1 _18533_ (.A1(_04267_),
    .A2(_04268_),
    .Y(_04270_),
    .B1(_04269_));
 sg13g2_a21o_1 _18534_ (.A2(net3200),
    .A1(net6391),
    .B1(_04270_),
    .X(_01100_));
 sg13g2_nand2_1 _18535_ (.Y(_04271_),
    .A(\soc_inst.cpu_core.if_funct3[1] ),
    .B(net5250));
 sg13g2_a21oi_1 _18536_ (.A1(_04268_),
    .A2(_04271_),
    .Y(_04272_),
    .B1(_04269_));
 sg13g2_a21o_1 _18537_ (.A2(net2906),
    .A1(net6388),
    .B1(_04272_),
    .X(_01101_));
 sg13g2_nand2_1 _18538_ (.Y(_04273_),
    .A(net2945),
    .B(net5250));
 sg13g2_a21oi_1 _18539_ (.A1(_04268_),
    .A2(_04273_),
    .Y(_04274_),
    .B1(_04269_));
 sg13g2_a21o_1 _18540_ (.A2(net3183),
    .A1(net6389),
    .B1(_04274_),
    .X(_01102_));
 sg13g2_nand2_1 _18541_ (.Y(_04275_),
    .A(net6450),
    .B(net5250));
 sg13g2_a21oi_1 _18542_ (.A1(_04268_),
    .A2(_04275_),
    .Y(_04276_),
    .B1(_04269_));
 sg13g2_a21o_1 _18543_ (.A2(net3241),
    .A1(net6391),
    .B1(_04276_),
    .X(_01103_));
 sg13g2_nand2_1 _18544_ (.Y(_04277_),
    .A(net6448),
    .B(net5250));
 sg13g2_a21oi_2 _18545_ (.B1(_04269_),
    .Y(_04278_),
    .A2(_04277_),
    .A1(_04268_));
 sg13g2_a21o_1 _18546_ (.A2(net3293),
    .A1(net6397),
    .B1(_04278_),
    .X(_01104_));
 sg13g2_nand2_1 _18547_ (.Y(_04279_),
    .A(net6445),
    .B(net5250));
 sg13g2_a21oi_2 _18548_ (.B1(_04269_),
    .Y(_04280_),
    .A2(_04279_),
    .A1(_04268_));
 sg13g2_a21o_1 _18549_ (.A2(net3234),
    .A1(net6386),
    .B1(_04280_),
    .X(_01105_));
 sg13g2_nand2_1 _18550_ (.Y(_04281_),
    .A(net6444),
    .B(net5250));
 sg13g2_a21oi_2 _18551_ (.B1(_04269_),
    .Y(_04282_),
    .A2(_04281_),
    .A1(_04268_));
 sg13g2_a21o_1 _18552_ (.A2(net3126),
    .A1(net6386),
    .B1(_04282_),
    .X(_01106_));
 sg13g2_nand2_1 _18553_ (.Y(_04283_),
    .A(net6443),
    .B(_04266_));
 sg13g2_a21oi_2 _18554_ (.B1(_04269_),
    .Y(_04284_),
    .A2(_04283_),
    .A1(_04268_));
 sg13g2_a21o_1 _18555_ (.A2(net3103),
    .A1(net6386),
    .B1(_04284_),
    .X(_01107_));
 sg13g2_o21ai_1 _18556_ (.B1(\soc_inst.cpu_core.if_funct7[6] ),
    .Y(_04285_),
    .A1(net5775),
    .A2(_04230_));
 sg13g2_nor2_1 _18557_ (.A(net6438),
    .B(net5466),
    .Y(_04286_));
 sg13g2_o21ai_1 _18558_ (.B1(net5250),
    .Y(_04287_),
    .A1(\soc_inst.cpu_core.if_funct7[6] ),
    .A2(_04258_));
 sg13g2_o21ai_1 _18559_ (.B1(net5101),
    .Y(_04288_),
    .A1(_04286_),
    .A2(net5099));
 sg13g2_a22oi_1 _18560_ (.Y(_04289_),
    .B1(net5302),
    .B2(_04288_),
    .A2(net3201),
    .A1(net6382));
 sg13g2_inv_1 _18561_ (.Y(_01108_),
    .A(_04289_));
 sg13g2_nor2_1 _18562_ (.A(net6436),
    .B(net5465),
    .Y(_04290_));
 sg13g2_o21ai_1 _18563_ (.B1(net5100),
    .Y(_04291_),
    .A1(net5098),
    .A2(_04290_));
 sg13g2_a22oi_1 _18564_ (.Y(_04292_),
    .B1(net5301),
    .B2(_04291_),
    .A2(net3277),
    .A1(net6385));
 sg13g2_inv_1 _18565_ (.Y(_01109_),
    .A(_04292_));
 sg13g2_nor2_1 _18566_ (.A(net6435),
    .B(net5465),
    .Y(_04293_));
 sg13g2_o21ai_1 _18567_ (.B1(net5100),
    .Y(_04294_),
    .A1(net5098),
    .A2(_04293_));
 sg13g2_a22oi_1 _18568_ (.Y(_04295_),
    .B1(net5301),
    .B2(_04294_),
    .A2(net3060),
    .A1(net6385));
 sg13g2_inv_1 _18569_ (.Y(_01110_),
    .A(_04295_));
 sg13g2_nor2_1 _18570_ (.A(net6433),
    .B(net5465),
    .Y(_04296_));
 sg13g2_o21ai_1 _18571_ (.B1(net5100),
    .Y(_04297_),
    .A1(net5098),
    .A2(_04296_));
 sg13g2_a22oi_1 _18572_ (.Y(_04298_),
    .B1(net5301),
    .B2(_04297_),
    .A2(net3202),
    .A1(net6398));
 sg13g2_inv_1 _18573_ (.Y(_01111_),
    .A(_04298_));
 sg13g2_nor2_1 _18574_ (.A(net6431),
    .B(net5465),
    .Y(_04299_));
 sg13g2_o21ai_1 _18575_ (.B1(net5100),
    .Y(_04300_),
    .A1(net5098),
    .A2(_04299_));
 sg13g2_a22oi_1 _18576_ (.Y(_04301_),
    .B1(net5301),
    .B2(_04300_),
    .A2(net3169),
    .A1(net6385));
 sg13g2_inv_1 _18577_ (.Y(_01112_),
    .A(_04301_));
 sg13g2_nor2_1 _18578_ (.A(\soc_inst.cpu_core.if_funct7[0] ),
    .B(net5465),
    .Y(_04302_));
 sg13g2_o21ai_1 _18579_ (.B1(net5100),
    .Y(_04303_),
    .A1(net5098),
    .A2(_04302_));
 sg13g2_a22oi_1 _18580_ (.Y(_04304_),
    .B1(net5301),
    .B2(_04303_),
    .A2(net3062),
    .A1(net6385));
 sg13g2_inv_1 _18581_ (.Y(_01113_),
    .A(_04304_));
 sg13g2_nor2_1 _18582_ (.A(\soc_inst.cpu_core.if_funct7[1] ),
    .B(net5465),
    .Y(_04305_));
 sg13g2_o21ai_1 _18583_ (.B1(net5100),
    .Y(_04306_),
    .A1(net5098),
    .A2(_04305_));
 sg13g2_a22oi_1 _18584_ (.Y(_04307_),
    .B1(net5301),
    .B2(_04306_),
    .A2(net3249),
    .A1(net6385));
 sg13g2_inv_1 _18585_ (.Y(_01114_),
    .A(_04307_));
 sg13g2_nor2_1 _18586_ (.A(\soc_inst.cpu_core.if_funct7[2] ),
    .B(net5465),
    .Y(_04308_));
 sg13g2_o21ai_1 _18587_ (.B1(net5100),
    .Y(_04309_),
    .A1(net5098),
    .A2(_04308_));
 sg13g2_a22oi_1 _18588_ (.Y(_04310_),
    .B1(net5301),
    .B2(_04309_),
    .A2(net3257),
    .A1(net6385));
 sg13g2_inv_1 _18589_ (.Y(_01115_),
    .A(net3258));
 sg13g2_nor2_1 _18590_ (.A(net3408),
    .B(net5465),
    .Y(_04311_));
 sg13g2_o21ai_1 _18591_ (.B1(net5100),
    .Y(_04312_),
    .A1(net5098),
    .A2(_04311_));
 sg13g2_a22oi_1 _18592_ (.Y(_04313_),
    .B1(net5302),
    .B2(_04312_),
    .A2(net3048),
    .A1(net6394));
 sg13g2_inv_1 _18593_ (.Y(_01116_),
    .A(_04313_));
 sg13g2_nor2_1 _18594_ (.A(\soc_inst.cpu_core.if_funct7[4] ),
    .B(net5466),
    .Y(_04314_));
 sg13g2_o21ai_1 _18595_ (.B1(net5101),
    .Y(_04315_),
    .A1(net5099),
    .A2(_04314_));
 sg13g2_a22oi_1 _18596_ (.Y(_04316_),
    .B1(net5302),
    .B2(_04315_),
    .A2(net3144),
    .A1(net6394));
 sg13g2_inv_1 _18597_ (.Y(_01117_),
    .A(_04316_));
 sg13g2_nor2_1 _18598_ (.A(\soc_inst.cpu_core.if_funct7[5] ),
    .B(net5466),
    .Y(_04317_));
 sg13g2_o21ai_1 _18599_ (.B1(net5101),
    .Y(_04318_),
    .A1(net5099),
    .A2(_04317_));
 sg13g2_a22oi_1 _18600_ (.Y(_04319_),
    .B1(net5302),
    .B2(_04318_),
    .A2(net2961),
    .A1(net6393));
 sg13g2_inv_1 _18601_ (.Y(_01118_),
    .A(net2962));
 sg13g2_a21oi_2 _18602_ (.B1(_02608_),
    .Y(_04320_),
    .A2(_04265_),
    .A1(_04248_));
 sg13g2_a21o_1 _18603_ (.A2(net2665),
    .A1(net6393),
    .B1(_04320_),
    .X(_01119_));
 sg13g2_nor2_1 _18604_ (.A(net6417),
    .B(_07933_),
    .Y(_04321_));
 sg13g2_a22oi_1 _18605_ (.Y(_04322_),
    .B1(net5007),
    .B2(_04321_),
    .A2(net3296),
    .A1(net6417));
 sg13g2_inv_1 _18606_ (.Y(_01120_),
    .A(_04322_));
 sg13g2_nand2_1 _18607_ (.Y(_04323_),
    .A(net6417),
    .B(net6288));
 sg13g2_nor2_2 _18608_ (.A(net2877),
    .B(net5779),
    .Y(_04324_));
 sg13g2_nor3_1 _18609_ (.A(net2877),
    .B(net3014),
    .C(net5779),
    .Y(_04325_));
 sg13g2_nand2_1 _18610_ (.Y(_04326_),
    .A(net2877),
    .B(_04223_));
 sg13g2_nand4_1 _18611_ (.B(_04228_),
    .C(_04265_),
    .A(net5309),
    .Y(_04327_),
    .D(_04326_));
 sg13g2_o21ai_1 _18612_ (.B1(_04323_),
    .Y(_01121_),
    .A1(_04325_),
    .A2(_04327_));
 sg13g2_a21oi_1 _18613_ (.A1(_08134_),
    .A2(_04324_),
    .Y(_04328_),
    .B1(_04327_));
 sg13g2_a21o_1 _18614_ (.A2(net3312),
    .A1(net6417),
    .B1(_04328_),
    .X(_01122_));
 sg13g2_nor3_1 _18615_ (.A(net2877),
    .B(net2945),
    .C(net5779),
    .Y(_04329_));
 sg13g2_nand2_1 _18616_ (.Y(_04330_),
    .A(net6417),
    .B(net3085));
 sg13g2_o21ai_1 _18617_ (.B1(_04330_),
    .Y(_01123_),
    .A1(_04327_),
    .A2(_04329_));
 sg13g2_nand2_2 _18618_ (.Y(_04331_),
    .A(net3174),
    .B(_04324_));
 sg13g2_nand4_1 _18619_ (.B(net3014),
    .C(_08134_),
    .A(net2743),
    .Y(_04332_),
    .D(net2945));
 sg13g2_a21oi_1 _18620_ (.A1(_04324_),
    .A2(_04332_),
    .Y(_04333_),
    .B1(_04327_));
 sg13g2_a21oi_1 _18621_ (.A1(net6417),
    .A2(net6285),
    .Y(_04334_),
    .B1(_04333_));
 sg13g2_o21ai_1 _18622_ (.B1(_04334_),
    .Y(_01124_),
    .A1(_11771_),
    .A2(net5248));
 sg13g2_o21ai_1 _18623_ (.B1(_04228_),
    .Y(_04335_),
    .A1(\soc_inst.cpu_core.if_instr[5] ),
    .A2(_04265_));
 sg13g2_nand2_1 _18624_ (.Y(_04336_),
    .A(net2809),
    .B(net5463));
 sg13g2_nand2_2 _18625_ (.Y(_04337_),
    .A(net5310),
    .B(net5779));
 sg13g2_a22oi_1 _18626_ (.Y(_04338_),
    .B1(net5097),
    .B2(_02677_),
    .A2(_04336_),
    .A1(net5780));
 sg13g2_a21o_1 _18627_ (.A2(net3136),
    .A1(net6423),
    .B1(_04338_),
    .X(_01125_));
 sg13g2_a21oi_1 _18628_ (.A1(net2093),
    .A2(net5464),
    .Y(_04339_),
    .B1(_04223_));
 sg13g2_nor2b_1 _18629_ (.A(_02701_),
    .B_N(net5097),
    .Y(_04340_));
 sg13g2_nand2_1 _18630_ (.Y(_04341_),
    .A(net6417),
    .B(net2926));
 sg13g2_o21ai_1 _18631_ (.B1(_04341_),
    .Y(_01126_),
    .A1(_04339_),
    .A2(_04340_));
 sg13g2_a21oi_1 _18632_ (.A1(net1316),
    .A2(net5464),
    .Y(_04342_),
    .B1(_04223_));
 sg13g2_nor2b_1 _18633_ (.A(_02725_),
    .B_N(net5097),
    .Y(_04343_));
 sg13g2_nand2_1 _18634_ (.Y(_04344_),
    .A(net6419),
    .B(net2035));
 sg13g2_o21ai_1 _18635_ (.B1(_04344_),
    .Y(_01127_),
    .A1(_04342_),
    .A2(_04343_));
 sg13g2_nand2_1 _18636_ (.Y(_04345_),
    .A(net2324),
    .B(net5463));
 sg13g2_a22oi_1 _18637_ (.Y(_04346_),
    .B1(_04345_),
    .B2(net5780),
    .A2(_04337_),
    .A1(_02749_));
 sg13g2_a21o_1 _18638_ (.A2(net2884),
    .A1(net6424),
    .B1(_04346_),
    .X(_01128_));
 sg13g2_nand2_1 _18639_ (.Y(_04347_),
    .A(net2046),
    .B(net5463));
 sg13g2_a22oi_1 _18640_ (.Y(_04348_),
    .B1(_04347_),
    .B2(net5779),
    .A2(_04337_),
    .A1(_02773_));
 sg13g2_a21o_1 _18641_ (.A2(net3019),
    .A1(net6422),
    .B1(_04348_),
    .X(_01129_));
 sg13g2_nand2_1 _18642_ (.Y(_04349_),
    .A(net1748),
    .B(net5463));
 sg13g2_a22oi_1 _18643_ (.Y(_04350_),
    .B1(_04349_),
    .B2(net5780),
    .A2(net5097),
    .A1(_02797_));
 sg13g2_a21o_1 _18644_ (.A2(net3088),
    .A1(net6418),
    .B1(_04350_),
    .X(_01130_));
 sg13g2_a21oi_1 _18645_ (.A1(net1946),
    .A2(net5464),
    .Y(_04351_),
    .B1(_04223_));
 sg13g2_a21o_1 _18646_ (.A2(net5097),
    .A1(_02821_),
    .B1(_04351_),
    .X(_04352_));
 sg13g2_o21ai_1 _18647_ (.B1(_04352_),
    .Y(_01131_),
    .A1(net6154),
    .A2(_08205_));
 sg13g2_nand2_1 _18648_ (.Y(_04353_),
    .A(net2271),
    .B(net5464));
 sg13g2_a22oi_1 _18649_ (.Y(_04354_),
    .B1(_04353_),
    .B2(net5779),
    .A2(_04337_),
    .A1(_02845_));
 sg13g2_a21o_1 _18650_ (.A2(net3145),
    .A1(net6419),
    .B1(_04354_),
    .X(_01132_));
 sg13g2_nand2_1 _18651_ (.Y(_04355_),
    .A(net2258),
    .B(net5463));
 sg13g2_a22oi_1 _18652_ (.Y(_04356_),
    .B1(_04355_),
    .B2(net5780),
    .A2(net5097),
    .A1(_02869_));
 sg13g2_a21o_1 _18653_ (.A2(net6284),
    .A1(net6409),
    .B1(_04356_),
    .X(_01133_));
 sg13g2_nor2b_1 _18654_ (.A(_11390_),
    .B_N(net5463),
    .Y(_04357_));
 sg13g2_nor2_2 _18655_ (.A(net6405),
    .B(_07918_),
    .Y(_04358_));
 sg13g2_a22oi_1 _18656_ (.Y(_04359_),
    .B1(net5244),
    .B2(_04358_),
    .A2(net3332),
    .A1(net6411));
 sg13g2_o21ai_1 _18657_ (.B1(_04359_),
    .Y(_01134_),
    .A1(_02893_),
    .A2(net5780));
 sg13g2_nor2_2 _18658_ (.A(net6409),
    .B(_07919_),
    .Y(_04360_));
 sg13g2_a22oi_1 _18659_ (.Y(_04361_),
    .B1(net5244),
    .B2(_04360_),
    .A2(net3309),
    .A1(net6410));
 sg13g2_o21ai_1 _18660_ (.B1(_04361_),
    .Y(_01135_),
    .A1(_02917_),
    .A2(net5780));
 sg13g2_nor2_2 _18661_ (.A(net6409),
    .B(_07920_),
    .Y(_04362_));
 sg13g2_a22oi_1 _18662_ (.Y(_04363_),
    .B1(net5244),
    .B2(_04362_),
    .A2(net3342),
    .A1(net6409));
 sg13g2_o21ai_1 _18663_ (.B1(_04363_),
    .Y(_01136_),
    .A1(_02941_),
    .A2(net5780));
 sg13g2_nor2_2 _18664_ (.A(net6351),
    .B(_07921_),
    .Y(_04364_));
 sg13g2_a22oi_1 _18665_ (.Y(_04365_),
    .B1(net5244),
    .B2(_04364_),
    .A2(net3290),
    .A1(net6396));
 sg13g2_o21ai_1 _18666_ (.B1(_04365_),
    .Y(_01137_),
    .A1(_02965_),
    .A2(net5778));
 sg13g2_nor2_2 _18667_ (.A(net6348),
    .B(_07922_),
    .Y(_04366_));
 sg13g2_a22oi_1 _18668_ (.Y(_04367_),
    .B1(net5243),
    .B2(_04366_),
    .A2(net3361),
    .A1(net6394));
 sg13g2_o21ai_1 _18669_ (.B1(_04367_),
    .Y(_01138_),
    .A1(_02989_),
    .A2(net5778));
 sg13g2_nor2_2 _18670_ (.A(net6348),
    .B(_07923_),
    .Y(_04368_));
 sg13g2_a22oi_1 _18671_ (.Y(_04369_),
    .B1(net5244),
    .B2(_04368_),
    .A2(net6283),
    .A1(net6393));
 sg13g2_o21ai_1 _18672_ (.B1(_04369_),
    .Y(_01139_),
    .A1(_03013_),
    .A2(net5778));
 sg13g2_nor2_2 _18673_ (.A(net6348),
    .B(_07924_),
    .Y(_04370_));
 sg13g2_a22oi_1 _18674_ (.Y(_04371_),
    .B1(net5243),
    .B2(_04370_),
    .A2(net3354),
    .A1(net6393));
 sg13g2_o21ai_1 _18675_ (.B1(_04371_),
    .Y(_01140_),
    .A1(_03037_),
    .A2(net5778));
 sg13g2_nor2_2 _18676_ (.A(net6343),
    .B(_07925_),
    .Y(_04372_));
 sg13g2_a22oi_1 _18677_ (.Y(_04373_),
    .B1(net5243),
    .B2(_04372_),
    .A2(net6282),
    .A1(net6397));
 sg13g2_o21ai_1 _18678_ (.B1(_04373_),
    .Y(_01141_),
    .A1(_03061_),
    .A2(net5776));
 sg13g2_nor2_2 _18679_ (.A(net6342),
    .B(_07926_),
    .Y(_04374_));
 sg13g2_a22oi_1 _18680_ (.Y(_04375_),
    .B1(net5243),
    .B2(_04374_),
    .A2(net6280),
    .A1(net6397));
 sg13g2_o21ai_1 _18681_ (.B1(_04375_),
    .Y(_01142_),
    .A1(_03085_),
    .A2(net5776));
 sg13g2_nor2_2 _18682_ (.A(net6343),
    .B(_07927_),
    .Y(_04376_));
 sg13g2_a22oi_1 _18683_ (.Y(_04377_),
    .B1(net5243),
    .B2(_04376_),
    .A2(net6278),
    .A1(net6397));
 sg13g2_o21ai_1 _18684_ (.B1(_04377_),
    .Y(_01143_),
    .A1(_03109_),
    .A2(net5776));
 sg13g2_nor2_2 _18685_ (.A(net6342),
    .B(_07928_),
    .Y(_04378_));
 sg13g2_a22oi_1 _18686_ (.Y(_04379_),
    .B1(net5243),
    .B2(_04378_),
    .A2(net6276),
    .A1(net6397));
 sg13g2_o21ai_1 _18687_ (.B1(_04379_),
    .Y(_01144_),
    .A1(_03133_),
    .A2(net5776));
 sg13g2_nor2_2 _18688_ (.A(net6345),
    .B(_07929_),
    .Y(_04380_));
 sg13g2_a22oi_1 _18689_ (.Y(_04381_),
    .B1(net5243),
    .B2(_04380_),
    .A2(net6274),
    .A1(net6399));
 sg13g2_o21ai_1 _18690_ (.B1(_04381_),
    .Y(_01145_),
    .A1(_03156_),
    .A2(net5776));
 sg13g2_a21oi_1 _18691_ (.A1(net2078),
    .A2(net5463),
    .Y(_04382_),
    .B1(_04223_));
 sg13g2_nor2b_1 _18692_ (.A(_03180_),
    .B_N(net5097),
    .Y(_04383_));
 sg13g2_nand2_1 _18693_ (.Y(_04384_),
    .A(net6396),
    .B(net6272));
 sg13g2_o21ai_1 _18694_ (.B1(_04384_),
    .Y(_01146_),
    .A1(_04382_),
    .A2(_04383_));
 sg13g2_nor2_2 _18695_ (.A(net6345),
    .B(_07931_),
    .Y(_04385_));
 sg13g2_a22oi_1 _18696_ (.Y(_04386_),
    .B1(net5243),
    .B2(_04385_),
    .A2(net6271),
    .A1(net6398));
 sg13g2_o21ai_1 _18697_ (.B1(_04386_),
    .Y(_01147_),
    .A1(_03204_),
    .A2(net5776));
 sg13g2_nand2_1 _18698_ (.Y(_04387_),
    .A(net2947),
    .B(net5463));
 sg13g2_a22oi_1 _18699_ (.Y(_04388_),
    .B1(_04387_),
    .B2(net5778),
    .A2(net5097),
    .A1(_03228_));
 sg13g2_a21o_1 _18700_ (.A2(net6270),
    .A1(net6402),
    .B1(_04388_),
    .X(_01148_));
 sg13g2_nand2_1 _18701_ (.Y(_04389_),
    .A(net6400),
    .B(net6269));
 sg13g2_o21ai_1 _18702_ (.B1(_04389_),
    .Y(_01149_),
    .A1(_03252_),
    .A2(net5776));
 sg13g2_nand2_1 _18703_ (.Y(_04390_),
    .A(net6400),
    .B(net6268));
 sg13g2_o21ai_1 _18704_ (.B1(_04390_),
    .Y(_01150_),
    .A1(_03276_),
    .A2(net5777));
 sg13g2_nand2_1 _18705_ (.Y(_04391_),
    .A(net6400),
    .B(net6266));
 sg13g2_o21ai_1 _18706_ (.B1(_04391_),
    .Y(_01151_),
    .A1(_03300_),
    .A2(net5777));
 sg13g2_nand2_1 _18707_ (.Y(_04392_),
    .A(net6401),
    .B(net6265));
 sg13g2_o21ai_1 _18708_ (.B1(_04392_),
    .Y(_01152_),
    .A1(_03324_),
    .A2(net5777));
 sg13g2_nand2_1 _18709_ (.Y(_04393_),
    .A(net6401),
    .B(net6264));
 sg13g2_o21ai_1 _18710_ (.B1(_04393_),
    .Y(_01153_),
    .A1(_03348_),
    .A2(net5777));
 sg13g2_a22oi_1 _18711_ (.Y(_04394_),
    .B1(_03372_),
    .B2(_04223_),
    .A2(net3077),
    .A1(net6426));
 sg13g2_inv_1 _18712_ (.Y(_01154_),
    .A(_04394_));
 sg13g2_nand2_1 _18713_ (.Y(_04395_),
    .A(net6425),
    .B(net3294));
 sg13g2_o21ai_1 _18714_ (.B1(_04395_),
    .Y(_01155_),
    .A1(_03396_),
    .A2(_04224_));
 sg13g2_nand2_1 _18715_ (.Y(_04396_),
    .A(net6400),
    .B(net6262));
 sg13g2_o21ai_1 _18716_ (.B1(_04396_),
    .Y(_01156_),
    .A1(_03419_),
    .A2(net5776));
 sg13g2_and2_1 _18717_ (.A(net5301),
    .B(net5245),
    .X(_04397_));
 sg13g2_o21ai_1 _18718_ (.B1(net5248),
    .Y(_04398_),
    .A1(net2936),
    .A2(_04232_));
 sg13g2_o21ai_1 _18719_ (.B1(_04398_),
    .Y(_04399_),
    .A1(_03493_),
    .A2(net5096));
 sg13g2_o21ai_1 _18720_ (.B1(_04399_),
    .Y(_01157_),
    .A1(net6157),
    .A2(net6112));
 sg13g2_o21ai_1 _18721_ (.B1(_04326_),
    .Y(_04400_),
    .A1(\soc_inst.cpu_core.if_instr[5] ),
    .A2(net5779));
 sg13g2_a22oi_1 _18722_ (.Y(_04401_),
    .B1(_04236_),
    .B2(_04400_),
    .A2(_04227_),
    .A1(net2451));
 sg13g2_nand2_1 _18723_ (.Y(_04402_),
    .A(net5248),
    .B(_04401_));
 sg13g2_o21ai_1 _18724_ (.B1(_04402_),
    .Y(_04403_),
    .A1(_03516_),
    .A2(net5096));
 sg13g2_o21ai_1 _18725_ (.B1(_04403_),
    .Y(_01158_),
    .A1(net6157),
    .A2(net6118));
 sg13g2_nand2_1 _18726_ (.Y(_04404_),
    .A(net6422),
    .B(net6238));
 sg13g2_nor2_1 _18727_ (.A(_03540_),
    .B(net5096),
    .Y(_04405_));
 sg13g2_o21ai_1 _18728_ (.B1(net5249),
    .Y(_04406_),
    .A1(net2451),
    .A2(_04228_));
 sg13g2_a21oi_1 _18729_ (.A1(_04239_),
    .A2(_04400_),
    .Y(_04407_),
    .B1(_04406_));
 sg13g2_o21ai_1 _18730_ (.B1(_04404_),
    .Y(_01159_),
    .A1(_04405_),
    .A2(_04407_));
 sg13g2_nor2_1 _18731_ (.A(net3236),
    .B(_04243_),
    .Y(_04408_));
 sg13g2_a21oi_1 _18732_ (.A1(net6425),
    .A2(net6231),
    .Y(_04409_),
    .B1(_04408_));
 sg13g2_o21ai_1 _18733_ (.B1(_04409_),
    .Y(_01160_),
    .A1(_03563_),
    .A2(net5249));
 sg13g2_nor2_1 _18734_ (.A(net6452),
    .B(_04246_),
    .Y(_04410_));
 sg13g2_a21oi_1 _18735_ (.A1(net6422),
    .A2(net6222),
    .Y(_04411_),
    .B1(_04410_));
 sg13g2_o21ai_1 _18736_ (.B1(_04411_),
    .Y(_01161_),
    .A1(_03586_),
    .A2(net5249));
 sg13g2_nor2_1 _18737_ (.A(net6451),
    .B(_04249_),
    .Y(_04412_));
 sg13g2_a21oi_1 _18738_ (.A1(net6418),
    .A2(net3063),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_o21ai_1 _18739_ (.B1(_04413_),
    .Y(_01162_),
    .A1(_03609_),
    .A2(net5248));
 sg13g2_nor2_1 _18740_ (.A(net6451),
    .B(_04250_),
    .Y(_04414_));
 sg13g2_a21oi_1 _18741_ (.A1(net6418),
    .A2(net2972),
    .Y(_04415_),
    .B1(_04414_));
 sg13g2_o21ai_1 _18742_ (.B1(net2973),
    .Y(_01163_),
    .A1(_03632_),
    .A2(net5249));
 sg13g2_nor2_1 _18743_ (.A(net6452),
    .B(_04251_),
    .Y(_04416_));
 sg13g2_a21oi_1 _18744_ (.A1(net6419),
    .A2(net2943),
    .Y(_04417_),
    .B1(_04416_));
 sg13g2_o21ai_1 _18745_ (.B1(net2944),
    .Y(_01164_),
    .A1(_03655_),
    .A2(net5248));
 sg13g2_nor2_1 _18746_ (.A(net6452),
    .B(_04252_),
    .Y(_04418_));
 sg13g2_a21oi_1 _18747_ (.A1(net6411),
    .A2(net3272),
    .Y(_04419_),
    .B1(_04418_));
 sg13g2_o21ai_1 _18748_ (.B1(_04419_),
    .Y(_01165_),
    .A1(_03678_),
    .A2(net5248));
 sg13g2_nor2_1 _18749_ (.A(net6452),
    .B(_04253_),
    .Y(_04420_));
 sg13g2_a21oi_1 _18750_ (.A1(net6411),
    .A2(net3178),
    .Y(_04421_),
    .B1(_04420_));
 sg13g2_o21ai_1 _18751_ (.B1(net3179),
    .Y(_01166_),
    .A1(_03701_),
    .A2(net5248));
 sg13g2_nor2_1 _18752_ (.A(net6452),
    .B(_04254_),
    .Y(_04422_));
 sg13g2_a21oi_1 _18753_ (.A1(net6409),
    .A2(net2998),
    .Y(_04423_),
    .B1(_04422_));
 sg13g2_o21ai_1 _18754_ (.B1(net2999),
    .Y(_01167_),
    .A1(_03724_),
    .A2(net5248));
 sg13g2_o21ai_1 _18755_ (.B1(net5249),
    .Y(_04424_),
    .A1(net6451),
    .A2(_04262_));
 sg13g2_o21ai_1 _18756_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_03748_),
    .A2(net5096));
 sg13g2_o21ai_1 _18757_ (.B1(_04425_),
    .Y(_01168_),
    .A1(net6156),
    .A2(_08202_));
 sg13g2_a22oi_1 _18758_ (.Y(_04426_),
    .B1(_04270_),
    .B2(net6139),
    .A2(net3040),
    .A1(net6391));
 sg13g2_o21ai_1 _18759_ (.B1(_04426_),
    .Y(_01169_),
    .A1(_03771_),
    .A2(net5247));
 sg13g2_a22oi_1 _18760_ (.Y(_04427_),
    .B1(_04272_),
    .B2(net6139),
    .A2(net3285),
    .A1(net6388));
 sg13g2_o21ai_1 _18761_ (.B1(net3286),
    .Y(_01170_),
    .A1(_03794_),
    .A2(net5247));
 sg13g2_a22oi_1 _18762_ (.Y(_04428_),
    .B1(_04274_),
    .B2(net6139),
    .A2(net3254),
    .A1(net6393));
 sg13g2_o21ai_1 _18763_ (.B1(_04428_),
    .Y(_01171_),
    .A1(_03817_),
    .A2(net5247));
 sg13g2_a22oi_1 _18764_ (.Y(_04429_),
    .B1(_04276_),
    .B2(net6139),
    .A2(net3203),
    .A1(net6395));
 sg13g2_o21ai_1 _18765_ (.B1(_04429_),
    .Y(_01172_),
    .A1(_03840_),
    .A2(net5247));
 sg13g2_a22oi_1 _18766_ (.Y(_04430_),
    .B1(_04278_),
    .B2(net6137),
    .A2(net3351),
    .A1(net6398));
 sg13g2_o21ai_1 _18767_ (.B1(_04430_),
    .Y(_01173_),
    .A1(_03863_),
    .A2(net5245));
 sg13g2_a22oi_1 _18768_ (.Y(_04431_),
    .B1(_04280_),
    .B2(net6137),
    .A2(net3316),
    .A1(net6398));
 sg13g2_o21ai_1 _18769_ (.B1(_04431_),
    .Y(_01174_),
    .A1(_03886_),
    .A2(net5245));
 sg13g2_a22oi_1 _18770_ (.Y(_04432_),
    .B1(_04282_),
    .B2(net6137),
    .A2(net3156),
    .A1(net6398));
 sg13g2_o21ai_1 _18771_ (.B1(_04432_),
    .Y(_01175_),
    .A1(_03909_),
    .A2(net5247));
 sg13g2_a22oi_1 _18772_ (.Y(_04433_),
    .B1(_04284_),
    .B2(net6138),
    .A2(net3320),
    .A1(net6385));
 sg13g2_o21ai_1 _18773_ (.B1(_04433_),
    .Y(_01176_),
    .A1(_03932_),
    .A2(net5247));
 sg13g2_a22oi_1 _18774_ (.Y(_04434_),
    .B1(_04324_),
    .B2(\soc_inst.cpu_core.if_instr[5] ),
    .A2(_04288_),
    .A1(net6140));
 sg13g2_nor2_2 _18775_ (.A(_03956_),
    .B(net5095),
    .Y(_04435_));
 sg13g2_nand2_1 _18776_ (.Y(_04436_),
    .A(net6426),
    .B(net2951));
 sg13g2_o21ai_1 _18777_ (.B1(_04436_),
    .Y(_01177_),
    .A1(_04434_),
    .A2(_04435_));
 sg13g2_nand2_1 _18778_ (.Y(_04437_),
    .A(net6137),
    .B(_04291_));
 sg13g2_nor2_1 _18779_ (.A(_03980_),
    .B(net5095),
    .Y(_04438_));
 sg13g2_a21o_1 _18780_ (.A2(_04437_),
    .A1(net5245),
    .B1(_04438_),
    .X(_04439_));
 sg13g2_o21ai_1 _18781_ (.B1(_04439_),
    .Y(_01178_),
    .A1(net6149),
    .A2(_08194_));
 sg13g2_nand2_1 _18782_ (.Y(_04440_),
    .A(net6137),
    .B(_04294_));
 sg13g2_nor2_1 _18783_ (.A(_04004_),
    .B(net5095),
    .Y(_04441_));
 sg13g2_a21o_1 _18784_ (.A2(_04440_),
    .A1(net5245),
    .B1(_04441_),
    .X(_04442_));
 sg13g2_o21ai_1 _18785_ (.B1(_04442_),
    .Y(_01179_),
    .A1(net6151),
    .A2(_08193_));
 sg13g2_nand2_1 _18786_ (.Y(_04443_),
    .A(net6137),
    .B(_04297_));
 sg13g2_nor2_1 _18787_ (.A(_04028_),
    .B(net5096),
    .Y(_04444_));
 sg13g2_a21o_1 _18788_ (.A2(_04443_),
    .A1(net5246),
    .B1(_04444_),
    .X(_04445_));
 sg13g2_o21ai_1 _18789_ (.B1(_04445_),
    .Y(_01180_),
    .A1(net6151),
    .A2(_08192_));
 sg13g2_nand2_1 _18790_ (.Y(_04446_),
    .A(net6137),
    .B(_04300_));
 sg13g2_nor2_1 _18791_ (.A(_04052_),
    .B(net5095),
    .Y(_04447_));
 sg13g2_a21o_1 _18792_ (.A2(_04446_),
    .A1(net5245),
    .B1(_04447_),
    .X(_04448_));
 sg13g2_o21ai_1 _18793_ (.B1(_04448_),
    .Y(_01181_),
    .A1(net6149),
    .A2(_08191_));
 sg13g2_nand2_1 _18794_ (.Y(_04449_),
    .A(net6137),
    .B(_04303_));
 sg13g2_nor2_1 _18795_ (.A(_04076_),
    .B(net5095),
    .Y(_04450_));
 sg13g2_a21o_1 _18796_ (.A2(_04449_),
    .A1(net5245),
    .B1(_04450_),
    .X(_04451_));
 sg13g2_o21ai_1 _18797_ (.B1(_04451_),
    .Y(_01182_),
    .A1(net6149),
    .A2(_08190_));
 sg13g2_nand2_1 _18798_ (.Y(_04452_),
    .A(net6138),
    .B(_04306_));
 sg13g2_nor2_1 _18799_ (.A(_04100_),
    .B(net5095),
    .Y(_04453_));
 sg13g2_a21o_1 _18800_ (.A2(_04452_),
    .A1(net5245),
    .B1(_04453_),
    .X(_04454_));
 sg13g2_o21ai_1 _18801_ (.B1(_04454_),
    .Y(_01183_),
    .A1(net6149),
    .A2(_08189_));
 sg13g2_nand2_1 _18802_ (.Y(_04455_),
    .A(net6138),
    .B(_04309_));
 sg13g2_nor2_1 _18803_ (.A(_04124_),
    .B(net5095),
    .Y(_04456_));
 sg13g2_a21oi_1 _18804_ (.A1(net5246),
    .A2(_04455_),
    .Y(_04457_),
    .B1(_04456_));
 sg13g2_a21o_1 _18805_ (.A2(net2942),
    .A1(net6401),
    .B1(_04457_),
    .X(_01184_));
 sg13g2_nand2_1 _18806_ (.Y(_04458_),
    .A(net6138),
    .B(_04312_));
 sg13g2_nor2_1 _18807_ (.A(_04148_),
    .B(net5096),
    .Y(_04459_));
 sg13g2_a21oi_1 _18808_ (.A1(net5246),
    .A2(_04458_),
    .Y(_04460_),
    .B1(_04459_));
 sg13g2_a21o_1 _18809_ (.A2(net3061),
    .A1(net6402),
    .B1(_04460_),
    .X(_01185_));
 sg13g2_nand2_1 _18810_ (.Y(_04461_),
    .A(net6139),
    .B(_04315_));
 sg13g2_nor2_1 _18811_ (.A(_04172_),
    .B(net5096),
    .Y(_04462_));
 sg13g2_a21oi_1 _18812_ (.A1(net5246),
    .A2(_04461_),
    .Y(_04463_),
    .B1(_04462_));
 sg13g2_a21o_1 _18813_ (.A2(net3162),
    .A1(net6402),
    .B1(_04463_),
    .X(_01186_));
 sg13g2_nand2_1 _18814_ (.Y(_04464_),
    .A(net6139),
    .B(_04318_));
 sg13g2_nor2_1 _18815_ (.A(_04196_),
    .B(net5095),
    .Y(_04465_));
 sg13g2_a21o_1 _18816_ (.A2(_04464_),
    .A1(net5246),
    .B1(_04465_),
    .X(_04466_));
 sg13g2_o21ai_1 _18817_ (.B1(_04466_),
    .Y(_01187_),
    .A1(net6149),
    .A2(_08187_));
 sg13g2_a22oi_1 _18818_ (.Y(_04467_),
    .B1(_04320_),
    .B2(net6140),
    .A2(net3242),
    .A1(net6426));
 sg13g2_o21ai_1 _18819_ (.B1(net3243),
    .Y(_01188_),
    .A1(_04219_),
    .A2(net5247));
 sg13g2_mux2_1 _18820_ (.A0(net3196),
    .A1(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .S(net6422),
    .X(_01189_));
 sg13g2_mux2_1 _18821_ (.A0(net2528),
    .A1(net3248),
    .S(net6418),
    .X(_01190_));
 sg13g2_mux2_1 _18822_ (.A0(\soc_inst.cpu_core.ex_instr[9] ),
    .A1(net1593),
    .S(net6418),
    .X(_01191_));
 sg13g2_mux2_1 _18823_ (.A0(net2022),
    .A1(net2543),
    .S(net6422),
    .X(_01192_));
 sg13g2_a22oi_1 _18824_ (.Y(_04468_),
    .B1(net2451),
    .B2(net5309),
    .A2(\soc_inst.cpu_core.id_is_compressed ),
    .A1(net6416));
 sg13g2_inv_1 _18825_ (.Y(_01193_),
    .A(net2452));
 sg13g2_mux2_1 _18826_ (.A0(net2480),
    .A1(net2762),
    .S(net6371),
    .X(_01194_));
 sg13g2_mux2_1 _18827_ (.A0(net2833),
    .A1(net2888),
    .S(net6365),
    .X(_01195_));
 sg13g2_mux2_1 _18828_ (.A0(net3016),
    .A1(net3017),
    .S(net6365),
    .X(_01196_));
 sg13g2_mux2_1 _18829_ (.A0(net3051),
    .A1(\soc_inst.cpu_core.ex_instr[3] ),
    .S(net6371),
    .X(_01197_));
 sg13g2_nor2_1 _18830_ (.A(_00257_),
    .B(net6365),
    .Y(_04469_));
 sg13g2_a21oi_1 _18831_ (.A1(_07791_),
    .A2(net6364),
    .Y(_01198_),
    .B1(_04469_));
 sg13g2_mux2_1 _18832_ (.A0(net3182),
    .A1(net6213),
    .S(net6407),
    .X(_01199_));
 sg13g2_mux2_1 _18833_ (.A0(net2587),
    .A1(\soc_inst.cpu_core.ex_instr[6] ),
    .S(net6412),
    .X(_01200_));
 sg13g2_mux2_1 _18834_ (.A0(net2416),
    .A1(\soc_inst.cpu_core.ex_instr[7] ),
    .S(net6415),
    .X(_01201_));
 sg13g2_mux2_1 _18835_ (.A0(net2345),
    .A1(net2528),
    .S(net6377),
    .X(_01202_));
 sg13g2_mux2_1 _18836_ (.A0(net2153),
    .A1(\soc_inst.cpu_core.ex_instr[9] ),
    .S(net6377),
    .X(_01203_));
 sg13g2_mux2_1 _18837_ (.A0(net1652),
    .A1(net2022),
    .S(net6377),
    .X(_01204_));
 sg13g2_mux2_1 _18838_ (.A0(net1835),
    .A1(net2130),
    .S(net6415),
    .X(_01205_));
 sg13g2_mux2_1 _18839_ (.A0(\soc_inst.cpu_core.id_funct3[0] ),
    .A1(net2978),
    .S(net6368),
    .X(_01206_));
 sg13g2_mux2_1 _18840_ (.A0(\soc_inst.cpu_core.id_funct3[1] ),
    .A1(net3028),
    .S(net6405),
    .X(_01207_));
 sg13g2_nor2_1 _18841_ (.A(net6366),
    .B(net2234),
    .Y(_04470_));
 sg13g2_a21oi_1 _18842_ (.A1(_07869_),
    .A2(net6366),
    .Y(_01208_),
    .B1(_04470_));
 sg13g2_nor2_1 _18843_ (.A(net6395),
    .B(net360),
    .Y(_04471_));
 sg13g2_a21oi_1 _18844_ (.A1(net6389),
    .A2(_08173_),
    .Y(_01209_),
    .B1(_04471_));
 sg13g2_mux2_1 _18845_ (.A0(net1350),
    .A1(\soc_inst.cpu_core.ex_instr[16] ),
    .S(net6360),
    .X(_01210_));
 sg13g2_nor2_1 _18846_ (.A(net6355),
    .B(net1545),
    .Y(_04472_));
 sg13g2_a21oi_1 _18847_ (.A1(net6354),
    .A2(_08175_),
    .Y(_01211_),
    .B1(_04472_));
 sg13g2_mux2_1 _18848_ (.A0(net1363),
    .A1(\soc_inst.cpu_core.ex_instr[18] ),
    .S(net6367),
    .X(_01212_));
 sg13g2_mux2_1 _18849_ (.A0(net1864),
    .A1(\soc_inst.cpu_core.ex_instr[19] ),
    .S(net6371),
    .X(_01213_));
 sg13g2_nor2_1 _18850_ (.A(net6345),
    .B(net630),
    .Y(_04473_));
 sg13g2_a21oi_1 _18851_ (.A1(net6345),
    .A2(_08176_),
    .Y(_01214_),
    .B1(_04473_));
 sg13g2_mux2_1 _18852_ (.A0(net2501),
    .A1(net2487),
    .S(net6390),
    .X(_01215_));
 sg13g2_a21oi_1 _18853_ (.A1(net6348),
    .A2(_08177_),
    .Y(_01216_),
    .B1(_11413_));
 sg13g2_mux2_1 _18854_ (.A0(net2885),
    .A1(net2715),
    .S(net6388),
    .X(_01217_));
 sg13g2_mux2_1 _18855_ (.A0(net2286),
    .A1(\soc_inst.cpu_core.ex_instr[24] ),
    .S(net6351),
    .X(_01218_));
 sg13g2_nor2_1 _18856_ (.A(net6349),
    .B(net1121),
    .Y(_04474_));
 sg13g2_a21oi_1 _18857_ (.A1(net6349),
    .A2(_08179_),
    .Y(_01219_),
    .B1(_04474_));
 sg13g2_mux2_1 _18858_ (.A0(\soc_inst.cpu_core.id_imm12[6] ),
    .A1(net2338),
    .S(net6348),
    .X(_01220_));
 sg13g2_mux2_1 _18859_ (.A0(net2613),
    .A1(net2393),
    .S(net6349),
    .X(_01221_));
 sg13g2_mux2_1 _18860_ (.A0(\soc_inst.cpu_core.id_imm12[8] ),
    .A1(net2841),
    .S(net6355),
    .X(_01222_));
 sg13g2_mux2_1 _18861_ (.A0(\soc_inst.cpu_core.id_imm12[9] ),
    .A1(net2371),
    .S(net6354),
    .X(_01223_));
 sg13g2_mux2_1 _18862_ (.A0(net2566),
    .A1(net2098),
    .S(net6349),
    .X(_01224_));
 sg13g2_mux2_1 _18863_ (.A0(net2726),
    .A1(net2785),
    .S(net6354),
    .X(_01225_));
 sg13g2_nor2_2 _18864_ (.A(net6478),
    .B(net6344),
    .Y(_04475_));
 sg13g2_a22oi_1 _18865_ (.Y(_01226_),
    .B1(net6074),
    .B2(_08082_),
    .A2(_08136_),
    .A1(net6365));
 sg13g2_a22oi_1 _18866_ (.Y(_01227_),
    .B1(net6075),
    .B2(_08083_),
    .A2(_08137_),
    .A1(net6406));
 sg13g2_a22oi_1 _18867_ (.Y(_01228_),
    .B1(net6075),
    .B2(_08084_),
    .A2(_08138_),
    .A1(net6370));
 sg13g2_a22oi_1 _18868_ (.Y(_01229_),
    .B1(net6075),
    .B2(_08085_),
    .A2(_08139_),
    .A1(net6369));
 sg13g2_a22oi_1 _18869_ (.Y(_01230_),
    .B1(net6075),
    .B2(_08087_),
    .A2(_08140_),
    .A1(net6406));
 sg13g2_a22oi_1 _18870_ (.Y(_01231_),
    .B1(net6074),
    .B2(_08089_),
    .A2(_08141_),
    .A1(net6364));
 sg13g2_a22oi_1 _18871_ (.Y(_01232_),
    .B1(net6074),
    .B2(_08091_),
    .A2(_08142_),
    .A1(net6364));
 sg13g2_a22oi_1 _18872_ (.Y(_01233_),
    .B1(net6074),
    .B2(_08093_),
    .A2(_08143_),
    .A1(net6371));
 sg13g2_a22oi_1 _18873_ (.Y(_01234_),
    .B1(net6074),
    .B2(_08095_),
    .A2(_08144_),
    .A1(net6367));
 sg13g2_a22oi_1 _18874_ (.Y(_01235_),
    .B1(net6074),
    .B2(_08097_),
    .A2(_08145_),
    .A1(net6366));
 sg13g2_a22oi_1 _18875_ (.Y(_01236_),
    .B1(net6074),
    .B2(_08099_),
    .A2(_08146_),
    .A1(net6357));
 sg13g2_a22oi_1 _18876_ (.Y(_01237_),
    .B1(net6075),
    .B2(_08101_),
    .A2(_08147_),
    .A1(net6367));
 sg13g2_a22oi_1 _18877_ (.Y(_01238_),
    .B1(net6074),
    .B2(_08103_),
    .A2(_08148_),
    .A1(net6354));
 sg13g2_a22oi_1 _18878_ (.Y(_01239_),
    .B1(net6073),
    .B2(_08105_),
    .A2(_08149_),
    .A1(net6349));
 sg13g2_a22oi_1 _18879_ (.Y(_01240_),
    .B1(net6072),
    .B2(_08106_),
    .A2(_08150_),
    .A1(net6344));
 sg13g2_a22oi_1 _18880_ (.Y(_01241_),
    .B1(net6072),
    .B2(_08107_),
    .A2(_08151_),
    .A1(net6339));
 sg13g2_a22oi_1 _18881_ (.Y(_01242_),
    .B1(net6072),
    .B2(_08108_),
    .A2(_08152_),
    .A1(net6340));
 sg13g2_a22oi_1 _18882_ (.Y(_01243_),
    .B1(net6073),
    .B2(_08109_),
    .A2(_08153_),
    .A1(net6344));
 sg13g2_a22oi_1 _18883_ (.Y(_01244_),
    .B1(net6072),
    .B2(_08110_),
    .A2(_08154_),
    .A1(net6340));
 sg13g2_a22oi_1 _18884_ (.Y(_01245_),
    .B1(net6072),
    .B2(_08111_),
    .A2(_08155_),
    .A1(net6340));
 sg13g2_a22oi_1 _18885_ (.Y(_01246_),
    .B1(net6072),
    .B2(_08112_),
    .A2(_08156_),
    .A1(net6339));
 sg13g2_a22oi_1 _18886_ (.Y(_01247_),
    .B1(net6072),
    .B2(_08113_),
    .A2(_08157_),
    .A1(net6339));
 sg13g2_a22oi_1 _18887_ (.Y(_01248_),
    .B1(net6073),
    .B2(_08115_),
    .A2(_08158_),
    .A1(net6344));
 sg13g2_a22oi_1 _18888_ (.Y(_01249_),
    .B1(net6072),
    .B2(_08116_),
    .A2(_08159_),
    .A1(net6339));
 sg13g2_nand2_1 _18889_ (.Y(_04476_),
    .A(net6373),
    .B(net644));
 sg13g2_o21ai_1 _18890_ (.B1(_04476_),
    .Y(_01250_),
    .A1(net6373),
    .A2(_08029_));
 sg13g2_nand2_1 _18891_ (.Y(_04477_),
    .A(net6371),
    .B(net394));
 sg13g2_o21ai_1 _18892_ (.B1(_04477_),
    .Y(_01251_),
    .A1(net6371),
    .A2(_08030_));
 sg13g2_mux2_1 _18893_ (.A0(\soc_inst.cpu_core.id_rs1_data[2] ),
    .A1(net2043),
    .S(net6363),
    .X(_01252_));
 sg13g2_nand2_1 _18894_ (.Y(_04478_),
    .A(net6374),
    .B(net316));
 sg13g2_o21ai_1 _18895_ (.B1(_04478_),
    .Y(_01253_),
    .A1(net6374),
    .A2(_08031_));
 sg13g2_nand2_1 _18896_ (.Y(_04479_),
    .A(net6364),
    .B(net257));
 sg13g2_o21ai_1 _18897_ (.B1(_04479_),
    .Y(_01254_),
    .A1(net6359),
    .A2(_08039_));
 sg13g2_nand2_1 _18898_ (.Y(_04480_),
    .A(net6378),
    .B(net519));
 sg13g2_o21ai_1 _18899_ (.B1(_04480_),
    .Y(_01255_),
    .A1(net6378),
    .A2(_08037_));
 sg13g2_nand2_1 _18900_ (.Y(_04481_),
    .A(net6330),
    .B(net455));
 sg13g2_o21ai_1 _18901_ (.B1(_04481_),
    .Y(_01256_),
    .A1(net6330),
    .A2(_08035_));
 sg13g2_nand2_1 _18902_ (.Y(_04482_),
    .A(net6361),
    .B(net1197));
 sg13g2_o21ai_1 _18903_ (.B1(_04482_),
    .Y(_01257_),
    .A1(net6362),
    .A2(_08033_));
 sg13g2_nand2_1 _18904_ (.Y(_04483_),
    .A(net6334),
    .B(net260));
 sg13g2_o21ai_1 _18905_ (.B1(_04483_),
    .Y(_01258_),
    .A1(net6334),
    .A2(_08054_));
 sg13g2_nand2_1 _18906_ (.Y(_04484_),
    .A(net6362),
    .B(net206));
 sg13g2_o21ai_1 _18907_ (.B1(_04484_),
    .Y(_01259_),
    .A1(net6361),
    .A2(_08052_));
 sg13g2_nand2_1 _18908_ (.Y(_04485_),
    .A(net6334),
    .B(net243));
 sg13g2_o21ai_1 _18909_ (.B1(_04485_),
    .Y(_01260_),
    .A1(net6333),
    .A2(_08050_));
 sg13g2_nand2_1 _18910_ (.Y(_04486_),
    .A(net6334),
    .B(net326));
 sg13g2_o21ai_1 _18911_ (.B1(_04486_),
    .Y(_01261_),
    .A1(net6334),
    .A2(_08049_));
 sg13g2_nand2_1 _18912_ (.Y(_04487_),
    .A(net6323),
    .B(net231));
 sg13g2_o21ai_1 _18913_ (.B1(_04487_),
    .Y(_01262_),
    .A1(net6323),
    .A2(_08047_));
 sg13g2_nand2_1 _18914_ (.Y(_04488_),
    .A(net6324),
    .B(net288));
 sg13g2_o21ai_1 _18915_ (.B1(_04488_),
    .Y(_01263_),
    .A1(net6324),
    .A2(_08045_));
 sg13g2_nand2_1 _18916_ (.Y(_04489_),
    .A(net6336),
    .B(net367));
 sg13g2_o21ai_1 _18917_ (.B1(_04489_),
    .Y(_01264_),
    .A1(net6336),
    .A2(_08043_));
 sg13g2_nand2_1 _18918_ (.Y(_04490_),
    .A(net6335),
    .B(net729));
 sg13g2_o21ai_1 _18919_ (.B1(_04490_),
    .Y(_01265_),
    .A1(net6335),
    .A2(_08041_));
 sg13g2_nand2_1 _18920_ (.Y(_04491_),
    .A(net6343),
    .B(net275));
 sg13g2_o21ai_1 _18921_ (.B1(_04491_),
    .Y(_01266_),
    .A1(net6343),
    .A2(_08080_));
 sg13g2_nand2_1 _18922_ (.Y(_04492_),
    .A(net6338),
    .B(net217));
 sg13g2_o21ai_1 _18923_ (.B1(_04492_),
    .Y(_01267_),
    .A1(net6338),
    .A2(_08078_));
 sg13g2_nand2_1 _18924_ (.Y(_04493_),
    .A(net6343),
    .B(net1033));
 sg13g2_o21ai_1 _18925_ (.B1(_04493_),
    .Y(_01268_),
    .A1(net6341),
    .A2(_08076_));
 sg13g2_nand2_1 _18926_ (.Y(_04494_),
    .A(net6337),
    .B(net524));
 sg13g2_o21ai_1 _18927_ (.B1(_04494_),
    .Y(_01269_),
    .A1(net6337),
    .A2(_08074_));
 sg13g2_nand2_1 _18928_ (.Y(_04495_),
    .A(net6341),
    .B(net891));
 sg13g2_o21ai_1 _18929_ (.B1(_04495_),
    .Y(_01270_),
    .A1(net6341),
    .A2(_08073_));
 sg13g2_mux2_1 _18930_ (.A0(\soc_inst.cpu_core.id_rs1_data[21] ),
    .A1(net2223),
    .S(net6341),
    .X(_01271_));
 sg13g2_nand2_1 _18931_ (.Y(_04496_),
    .A(net6342),
    .B(net885));
 sg13g2_o21ai_1 _18932_ (.B1(_04496_),
    .Y(_01272_),
    .A1(net6342),
    .A2(_08070_));
 sg13g2_nand2_1 _18933_ (.Y(_04497_),
    .A(net6341),
    .B(net1368));
 sg13g2_o21ai_1 _18934_ (.B1(_04497_),
    .Y(_01273_),
    .A1(net6341),
    .A2(_08068_));
 sg13g2_nand2_1 _18935_ (.Y(_04498_),
    .A(net6381),
    .B(net1279));
 sg13g2_o21ai_1 _18936_ (.B1(_04498_),
    .Y(_01274_),
    .A1(net6381),
    .A2(_08066_));
 sg13g2_nand2_1 _18937_ (.Y(_04499_),
    .A(net6340),
    .B(net732));
 sg13g2_o21ai_1 _18938_ (.B1(_04499_),
    .Y(_01275_),
    .A1(net6340),
    .A2(_08065_));
 sg13g2_nand2_1 _18939_ (.Y(_04500_),
    .A(net6397),
    .B(net214));
 sg13g2_o21ai_1 _18940_ (.B1(_04500_),
    .Y(_01276_),
    .A1(net6386),
    .A2(_08063_));
 sg13g2_nand2_1 _18941_ (.Y(_04501_),
    .A(net6339),
    .B(net320));
 sg13g2_o21ai_1 _18942_ (.B1(_04501_),
    .Y(_01277_),
    .A1(net6339),
    .A2(_08061_));
 sg13g2_nand2_1 _18943_ (.Y(_04502_),
    .A(net6341),
    .B(net328));
 sg13g2_o21ai_1 _18944_ (.B1(_04502_),
    .Y(_01278_),
    .A1(net6343),
    .A2(_08060_));
 sg13g2_nand2_1 _18945_ (.Y(_04503_),
    .A(net6342),
    .B(net2822));
 sg13g2_o21ai_1 _18946_ (.B1(_04503_),
    .Y(_01279_),
    .A1(net6344),
    .A2(_08059_));
 sg13g2_nand2_1 _18947_ (.Y(_04504_),
    .A(net6340),
    .B(net374));
 sg13g2_o21ai_1 _18948_ (.B1(_04504_),
    .Y(_01280_),
    .A1(net6339),
    .A2(_08058_));
 sg13g2_nand2_1 _18949_ (.Y(_04505_),
    .A(net6353),
    .B(net381));
 sg13g2_o21ai_1 _18950_ (.B1(_04505_),
    .Y(_01281_),
    .A1(net6352),
    .A2(_08057_));
 sg13g2_nor2_2 _18951_ (.A(net2814),
    .B(net6359),
    .Y(_04506_));
 sg13g2_a21oi_1 _18952_ (.A1(net6327),
    .A2(_07886_),
    .Y(_01282_),
    .B1(_04506_));
 sg13g2_nor2_2 _18953_ (.A(net3205),
    .B(net6359),
    .Y(_04507_));
 sg13g2_a21oi_1 _18954_ (.A1(net6327),
    .A2(_07885_),
    .Y(_01283_),
    .B1(_04507_));
 sg13g2_nor2_1 _18955_ (.A(net6326),
    .B(net3266),
    .Y(_04508_));
 sg13g2_a21oi_1 _18956_ (.A1(net6330),
    .A2(_07887_),
    .Y(_01284_),
    .B1(_04508_));
 sg13g2_nor2_1 _18957_ (.A(net6326),
    .B(net3279),
    .Y(_04509_));
 sg13g2_a21oi_1 _18958_ (.A1(net6326),
    .A2(_07888_),
    .Y(_01285_),
    .B1(_04509_));
 sg13g2_nor2_2 _18959_ (.A(net6359),
    .B(\soc_inst.cpu_core.ex_alu_result[4] ),
    .Y(_04510_));
 sg13g2_a21oi_1 _18960_ (.A1(net6327),
    .A2(_07889_),
    .Y(_01286_),
    .B1(_04510_));
 sg13g2_nor2_1 _18961_ (.A(net6327),
    .B(net2938),
    .Y(_04511_));
 sg13g2_a21oi_1 _18962_ (.A1(net6327),
    .A2(_07890_),
    .Y(_01287_),
    .B1(_04511_));
 sg13g2_nor2_1 _18963_ (.A(net6327),
    .B(net2900),
    .Y(_04512_));
 sg13g2_a21oi_1 _18964_ (.A1(net6326),
    .A2(_07892_),
    .Y(_01288_),
    .B1(_04512_));
 sg13g2_nor2_2 _18965_ (.A(net6411),
    .B(net2656),
    .Y(_04513_));
 sg13g2_a21oi_1 _18966_ (.A1(net6327),
    .A2(_07891_),
    .Y(_01289_),
    .B1(_04513_));
 sg13g2_nand2_1 _18967_ (.Y(_04514_),
    .A(net1051),
    .B(net6326));
 sg13g2_o21ai_1 _18968_ (.B1(_04514_),
    .Y(_01290_),
    .A1(net6326),
    .A2(_08166_));
 sg13g2_nand2_1 _18969_ (.Y(_04515_),
    .A(net1927),
    .B(net6329));
 sg13g2_o21ai_1 _18970_ (.B1(_04515_),
    .Y(_01291_),
    .A1(net6329),
    .A2(_08167_));
 sg13g2_nand2_1 _18971_ (.Y(_04516_),
    .A(net1110),
    .B(net6324));
 sg13g2_o21ai_1 _18972_ (.B1(_04516_),
    .Y(_01292_),
    .A1(net6329),
    .A2(_08168_));
 sg13g2_nor2_1 _18973_ (.A(net6326),
    .B(\soc_inst.cpu_core.ex_alu_result[11] ),
    .Y(_04517_));
 sg13g2_a21oi_1 _18974_ (.A1(_07812_),
    .A2(net6324),
    .Y(_01293_),
    .B1(_04517_));
 sg13g2_nand2_1 _18975_ (.Y(_04518_),
    .A(\soc_inst.core_mem_addr[12] ),
    .B(net6392));
 sg13g2_o21ai_1 _18976_ (.B1(_04518_),
    .Y(_01294_),
    .A1(net6392),
    .A2(_08170_));
 sg13g2_nor2_1 _18977_ (.A(net6323),
    .B(net3287),
    .Y(_04519_));
 sg13g2_a21oi_1 _18978_ (.A1(_07813_),
    .A2(net6320),
    .Y(_01295_),
    .B1(_04519_));
 sg13g2_nor2_1 _18979_ (.A(net6323),
    .B(\soc_inst.cpu_core.ex_alu_result[14] ),
    .Y(_04520_));
 sg13g2_a21oi_1 _18980_ (.A1(_07815_),
    .A2(net6320),
    .Y(_01296_),
    .B1(_04520_));
 sg13g2_nor2_1 _18981_ (.A(net6324),
    .B(\soc_inst.cpu_core.ex_alu_result[15] ),
    .Y(_04521_));
 sg13g2_a21oi_1 _18982_ (.A1(_07814_),
    .A2(net6324),
    .Y(_01297_),
    .B1(_04521_));
 sg13g2_mux2_1 _18983_ (.A0(net2299),
    .A1(net3105),
    .S(net6348),
    .X(_01298_));
 sg13g2_mux2_1 _18984_ (.A0(\soc_inst.cpu_core.ex_alu_result[17] ),
    .A1(net2856),
    .S(net6323),
    .X(_01299_));
 sg13g2_mux2_1 _18985_ (.A0(\soc_inst.cpu_core.ex_alu_result[18] ),
    .A1(net2836),
    .S(net6320),
    .X(_01300_));
 sg13g2_mux2_1 _18986_ (.A0(\soc_inst.cpu_core.ex_alu_result[19] ),
    .A1(net2687),
    .S(net6317),
    .X(_01301_));
 sg13g2_mux2_1 _18987_ (.A0(\soc_inst.cpu_core.ex_alu_result[20] ),
    .A1(net2805),
    .S(net6323),
    .X(_01302_));
 sg13g2_mux2_1 _18988_ (.A0(net2879),
    .A1(net2889),
    .S(net6323),
    .X(_01303_));
 sg13g2_mux2_1 _18989_ (.A0(\soc_inst.cpu_core.ex_alu_result[22] ),
    .A1(net2694),
    .S(net6320),
    .X(_01304_));
 sg13g2_mux2_1 _18990_ (.A0(\soc_inst.cpu_core.ex_alu_result[23] ),
    .A1(net2902),
    .S(net6323),
    .X(_01305_));
 sg13g2_mux2_1 _18991_ (.A0(\soc_inst.cpu_core.ex_alu_result[24] ),
    .A1(net2731),
    .S(net6331),
    .X(_01306_));
 sg13g2_mux2_1 _18992_ (.A0(\soc_inst.cpu_core.ex_alu_result[25] ),
    .A1(net2847),
    .S(net6331),
    .X(_01307_));
 sg13g2_mux2_1 _18993_ (.A0(\soc_inst.cpu_core.ex_alu_result[26] ),
    .A1(net2733),
    .S(net6331),
    .X(_01308_));
 sg13g2_mux2_1 _18994_ (.A0(\soc_inst.cpu_core.ex_alu_result[27] ),
    .A1(net2757),
    .S(net6331),
    .X(_01309_));
 sg13g2_mux2_1 _18995_ (.A0(\soc_inst.cpu_core.ex_alu_result[28] ),
    .A1(net2630),
    .S(net6325),
    .X(_01310_));
 sg13g2_mux2_1 _18996_ (.A0(\soc_inst.cpu_core.ex_alu_result[29] ),
    .A1(net2545),
    .S(net6329),
    .X(_01311_));
 sg13g2_mux2_1 _18997_ (.A0(\soc_inst.cpu_core.ex_alu_result[30] ),
    .A1(net2701),
    .S(net6326),
    .X(_01312_));
 sg13g2_nand2_1 _18998_ (.Y(_04522_),
    .A(net403),
    .B(net6329));
 sg13g2_o21ai_1 _18999_ (.B1(_04522_),
    .Y(_01313_),
    .A1(net6329),
    .A2(_08184_));
 sg13g2_mux2_1 _19000_ (.A0(net1491),
    .A1(net377),
    .S(net6312),
    .X(_01314_));
 sg13g2_mux2_1 _19001_ (.A0(net1466),
    .A1(net299),
    .S(net6310),
    .X(_01315_));
 sg13g2_mux2_1 _19002_ (.A0(net1291),
    .A1(net791),
    .S(net6330),
    .X(_01316_));
 sg13g2_nand2_1 _19003_ (.Y(_04523_),
    .A(net6312),
    .B(net398));
 sg13g2_o21ai_1 _19004_ (.B1(_04523_),
    .Y(_01317_),
    .A1(net6312),
    .A2(_08032_));
 sg13g2_nand2_1 _19005_ (.Y(_04524_),
    .A(net6310),
    .B(net251));
 sg13g2_o21ai_1 _19006_ (.B1(_04524_),
    .Y(_01318_),
    .A1(net6310),
    .A2(_08040_));
 sg13g2_nand2_1 _19007_ (.Y(_04525_),
    .A(net6311),
    .B(net638));
 sg13g2_o21ai_1 _19008_ (.B1(_04525_),
    .Y(_01319_),
    .A1(net6311),
    .A2(_08038_));
 sg13g2_nand2_1 _19009_ (.Y(_04526_),
    .A(net6310),
    .B(net297));
 sg13g2_o21ai_1 _19010_ (.B1(_04526_),
    .Y(_01320_),
    .A1(net6310),
    .A2(_08036_));
 sg13g2_nand2_1 _19011_ (.Y(_04527_),
    .A(net6313),
    .B(net856));
 sg13g2_o21ai_1 _19012_ (.B1(net857),
    .Y(_01321_),
    .A1(net6313),
    .A2(_08034_));
 sg13g2_nand2_1 _19013_ (.Y(_04528_),
    .A(net6321),
    .B(net255));
 sg13g2_o21ai_1 _19014_ (.B1(_04528_),
    .Y(_01322_),
    .A1(net6321),
    .A2(_08055_));
 sg13g2_nand2_1 _19015_ (.Y(_04529_),
    .A(net6308),
    .B(net926));
 sg13g2_o21ai_1 _19016_ (.B1(_04529_),
    .Y(_01323_),
    .A1(net6308),
    .A2(_08053_));
 sg13g2_nand2_1 _19017_ (.Y(_04530_),
    .A(net6321),
    .B(net293));
 sg13g2_o21ai_1 _19018_ (.B1(_04530_),
    .Y(_01324_),
    .A1(net6320),
    .A2(_08051_));
 sg13g2_mux2_1 _19019_ (.A0(net1726),
    .A1(net1396),
    .S(net6307),
    .X(_01325_));
 sg13g2_nand2_1 _19020_ (.Y(_04531_),
    .A(net6320),
    .B(net1799));
 sg13g2_o21ai_1 _19021_ (.B1(_04531_),
    .Y(_01326_),
    .A1(net6320),
    .A2(_08048_));
 sg13g2_nand2_1 _19022_ (.Y(_04532_),
    .A(net6309),
    .B(net238));
 sg13g2_o21ai_1 _19023_ (.B1(net239),
    .Y(_01327_),
    .A1(net6309),
    .A2(_08046_));
 sg13g2_nand2_1 _19024_ (.Y(_04533_),
    .A(net6309),
    .B(net335));
 sg13g2_o21ai_1 _19025_ (.B1(net336),
    .Y(_01328_),
    .A1(net6309),
    .A2(_08044_));
 sg13g2_nand2_1 _19026_ (.Y(_04534_),
    .A(net6325),
    .B(net1548));
 sg13g2_o21ai_1 _19027_ (.B1(_04534_),
    .Y(_01329_),
    .A1(net6322),
    .A2(_08042_));
 sg13g2_nand2_1 _19028_ (.Y(_04535_),
    .A(net6314),
    .B(net324));
 sg13g2_o21ai_1 _19029_ (.B1(_04535_),
    .Y(_01330_),
    .A1(net6314),
    .A2(_08081_));
 sg13g2_nand2_1 _19030_ (.Y(_04536_),
    .A(net6315),
    .B(net566));
 sg13g2_o21ai_1 _19031_ (.B1(_04536_),
    .Y(_01331_),
    .A1(net6315),
    .A2(_08079_));
 sg13g2_nand2_1 _19032_ (.Y(_04537_),
    .A(net6322),
    .B(net510));
 sg13g2_o21ai_1 _19033_ (.B1(_04537_),
    .Y(_01332_),
    .A1(net6322),
    .A2(_08077_));
 sg13g2_nand2_1 _19034_ (.Y(_04538_),
    .A(net6315),
    .B(net687));
 sg13g2_o21ai_1 _19035_ (.B1(_04538_),
    .Y(_01333_),
    .A1(net6315),
    .A2(_08075_));
 sg13g2_mux2_1 _19036_ (.A0(\soc_inst.cpu_core.id_rs2_data[20] ),
    .A1(net1976),
    .S(net6315),
    .X(_01334_));
 sg13g2_nand2_1 _19037_ (.Y(_04539_),
    .A(net6322),
    .B(net522));
 sg13g2_o21ai_1 _19038_ (.B1(_04539_),
    .Y(_01335_),
    .A1(net6322),
    .A2(_08072_));
 sg13g2_nand2_1 _19039_ (.Y(_04540_),
    .A(net6316),
    .B(net586));
 sg13g2_o21ai_1 _19040_ (.B1(_04540_),
    .Y(_01336_),
    .A1(net6316),
    .A2(_08071_));
 sg13g2_nand2_1 _19041_ (.Y(_04541_),
    .A(net6322),
    .B(net273));
 sg13g2_o21ai_1 _19042_ (.B1(_04541_),
    .Y(_01337_),
    .A1(net6322),
    .A2(_08069_));
 sg13g2_nand2_1 _19043_ (.Y(_04542_),
    .A(net6319),
    .B(net347));
 sg13g2_o21ai_1 _19044_ (.B1(_04542_),
    .Y(_01338_),
    .A1(net6319),
    .A2(_08067_));
 sg13g2_mux2_1 _19045_ (.A0(\soc_inst.cpu_core.id_rs2_data[25] ),
    .A1(net2573),
    .S(net6314),
    .X(_01339_));
 sg13g2_nand2_1 _19046_ (.Y(_04543_),
    .A(net6318),
    .B(net208));
 sg13g2_o21ai_1 _19047_ (.B1(_04543_),
    .Y(_01340_),
    .A1(net6317),
    .A2(_08064_));
 sg13g2_nand2_1 _19048_ (.Y(_04544_),
    .A(net6318),
    .B(net472));
 sg13g2_o21ai_1 _19049_ (.B1(_04544_),
    .Y(_01341_),
    .A1(net6317),
    .A2(_08062_));
 sg13g2_mux2_1 _19050_ (.A0(net1318),
    .A1(net1089),
    .S(net6307),
    .X(_01342_));
 sg13g2_mux2_1 _19051_ (.A0(net1343),
    .A1(net852),
    .S(net6307),
    .X(_01343_));
 sg13g2_mux2_1 _19052_ (.A0(\soc_inst.cpu_core.id_rs2_data[30] ),
    .A1(net1795),
    .S(net6318),
    .X(_01344_));
 sg13g2_nand2_1 _19053_ (.Y(_04545_),
    .A(net6317),
    .B(net426));
 sg13g2_o21ai_1 _19054_ (.B1(_04545_),
    .Y(_01345_),
    .A1(net6317),
    .A2(_08056_));
 sg13g2_nand2_1 _19055_ (.Y(_04546_),
    .A(net2814),
    .B(net6410));
 sg13g2_nor2_2 _19056_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B(net6288),
    .Y(_04547_));
 sg13g2_nor3_1 _19057_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B(net6288),
    .C(\soc_inst.cpu_core.alu.op[2] ),
    .Y(_04548_));
 sg13g2_nor2b_2 _19058_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B_N(net6287),
    .Y(_04549_));
 sg13g2_and2_1 _19059_ (.A(\soc_inst.cpu_core.alu.op[2] ),
    .B(_04549_),
    .X(_04550_));
 sg13g2_nand2_2 _19060_ (.Y(_04551_),
    .A(\soc_inst.cpu_core.alu.op[2] ),
    .B(_04549_));
 sg13g2_and2_1 _19061_ (.A(net6285),
    .B(_04548_),
    .X(_04552_));
 sg13g2_nand2_1 _19062_ (.Y(_04553_),
    .A(net6285),
    .B(_04548_));
 sg13g2_nand3_1 _19063_ (.B(_04551_),
    .C(net5771),
    .A(net3400),
    .Y(_04554_));
 sg13g2_and2_1 _19064_ (.A(net6156),
    .B(_04554_),
    .X(_04555_));
 sg13g2_nand2_2 _19065_ (.Y(_04556_),
    .A(net6156),
    .B(_04554_));
 sg13g2_nand2b_1 _19066_ (.Y(_04557_),
    .B(net6261),
    .A_N(\soc_inst.cpu_core.alu.b[31] ));
 sg13g2_xor2_1 _19067_ (.B(net6261),
    .A(\soc_inst.cpu_core.alu.b[31] ),
    .X(_04558_));
 sg13g2_xnor2_1 _19068_ (.Y(_04559_),
    .A(\soc_inst.cpu_core.alu.b[29] ),
    .B(net6263));
 sg13g2_nor2_2 _19069_ (.A(\soc_inst.cpu_core.alu.b[15] ),
    .B(\soc_inst.cpu_core.alu.a[15] ),
    .Y(_04560_));
 sg13g2_nand2_1 _19070_ (.Y(_04561_),
    .A(\soc_inst.cpu_core.alu.b[15] ),
    .B(\soc_inst.cpu_core.alu.a[15] ));
 sg13g2_nor2b_2 _19071_ (.A(_04560_),
    .B_N(_04561_),
    .Y(_04562_));
 sg13g2_and2_1 _19072_ (.A(\soc_inst.cpu_core.alu.b[14] ),
    .B(net6283),
    .X(_04563_));
 sg13g2_nand2_1 _19073_ (.Y(_04564_),
    .A(\soc_inst.cpu_core.alu.b[14] ),
    .B(net6283));
 sg13g2_nor2_1 _19074_ (.A(\soc_inst.cpu_core.alu.b[14] ),
    .B(net6283),
    .Y(_04565_));
 sg13g2_nor2_2 _19075_ (.A(_04563_),
    .B(_04565_),
    .Y(_04566_));
 sg13g2_nor2_1 _19076_ (.A(_04562_),
    .B(_04566_),
    .Y(_04567_));
 sg13g2_nand2b_1 _19077_ (.Y(_04568_),
    .B(net6283),
    .A_N(\soc_inst.cpu_core.alu.b[14] ));
 sg13g2_nor2_1 _19078_ (.A(\soc_inst.cpu_core.alu.b[13] ),
    .B(\soc_inst.cpu_core.alu.a[13] ),
    .Y(_04569_));
 sg13g2_nand2_2 _19079_ (.Y(_04570_),
    .A(\soc_inst.cpu_core.alu.b[13] ),
    .B(\soc_inst.cpu_core.alu.a[13] ));
 sg13g2_nor2b_1 _19080_ (.A(_04569_),
    .B_N(_04570_),
    .Y(_04571_));
 sg13g2_nand2b_2 _19081_ (.Y(_04572_),
    .B(_04570_),
    .A_N(_04569_));
 sg13g2_nand2_1 _19082_ (.Y(_04573_),
    .A(_08202_),
    .B(\soc_inst.cpu_core.alu.a[11] ));
 sg13g2_or2_1 _19083_ (.X(_04574_),
    .B(\soc_inst.cpu_core.alu.a[11] ),
    .A(\soc_inst.cpu_core.alu.b[11] ));
 sg13g2_xor2_1 _19084_ (.B(\soc_inst.cpu_core.alu.a[11] ),
    .A(\soc_inst.cpu_core.alu.b[11] ),
    .X(_04575_));
 sg13g2_nand2b_1 _19085_ (.Y(_04576_),
    .B(\soc_inst.cpu_core.alu.a[10] ),
    .A_N(net2998));
 sg13g2_o21ai_1 _19086_ (.B1(_04573_),
    .Y(_04577_),
    .A1(_04575_),
    .A2(_04576_));
 sg13g2_nor2_1 _19087_ (.A(\soc_inst.cpu_core.alu.b[10] ),
    .B(\soc_inst.cpu_core.alu.a[10] ),
    .Y(_04578_));
 sg13g2_nand2_2 _19088_ (.Y(_04579_),
    .A(\soc_inst.cpu_core.alu.b[10] ),
    .B(\soc_inst.cpu_core.alu.a[10] ));
 sg13g2_nor2b_2 _19089_ (.A(_04578_),
    .B_N(_04579_),
    .Y(_04580_));
 sg13g2_or2_1 _19090_ (.X(_04581_),
    .B(_04580_),
    .A(_04575_));
 sg13g2_nor2_1 _19091_ (.A(\soc_inst.cpu_core.alu.b[9] ),
    .B(\soc_inst.cpu_core.alu.a[9] ),
    .Y(_04582_));
 sg13g2_nand2_2 _19092_ (.Y(_04583_),
    .A(\soc_inst.cpu_core.alu.b[9] ),
    .B(\soc_inst.cpu_core.alu.a[9] ));
 sg13g2_nor2b_2 _19093_ (.A(_04582_),
    .B_N(_04583_),
    .Y(_04584_));
 sg13g2_nand2b_2 _19094_ (.Y(_04585_),
    .B(_04583_),
    .A_N(_04582_));
 sg13g2_nand2b_1 _19095_ (.Y(_04586_),
    .B(net6284),
    .A_N(\soc_inst.cpu_core.alu.b[8] ));
 sg13g2_nand2b_1 _19096_ (.Y(_04587_),
    .B(_04585_),
    .A_N(_04586_));
 sg13g2_o21ai_1 _19097_ (.B1(_04587_),
    .Y(_04588_),
    .A1(\soc_inst.cpu_core.alu.b[9] ),
    .A2(_08204_));
 sg13g2_nor2b_1 _19098_ (.A(\soc_inst.cpu_core.alu.b[7] ),
    .B_N(\soc_inst.cpu_core.alu.a[7] ),
    .Y(_04589_));
 sg13g2_and2_1 _19099_ (.A(\soc_inst.cpu_core.alu.b[7] ),
    .B(\soc_inst.cpu_core.alu.a[7] ),
    .X(_04590_));
 sg13g2_nand2_1 _19100_ (.Y(_04591_),
    .A(\soc_inst.cpu_core.alu.b[7] ),
    .B(\soc_inst.cpu_core.alu.a[7] ));
 sg13g2_or2_1 _19101_ (.X(_04592_),
    .B(\soc_inst.cpu_core.alu.a[7] ),
    .A(\soc_inst.cpu_core.alu.b[7] ));
 sg13g2_nand2_2 _19102_ (.Y(_04593_),
    .A(_04591_),
    .B(_04592_));
 sg13g2_nand2b_1 _19103_ (.Y(_04594_),
    .B(\soc_inst.cpu_core.alu.a[6] ),
    .A_N(\soc_inst.cpu_core.alu.b[6] ));
 sg13g2_nor2_1 _19104_ (.A(\soc_inst.cpu_core.alu.b[6] ),
    .B(\soc_inst.cpu_core.alu.a[6] ),
    .Y(_04595_));
 sg13g2_nand2_1 _19105_ (.Y(_04596_),
    .A(\soc_inst.cpu_core.alu.b[6] ),
    .B(\soc_inst.cpu_core.alu.a[6] ));
 sg13g2_nand2b_2 _19106_ (.Y(_04597_),
    .B(_04596_),
    .A_N(_04595_));
 sg13g2_inv_1 _19107_ (.Y(_04598_),
    .A(_04597_));
 sg13g2_nor2b_1 _19108_ (.A(\soc_inst.cpu_core.alu.b[5] ),
    .B_N(\soc_inst.cpu_core.alu.a[5] ),
    .Y(_04599_));
 sg13g2_or2_1 _19109_ (.X(_04600_),
    .B(\soc_inst.cpu_core.alu.a[5] ),
    .A(\soc_inst.cpu_core.alu.b[5] ));
 sg13g2_and2_1 _19110_ (.A(\soc_inst.cpu_core.alu.b[5] ),
    .B(\soc_inst.cpu_core.alu.a[5] ),
    .X(_04601_));
 sg13g2_xnor2_1 _19111_ (.Y(_04602_),
    .A(\soc_inst.cpu_core.alu.b[5] ),
    .B(\soc_inst.cpu_core.alu.a[5] ));
 sg13g2_nand2_1 _19112_ (.Y(_04603_),
    .A(net6136),
    .B(\soc_inst.cpu_core.alu.a[4] ));
 sg13g2_nor2_1 _19113_ (.A(net6222),
    .B(\soc_inst.cpu_core.alu.a[4] ),
    .Y(_04604_));
 sg13g2_nand2_1 _19114_ (.Y(_04605_),
    .A(net6222),
    .B(\soc_inst.cpu_core.alu.a[4] ));
 sg13g2_nor2b_2 _19115_ (.A(_04604_),
    .B_N(_04605_),
    .Y(_04606_));
 sg13g2_nand2b_1 _19116_ (.Y(_04607_),
    .B(_04605_),
    .A_N(_04604_));
 sg13g2_nor2b_1 _19117_ (.A(net6230),
    .B_N(\soc_inst.cpu_core.alu.a[3] ),
    .Y(_04608_));
 sg13g2_or2_1 _19118_ (.X(_04609_),
    .B(\soc_inst.cpu_core.alu.a[3] ),
    .A(net6230));
 sg13g2_nand2_1 _19119_ (.Y(_04610_),
    .A(net6230),
    .B(\soc_inst.cpu_core.alu.a[3] ));
 sg13g2_inv_1 _19120_ (.Y(_04611_),
    .A(_04610_));
 sg13g2_and2_1 _19121_ (.A(_04609_),
    .B(_04610_),
    .X(_04612_));
 sg13g2_nand2_1 _19122_ (.Y(_04613_),
    .A(_04609_),
    .B(_04610_));
 sg13g2_nand2_1 _19123_ (.Y(_04614_),
    .A(net6123),
    .B(\soc_inst.cpu_core.alu.a[2] ));
 sg13g2_nor2_1 _19124_ (.A(net6238),
    .B(net3271),
    .Y(_04615_));
 sg13g2_and2_1 _19125_ (.A(net6238),
    .B(\soc_inst.cpu_core.alu.a[2] ),
    .X(_04616_));
 sg13g2_nor2_2 _19126_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sg13g2_nor2b_1 _19127_ (.A(net6241),
    .B_N(\soc_inst.cpu_core.alu.a[1] ),
    .Y(_04618_));
 sg13g2_nand2_1 _19128_ (.Y(_04619_),
    .A(net6241),
    .B(\soc_inst.cpu_core.alu.a[1] ));
 sg13g2_xnor2_1 _19129_ (.Y(_04620_),
    .A(net6241),
    .B(\soc_inst.cpu_core.alu.a[1] ));
 sg13g2_nand2b_1 _19130_ (.Y(_04621_),
    .B(net6252),
    .A_N(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_a21oi_1 _19131_ (.A1(_04620_),
    .A2(_04621_),
    .Y(_04622_),
    .B1(_04618_));
 sg13g2_o21ai_1 _19132_ (.B1(_04614_),
    .Y(_04623_),
    .A1(_04617_),
    .A2(_04622_));
 sg13g2_a21oi_1 _19133_ (.A1(_04613_),
    .A2(_04623_),
    .Y(_04624_),
    .B1(_04608_));
 sg13g2_o21ai_1 _19134_ (.B1(_04603_),
    .Y(_04625_),
    .A1(_04606_),
    .A2(_04624_));
 sg13g2_a21oi_1 _19135_ (.A1(_04602_),
    .A2(_04625_),
    .Y(_04626_),
    .B1(_04599_));
 sg13g2_o21ai_1 _19136_ (.B1(_04594_),
    .Y(_04627_),
    .A1(_04598_),
    .A2(_04626_));
 sg13g2_a21oi_1 _19137_ (.A1(_04593_),
    .A2(_04627_),
    .Y(_04628_),
    .B1(_04589_));
 sg13g2_nand2_1 _19138_ (.Y(_04629_),
    .A(\soc_inst.cpu_core.alu.b[8] ),
    .B(net6284));
 sg13g2_xor2_1 _19139_ (.B(net6284),
    .A(\soc_inst.cpu_core.alu.b[8] ),
    .X(_04630_));
 sg13g2_xnor2_1 _19140_ (.Y(_04631_),
    .A(\soc_inst.cpu_core.alu.b[8] ),
    .B(net6284));
 sg13g2_nand2b_1 _19141_ (.Y(_04632_),
    .B(_04631_),
    .A_N(_04628_));
 sg13g2_nand2b_1 _19142_ (.Y(_04633_),
    .B(_04585_),
    .A_N(_04632_));
 sg13g2_nor2b_1 _19143_ (.A(_04588_),
    .B_N(_04633_),
    .Y(_04634_));
 sg13g2_nor2b_1 _19144_ (.A(_04581_),
    .B_N(_04588_),
    .Y(_04635_));
 sg13g2_nor4_1 _19145_ (.A(_04581_),
    .B(_04584_),
    .C(_04628_),
    .D(_04630_),
    .Y(_04636_));
 sg13g2_nor3_2 _19146_ (.A(_04577_),
    .B(_04635_),
    .C(_04636_),
    .Y(_04637_));
 sg13g2_inv_1 _19147_ (.Y(_04638_),
    .A(_04637_));
 sg13g2_nor2_1 _19148_ (.A(\soc_inst.cpu_core.alu.b[12] ),
    .B(\soc_inst.cpu_core.alu.a[12] ),
    .Y(_04639_));
 sg13g2_nand2_2 _19149_ (.Y(_04640_),
    .A(net3040),
    .B(\soc_inst.cpu_core.alu.a[12] ));
 sg13g2_nand2b_2 _19150_ (.Y(_04641_),
    .B(_04640_),
    .A_N(_04639_));
 sg13g2_nor2b_1 _19151_ (.A(_04637_),
    .B_N(_04641_),
    .Y(_04642_));
 sg13g2_nand2_1 _19152_ (.Y(_04643_),
    .A(_04572_),
    .B(_04642_));
 sg13g2_nor3_1 _19153_ (.A(\soc_inst.cpu_core.alu.b[12] ),
    .B(_08201_),
    .C(_04571_),
    .Y(_04644_));
 sg13g2_a21oi_1 _19154_ (.A1(_08199_),
    .A2(\soc_inst.cpu_core.alu.a[13] ),
    .Y(_04645_),
    .B1(_04644_));
 sg13g2_o21ai_1 _19155_ (.B1(_04568_),
    .Y(_04646_),
    .A1(_04566_),
    .A2(_04645_));
 sg13g2_nor2b_1 _19156_ (.A(_04562_),
    .B_N(_04646_),
    .Y(_04647_));
 sg13g2_a21oi_1 _19157_ (.A1(_08197_),
    .A2(\soc_inst.cpu_core.alu.a[15] ),
    .Y(_04648_),
    .B1(_04647_));
 sg13g2_nand3_1 _19158_ (.B(_04572_),
    .C(_04641_),
    .A(_04567_),
    .Y(_04649_));
 sg13g2_o21ai_1 _19159_ (.B1(_04648_),
    .Y(_04650_),
    .A1(_04637_),
    .A2(_04649_));
 sg13g2_or2_1 _19160_ (.X(_04651_),
    .B(net6279),
    .A(\soc_inst.cpu_core.alu.b[17] ));
 sg13g2_and2_1 _19161_ (.A(\soc_inst.cpu_core.alu.b[17] ),
    .B(net6279),
    .X(_04652_));
 sg13g2_xor2_1 _19162_ (.B(net6279),
    .A(\soc_inst.cpu_core.alu.b[17] ),
    .X(_04653_));
 sg13g2_xnor2_1 _19163_ (.Y(_04654_),
    .A(\soc_inst.cpu_core.alu.b[17] ),
    .B(net6279));
 sg13g2_nand2_1 _19164_ (.Y(_04655_),
    .A(\soc_inst.cpu_core.alu.b[16] ),
    .B(net6281));
 sg13g2_xor2_1 _19165_ (.B(net6281),
    .A(\soc_inst.cpu_core.alu.b[16] ),
    .X(_04656_));
 sg13g2_xnor2_1 _19166_ (.Y(_04657_),
    .A(\soc_inst.cpu_core.alu.b[16] ),
    .B(net6281));
 sg13g2_nor2_2 _19167_ (.A(_04653_),
    .B(_04656_),
    .Y(_04658_));
 sg13g2_nand2_1 _19168_ (.Y(_04659_),
    .A(_04650_),
    .B(_04658_));
 sg13g2_nand2_1 _19169_ (.Y(_04660_),
    .A(\soc_inst.cpu_core.alu.b[21] ),
    .B(net6272));
 sg13g2_xor2_1 _19170_ (.B(net6272),
    .A(\soc_inst.cpu_core.alu.b[21] ),
    .X(_04661_));
 sg13g2_xnor2_1 _19171_ (.Y(_04662_),
    .A(\soc_inst.cpu_core.alu.b[21] ),
    .B(net6272));
 sg13g2_nor2_2 _19172_ (.A(\soc_inst.cpu_core.alu.b[22] ),
    .B(net6271),
    .Y(_04663_));
 sg13g2_nand2_2 _19173_ (.Y(_04664_),
    .A(\soc_inst.cpu_core.alu.b[22] ),
    .B(net6271));
 sg13g2_nor2b_2 _19174_ (.A(_04663_),
    .B_N(_04664_),
    .Y(_04665_));
 sg13g2_nand2b_2 _19175_ (.Y(_04666_),
    .B(_04664_),
    .A_N(_04663_));
 sg13g2_nand2_1 _19176_ (.Y(_04667_),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .B(net6275));
 sg13g2_xor2_1 _19177_ (.B(net6274),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .X(_04668_));
 sg13g2_xnor2_1 _19178_ (.Y(_04669_),
    .A(\soc_inst.cpu_core.alu.b[20] ),
    .B(net6274));
 sg13g2_nor2_1 _19179_ (.A(\soc_inst.cpu_core.alu.b[23] ),
    .B(net6270),
    .Y(_04670_));
 sg13g2_nand2_2 _19180_ (.Y(_04671_),
    .A(\soc_inst.cpu_core.alu.b[23] ),
    .B(net6270));
 sg13g2_nand2b_2 _19181_ (.Y(_04672_),
    .B(_04671_),
    .A_N(_04670_));
 sg13g2_nand3_1 _19182_ (.B(_04669_),
    .C(_04672_),
    .A(_04666_),
    .Y(_04673_));
 sg13g2_or2_1 _19183_ (.X(_04674_),
    .B(net6276),
    .A(\soc_inst.cpu_core.alu.b[19] ));
 sg13g2_and2_1 _19184_ (.A(\soc_inst.cpu_core.alu.b[19] ),
    .B(net6276),
    .X(_04675_));
 sg13g2_xor2_1 _19185_ (.B(net6276),
    .A(\soc_inst.cpu_core.alu.b[19] ),
    .X(_04676_));
 sg13g2_xnor2_1 _19186_ (.Y(_04677_),
    .A(\soc_inst.cpu_core.alu.b[19] ),
    .B(net6276));
 sg13g2_or2_1 _19187_ (.X(_04678_),
    .B(net6278),
    .A(\soc_inst.cpu_core.alu.b[18] ));
 sg13g2_and2_1 _19188_ (.A(\soc_inst.cpu_core.alu.b[18] ),
    .B(net6278),
    .X(_04679_));
 sg13g2_nand2_1 _19189_ (.Y(_04680_),
    .A(\soc_inst.cpu_core.alu.b[18] ),
    .B(net6278));
 sg13g2_and2_1 _19190_ (.A(_04678_),
    .B(_04680_),
    .X(_04681_));
 sg13g2_nor2_1 _19191_ (.A(_04676_),
    .B(_04681_),
    .Y(_04682_));
 sg13g2_nand2_1 _19192_ (.Y(_04683_),
    .A(_04658_),
    .B(_04682_));
 sg13g2_nor3_1 _19193_ (.A(_04661_),
    .B(_04673_),
    .C(_04683_),
    .Y(_04684_));
 sg13g2_nand2_1 _19194_ (.Y(_04685_),
    .A(_08193_),
    .B(net6271));
 sg13g2_nand2_1 _19195_ (.Y(_04686_),
    .A(_08194_),
    .B(net6272));
 sg13g2_nand3b_1 _19196_ (.B(net6281),
    .C(_04654_),
    .Y(_04687_),
    .A_N(\soc_inst.cpu_core.alu.b[16] ));
 sg13g2_o21ai_1 _19197_ (.B1(_04687_),
    .Y(_04688_),
    .A1(\soc_inst.cpu_core.alu.b[17] ),
    .A2(_08195_));
 sg13g2_nand2b_1 _19198_ (.Y(_04689_),
    .B(net6276),
    .A_N(\soc_inst.cpu_core.alu.b[19] ));
 sg13g2_nand2b_1 _19199_ (.Y(_04690_),
    .B(net6278),
    .A_N(\soc_inst.cpu_core.alu.b[18] ));
 sg13g2_o21ai_1 _19200_ (.B1(_04689_),
    .Y(_04691_),
    .A1(_04676_),
    .A2(_04690_));
 sg13g2_a21oi_1 _19201_ (.A1(_04682_),
    .A2(_04688_),
    .Y(_04692_),
    .B1(_04691_));
 sg13g2_nor2_1 _19202_ (.A(_04668_),
    .B(_04692_),
    .Y(_04693_));
 sg13g2_nor2b_1 _19203_ (.A(\soc_inst.cpu_core.alu.b[20] ),
    .B_N(net6274),
    .Y(_04694_));
 sg13g2_o21ai_1 _19204_ (.B1(_04662_),
    .Y(_04695_),
    .A1(_04693_),
    .A2(_04694_));
 sg13g2_and2_1 _19205_ (.A(_04686_),
    .B(_04695_),
    .X(_04696_));
 sg13g2_o21ai_1 _19206_ (.B1(_04685_),
    .Y(_04697_),
    .A1(_04665_),
    .A2(_04696_));
 sg13g2_and2_1 _19207_ (.A(_04672_),
    .B(_04697_),
    .X(_04698_));
 sg13g2_a221oi_1 _19208_ (.B2(_04684_),
    .C1(_04698_),
    .B1(_04650_),
    .A1(_08192_),
    .Y(_04699_),
    .A2(net6270));
 sg13g2_or2_1 _19209_ (.X(_04700_),
    .B(net6265),
    .A(\soc_inst.cpu_core.alu.b[27] ));
 sg13g2_and2_1 _19210_ (.A(\soc_inst.cpu_core.alu.b[27] ),
    .B(net6265),
    .X(_04701_));
 sg13g2_xnor2_1 _19211_ (.Y(_04702_),
    .A(\soc_inst.cpu_core.alu.b[27] ),
    .B(net6265));
 sg13g2_nand2_2 _19212_ (.Y(_04703_),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .B(net6266));
 sg13g2_nor2_1 _19213_ (.A(\soc_inst.cpu_core.alu.b[26] ),
    .B(net6266),
    .Y(_04704_));
 sg13g2_xor2_1 _19214_ (.B(net6266),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .X(_04705_));
 sg13g2_xnor2_1 _19215_ (.Y(_04706_),
    .A(\soc_inst.cpu_core.alu.b[26] ),
    .B(net6266));
 sg13g2_and2_1 _19216_ (.A(\soc_inst.cpu_core.alu.b[24] ),
    .B(net6269),
    .X(_04707_));
 sg13g2_or2_1 _19217_ (.X(_04708_),
    .B(net6269),
    .A(\soc_inst.cpu_core.alu.b[24] ));
 sg13g2_nor2b_1 _19218_ (.A(_04707_),
    .B_N(_04708_),
    .Y(_04709_));
 sg13g2_nand2b_2 _19219_ (.Y(_04710_),
    .B(_04708_),
    .A_N(_04707_));
 sg13g2_or2_1 _19220_ (.X(_04711_),
    .B(net6268),
    .A(\soc_inst.cpu_core.alu.b[25] ));
 sg13g2_and2_1 _19221_ (.A(\soc_inst.cpu_core.alu.b[25] ),
    .B(net6268),
    .X(_04712_));
 sg13g2_nand2_1 _19222_ (.Y(_04713_),
    .A(\soc_inst.cpu_core.alu.b[25] ),
    .B(net6268));
 sg13g2_and2_1 _19223_ (.A(_04711_),
    .B(_04713_),
    .X(_04714_));
 sg13g2_nand2_1 _19224_ (.Y(_04715_),
    .A(_04711_),
    .B(_04713_));
 sg13g2_nand4_1 _19225_ (.B(_04706_),
    .C(_04710_),
    .A(_04702_),
    .Y(_04716_),
    .D(_04715_));
 sg13g2_nand2_1 _19226_ (.Y(_04717_),
    .A(_08191_),
    .B(net6269));
 sg13g2_nor2_1 _19227_ (.A(_04714_),
    .B(_04717_),
    .Y(_04718_));
 sg13g2_a21oi_1 _19228_ (.A1(_08190_),
    .A2(net6268),
    .Y(_04719_),
    .B1(_04718_));
 sg13g2_nor2b_1 _19229_ (.A(\soc_inst.cpu_core.alu.b[27] ),
    .B_N(net6265),
    .Y(_04720_));
 sg13g2_nand2_1 _19230_ (.Y(_04721_),
    .A(_08189_),
    .B(net6266));
 sg13g2_o21ai_1 _19231_ (.B1(_04721_),
    .Y(_04722_),
    .A1(_04705_),
    .A2(_04719_));
 sg13g2_a21oi_1 _19232_ (.A1(_04702_),
    .A2(_04722_),
    .Y(_04723_),
    .B1(_04720_));
 sg13g2_o21ai_1 _19233_ (.B1(_04723_),
    .Y(_04724_),
    .A1(_04699_),
    .A2(_04716_));
 sg13g2_nand2_1 _19234_ (.Y(_04725_),
    .A(\soc_inst.cpu_core.alu.b[28] ),
    .B(net6264));
 sg13g2_xnor2_1 _19235_ (.Y(_04726_),
    .A(\soc_inst.cpu_core.alu.b[28] ),
    .B(net6264));
 sg13g2_nand2_1 _19236_ (.Y(_04727_),
    .A(_04724_),
    .B(_04726_));
 sg13g2_nand3_1 _19237_ (.B(_04724_),
    .C(_04726_),
    .A(_04559_),
    .Y(_04728_));
 sg13g2_nor2b_1 _19238_ (.A(\soc_inst.cpu_core.alu.b[29] ),
    .B_N(net6263),
    .Y(_04729_));
 sg13g2_nor2b_1 _19239_ (.A(\soc_inst.cpu_core.alu.b[28] ),
    .B_N(net6264),
    .Y(_04730_));
 sg13g2_a21oi_1 _19240_ (.A1(_04559_),
    .A2(_04730_),
    .Y(_04731_),
    .B1(_04729_));
 sg13g2_nor2_2 _19241_ (.A(_08187_),
    .B(_08188_),
    .Y(_04732_));
 sg13g2_xor2_1 _19242_ (.B(\soc_inst.cpu_core.alu.a[30] ),
    .A(\soc_inst.cpu_core.alu.b[30] ),
    .X(_04733_));
 sg13g2_inv_1 _19243_ (.Y(_04734_),
    .A(_04733_));
 sg13g2_a21o_1 _19244_ (.A2(_04731_),
    .A1(_04728_),
    .B1(_04733_),
    .X(_04735_));
 sg13g2_o21ai_1 _19245_ (.B1(_04735_),
    .Y(_04736_),
    .A1(\soc_inst.cpu_core.alu.b[30] ),
    .A2(_08188_));
 sg13g2_o21ai_1 _19246_ (.B1(_04557_),
    .Y(_04737_),
    .A1(_04558_),
    .A2(_04736_));
 sg13g2_nor2_2 _19247_ (.A(\soc_inst.cpu_core.alu.op[2] ),
    .B(\soc_inst.cpu_core.alu.op[3] ),
    .Y(_04738_));
 sg13g2_nand2_1 _19248_ (.Y(_04739_),
    .A(\soc_inst.cpu_core.alu.op[1] ),
    .B(_04738_));
 sg13g2_nor2_1 _19249_ (.A(net6287),
    .B(_04739_),
    .Y(_04740_));
 sg13g2_nand2b_1 _19250_ (.Y(_04741_),
    .B(_04736_),
    .A_N(_04558_));
 sg13g2_and4_1 _19251_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B(net6287),
    .C(_04557_),
    .D(_04738_),
    .X(_04742_));
 sg13g2_mux4_1 _19252_ (.S0(net6256),
    .A0(net6274),
    .A1(net6273),
    .A2(net6271),
    .A3(net6270),
    .S1(net6245),
    .X(_04743_));
 sg13g2_and2_1 _19253_ (.A(net6233),
    .B(_04743_),
    .X(_04744_));
 sg13g2_mux4_1 _19254_ (.S0(net6250),
    .A0(net6281),
    .A1(net6279),
    .A2(net6278),
    .A3(net6276),
    .S1(net6240),
    .X(_04745_));
 sg13g2_a21oi_1 _19255_ (.A1(net6122),
    .A2(_04745_),
    .Y(_04746_),
    .B1(_04744_));
 sg13g2_nor2b_1 _19256_ (.A(net6257),
    .B_N(net6264),
    .Y(_04747_));
 sg13g2_a21oi_1 _19257_ (.A1(net6263),
    .A2(net6257),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_mux2_1 _19258_ (.A0(\soc_inst.cpu_core.alu.a[30] ),
    .A1(net6262),
    .S(net6255),
    .X(_04749_));
 sg13g2_nand2_1 _19259_ (.Y(_04750_),
    .A(net6245),
    .B(_04749_));
 sg13g2_o21ai_1 _19260_ (.B1(_04750_),
    .Y(_04751_),
    .A1(net6245),
    .A2(_04748_));
 sg13g2_mux4_1 _19261_ (.S0(net6256),
    .A0(net6269),
    .A1(net6268),
    .A2(net6267),
    .A3(\soc_inst.cpu_core.alu.a[27] ),
    .S1(net6245),
    .X(_04752_));
 sg13g2_mux2_1 _19262_ (.A0(_04751_),
    .A1(_04752_),
    .S(net6121),
    .X(_04753_));
 sg13g2_nor2_1 _19263_ (.A(net6129),
    .B(_04753_),
    .Y(_04754_));
 sg13g2_a21oi_1 _19264_ (.A1(net6129),
    .A2(_04746_),
    .Y(_04755_),
    .B1(_04754_));
 sg13g2_nand3_1 _19265_ (.B(_04550_),
    .C(_04755_),
    .A(net6219),
    .Y(_04756_));
 sg13g2_nor2_1 _19266_ (.A(_08201_),
    .B(net6249),
    .Y(_04757_));
 sg13g2_a21oi_1 _19267_ (.A1(\soc_inst.cpu_core.alu.a[13] ),
    .A2(net6249),
    .Y(_04758_),
    .B1(_04757_));
 sg13g2_nand2_1 _19268_ (.Y(_04759_),
    .A(net6283),
    .B(net6111));
 sg13g2_nand2_1 _19269_ (.Y(_04760_),
    .A(\soc_inst.cpu_core.alu.a[15] ),
    .B(net6249));
 sg13g2_and3_1 _19270_ (.X(_04761_),
    .A(net6240),
    .B(_04759_),
    .C(_04760_));
 sg13g2_a21oi_1 _19271_ (.A1(net6115),
    .A2(_04758_),
    .Y(_04762_),
    .B1(_04761_));
 sg13g2_nand2_1 _19272_ (.Y(_04763_),
    .A(net6236),
    .B(_04762_));
 sg13g2_nor2b_1 _19273_ (.A(net6253),
    .B_N(net6284),
    .Y(_04764_));
 sg13g2_a21oi_1 _19274_ (.A1(\soc_inst.cpu_core.alu.a[9] ),
    .A2(net6253),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nand2_1 _19275_ (.Y(_04766_),
    .A(\soc_inst.cpu_core.alu.a[10] ),
    .B(net6111));
 sg13g2_nand2_1 _19276_ (.Y(_04767_),
    .A(\soc_inst.cpu_core.alu.a[11] ),
    .B(net6249));
 sg13g2_nand2_1 _19277_ (.Y(_04768_),
    .A(_04766_),
    .B(_04767_));
 sg13g2_nor2_1 _19278_ (.A(net6116),
    .B(_04768_),
    .Y(_04769_));
 sg13g2_a21oi_1 _19279_ (.A1(net6116),
    .A2(_04765_),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_inv_1 _19280_ (.Y(_04771_),
    .A(_04770_));
 sg13g2_o21ai_1 _19281_ (.B1(_04763_),
    .Y(_04772_),
    .A1(net6236),
    .A2(_04771_));
 sg13g2_nor2_2 _19282_ (.A(net6219),
    .B(_04551_),
    .Y(_04773_));
 sg13g2_nand2_2 _19283_ (.Y(_04774_),
    .A(net6136),
    .B(_04550_));
 sg13g2_nor2b_1 _19284_ (.A(net6251),
    .B_N(\soc_inst.cpu_core.alu.a[4] ),
    .Y(_04775_));
 sg13g2_nand2_1 _19285_ (.Y(_04776_),
    .A(\soc_inst.cpu_core.alu.a[5] ),
    .B(net6252));
 sg13g2_nand2b_1 _19286_ (.Y(_04777_),
    .B(_04776_),
    .A_N(_04775_));
 sg13g2_nand2_1 _19287_ (.Y(_04778_),
    .A(\soc_inst.cpu_core.alu.a[7] ),
    .B(net6253));
 sg13g2_o21ai_1 _19288_ (.B1(_04778_),
    .Y(_04779_),
    .A1(_08205_),
    .A2(net6252));
 sg13g2_mux2_1 _19289_ (.A0(_04777_),
    .A1(_04779_),
    .S(net6243),
    .X(_04780_));
 sg13g2_nand2_1 _19290_ (.Y(_04781_),
    .A(\soc_inst.cpu_core.alu.a[3] ),
    .B(net6251));
 sg13g2_o21ai_1 _19291_ (.B1(_04781_),
    .Y(_04782_),
    .A1(_08209_),
    .A2(net6251));
 sg13g2_nor2_2 _19292_ (.A(net6237),
    .B(net6116),
    .Y(_04783_));
 sg13g2_nand2_1 _19293_ (.Y(_04784_),
    .A(\soc_inst.cpu_core.alu.a[1] ),
    .B(net6252));
 sg13g2_nor2_2 _19294_ (.A(net6239),
    .B(net6248),
    .Y(_04785_));
 sg13g2_nand2_2 _19295_ (.Y(_04786_),
    .A(net6123),
    .B(net6116));
 sg13g2_nand2_2 _19296_ (.Y(_04787_),
    .A(net6112),
    .B(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_nor2_1 _19297_ (.A(net5769),
    .B(_04787_),
    .Y(_04788_));
 sg13g2_nor2_1 _19298_ (.A(net6227),
    .B(_04788_),
    .Y(_04789_));
 sg13g2_o21ai_1 _19299_ (.B1(_04789_),
    .Y(_04790_),
    .A1(_04784_),
    .A2(net5769));
 sg13g2_a221oi_1 _19300_ (.B2(_04783_),
    .C1(_04790_),
    .B1(_04782_),
    .A1(net6237),
    .Y(_04791_),
    .A2(_04780_));
 sg13g2_nor2_1 _19301_ (.A(_04774_),
    .B(_04791_),
    .Y(_04792_));
 sg13g2_o21ai_1 _19302_ (.B1(_04792_),
    .Y(_04793_),
    .A1(net6127),
    .A2(_04772_));
 sg13g2_nor2b_1 _19303_ (.A(net6285),
    .B_N(\soc_inst.cpu_core.alu.op[2] ),
    .Y(_04794_));
 sg13g2_and2_1 _19304_ (.A(\soc_inst.cpu_core.alu.op[1] ),
    .B(_04794_),
    .X(_04795_));
 sg13g2_nor2b_2 _19305_ (.A(net6286),
    .B_N(net5766),
    .Y(_04796_));
 sg13g2_nand2b_2 _19306_ (.Y(_04797_),
    .B(net5766),
    .A_N(net6286));
 sg13g2_and2_1 _19307_ (.A(net6251),
    .B(\soc_inst.cpu_core.alu.a[0] ),
    .X(_04798_));
 sg13g2_nand2_2 _19308_ (.Y(_04799_),
    .A(net6252),
    .B(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_nand2_1 _19309_ (.Y(_04800_),
    .A(\soc_inst.cpu_core.alu.op[2] ),
    .B(net6285));
 sg13g2_nand3_1 _19310_ (.B(_04799_),
    .C(_04800_),
    .A(_04547_),
    .Y(_04801_));
 sg13g2_nand2_1 _19311_ (.Y(_04802_),
    .A(_04797_),
    .B(_04801_));
 sg13g2_o21ai_1 _19312_ (.B1(_04802_),
    .Y(_04803_),
    .A1(net6251),
    .A2(\soc_inst.cpu_core.alu.a[0] ));
 sg13g2_and2_1 _19313_ (.A(net6286),
    .B(net5766),
    .X(_04804_));
 sg13g2_nand2_2 _19314_ (.Y(_04805_),
    .A(net6286),
    .B(net5766));
 sg13g2_nor3_2 _19315_ (.A(net6228),
    .B(net5769),
    .C(_04787_),
    .Y(_04806_));
 sg13g2_and2_1 _19316_ (.A(_04549_),
    .B(_04738_),
    .X(_04807_));
 sg13g2_nand2_2 _19317_ (.Y(_04808_),
    .A(_04549_),
    .B(_04738_));
 sg13g2_nor2_1 _19318_ (.A(net6221),
    .B(_04808_),
    .Y(_04809_));
 sg13g2_nand2_2 _19319_ (.Y(_04810_),
    .A(net6135),
    .B(_04807_));
 sg13g2_a22oi_1 _19320_ (.Y(_04811_),
    .B1(_04806_),
    .B2(net5457),
    .A2(net5459),
    .A1(_04798_));
 sg13g2_nand4_1 _19321_ (.B(_04793_),
    .C(_04803_),
    .A(_04756_),
    .Y(_04812_),
    .D(_04811_));
 sg13g2_a221oi_1 _19322_ (.B2(_04742_),
    .C1(_04812_),
    .B1(_04741_),
    .A1(_04737_),
    .Y(_04813_),
    .A2(_04740_));
 sg13g2_o21ai_1 _19323_ (.B1(_04546_),
    .Y(_01346_),
    .A1(_04556_),
    .A2(_04813_));
 sg13g2_and2_1 _19324_ (.A(net6285),
    .B(_04550_),
    .X(_04814_));
 sg13g2_mux4_1 _19325_ (.S0(net6258),
    .A0(net6273),
    .A1(net6271),
    .A2(net6270),
    .A3(net6269),
    .S1(net6246),
    .X(_04815_));
 sg13g2_mux4_1 _19326_ (.S0(net6256),
    .A0(net6279),
    .A1(net6278),
    .A2(net6276),
    .A3(net6274),
    .S1(net6245),
    .X(_04816_));
 sg13g2_mux2_1 _19327_ (.A0(_04815_),
    .A1(_04816_),
    .S(net6126),
    .X(_04817_));
 sg13g2_nand2_1 _19328_ (.Y(_04818_),
    .A(net6131),
    .B(_04817_));
 sg13g2_nor2b_1 _19329_ (.A(net6255),
    .B_N(net6265),
    .Y(_04819_));
 sg13g2_and2_1 _19330_ (.A(net6264),
    .B(net6255),
    .X(_04820_));
 sg13g2_mux4_1 _19331_ (.S0(net6255),
    .A0(net6268),
    .A1(net6266),
    .A2(net6265),
    .A3(\soc_inst.cpu_core.alu.a[28] ),
    .S1(net6246),
    .X(_04821_));
 sg13g2_and2_1 _19332_ (.A(net6120),
    .B(_04821_),
    .X(_04822_));
 sg13g2_nor2b_1 _19333_ (.A(net6255),
    .B_N(net6263),
    .Y(_04823_));
 sg13g2_a21oi_1 _19334_ (.A1(\soc_inst.cpu_core.alu.a[30] ),
    .A2(net6258),
    .Y(_04824_),
    .B1(_04823_));
 sg13g2_nor2_1 _19335_ (.A(net6247),
    .B(_04824_),
    .Y(_04825_));
 sg13g2_and2_1 _19336_ (.A(net6261),
    .B(net6234),
    .X(_04826_));
 sg13g2_nand2_1 _19337_ (.Y(_04827_),
    .A(net6261),
    .B(net6234));
 sg13g2_a21oi_1 _19338_ (.A1(net6261),
    .A2(net6247),
    .Y(_04828_),
    .B1(_04825_));
 sg13g2_a221oi_1 _19339_ (.B2(net6247),
    .C1(_04822_),
    .B1(_04826_),
    .A1(net6234),
    .Y(_04829_),
    .A2(_04825_));
 sg13g2_o21ai_1 _19340_ (.B1(_04818_),
    .Y(_04830_),
    .A1(net6131),
    .A2(_04829_));
 sg13g2_nor2_2 _19341_ (.A(net6285),
    .B(_04551_),
    .Y(_04831_));
 sg13g2_nand2_2 _19342_ (.Y(_04832_),
    .A(net6262),
    .B(net6111));
 sg13g2_nor2_1 _19343_ (.A(net6113),
    .B(_04832_),
    .Y(_04833_));
 sg13g2_or2_1 _19344_ (.X(_04834_),
    .B(_04833_),
    .A(_04825_));
 sg13g2_a21oi_1 _19345_ (.A1(net6234),
    .A2(_04834_),
    .Y(_04835_),
    .B1(_04822_));
 sg13g2_inv_1 _19346_ (.Y(_04836_),
    .A(_04835_));
 sg13g2_o21ai_1 _19347_ (.B1(_04818_),
    .Y(_04837_),
    .A1(net6131),
    .A2(_04835_));
 sg13g2_a22oi_1 _19348_ (.Y(_04838_),
    .B1(_04831_),
    .B2(_04837_),
    .A2(_04830_),
    .A1(net5455));
 sg13g2_nand2b_1 _19349_ (.Y(_04839_),
    .B(net6221),
    .A_N(_04838_));
 sg13g2_o21ai_1 _19350_ (.B1(net5461),
    .Y(_04840_),
    .A1(net6241),
    .A2(net2926));
 sg13g2_nor2_1 _19351_ (.A(_04619_),
    .B(_04805_),
    .Y(_04841_));
 sg13g2_and2_1 _19352_ (.A(_04547_),
    .B(_04794_),
    .X(_04842_));
 sg13g2_nand2_1 _19353_ (.Y(_04843_),
    .A(_04547_),
    .B(_04794_));
 sg13g2_o21ai_1 _19354_ (.B1(net6156),
    .Y(_04844_),
    .A1(_04620_),
    .A2(net5762));
 sg13g2_nor2_1 _19355_ (.A(_04841_),
    .B(_04844_),
    .Y(_04845_));
 sg13g2_a21oi_1 _19356_ (.A1(_04620_),
    .A2(_04621_),
    .Y(_04846_),
    .B1(net5771));
 sg13g2_o21ai_1 _19357_ (.B1(_04846_),
    .Y(_04847_),
    .A1(_04620_),
    .A2(_04621_));
 sg13g2_nor2_2 _19358_ (.A(net6229),
    .B(_04808_),
    .Y(_04848_));
 sg13g2_nand2_1 _19359_ (.Y(_04849_),
    .A(\soc_inst.cpu_core.alu.a[1] ),
    .B(net6112));
 sg13g2_a21oi_1 _19360_ (.A1(\soc_inst.cpu_core.alu.a[1] ),
    .A2(net6112),
    .Y(_04850_),
    .B1(_04798_));
 sg13g2_nand2b_1 _19361_ (.Y(_04851_),
    .B(_04785_),
    .A_N(_04850_));
 sg13g2_nor3_1 _19362_ (.A(net6229),
    .B(_04808_),
    .C(_04851_),
    .Y(_04852_));
 sg13g2_and2_1 _19363_ (.A(_04547_),
    .B(_04738_),
    .X(_04853_));
 sg13g2_nand2_1 _19364_ (.Y(_04854_),
    .A(_04547_),
    .B(_04738_));
 sg13g2_a21oi_1 _19365_ (.A1(_04620_),
    .A2(_04799_),
    .Y(_04855_),
    .B1(net5758));
 sg13g2_o21ai_1 _19366_ (.B1(_04855_),
    .Y(_04856_),
    .A1(_04620_),
    .A2(_04799_));
 sg13g2_nand4_1 _19367_ (.B(_04845_),
    .C(_04847_),
    .A(_04840_),
    .Y(_04857_),
    .D(_04856_));
 sg13g2_nor2_1 _19368_ (.A(_08200_),
    .B(net6250),
    .Y(_04858_));
 sg13g2_a21oi_1 _19369_ (.A1(net6283),
    .A2(net6250),
    .Y(_04859_),
    .B1(_04858_));
 sg13g2_nand2_1 _19370_ (.Y(_04860_),
    .A(net6281),
    .B(net6250));
 sg13g2_nand2_1 _19371_ (.Y(_04861_),
    .A(\soc_inst.cpu_core.alu.a[15] ),
    .B(net6111));
 sg13g2_and3_1 _19372_ (.X(_04862_),
    .A(net6244),
    .B(_04860_),
    .C(_04861_));
 sg13g2_a21oi_1 _19373_ (.A1(net6115),
    .A2(_04859_),
    .Y(_04863_),
    .B1(_04862_));
 sg13g2_nor2_1 _19374_ (.A(_08204_),
    .B(net6253),
    .Y(_04864_));
 sg13g2_a21oi_1 _19375_ (.A1(\soc_inst.cpu_core.alu.a[10] ),
    .A2(net6253),
    .Y(_04865_),
    .B1(_04864_));
 sg13g2_nand2_1 _19376_ (.Y(_04866_),
    .A(\soc_inst.cpu_core.alu.a[12] ),
    .B(net6249));
 sg13g2_nand2_1 _19377_ (.Y(_04867_),
    .A(\soc_inst.cpu_core.alu.a[11] ),
    .B(net6111));
 sg13g2_nand2_1 _19378_ (.Y(_04868_),
    .A(_04866_),
    .B(_04867_));
 sg13g2_nor2_1 _19379_ (.A(net6116),
    .B(_04868_),
    .Y(_04869_));
 sg13g2_a21oi_1 _19380_ (.A1(net6116),
    .A2(_04865_),
    .Y(_04870_),
    .B1(_04869_));
 sg13g2_mux2_1 _19381_ (.A0(_04863_),
    .A1(_04870_),
    .S(net6124),
    .X(_04871_));
 sg13g2_inv_1 _19382_ (.Y(_04872_),
    .A(_04871_));
 sg13g2_nand2_1 _19383_ (.Y(_04873_),
    .A(net6229),
    .B(_04872_));
 sg13g2_nor2b_1 _19384_ (.A(net6254),
    .B_N(\soc_inst.cpu_core.alu.a[5] ),
    .Y(_04874_));
 sg13g2_a21oi_1 _19385_ (.A1(\soc_inst.cpu_core.alu.a[6] ),
    .A2(net6251),
    .Y(_04875_),
    .B1(_04874_));
 sg13g2_mux2_1 _19386_ (.A0(\soc_inst.cpu_core.alu.a[7] ),
    .A1(net6284),
    .S(net6253),
    .X(_04876_));
 sg13g2_nor2_1 _19387_ (.A(net6117),
    .B(_04876_),
    .Y(_04877_));
 sg13g2_a21oi_1 _19388_ (.A1(net6118),
    .A2(_04875_),
    .Y(_04878_),
    .B1(_04877_));
 sg13g2_nand2_1 _19389_ (.Y(_04879_),
    .A(\soc_inst.cpu_core.alu.a[2] ),
    .B(net6251));
 sg13g2_a21oi_1 _19390_ (.A1(_04849_),
    .A2(_04879_),
    .Y(_04880_),
    .B1(net5769));
 sg13g2_nand2_1 _19391_ (.Y(_04881_),
    .A(\soc_inst.cpu_core.alu.a[4] ),
    .B(net6251));
 sg13g2_nand2_1 _19392_ (.Y(_04882_),
    .A(\soc_inst.cpu_core.alu.a[3] ),
    .B(net6112));
 sg13g2_nand2_1 _19393_ (.Y(_04883_),
    .A(_04881_),
    .B(_04882_));
 sg13g2_a221oi_1 _19394_ (.B2(_04783_),
    .C1(_04880_),
    .B1(_04883_),
    .A1(net6238),
    .Y(_04884_),
    .A2(_04878_));
 sg13g2_a21oi_1 _19395_ (.A1(net6127),
    .A2(_04884_),
    .Y(_04885_),
    .B1(_04774_));
 sg13g2_a221oi_1 _19396_ (.B2(_04885_),
    .C1(_04857_),
    .B1(_04873_),
    .A1(net6136),
    .Y(_04886_),
    .A2(_04852_));
 sg13g2_a22oi_1 _19397_ (.Y(_01347_),
    .B1(_04839_),
    .B2(_04886_),
    .A2(net6424),
    .A1(_07870_));
 sg13g2_mux4_1 _19398_ (.S0(net6256),
    .A0(net6278),
    .A1(net6277),
    .A2(net6274),
    .A3(net6273),
    .S1(net6245),
    .X(_04887_));
 sg13g2_mux4_1 _19399_ (.S0(net6255),
    .A0(net6271),
    .A1(net6270),
    .A2(net6269),
    .A3(net6268),
    .S1(net6246),
    .X(_04888_));
 sg13g2_mux2_1 _19400_ (.A0(_04887_),
    .A1(_04888_),
    .S(net6236),
    .X(_04889_));
 sg13g2_inv_1 _19401_ (.Y(_04890_),
    .A(_04889_));
 sg13g2_nand2_1 _19402_ (.Y(_04891_),
    .A(net6134),
    .B(_04889_));
 sg13g2_nand2_2 _19403_ (.Y(_04892_),
    .A(net6237),
    .B(net6117));
 sg13g2_nand2_1 _19404_ (.Y(_04893_),
    .A(net6113),
    .B(_04749_));
 sg13g2_nor2_1 _19405_ (.A(net6120),
    .B(_04893_),
    .Y(_04894_));
 sg13g2_mux4_1 _19406_ (.S0(net6255),
    .A0(net6266),
    .A1(net6265),
    .A2(\soc_inst.cpu_core.alu.a[28] ),
    .A3(\soc_inst.cpu_core.alu.a[29] ),
    .S1(net6245),
    .X(_04895_));
 sg13g2_a21oi_2 _19407_ (.B1(_04894_),
    .Y(_04896_),
    .A2(_04895_),
    .A1(net6120));
 sg13g2_o21ai_1 _19408_ (.B1(_04891_),
    .Y(_04897_),
    .A1(net6131),
    .A2(_04896_));
 sg13g2_o21ai_1 _19409_ (.B1(_04896_),
    .Y(_04898_),
    .A1(net6113),
    .A2(_04827_));
 sg13g2_nand2_1 _19410_ (.Y(_04899_),
    .A(net6225),
    .B(_04898_));
 sg13g2_nand2_1 _19411_ (.Y(_04900_),
    .A(_04891_),
    .B(_04899_));
 sg13g2_a22oi_1 _19412_ (.Y(_04901_),
    .B1(_04900_),
    .B2(net5455),
    .A2(_04897_),
    .A1(_04831_));
 sg13g2_nor2_1 _19413_ (.A(net6136),
    .B(_04901_),
    .Y(_04902_));
 sg13g2_mux4_1 _19414_ (.S0(net6249),
    .A0(\soc_inst.cpu_core.alu.a[14] ),
    .A1(\soc_inst.cpu_core.alu.a[15] ),
    .A2(net6282),
    .A3(net6279),
    .S1(net6240),
    .X(_04903_));
 sg13g2_nor2_1 _19415_ (.A(net6240),
    .B(_04768_),
    .Y(_04904_));
 sg13g2_a21oi_1 _19416_ (.A1(net6240),
    .A2(_04758_),
    .Y(_04905_),
    .B1(_04904_));
 sg13g2_mux2_1 _19417_ (.A0(_04903_),
    .A1(_04905_),
    .S(net6122),
    .X(_04906_));
 sg13g2_nor2_1 _19418_ (.A(net6242),
    .B(_04779_),
    .Y(_04907_));
 sg13g2_a21oi_1 _19419_ (.A1(net6242),
    .A2(_04765_),
    .Y(_04908_),
    .B1(_04907_));
 sg13g2_a22oi_1 _19420_ (.Y(_04909_),
    .B1(_04785_),
    .B2(_04782_),
    .A2(_04783_),
    .A1(_04777_));
 sg13g2_a21oi_1 _19421_ (.A1(net6237),
    .A2(_04908_),
    .Y(_04910_),
    .B1(net6228));
 sg13g2_o21ai_1 _19422_ (.B1(net5462),
    .Y(_04911_),
    .A1(net6127),
    .A2(_04906_));
 sg13g2_a21oi_1 _19423_ (.A1(_04909_),
    .A2(_04910_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_o21ai_1 _19424_ (.B1(_04784_),
    .Y(_04913_),
    .A1(_08209_),
    .A2(net6252));
 sg13g2_nand2_1 _19425_ (.Y(_04914_),
    .A(net6241),
    .B(_04787_));
 sg13g2_o21ai_1 _19426_ (.B1(_04914_),
    .Y(_04915_),
    .A1(net6241),
    .A2(_04913_));
 sg13g2_nand2b_2 _19427_ (.Y(_04916_),
    .B(net6123),
    .A_N(_04915_));
 sg13g2_nor3_1 _19428_ (.A(net6230),
    .B(_04810_),
    .C(_04916_),
    .Y(_04917_));
 sg13g2_o21ai_1 _19429_ (.B1(_04619_),
    .Y(_04918_),
    .A1(_04620_),
    .A2(_04799_));
 sg13g2_xor2_1 _19430_ (.B(_04918_),
    .A(_04617_),
    .X(_04919_));
 sg13g2_a21o_1 _19431_ (.A2(_04919_),
    .A1(net5760),
    .B1(_04917_),
    .X(_04920_));
 sg13g2_o21ai_1 _19432_ (.B1(net5774),
    .Y(_04921_),
    .A1(_04617_),
    .A2(_04622_));
 sg13g2_a21o_1 _19433_ (.A2(_04622_),
    .A1(_04617_),
    .B1(_04921_),
    .X(_04922_));
 sg13g2_nor2_1 _19434_ (.A(_04616_),
    .B(net5762),
    .Y(_04923_));
 sg13g2_nor2_1 _19435_ (.A(net5461),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_a21oi_1 _19436_ (.A1(_04616_),
    .A2(net5459),
    .Y(_04925_),
    .B1(net6422));
 sg13g2_o21ai_1 _19437_ (.B1(_04925_),
    .Y(_04926_),
    .A1(_04615_),
    .A2(_04924_));
 sg13g2_nor4_1 _19438_ (.A(_04902_),
    .B(_04912_),
    .C(_04920_),
    .D(_04926_),
    .Y(_04927_));
 sg13g2_a22oi_1 _19439_ (.Y(_01348_),
    .B1(_04922_),
    .B2(_04927_),
    .A2(_08160_),
    .A1(net6424));
 sg13g2_mux4_1 _19440_ (.S0(net6255),
    .A0(net6270),
    .A1(net6269),
    .A2(\soc_inst.cpu_core.alu.a[25] ),
    .A3(net6267),
    .S1(net6245),
    .X(_04928_));
 sg13g2_mux4_1 _19441_ (.S0(net6259),
    .A0(net6277),
    .A1(net6275),
    .A2(net6272),
    .A3(net6271),
    .S1(net6247),
    .X(_04929_));
 sg13g2_mux2_1 _19442_ (.A0(_04928_),
    .A1(_04929_),
    .S(net6121),
    .X(_04930_));
 sg13g2_nand2_1 _19443_ (.Y(_04931_),
    .A(net6131),
    .B(_04930_));
 sg13g2_nor3_1 _19444_ (.A(net6247),
    .B(_04819_),
    .C(_04820_),
    .Y(_04932_));
 sg13g2_a21oi_2 _19445_ (.B1(_04932_),
    .Y(_04933_),
    .A2(_04824_),
    .A1(net6247));
 sg13g2_nand2_1 _19446_ (.Y(_04934_),
    .A(net6120),
    .B(_04933_));
 sg13g2_o21ai_1 _19447_ (.B1(_04934_),
    .Y(_04935_),
    .A1(_04832_),
    .A2(_04892_));
 sg13g2_nand2_1 _19448_ (.Y(_04936_),
    .A(net6231),
    .B(_04935_));
 sg13g2_nand2_1 _19449_ (.Y(_04937_),
    .A(_04931_),
    .B(_04936_));
 sg13g2_a21oi_1 _19450_ (.A1(net6120),
    .A2(_04933_),
    .Y(_04938_),
    .B1(_04826_));
 sg13g2_o21ai_1 _19451_ (.B1(_04931_),
    .Y(_04939_),
    .A1(net6131),
    .A2(_04938_));
 sg13g2_a22oi_1 _19452_ (.Y(_04940_),
    .B1(_04939_),
    .B2(_04814_),
    .A2(_04937_),
    .A1(_04831_));
 sg13g2_nand2b_1 _19453_ (.Y(_04941_),
    .B(net6222),
    .A_N(_04940_));
 sg13g2_xnor2_1 _19454_ (.Y(_04942_),
    .A(_04612_),
    .B(_04623_));
 sg13g2_a21o_1 _19455_ (.A2(_04918_),
    .A1(_04617_),
    .B1(_04616_),
    .X(_04943_));
 sg13g2_xnor2_1 _19456_ (.Y(_04944_),
    .A(_04612_),
    .B(_04943_));
 sg13g2_nor2_1 _19457_ (.A(net6240),
    .B(_04868_),
    .Y(_04945_));
 sg13g2_a21oi_1 _19458_ (.A1(net6244),
    .A2(_04859_),
    .Y(_04946_),
    .B1(_04945_));
 sg13g2_mux4_1 _19459_ (.S0(net6249),
    .A0(\soc_inst.cpu_core.alu.a[15] ),
    .A1(net6282),
    .A2(net6280),
    .A3(\soc_inst.cpu_core.alu.a[18] ),
    .S1(net6240),
    .X(_04947_));
 sg13g2_mux2_1 _19460_ (.A0(_04946_),
    .A1(_04947_),
    .S(net6236),
    .X(_04948_));
 sg13g2_nor2_1 _19461_ (.A(net6242),
    .B(_04876_),
    .Y(_04949_));
 sg13g2_a21oi_1 _19462_ (.A1(net6242),
    .A2(_04865_),
    .Y(_04950_),
    .B1(_04949_));
 sg13g2_nand2_1 _19463_ (.Y(_04951_),
    .A(net6237),
    .B(_04950_));
 sg13g2_nor2b_1 _19464_ (.A(_04875_),
    .B_N(_04783_),
    .Y(_04952_));
 sg13g2_a21oi_1 _19465_ (.A1(_04881_),
    .A2(_04882_),
    .Y(_04953_),
    .B1(net5769));
 sg13g2_nor3_1 _19466_ (.A(net6230),
    .B(_04952_),
    .C(_04953_),
    .Y(_04954_));
 sg13g2_o21ai_1 _19467_ (.B1(net5462),
    .Y(_04955_),
    .A1(net6127),
    .A2(_04948_));
 sg13g2_a21oi_1 _19468_ (.A1(_04951_),
    .A2(_04954_),
    .Y(_04956_),
    .B1(_04955_));
 sg13g2_nand2_1 _19469_ (.Y(_04957_),
    .A(_04879_),
    .B(_04882_));
 sg13g2_nor2_1 _19470_ (.A(net6243),
    .B(_04957_),
    .Y(_04958_));
 sg13g2_a21oi_1 _19471_ (.A1(net6243),
    .A2(_04850_),
    .Y(_04959_),
    .B1(_04958_));
 sg13g2_nand2_2 _19472_ (.Y(_04960_),
    .A(net6123),
    .B(_04959_));
 sg13g2_nor3_1 _19473_ (.A(net6230),
    .B(_04810_),
    .C(_04960_),
    .Y(_04961_));
 sg13g2_a221oi_1 _19474_ (.B2(_04612_),
    .C1(net6422),
    .B1(net5765),
    .A1(_04609_),
    .Y(_04962_),
    .A2(net5461));
 sg13g2_o21ai_1 _19475_ (.B1(_04962_),
    .Y(_04963_),
    .A1(_04610_),
    .A2(_04805_));
 sg13g2_nor3_1 _19476_ (.A(_04956_),
    .B(_04961_),
    .C(_04963_),
    .Y(_04964_));
 sg13g2_o21ai_1 _19477_ (.B1(_04964_),
    .Y(_04965_),
    .A1(net5758),
    .A2(_04944_));
 sg13g2_a21oi_1 _19478_ (.A1(net5774),
    .A2(_04942_),
    .Y(_04966_),
    .B1(_04965_));
 sg13g2_a22oi_1 _19479_ (.Y(_01349_),
    .B1(_04941_),
    .B2(_04966_),
    .A2(_08161_),
    .A1(net6425));
 sg13g2_a21oi_1 _19480_ (.A1(_04612_),
    .A2(_04943_),
    .Y(_04967_),
    .B1(_04611_));
 sg13g2_o21ai_1 _19481_ (.B1(net5760),
    .Y(_04968_),
    .A1(_04607_),
    .A2(_04967_));
 sg13g2_a21o_1 _19482_ (.A2(_04967_),
    .A1(_04607_),
    .B1(_04968_),
    .X(_04969_));
 sg13g2_xnor2_1 _19483_ (.Y(_04970_),
    .A(_04606_),
    .B(_04624_));
 sg13g2_o21ai_1 _19484_ (.B1(_04969_),
    .Y(_04971_),
    .A1(net5771),
    .A2(_04970_));
 sg13g2_mux2_1 _19485_ (.A0(_04743_),
    .A1(_04752_),
    .S(net6233),
    .X(_04972_));
 sg13g2_and2_1 _19486_ (.A(net6130),
    .B(_04972_),
    .X(_04973_));
 sg13g2_and2_1 _19487_ (.A(net6121),
    .B(_04751_),
    .X(_04974_));
 sg13g2_a21o_1 _19488_ (.A2(_04974_),
    .A1(net6226),
    .B1(_04973_),
    .X(_04975_));
 sg13g2_or2_1 _19489_ (.X(_04976_),
    .B(_04974_),
    .A(_04826_));
 sg13g2_a21o_1 _19490_ (.A2(_04976_),
    .A1(net6226),
    .B1(_04973_),
    .X(_04977_));
 sg13g2_a22oi_1 _19491_ (.Y(_04978_),
    .B1(_04977_),
    .B2(net5455),
    .A2(_04975_),
    .A1(_04831_));
 sg13g2_nand2b_1 _19492_ (.Y(_04979_),
    .B(net6221),
    .A_N(_04978_));
 sg13g2_mux2_1 _19493_ (.A0(_04745_),
    .A1(_04762_),
    .S(net6122),
    .X(_04980_));
 sg13g2_a21oi_1 _19494_ (.A1(net6237),
    .A2(_04771_),
    .Y(_04981_),
    .B1(net6228));
 sg13g2_o21ai_1 _19495_ (.B1(_04981_),
    .Y(_04982_),
    .A1(net6237),
    .A2(_04780_));
 sg13g2_nand2_1 _19496_ (.Y(_04983_),
    .A(net6227),
    .B(_04980_));
 sg13g2_a21oi_1 _19497_ (.A1(_04982_),
    .A2(_04983_),
    .Y(_04984_),
    .B1(_04774_));
 sg13g2_nor2_1 _19498_ (.A(_04787_),
    .B(_04892_),
    .Y(_04985_));
 sg13g2_nor2b_1 _19499_ (.A(_04775_),
    .B_N(_04781_),
    .Y(_04986_));
 sg13g2_nand2_1 _19500_ (.Y(_04987_),
    .A(net6241),
    .B(_04913_));
 sg13g2_o21ai_1 _19501_ (.B1(_04987_),
    .Y(_04988_),
    .A1(net6241),
    .A2(_04986_));
 sg13g2_a21oi_1 _19502_ (.A1(net6124),
    .A2(_04988_),
    .Y(_04989_),
    .B1(_04985_));
 sg13g2_or2_1 _19503_ (.X(_04990_),
    .B(_04989_),
    .A(net6227));
 sg13g2_nor2_1 _19504_ (.A(_04604_),
    .B(_04797_),
    .Y(_04991_));
 sg13g2_a21oi_1 _19505_ (.A1(_04606_),
    .A2(net5765),
    .Y(_04992_),
    .B1(net6419));
 sg13g2_o21ai_1 _19506_ (.B1(_04992_),
    .Y(_04993_),
    .A1(_04605_),
    .A2(_04805_));
 sg13g2_nor3_1 _19507_ (.A(_04984_),
    .B(_04991_),
    .C(_04993_),
    .Y(_04994_));
 sg13g2_o21ai_1 _19508_ (.B1(_04994_),
    .Y(_04995_),
    .A1(_04810_),
    .A2(_04990_));
 sg13g2_nor2_1 _19509_ (.A(_04971_),
    .B(_04995_),
    .Y(_04996_));
 sg13g2_a22oi_1 _19510_ (.Y(_01350_),
    .B1(_04979_),
    .B2(_04996_),
    .A2(_08162_),
    .A1(net6425));
 sg13g2_o21ai_1 _19511_ (.B1(_04605_),
    .Y(_04997_),
    .A1(_04607_),
    .A2(_04967_));
 sg13g2_xnor2_1 _19512_ (.Y(_04998_),
    .A(_04602_),
    .B(_04997_));
 sg13g2_xor2_1 _19513_ (.B(_04625_),
    .A(_04602_),
    .X(_04999_));
 sg13g2_mux2_1 _19514_ (.A0(_04815_),
    .A1(_04821_),
    .S(net6234),
    .X(_05000_));
 sg13g2_nand2_1 _19515_ (.Y(_05001_),
    .A(net6131),
    .B(_05000_));
 sg13g2_and2_1 _19516_ (.A(net6120),
    .B(_04834_),
    .X(_05002_));
 sg13g2_nand2_1 _19517_ (.Y(_05003_),
    .A(net6231),
    .B(_05002_));
 sg13g2_nand2_1 _19518_ (.Y(_05004_),
    .A(_05001_),
    .B(_05003_));
 sg13g2_o21ai_1 _19519_ (.B1(_04827_),
    .Y(_05005_),
    .A1(net6235),
    .A2(_04828_));
 sg13g2_nand2_1 _19520_ (.Y(_05006_),
    .A(net6231),
    .B(_05005_));
 sg13g2_nand2_1 _19521_ (.Y(_05007_),
    .A(_05001_),
    .B(_05006_));
 sg13g2_a22oi_1 _19522_ (.Y(_05008_),
    .B1(_05007_),
    .B2(net5455),
    .A2(_05004_),
    .A1(_04831_));
 sg13g2_nor2_1 _19523_ (.A(_04850_),
    .B(_04892_),
    .Y(_05009_));
 sg13g2_nor2b_1 _19524_ (.A(_04874_),
    .B_N(_04881_),
    .Y(_05010_));
 sg13g2_nand2_1 _19525_ (.Y(_05011_),
    .A(net6243),
    .B(_04957_));
 sg13g2_o21ai_1 _19526_ (.B1(_05011_),
    .Y(_05012_),
    .A1(net6243),
    .A2(_05010_));
 sg13g2_a21oi_1 _19527_ (.A1(net6123),
    .A2(_05012_),
    .Y(_05013_),
    .B1(_05009_));
 sg13g2_nor2_2 _19528_ (.A(net6228),
    .B(_05013_),
    .Y(_05014_));
 sg13g2_a221oi_1 _19529_ (.B2(_04601_),
    .C1(net6418),
    .B1(net5459),
    .A1(_04600_),
    .Y(_05015_),
    .A2(net5461));
 sg13g2_o21ai_1 _19530_ (.B1(_05015_),
    .Y(_05016_),
    .A1(_04602_),
    .A2(net5762));
 sg13g2_nor2_1 _19531_ (.A(net6237),
    .B(_04878_),
    .Y(_05017_));
 sg13g2_nor2_1 _19532_ (.A(net6124),
    .B(_04870_),
    .Y(_05018_));
 sg13g2_o21ai_1 _19533_ (.B1(net6127),
    .Y(_05019_),
    .A1(_05017_),
    .A2(_05018_));
 sg13g2_mux2_1 _19534_ (.A0(_04816_),
    .A1(_04863_),
    .S(net6120),
    .X(_05020_));
 sg13g2_inv_1 _19535_ (.Y(_05021_),
    .A(_05020_));
 sg13g2_a21oi_1 _19536_ (.A1(net6227),
    .A2(_05021_),
    .Y(_05022_),
    .B1(_04774_));
 sg13g2_a221oi_1 _19537_ (.B2(_05022_),
    .C1(_05016_),
    .B1(_05019_),
    .A1(net5457),
    .Y(_05023_),
    .A2(_05014_));
 sg13g2_o21ai_1 _19538_ (.B1(_05023_),
    .Y(_05024_),
    .A1(net6136),
    .A2(_05008_));
 sg13g2_a221oi_1 _19539_ (.B2(net5774),
    .C1(_05024_),
    .B1(_04999_),
    .A1(_04853_),
    .Y(_05025_),
    .A2(_04998_));
 sg13g2_a21oi_1 _19540_ (.A1(net6375),
    .A2(_08163_),
    .Y(_01351_),
    .B1(_05025_));
 sg13g2_a21oi_1 _19541_ (.A1(_04600_),
    .A2(_04997_),
    .Y(_05026_),
    .B1(_04601_));
 sg13g2_xnor2_1 _19542_ (.Y(_05027_),
    .A(_04598_),
    .B(_05026_));
 sg13g2_xnor2_1 _19543_ (.Y(_05028_),
    .A(_04597_),
    .B(_04626_));
 sg13g2_mux2_1 _19544_ (.A0(_04888_),
    .A1(_04895_),
    .S(net6233),
    .X(_05029_));
 sg13g2_nand2_1 _19545_ (.Y(_05030_),
    .A(net6130),
    .B(_05029_));
 sg13g2_nor2_1 _19546_ (.A(net6234),
    .B(_04893_),
    .Y(_05031_));
 sg13g2_nand2_1 _19547_ (.Y(_05032_),
    .A(net6225),
    .B(_05031_));
 sg13g2_nand2_1 _19548_ (.Y(_05033_),
    .A(_05030_),
    .B(_05032_));
 sg13g2_a21oi_1 _19549_ (.A1(net6261),
    .A2(net5769),
    .Y(_05034_),
    .B1(_05031_));
 sg13g2_o21ai_1 _19550_ (.B1(_05030_),
    .Y(_05035_),
    .A1(net6133),
    .A2(_05034_));
 sg13g2_a22oi_1 _19551_ (.Y(_05036_),
    .B1(_05035_),
    .B2(net5455),
    .A2(_05033_),
    .A1(_04831_));
 sg13g2_nor2_1 _19552_ (.A(net6136),
    .B(_05036_),
    .Y(_05037_));
 sg13g2_nand2_1 _19553_ (.Y(_05038_),
    .A(net6124),
    .B(_04908_));
 sg13g2_a21oi_1 _19554_ (.A1(net6236),
    .A2(_04905_),
    .Y(_05039_),
    .B1(net6227));
 sg13g2_mux2_1 _19555_ (.A0(_04887_),
    .A1(_04903_),
    .S(net6120),
    .X(_05040_));
 sg13g2_inv_2 _19556_ (.Y(_05041_),
    .A(_05040_));
 sg13g2_a221oi_1 _19557_ (.B2(net6227),
    .C1(_04774_),
    .B1(_05041_),
    .A1(_05038_),
    .Y(_05042_),
    .A2(_05039_));
 sg13g2_nand2_1 _19558_ (.Y(_05043_),
    .A(_04598_),
    .B(net5765));
 sg13g2_o21ai_1 _19559_ (.B1(_05043_),
    .Y(_05044_),
    .A1(_04595_),
    .A2(_04797_));
 sg13g2_o21ai_1 _19560_ (.B1(net6156),
    .Y(_05045_),
    .A1(_04596_),
    .A2(_04805_));
 sg13g2_nor2_1 _19561_ (.A(net6123),
    .B(_04915_),
    .Y(_05046_));
 sg13g2_o21ai_1 _19562_ (.B1(_04776_),
    .Y(_05047_),
    .A1(_08205_),
    .A2(net6252));
 sg13g2_nor2_1 _19563_ (.A(net6242),
    .B(_05047_),
    .Y(_05048_));
 sg13g2_a21oi_1 _19564_ (.A1(net6242),
    .A2(_04986_),
    .Y(_05049_),
    .B1(_05048_));
 sg13g2_a21oi_1 _19565_ (.A1(net6124),
    .A2(_05049_),
    .Y(_05050_),
    .B1(_05046_));
 sg13g2_nor2_1 _19566_ (.A(net6227),
    .B(_05050_),
    .Y(_05051_));
 sg13g2_a21o_1 _19567_ (.A2(_05051_),
    .A1(net5457),
    .B1(_05042_),
    .X(_05052_));
 sg13g2_or4_1 _19568_ (.A(_05037_),
    .B(_05044_),
    .C(_05045_),
    .D(_05052_),
    .X(_05053_));
 sg13g2_a221oi_1 _19569_ (.B2(net5774),
    .C1(_05053_),
    .B1(_05028_),
    .A1(_04853_),
    .Y(_05054_),
    .A2(_05027_));
 sg13g2_a21oi_1 _19570_ (.A1(net6375),
    .A2(_08164_),
    .Y(_01352_),
    .B1(_05054_));
 sg13g2_xor2_1 _19571_ (.B(_04627_),
    .A(_04593_),
    .X(_05055_));
 sg13g2_o21ai_1 _19572_ (.B1(_04596_),
    .Y(_05056_),
    .A1(_04597_),
    .A2(_05026_));
 sg13g2_nand2b_1 _19573_ (.Y(_05057_),
    .B(_04593_),
    .A_N(_05056_));
 sg13g2_nand2b_1 _19574_ (.Y(_05058_),
    .B(_05056_),
    .A_N(_04593_));
 sg13g2_and2_1 _19575_ (.A(_04853_),
    .B(_05057_),
    .X(_05059_));
 sg13g2_nand2_1 _19576_ (.Y(_05060_),
    .A(net6124),
    .B(_04950_));
 sg13g2_a21oi_1 _19577_ (.A1(net6236),
    .A2(_04946_),
    .Y(_05061_),
    .B1(net6223));
 sg13g2_mux2_1 _19578_ (.A0(_04929_),
    .A1(_04947_),
    .S(net6122),
    .X(_05062_));
 sg13g2_o21ai_1 _19579_ (.B1(net5462),
    .Y(_05063_),
    .A1(net6129),
    .A2(_05062_));
 sg13g2_a21oi_1 _19580_ (.A1(_05060_),
    .A2(_05061_),
    .Y(_05064_),
    .B1(_05063_));
 sg13g2_mux2_1 _19581_ (.A0(\soc_inst.cpu_core.alu.a[7] ),
    .A1(\soc_inst.cpu_core.alu.a[6] ),
    .S(net6252),
    .X(_05065_));
 sg13g2_nor2_1 _19582_ (.A(net6243),
    .B(_05065_),
    .Y(_05066_));
 sg13g2_a21oi_1 _19583_ (.A1(net6243),
    .A2(_05010_),
    .Y(_05067_),
    .B1(_05066_));
 sg13g2_mux2_1 _19584_ (.A0(_04959_),
    .A1(_05067_),
    .S(net6123),
    .X(_05068_));
 sg13g2_and2_1 _19585_ (.A(_08207_),
    .B(_05068_),
    .X(_05069_));
 sg13g2_a22oi_1 _19586_ (.Y(_05070_),
    .B1(net5459),
    .B2(_04590_),
    .A2(net5461),
    .A1(_04592_));
 sg13g2_o21ai_1 _19587_ (.B1(net6156),
    .Y(_05071_),
    .A1(_04593_),
    .A2(net5762));
 sg13g2_nand2b_1 _19588_ (.Y(_05072_),
    .B(_05070_),
    .A_N(_05071_));
 sg13g2_mux2_1 _19589_ (.A0(_04928_),
    .A1(_04933_),
    .S(net6234),
    .X(_05073_));
 sg13g2_inv_1 _19590_ (.Y(_05074_),
    .A(_05073_));
 sg13g2_and2_1 _19591_ (.A(net6262),
    .B(net5455),
    .X(_05075_));
 sg13g2_and2_1 _19592_ (.A(net6130),
    .B(net5455),
    .X(_05076_));
 sg13g2_nand2_1 _19593_ (.Y(_05077_),
    .A(net6133),
    .B(net5455));
 sg13g2_nor2_1 _19594_ (.A(_05075_),
    .B(_05076_),
    .Y(_05078_));
 sg13g2_o21ai_1 _19595_ (.B1(net6231),
    .Y(_05079_),
    .A1(net5769),
    .A2(_04832_));
 sg13g2_nand2_1 _19596_ (.Y(_05080_),
    .A(_04831_),
    .B(_05079_));
 sg13g2_and2_1 _19597_ (.A(net6226),
    .B(_05075_),
    .X(_05081_));
 sg13g2_a22oi_1 _19598_ (.Y(_05082_),
    .B1(_05078_),
    .B2(_05080_),
    .A2(_05074_),
    .A1(net6133));
 sg13g2_a221oi_1 _19599_ (.B2(net6221),
    .C1(_05072_),
    .B1(_05082_),
    .A1(net5457),
    .Y(_05083_),
    .A2(_05069_));
 sg13g2_nand2b_1 _19600_ (.Y(_05084_),
    .B(_05083_),
    .A_N(_05064_));
 sg13g2_a221oi_1 _19601_ (.B2(_05059_),
    .C1(_05084_),
    .B1(_05058_),
    .A1(net5774),
    .Y(_05085_),
    .A2(_05055_));
 sg13g2_a21oi_1 _19602_ (.A1(net6411),
    .A2(_08165_),
    .Y(_01353_),
    .B1(_05085_));
 sg13g2_a21oi_1 _19603_ (.A1(_04592_),
    .A2(_05056_),
    .Y(_05086_),
    .B1(_04590_));
 sg13g2_nand2_1 _19604_ (.Y(_05087_),
    .A(_04591_),
    .B(_05058_));
 sg13g2_nand2_1 _19605_ (.Y(_05088_),
    .A(_04631_),
    .B(_05086_));
 sg13g2_nand2_1 _19606_ (.Y(_05089_),
    .A(_04630_),
    .B(_05087_));
 sg13g2_nand3_1 _19607_ (.B(_05088_),
    .C(_05089_),
    .A(net5760),
    .Y(_05090_));
 sg13g2_a21oi_1 _19608_ (.A1(_04628_),
    .A2(_04630_),
    .Y(_05091_),
    .B1(net5771));
 sg13g2_nor2b_1 _19609_ (.A(_04764_),
    .B_N(_04778_),
    .Y(_05092_));
 sg13g2_nor2_1 _19610_ (.A(net6116),
    .B(_05047_),
    .Y(_05093_));
 sg13g2_a21oi_1 _19611_ (.A1(net6116),
    .A2(_05092_),
    .Y(_05094_),
    .B1(_05093_));
 sg13g2_mux2_1 _19612_ (.A0(_04988_),
    .A1(_05094_),
    .S(net6124),
    .X(_05095_));
 sg13g2_nor2_1 _19613_ (.A(net6127),
    .B(_04808_),
    .Y(_05096_));
 sg13g2_a22oi_1 _19614_ (.Y(_05097_),
    .B1(net5453),
    .B2(_04788_),
    .A2(_05095_),
    .A1(net5454));
 sg13g2_a21oi_1 _19615_ (.A1(net6223),
    .A2(_04746_),
    .Y(_05098_),
    .B1(_04551_));
 sg13g2_o21ai_1 _19616_ (.B1(_05098_),
    .Y(_05099_),
    .A1(net6223),
    .A2(_04772_));
 sg13g2_nand2_1 _19617_ (.Y(_05100_),
    .A(_05097_),
    .B(_05099_));
 sg13g2_a21o_1 _19618_ (.A2(_04753_),
    .A1(net6129),
    .B1(_05081_),
    .X(_05101_));
 sg13g2_nand3_1 _19619_ (.B(_04550_),
    .C(_05101_),
    .A(net6219),
    .Y(_05102_));
 sg13g2_nor2_1 _19620_ (.A(_04629_),
    .B(_04805_),
    .Y(_05103_));
 sg13g2_o21ai_1 _19621_ (.B1(_04796_),
    .Y(_05104_),
    .A1(\soc_inst.cpu_core.alu.b[8] ),
    .A2(net6284));
 sg13g2_a21oi_1 _19622_ (.A1(_04630_),
    .A2(net5765),
    .Y(_05105_),
    .B1(_05103_));
 sg13g2_nand4_1 _19623_ (.B(_05102_),
    .C(_05104_),
    .A(net6156),
    .Y(_05106_),
    .D(_05105_));
 sg13g2_a221oi_1 _19624_ (.B2(net6135),
    .C1(_05106_),
    .B1(_05100_),
    .A1(_04632_),
    .Y(_05107_),
    .A2(_05091_));
 sg13g2_a22oi_1 _19625_ (.Y(_01354_),
    .B1(_05090_),
    .B2(_05107_),
    .A2(_08166_),
    .A1(net6410));
 sg13g2_nand3_1 _19626_ (.B(_04629_),
    .C(_05089_),
    .A(_04585_),
    .Y(_05108_));
 sg13g2_nand3_1 _19627_ (.B(_04630_),
    .C(_05087_),
    .A(_04584_),
    .Y(_05109_));
 sg13g2_or2_1 _19628_ (.X(_05110_),
    .B(_04629_),
    .A(_04585_));
 sg13g2_nand4_1 _19629_ (.B(_05108_),
    .C(_05109_),
    .A(net5760),
    .Y(_05111_),
    .D(_05110_));
 sg13g2_nand3_1 _19630_ (.B(_04586_),
    .C(_04632_),
    .A(_04584_),
    .Y(_05112_));
 sg13g2_nand4_1 _19631_ (.B(_04587_),
    .C(_04633_),
    .A(net5774),
    .Y(_05113_),
    .D(_05112_));
 sg13g2_nor2_1 _19632_ (.A(net6132),
    .B(_04817_),
    .Y(_05114_));
 sg13g2_a21oi_1 _19633_ (.A1(net6128),
    .A2(_04872_),
    .Y(_05115_),
    .B1(_05114_));
 sg13g2_a21o_2 _19634_ (.A2(net6253),
    .A1(\soc_inst.cpu_core.alu.a[8] ),
    .B1(_04864_),
    .X(_05116_));
 sg13g2_mux2_1 _19635_ (.A0(_05065_),
    .A1(_05116_),
    .S(net6118),
    .X(_05117_));
 sg13g2_mux2_1 _19636_ (.A0(_05012_),
    .A1(_05117_),
    .S(net6123),
    .X(_05118_));
 sg13g2_nand2_1 _19637_ (.Y(_05119_),
    .A(net6128),
    .B(_05118_));
 sg13g2_o21ai_1 _19638_ (.B1(_05119_),
    .Y(_05120_),
    .A1(net6128),
    .A2(_04851_));
 sg13g2_nand2_1 _19639_ (.Y(_05121_),
    .A(net5456),
    .B(_05120_));
 sg13g2_o21ai_1 _19640_ (.B1(_04583_),
    .Y(_05122_),
    .A1(net6287),
    .A2(_04582_));
 sg13g2_a221oi_1 _19641_ (.B2(net5768),
    .C1(net6412),
    .B1(_05122_),
    .A1(_04584_),
    .Y(_05123_),
    .A2(net5765));
 sg13g2_nor3_2 _19642_ (.A(net6224),
    .B(net6285),
    .C(_04551_),
    .Y(_05124_));
 sg13g2_nand2_1 _19643_ (.Y(_05125_),
    .A(net6133),
    .B(_04831_));
 sg13g2_a21oi_1 _19644_ (.A1(_04836_),
    .A2(_05124_),
    .Y(_05126_),
    .B1(_05081_));
 sg13g2_o21ai_1 _19645_ (.B1(_05126_),
    .Y(_05127_),
    .A1(_04829_),
    .A2(_05077_));
 sg13g2_a22oi_1 _19646_ (.Y(_05128_),
    .B1(_05127_),
    .B2(net6220),
    .A2(_05115_),
    .A1(net5462));
 sg13g2_and4_1 _19647_ (.A(_05113_),
    .B(_05121_),
    .C(_05123_),
    .D(_05128_),
    .X(_05129_));
 sg13g2_a22oi_1 _19648_ (.Y(_01355_),
    .B1(_05111_),
    .B2(_05129_),
    .A2(_08167_),
    .A1(net6410));
 sg13g2_and2_1 _19649_ (.A(_04583_),
    .B(_05110_),
    .X(_05130_));
 sg13g2_nand2_1 _19650_ (.Y(_05131_),
    .A(_05109_),
    .B(_05130_));
 sg13g2_nand2_1 _19651_ (.Y(_05132_),
    .A(_04580_),
    .B(_05131_));
 sg13g2_o21ai_1 _19652_ (.B1(net5760),
    .Y(_05133_),
    .A1(_04580_),
    .A2(_05131_));
 sg13g2_nand2b_1 _19653_ (.Y(_05134_),
    .B(_05132_),
    .A_N(_05133_));
 sg13g2_or2_1 _19654_ (.X(_05135_),
    .B(_04634_),
    .A(_04580_));
 sg13g2_nand2_1 _19655_ (.Y(_05136_),
    .A(net5773),
    .B(_05135_));
 sg13g2_a21oi_1 _19656_ (.A1(_04580_),
    .A2(_04634_),
    .Y(_05137_),
    .B1(_05136_));
 sg13g2_o21ai_1 _19657_ (.B1(net5462),
    .Y(_05138_),
    .A1(net6223),
    .A2(_04906_));
 sg13g2_a21oi_1 _19658_ (.A1(net6223),
    .A2(_04890_),
    .Y(_05139_),
    .B1(_05138_));
 sg13g2_o21ai_1 _19659_ (.B1(_04766_),
    .Y(_05140_),
    .A1(_08204_),
    .A2(net6111));
 sg13g2_nor2_1 _19660_ (.A(net6240),
    .B(_05140_),
    .Y(_05141_));
 sg13g2_a21oi_1 _19661_ (.A1(net6242),
    .A2(_05092_),
    .Y(_05142_),
    .B1(_05141_));
 sg13g2_mux2_1 _19662_ (.A0(_05049_),
    .A1(_05142_),
    .S(net6124),
    .X(_05143_));
 sg13g2_nand2_1 _19663_ (.Y(_05144_),
    .A(net6224),
    .B(_04916_));
 sg13g2_o21ai_1 _19664_ (.B1(_05144_),
    .Y(_05145_),
    .A1(net6224),
    .A2(_05143_));
 sg13g2_o21ai_1 _19665_ (.B1(_04579_),
    .Y(_05146_),
    .A1(net6286),
    .A2(_04578_));
 sg13g2_a221oi_1 _19666_ (.B2(net5768),
    .C1(net6410),
    .B1(_05146_),
    .A1(_04580_),
    .Y(_05147_),
    .A2(net5764));
 sg13g2_o21ai_1 _19667_ (.B1(_05147_),
    .Y(_05148_),
    .A1(_04810_),
    .A2(_05145_));
 sg13g2_o21ai_1 _19668_ (.B1(_05077_),
    .Y(_05149_),
    .A1(_04896_),
    .A2(_05125_));
 sg13g2_a21oi_2 _19669_ (.B1(_05081_),
    .Y(_05150_),
    .A2(_05149_),
    .A1(_04898_));
 sg13g2_nor2_1 _19670_ (.A(net6135),
    .B(_05150_),
    .Y(_05151_));
 sg13g2_nor4_1 _19671_ (.A(_05137_),
    .B(_05139_),
    .C(_05148_),
    .D(_05151_),
    .Y(_05152_));
 sg13g2_a22oi_1 _19672_ (.Y(_01356_),
    .B1(_05134_),
    .B2(_05152_),
    .A2(_08168_),
    .A1(net6426));
 sg13g2_nand2_1 _19673_ (.Y(_05153_),
    .A(_04579_),
    .B(_05132_));
 sg13g2_xor2_1 _19674_ (.B(_05153_),
    .A(_04575_),
    .X(_05154_));
 sg13g2_nand3_1 _19675_ (.B(_04576_),
    .C(_05135_),
    .A(_04575_),
    .Y(_05155_));
 sg13g2_a21o_1 _19676_ (.A2(_05135_),
    .A1(_04576_),
    .B1(_04575_),
    .X(_05156_));
 sg13g2_nand3_1 _19677_ (.B(_05155_),
    .C(_05156_),
    .A(net5773),
    .Y(_05157_));
 sg13g2_nor2_1 _19678_ (.A(net6223),
    .B(_04948_),
    .Y(_05158_));
 sg13g2_o21ai_1 _19679_ (.B1(_04773_),
    .Y(_05159_),
    .A1(net6130),
    .A2(_04930_));
 sg13g2_o21ai_1 _19680_ (.B1(_04867_),
    .Y(_05160_),
    .A1(_08203_),
    .A2(net6111));
 sg13g2_mux2_1 _19681_ (.A0(_05116_),
    .A1(_05160_),
    .S(net6117),
    .X(_05161_));
 sg13g2_mux2_1 _19682_ (.A0(_05067_),
    .A1(_05161_),
    .S(net6125),
    .X(_05162_));
 sg13g2_nor2_1 _19683_ (.A(net6231),
    .B(_05162_),
    .Y(_05163_));
 sg13g2_a21oi_2 _19684_ (.B1(_05163_),
    .Y(_05164_),
    .A2(_04960_),
    .A1(net6230));
 sg13g2_nand3_1 _19685_ (.B(\soc_inst.cpu_core.alu.a[11] ),
    .C(net5459),
    .A(\soc_inst.cpu_core.alu.b[11] ),
    .Y(_05165_));
 sg13g2_a221oi_1 _19686_ (.B2(_04575_),
    .C1(net6412),
    .B1(net5765),
    .A1(_04574_),
    .Y(_05166_),
    .A2(net5461));
 sg13g2_nand2_1 _19687_ (.Y(_05167_),
    .A(_05165_),
    .B(_05166_));
 sg13g2_a21oi_1 _19688_ (.A1(net5456),
    .A2(_05164_),
    .Y(_05168_),
    .B1(_05167_));
 sg13g2_o21ai_1 _19689_ (.B1(_05168_),
    .Y(_05169_),
    .A1(_05158_),
    .A2(_05159_));
 sg13g2_a21oi_1 _19690_ (.A1(_04935_),
    .A2(_05124_),
    .Y(_05170_),
    .B1(_05081_));
 sg13g2_o21ai_1 _19691_ (.B1(_05170_),
    .Y(_05171_),
    .A1(_04938_),
    .A2(_05077_));
 sg13g2_a221oi_1 _19692_ (.B2(net6219),
    .C1(_05169_),
    .B1(_05171_),
    .A1(net5760),
    .Y(_05172_),
    .A2(_05154_));
 sg13g2_a22oi_1 _19693_ (.Y(_01357_),
    .B1(_05157_),
    .B2(_05172_),
    .A2(_08169_),
    .A1(net6426));
 sg13g2_nor2b_1 _19694_ (.A(_04579_),
    .B_N(_04574_),
    .Y(_05173_));
 sg13g2_a21oi_1 _19695_ (.A1(\soc_inst.cpu_core.alu.b[11] ),
    .A2(\soc_inst.cpu_core.alu.a[11] ),
    .Y(_05174_),
    .B1(_05173_));
 sg13g2_nand2_1 _19696_ (.Y(_05175_),
    .A(_04575_),
    .B(_04580_));
 sg13g2_nor4_1 _19697_ (.A(_04585_),
    .B(_04631_),
    .C(_05086_),
    .D(_05175_),
    .Y(_05176_));
 sg13g2_o21ai_1 _19698_ (.B1(_05174_),
    .Y(_05177_),
    .A1(_05130_),
    .A2(_05175_));
 sg13g2_nor2_1 _19699_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sg13g2_or2_1 _19700_ (.X(_05179_),
    .B(_05178_),
    .A(_04641_));
 sg13g2_a21oi_1 _19701_ (.A1(_04641_),
    .A2(_05178_),
    .Y(_05180_),
    .B1(net5757));
 sg13g2_o21ai_1 _19702_ (.B1(_04767_),
    .Y(_05181_),
    .A1(_08201_),
    .A2(net6249));
 sg13g2_mux2_1 _19703_ (.A0(_05140_),
    .A1(_05181_),
    .S(net6115),
    .X(_05182_));
 sg13g2_mux2_1 _19704_ (.A0(_05094_),
    .A1(_05182_),
    .S(net6122),
    .X(_05183_));
 sg13g2_nand2_1 _19705_ (.Y(_05184_),
    .A(net6127),
    .B(_05183_));
 sg13g2_o21ai_1 _19706_ (.B1(_05184_),
    .Y(_05185_),
    .A1(net6127),
    .A2(_04989_));
 sg13g2_nor2_1 _19707_ (.A(_04640_),
    .B(_04805_),
    .Y(_05186_));
 sg13g2_nor2_1 _19708_ (.A(_04641_),
    .B(net5762),
    .Y(_05187_));
 sg13g2_o21ai_1 _19709_ (.B1(net6149),
    .Y(_05188_),
    .A1(_04639_),
    .A2(_04797_));
 sg13g2_nor2_1 _19710_ (.A(net6223),
    .B(_04980_),
    .Y(_05189_));
 sg13g2_o21ai_1 _19711_ (.B1(_04773_),
    .Y(_05190_),
    .A1(net6130),
    .A2(_04972_));
 sg13g2_nor2_1 _19712_ (.A(_05189_),
    .B(_05190_),
    .Y(_05191_));
 sg13g2_a221oi_1 _19713_ (.B2(_04974_),
    .C1(_05081_),
    .B1(_05124_),
    .A1(_04976_),
    .Y(_05192_),
    .A2(_05076_));
 sg13g2_nor4_1 _19714_ (.A(_05186_),
    .B(_05187_),
    .C(_05188_),
    .D(_05191_),
    .Y(_05193_));
 sg13g2_o21ai_1 _19715_ (.B1(_05193_),
    .Y(_05194_),
    .A1(net6135),
    .A2(_05192_));
 sg13g2_a21oi_1 _19716_ (.A1(net5456),
    .A2(_05185_),
    .Y(_05195_),
    .B1(_05194_));
 sg13g2_o21ai_1 _19717_ (.B1(net5772),
    .Y(_05196_),
    .A1(_04638_),
    .A2(_04641_));
 sg13g2_nor2_1 _19718_ (.A(_04642_),
    .B(_05196_),
    .Y(_05197_));
 sg13g2_a21oi_1 _19719_ (.A1(_05179_),
    .A2(_05180_),
    .Y(_05198_),
    .B1(_05197_));
 sg13g2_a22oi_1 _19720_ (.Y(_01358_),
    .B1(_05195_),
    .B2(_05198_),
    .A2(_08170_),
    .A1(net6395));
 sg13g2_nand3_1 _19721_ (.B(_04640_),
    .C(_05179_),
    .A(_04572_),
    .Y(_05199_));
 sg13g2_nor2_1 _19722_ (.A(_04572_),
    .B(_04641_),
    .Y(_05200_));
 sg13g2_o21ai_1 _19723_ (.B1(_05200_),
    .Y(_05201_),
    .A1(_05176_),
    .A2(_05177_));
 sg13g2_o21ai_1 _19724_ (.B1(_05201_),
    .Y(_05202_),
    .A1(_04572_),
    .A2(_04640_));
 sg13g2_nor2_1 _19725_ (.A(net5757),
    .B(_05202_),
    .Y(_05203_));
 sg13g2_nor2_1 _19726_ (.A(_04572_),
    .B(_04642_),
    .Y(_05204_));
 sg13g2_o21ai_1 _19727_ (.B1(_05204_),
    .Y(_05205_),
    .A1(net3040),
    .A2(_08201_));
 sg13g2_nor2_1 _19728_ (.A(net5770),
    .B(_04644_),
    .Y(_05206_));
 sg13g2_nand3_1 _19729_ (.B(_05205_),
    .C(_05206_),
    .A(_04643_),
    .Y(_05207_));
 sg13g2_o21ai_1 _19730_ (.B1(_04570_),
    .Y(_05208_),
    .A1(net6286),
    .A2(_04569_));
 sg13g2_a22oi_1 _19731_ (.Y(_05209_),
    .B1(_05208_),
    .B2(net5766),
    .A2(net5763),
    .A1(_04571_));
 sg13g2_a221oi_1 _19732_ (.B2(_05002_),
    .C1(_05081_),
    .B1(_05124_),
    .A1(_05005_),
    .Y(_05210_),
    .A2(_05076_));
 sg13g2_nand2b_1 _19733_ (.Y(_05211_),
    .B(net6218),
    .A_N(_05210_));
 sg13g2_nor2_1 _19734_ (.A(net6131),
    .B(_05000_),
    .Y(_05212_));
 sg13g2_a21oi_1 _19735_ (.A1(net6128),
    .A2(_05021_),
    .Y(_05213_),
    .B1(_05212_));
 sg13g2_nand2b_2 _19736_ (.Y(_05214_),
    .B(_04866_),
    .A_N(_04858_));
 sg13g2_mux2_1 _19737_ (.A0(_05160_),
    .A1(_05214_),
    .S(net6117),
    .X(_05215_));
 sg13g2_mux2_1 _19738_ (.A0(_05117_),
    .A1(_05215_),
    .S(net6125),
    .X(_05216_));
 sg13g2_nand2_1 _19739_ (.Y(_05217_),
    .A(net6128),
    .B(_05216_));
 sg13g2_o21ai_1 _19740_ (.B1(_05217_),
    .Y(_05218_),
    .A1(net6128),
    .A2(_05013_));
 sg13g2_a22oi_1 _19741_ (.Y(_05219_),
    .B1(_05218_),
    .B2(net5456),
    .A2(_05213_),
    .A1(net5462));
 sg13g2_nand4_1 _19742_ (.B(_05209_),
    .C(_05211_),
    .A(net6149),
    .Y(_05220_),
    .D(_05219_));
 sg13g2_a21oi_1 _19743_ (.A1(_05199_),
    .A2(_05203_),
    .Y(_05221_),
    .B1(_05220_));
 sg13g2_a22oi_1 _19744_ (.Y(_01359_),
    .B1(net3291),
    .B2(_05221_),
    .A2(_08171_),
    .A1(net6395));
 sg13g2_nand3_1 _19745_ (.B(_04643_),
    .C(_04645_),
    .A(_04566_),
    .Y(_05222_));
 sg13g2_a21o_1 _19746_ (.A2(_04645_),
    .A1(_04643_),
    .B1(_04566_),
    .X(_05223_));
 sg13g2_nand3_1 _19747_ (.B(_05222_),
    .C(_05223_),
    .A(net5772),
    .Y(_05224_));
 sg13g2_o21ai_1 _19748_ (.B1(_04570_),
    .Y(_05225_),
    .A1(_04569_),
    .A2(_04640_));
 sg13g2_nor2b_1 _19749_ (.A(_05225_),
    .B_N(_05201_),
    .Y(_05226_));
 sg13g2_nor2b_1 _19750_ (.A(_05226_),
    .B_N(_04566_),
    .Y(_05227_));
 sg13g2_xnor2_1 _19751_ (.Y(_05228_),
    .A(_04566_),
    .B(_05226_));
 sg13g2_o21ai_1 _19752_ (.B1(_04773_),
    .Y(_05229_),
    .A1(net6130),
    .A2(_05029_));
 sg13g2_a21oi_1 _19753_ (.A1(net6129),
    .A2(_05041_),
    .Y(_05230_),
    .B1(_05229_));
 sg13g2_o21ai_1 _19754_ (.B1(_04564_),
    .Y(_05231_),
    .A1(net6286),
    .A2(_04565_));
 sg13g2_a221oi_1 _19755_ (.B2(net5766),
    .C1(net6395),
    .B1(_05231_),
    .A1(_04566_),
    .Y(_05232_),
    .A2(net5763));
 sg13g2_a21oi_1 _19756_ (.A1(net6130),
    .A2(_05034_),
    .Y(_05233_),
    .B1(_05078_));
 sg13g2_a21o_1 _19757_ (.A2(_05124_),
    .A1(_05031_),
    .B1(_05233_),
    .X(_05234_));
 sg13g2_a21oi_1 _19758_ (.A1(net6219),
    .A2(_05234_),
    .Y(_05235_),
    .B1(_05230_));
 sg13g2_and2_1 _19759_ (.A(_05232_),
    .B(_05235_),
    .X(_05236_));
 sg13g2_o21ai_1 _19760_ (.B1(_04759_),
    .Y(_05237_),
    .A1(_08200_),
    .A2(net6111));
 sg13g2_mux2_1 _19761_ (.A0(_05181_),
    .A1(_05237_),
    .S(net6115),
    .X(_05238_));
 sg13g2_mux2_1 _19762_ (.A0(_05142_),
    .A1(_05238_),
    .S(net6122),
    .X(_05239_));
 sg13g2_nand2_1 _19763_ (.Y(_05240_),
    .A(net6227),
    .B(_05050_));
 sg13g2_o21ai_1 _19764_ (.B1(_05240_),
    .Y(_05241_),
    .A1(net6224),
    .A2(_05239_));
 sg13g2_o21ai_1 _19765_ (.B1(_05236_),
    .Y(_05242_),
    .A1(_04810_),
    .A2(_05241_));
 sg13g2_a21oi_1 _19766_ (.A1(net5759),
    .A2(_05228_),
    .Y(_05243_),
    .B1(_05242_));
 sg13g2_a22oi_1 _19767_ (.Y(_01360_),
    .B1(_05224_),
    .B2(_05243_),
    .A2(_08172_),
    .A1(net6394));
 sg13g2_nand2_1 _19768_ (.Y(_05244_),
    .A(_04568_),
    .B(_05223_));
 sg13g2_xnor2_1 _19769_ (.Y(_05245_),
    .A(_04562_),
    .B(_05244_));
 sg13g2_nor2_1 _19770_ (.A(_04563_),
    .B(_05227_),
    .Y(_05246_));
 sg13g2_xnor2_1 _19771_ (.Y(_05247_),
    .A(_04562_),
    .B(_05246_));
 sg13g2_a21oi_1 _19772_ (.A1(net6224),
    .A2(_05074_),
    .Y(_05248_),
    .B1(_04774_));
 sg13g2_o21ai_1 _19773_ (.B1(_05248_),
    .Y(_05249_),
    .A1(net6223),
    .A2(_05062_));
 sg13g2_nand2_1 _19774_ (.Y(_05250_),
    .A(net6286),
    .B(_04561_));
 sg13g2_a22oi_1 _19775_ (.Y(_05251_),
    .B1(_05250_),
    .B2(net5766),
    .A2(net5763),
    .A1(_04561_));
 sg13g2_nor3_1 _19776_ (.A(_04786_),
    .B(_04832_),
    .C(_05125_),
    .Y(_05252_));
 sg13g2_nand2_1 _19777_ (.Y(_05253_),
    .A(net6219),
    .B(_05252_));
 sg13g2_and2_1 _19778_ (.A(net6218),
    .B(_05075_),
    .X(_05254_));
 sg13g2_nand2_2 _19779_ (.Y(_05255_),
    .A(net6220),
    .B(_05075_));
 sg13g2_o21ai_1 _19780_ (.B1(net6149),
    .Y(_05256_),
    .A1(_04560_),
    .A2(_05251_));
 sg13g2_nor2_1 _19781_ (.A(net5094),
    .B(_05256_),
    .Y(_05257_));
 sg13g2_o21ai_1 _19782_ (.B1(_04861_),
    .Y(_05258_),
    .A1(_08198_),
    .A2(net6112));
 sg13g2_mux2_1 _19783_ (.A0(_05214_),
    .A1(_05258_),
    .S(net6119),
    .X(_05259_));
 sg13g2_mux2_1 _19784_ (.A0(_05161_),
    .A1(_05259_),
    .S(net6126),
    .X(_05260_));
 sg13g2_mux2_1 _19785_ (.A0(_05068_),
    .A1(_05260_),
    .S(net6128),
    .X(_05261_));
 sg13g2_a22oi_1 _19786_ (.Y(_05262_),
    .B1(_05261_),
    .B2(net5456),
    .A2(_05245_),
    .A1(net5773));
 sg13g2_nand4_1 _19787_ (.B(_05253_),
    .C(_05257_),
    .A(_05249_),
    .Y(_05263_),
    .D(_05262_));
 sg13g2_a21oi_1 _19788_ (.A1(net5759),
    .A2(_05247_),
    .Y(_05264_),
    .B1(_05263_));
 sg13g2_a21oi_1 _19789_ (.A1(net6355),
    .A2(_08174_),
    .Y(_01361_),
    .B1(_05264_));
 sg13g2_xnor2_1 _19790_ (.Y(_05265_),
    .A(_04650_),
    .B(_04656_));
 sg13g2_o21ai_1 _19791_ (.B1(_04561_),
    .Y(_05266_),
    .A1(_04560_),
    .A2(_04564_));
 sg13g2_inv_1 _19792_ (.Y(_05267_),
    .A(_05266_));
 sg13g2_nor2_1 _19793_ (.A(_05225_),
    .B(_05266_),
    .Y(_05268_));
 sg13g2_nand2_1 _19794_ (.Y(_05269_),
    .A(_05201_),
    .B(_05268_));
 sg13g2_nand2_1 _19795_ (.Y(_05270_),
    .A(_04562_),
    .B(_04566_));
 sg13g2_nand2_1 _19796_ (.Y(_05271_),
    .A(_05267_),
    .B(_05270_));
 sg13g2_nand3_1 _19797_ (.B(_05269_),
    .C(_05271_),
    .A(_04656_),
    .Y(_05272_));
 sg13g2_a21oi_1 _19798_ (.A1(_05269_),
    .A2(_05271_),
    .Y(_05273_),
    .B1(_04656_));
 sg13g2_nor2_1 _19799_ (.A(net5757),
    .B(_05273_),
    .Y(_05274_));
 sg13g2_or2_1 _19800_ (.X(_05275_),
    .B(_05075_),
    .A(net5462));
 sg13g2_o21ai_1 _19801_ (.B1(_05275_),
    .Y(_05276_),
    .A1(net6218),
    .A2(_04755_));
 sg13g2_o21ai_1 _19802_ (.B1(_04760_),
    .Y(_05277_),
    .A1(_08196_),
    .A2(net6250));
 sg13g2_mux2_1 _19803_ (.A0(_05237_),
    .A1(_05277_),
    .S(net6115),
    .X(_05278_));
 sg13g2_mux2_1 _19804_ (.A0(_05182_),
    .A1(_05278_),
    .S(net6122),
    .X(_05279_));
 sg13g2_inv_1 _19805_ (.Y(_05280_),
    .A(_05279_));
 sg13g2_a21oi_1 _19806_ (.A1(net6129),
    .A2(_05280_),
    .Y(_05281_),
    .B1(_04810_));
 sg13g2_o21ai_1 _19807_ (.B1(_05281_),
    .Y(_05282_),
    .A1(net6129),
    .A2(_05095_));
 sg13g2_nor2_2 _19808_ (.A(net6135),
    .B(_04808_),
    .Y(_05283_));
 sg13g2_nand2_2 _19809_ (.Y(_05284_),
    .A(net6218),
    .B(_04807_));
 sg13g2_o21ai_1 _19810_ (.B1(net5766),
    .Y(_05285_),
    .A1(\soc_inst.cpu_core.alu.b[16] ),
    .A2(net6281));
 sg13g2_a21oi_1 _19811_ (.A1(net6288),
    .A2(_04655_),
    .Y(_05286_),
    .B1(_05285_));
 sg13g2_a221oi_1 _19812_ (.B2(_04806_),
    .C1(_05286_),
    .B1(net5452),
    .A1(_04656_),
    .Y(_05287_),
    .A2(net5763));
 sg13g2_nand3_1 _19813_ (.B(_05282_),
    .C(_05287_),
    .A(_05276_),
    .Y(_05288_));
 sg13g2_a221oi_1 _19814_ (.B2(_05274_),
    .C1(_05288_),
    .B1(_05272_),
    .A1(net5772),
    .Y(_05289_),
    .A2(_05265_));
 sg13g2_nand2_1 _19815_ (.Y(_05290_),
    .A(net6396),
    .B(net2299));
 sg13g2_o21ai_1 _19816_ (.B1(_05290_),
    .Y(_01362_),
    .A1(net5241),
    .A2(_05289_));
 sg13g2_nand2_1 _19817_ (.Y(_05291_),
    .A(net6394),
    .B(net3152));
 sg13g2_nand2_1 _19818_ (.Y(_05292_),
    .A(_04655_),
    .B(_05272_));
 sg13g2_xnor2_1 _19819_ (.Y(_05293_),
    .A(_04654_),
    .B(_05292_));
 sg13g2_a21oi_1 _19820_ (.A1(_04650_),
    .A2(_04657_),
    .Y(_05294_),
    .B1(_04654_));
 sg13g2_o21ai_1 _19821_ (.B1(_05294_),
    .Y(_05295_),
    .A1(\soc_inst.cpu_core.alu.b[16] ),
    .A2(_08196_));
 sg13g2_nand4_1 _19822_ (.B(_04659_),
    .C(_04687_),
    .A(net5772),
    .Y(_05296_),
    .D(_05295_));
 sg13g2_o21ai_1 _19823_ (.B1(_04860_),
    .Y(_05297_),
    .A1(_08195_),
    .A2(net6250));
 sg13g2_mux2_1 _19824_ (.A0(_05258_),
    .A1(_05297_),
    .S(net6119),
    .X(_05298_));
 sg13g2_mux2_1 _19825_ (.A0(_05215_),
    .A1(_05298_),
    .S(net6125),
    .X(_05299_));
 sg13g2_a22oi_1 _19826_ (.Y(_05300_),
    .B1(_05299_),
    .B2(net5454),
    .A2(_05118_),
    .A1(net5453));
 sg13g2_a21oi_1 _19827_ (.A1(_04838_),
    .A2(_05300_),
    .Y(_05301_),
    .B1(net6221));
 sg13g2_a22oi_1 _19828_ (.Y(_05302_),
    .B1(net5458),
    .B2(_04652_),
    .A2(net5460),
    .A1(_04651_));
 sg13g2_a21oi_1 _19829_ (.A1(_04653_),
    .A2(net5764),
    .Y(_05303_),
    .B1(net5094));
 sg13g2_a21oi_2 _19830_ (.B1(_05301_),
    .Y(_05304_),
    .A2(_04852_),
    .A1(net6221));
 sg13g2_nand4_1 _19831_ (.B(_05302_),
    .C(_05303_),
    .A(_05296_),
    .Y(_05305_),
    .D(_05304_));
 sg13g2_a21oi_1 _19832_ (.A1(net5759),
    .A2(_05293_),
    .Y(_05306_),
    .B1(_05305_));
 sg13g2_o21ai_1 _19833_ (.B1(_05291_),
    .Y(_01363_),
    .A1(net5241),
    .A2(_05306_));
 sg13g2_a21oi_1 _19834_ (.A1(_04650_),
    .A2(_04658_),
    .Y(_05307_),
    .B1(_04688_));
 sg13g2_or2_1 _19835_ (.X(_05308_),
    .B(_05307_),
    .A(_04681_));
 sg13g2_a21oi_1 _19836_ (.A1(_04681_),
    .A2(_05307_),
    .Y(_05309_),
    .B1(net5770));
 sg13g2_nor2_1 _19837_ (.A(_04654_),
    .B(_05272_),
    .Y(_05310_));
 sg13g2_nand2b_1 _19838_ (.Y(_05311_),
    .B(_04651_),
    .A_N(_04655_));
 sg13g2_nand2b_1 _19839_ (.Y(_05312_),
    .B(_05311_),
    .A_N(_04652_));
 sg13g2_o21ai_1 _19840_ (.B1(_04681_),
    .Y(_05313_),
    .A1(_05310_),
    .A2(_05312_));
 sg13g2_nor3_1 _19841_ (.A(_04681_),
    .B(_05310_),
    .C(_05312_),
    .Y(_05314_));
 sg13g2_nand2_1 _19842_ (.Y(_05315_),
    .A(net5759),
    .B(_05313_));
 sg13g2_mux2_1 _19843_ (.A0(\soc_inst.cpu_core.alu.a[18] ),
    .A1(net6280),
    .S(net6256),
    .X(_05316_));
 sg13g2_mux2_1 _19844_ (.A0(_05277_),
    .A1(_05316_),
    .S(net6113),
    .X(_05317_));
 sg13g2_mux2_1 _19845_ (.A0(_05238_),
    .A1(_05317_),
    .S(net6121),
    .X(_05318_));
 sg13g2_a22oi_1 _19846_ (.Y(_05319_),
    .B1(_05318_),
    .B2(net5454),
    .A2(_05143_),
    .A1(net5453));
 sg13g2_a21oi_1 _19847_ (.A1(_04901_),
    .A2(_05319_),
    .Y(_05320_),
    .B1(net6219));
 sg13g2_nor3_1 _19848_ (.A(net6224),
    .B(_04916_),
    .C(_05284_),
    .Y(_05321_));
 sg13g2_nand2_1 _19849_ (.Y(_05322_),
    .A(_04678_),
    .B(net5460));
 sg13g2_a22oi_1 _19850_ (.Y(_05323_),
    .B1(net5764),
    .B2(_04681_),
    .A2(net5458),
    .A1(_04679_));
 sg13g2_nand2_1 _19851_ (.Y(_05324_),
    .A(_05322_),
    .B(_05323_));
 sg13g2_nor4_1 _19852_ (.A(net5094),
    .B(_05320_),
    .C(_05321_),
    .D(_05324_),
    .Y(_05325_));
 sg13g2_o21ai_1 _19853_ (.B1(_05325_),
    .Y(_05326_),
    .A1(_05314_),
    .A2(_05315_));
 sg13g2_a21oi_1 _19854_ (.A1(_05308_),
    .A2(_05309_),
    .Y(_05327_),
    .B1(_05326_));
 sg13g2_nand2_1 _19855_ (.Y(_05328_),
    .A(net6389),
    .B(net3033));
 sg13g2_o21ai_1 _19856_ (.B1(_05328_),
    .Y(_01364_),
    .A1(net5242),
    .A2(_05327_));
 sg13g2_a21oi_1 _19857_ (.A1(_04680_),
    .A2(_05313_),
    .Y(_05329_),
    .B1(_04677_));
 sg13g2_nand3_1 _19858_ (.B(_04680_),
    .C(_05313_),
    .A(_04677_),
    .Y(_05330_));
 sg13g2_nand2_1 _19859_ (.Y(_05331_),
    .A(net5759),
    .B(_05330_));
 sg13g2_nand3_1 _19860_ (.B(_04690_),
    .C(_05308_),
    .A(_04676_),
    .Y(_05332_));
 sg13g2_a21oi_1 _19861_ (.A1(_04690_),
    .A2(_05308_),
    .Y(_05333_),
    .B1(_04676_));
 sg13g2_nor2_1 _19862_ (.A(net5770),
    .B(_05333_),
    .Y(_05334_));
 sg13g2_mux2_1 _19863_ (.A0(net6277),
    .A1(\soc_inst.cpu_core.alu.a[18] ),
    .S(net6259),
    .X(_05335_));
 sg13g2_mux2_1 _19864_ (.A0(_05297_),
    .A1(_05335_),
    .S(net6119),
    .X(_05336_));
 sg13g2_mux2_1 _19865_ (.A0(_05259_),
    .A1(_05336_),
    .S(net6126),
    .X(_05337_));
 sg13g2_a22oi_1 _19866_ (.Y(_05338_),
    .B1(_05337_),
    .B2(net5454),
    .A2(_05162_),
    .A1(net5453));
 sg13g2_a21oi_1 _19867_ (.A1(_04940_),
    .A2(_05338_),
    .Y(_05339_),
    .B1(net6221));
 sg13g2_nor3_1 _19868_ (.A(net6224),
    .B(_04960_),
    .C(_05284_),
    .Y(_05340_));
 sg13g2_a22oi_1 _19869_ (.Y(_05341_),
    .B1(net5458),
    .B2(_04675_),
    .A2(net5460),
    .A1(_04674_));
 sg13g2_o21ai_1 _19870_ (.B1(_05341_),
    .Y(_05342_),
    .A1(_04677_),
    .A2(net5761));
 sg13g2_nor4_1 _19871_ (.A(_05254_),
    .B(_05339_),
    .C(_05340_),
    .D(_05342_),
    .Y(_05343_));
 sg13g2_o21ai_1 _19872_ (.B1(_05343_),
    .Y(_05344_),
    .A1(_05329_),
    .A2(_05331_));
 sg13g2_a21oi_1 _19873_ (.A1(_05332_),
    .A2(_05334_),
    .Y(_05345_),
    .B1(_05344_));
 sg13g2_nand2_1 _19874_ (.Y(_05346_),
    .A(net6396),
    .B(net3244));
 sg13g2_o21ai_1 _19875_ (.B1(_05346_),
    .Y(_01365_),
    .A1(net5241),
    .A2(_05345_));
 sg13g2_nand3_1 _19876_ (.B(_04658_),
    .C(_04682_),
    .A(_04650_),
    .Y(_05347_));
 sg13g2_nand3_1 _19877_ (.B(_04692_),
    .C(_05347_),
    .A(_04668_),
    .Y(_05348_));
 sg13g2_a21oi_1 _19878_ (.A1(_04692_),
    .A2(_05347_),
    .Y(_05349_),
    .B1(_04668_));
 sg13g2_nor2_1 _19879_ (.A(net5770),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_and2_1 _19880_ (.A(_04676_),
    .B(_04681_),
    .X(_05351_));
 sg13g2_nand3_1 _19881_ (.B(_04656_),
    .C(_05351_),
    .A(_04653_),
    .Y(_05352_));
 sg13g2_a221oi_1 _19882_ (.B2(_05267_),
    .C1(_05352_),
    .B1(_05270_),
    .A1(_05201_),
    .Y(_05353_),
    .A2(_05268_));
 sg13g2_a21oi_1 _19883_ (.A1(_04674_),
    .A2(_04679_),
    .Y(_05354_),
    .B1(_04675_));
 sg13g2_nand2_1 _19884_ (.Y(_05355_),
    .A(_05312_),
    .B(_05351_));
 sg13g2_nand2_1 _19885_ (.Y(_05356_),
    .A(_05354_),
    .B(_05355_));
 sg13g2_or2_1 _19886_ (.X(_05357_),
    .B(_05356_),
    .A(_05353_));
 sg13g2_and2_1 _19887_ (.A(_04668_),
    .B(_05357_),
    .X(_05358_));
 sg13g2_xnor2_1 _19888_ (.Y(_05359_),
    .A(_04669_),
    .B(_05357_));
 sg13g2_mux2_1 _19889_ (.A0(net6275),
    .A1(net6277),
    .S(net6257),
    .X(_05360_));
 sg13g2_mux2_1 _19890_ (.A0(_05316_),
    .A1(_05360_),
    .S(net6113),
    .X(_05361_));
 sg13g2_and2_1 _19891_ (.A(net6121),
    .B(_05361_),
    .X(_05362_));
 sg13g2_a21oi_1 _19892_ (.A1(net6233),
    .A2(_05278_),
    .Y(_05363_),
    .B1(_05362_));
 sg13g2_inv_1 _19893_ (.Y(_05364_),
    .A(_05363_));
 sg13g2_a22oi_1 _19894_ (.Y(_05365_),
    .B1(_05364_),
    .B2(net5454),
    .A2(_05183_),
    .A1(net5453));
 sg13g2_a21oi_1 _19895_ (.A1(_04978_),
    .A2(_05365_),
    .Y(_05366_),
    .B1(net6220));
 sg13g2_nor2_1 _19896_ (.A(_04990_),
    .B(_05284_),
    .Y(_05367_));
 sg13g2_o21ai_1 _19897_ (.B1(net5460),
    .Y(_05368_),
    .A1(\soc_inst.cpu_core.alu.b[20] ),
    .A2(net6274));
 sg13g2_o21ai_1 _19898_ (.B1(_05368_),
    .Y(_05369_),
    .A1(_04667_),
    .A2(_04805_));
 sg13g2_nor4_1 _19899_ (.A(net5094),
    .B(_05366_),
    .C(_05367_),
    .D(_05369_),
    .Y(_05370_));
 sg13g2_o21ai_1 _19900_ (.B1(_05370_),
    .Y(_05371_),
    .A1(_04669_),
    .A2(net5761));
 sg13g2_a221oi_1 _19901_ (.B2(net5759),
    .C1(_05371_),
    .B1(_05359_),
    .A1(_05348_),
    .Y(_05372_),
    .A2(_05350_));
 sg13g2_nand2_1 _19902_ (.Y(_05373_),
    .A(net6388),
    .B(net3001));
 sg13g2_o21ai_1 _19903_ (.B1(_05373_),
    .Y(_01366_),
    .A1(net5242),
    .A2(_05372_));
 sg13g2_nand2_1 _19904_ (.Y(_05374_),
    .A(net6390),
    .B(net2879));
 sg13g2_nor3_1 _19905_ (.A(_04662_),
    .B(_04694_),
    .C(_05349_),
    .Y(_05375_));
 sg13g2_o21ai_1 _19906_ (.B1(_04662_),
    .Y(_05376_),
    .A1(_04694_),
    .A2(_05349_));
 sg13g2_nor2_1 _19907_ (.A(net5770),
    .B(_05375_),
    .Y(_05377_));
 sg13g2_nand2_1 _19908_ (.Y(_05378_),
    .A(_04662_),
    .B(_04667_));
 sg13g2_nor2_1 _19909_ (.A(_05358_),
    .B(_05378_),
    .Y(_05379_));
 sg13g2_nand2_1 _19910_ (.Y(_05380_),
    .A(_04661_),
    .B(_05358_));
 sg13g2_nor2_1 _19911_ (.A(_04662_),
    .B(_04667_),
    .Y(_05381_));
 sg13g2_nor3_1 _19912_ (.A(net5757),
    .B(_05379_),
    .C(_05381_),
    .Y(_05382_));
 sg13g2_mux2_1 _19913_ (.A0(net6273),
    .A1(net6275),
    .S(net6258),
    .X(_05383_));
 sg13g2_mux2_1 _19914_ (.A0(_05335_),
    .A1(_05383_),
    .S(net6114),
    .X(_05384_));
 sg13g2_mux2_1 _19915_ (.A0(_05298_),
    .A1(_05384_),
    .S(net6125),
    .X(_05385_));
 sg13g2_a22oi_1 _19916_ (.Y(_05386_),
    .B1(_05385_),
    .B2(net5454),
    .A2(_05216_),
    .A1(net5453));
 sg13g2_a21o_1 _19917_ (.A2(_05386_),
    .A1(_05008_),
    .B1(net6221),
    .X(_05387_));
 sg13g2_o21ai_1 _19918_ (.B1(net5767),
    .Y(_05388_),
    .A1(\soc_inst.cpu_core.alu.b[21] ),
    .A2(net6272));
 sg13g2_a21oi_1 _19919_ (.A1(net6287),
    .A2(_04660_),
    .Y(_05389_),
    .B1(_05388_));
 sg13g2_a221oi_1 _19920_ (.B2(net5452),
    .C1(_05389_),
    .B1(_05014_),
    .A1(_04661_),
    .Y(_05390_),
    .A2(net5763));
 sg13g2_nand3_1 _19921_ (.B(_05387_),
    .C(_05390_),
    .A(_05255_),
    .Y(_05391_));
 sg13g2_a221oi_1 _19922_ (.B2(_05382_),
    .C1(_05391_),
    .B1(_05380_),
    .A1(_05376_),
    .Y(_05392_),
    .A2(_05377_));
 sg13g2_o21ai_1 _19923_ (.B1(_05374_),
    .Y(_01367_),
    .A1(net5242),
    .A2(_05392_));
 sg13g2_nand2_1 _19924_ (.Y(_05393_),
    .A(net6388),
    .B(net3064));
 sg13g2_a21o_1 _19925_ (.A2(_05376_),
    .A1(_04686_),
    .B1(_04665_),
    .X(_05394_));
 sg13g2_nand3_1 _19926_ (.B(_04686_),
    .C(_05376_),
    .A(_04665_),
    .Y(_05395_));
 sg13g2_and2_1 _19927_ (.A(net5772),
    .B(_05395_),
    .X(_05396_));
 sg13g2_a21oi_1 _19928_ (.A1(\soc_inst.cpu_core.alu.b[21] ),
    .A2(net6272),
    .Y(_05397_),
    .B1(_05381_));
 sg13g2_a21o_1 _19929_ (.A2(_05397_),
    .A1(_05380_),
    .B1(_04666_),
    .X(_05398_));
 sg13g2_nand3_1 _19930_ (.B(_05380_),
    .C(_05397_),
    .A(_04666_),
    .Y(_05399_));
 sg13g2_nand3_1 _19931_ (.B(_05398_),
    .C(_05399_),
    .A(net5759),
    .Y(_05400_));
 sg13g2_mux2_1 _19932_ (.A0(\soc_inst.cpu_core.alu.a[22] ),
    .A1(net6273),
    .S(net6257),
    .X(_05401_));
 sg13g2_mux2_1 _19933_ (.A0(_05360_),
    .A1(_05401_),
    .S(net6113),
    .X(_05402_));
 sg13g2_mux2_1 _19934_ (.A0(_05317_),
    .A1(_05402_),
    .S(net6121),
    .X(_05403_));
 sg13g2_a22oi_1 _19935_ (.Y(_05404_),
    .B1(_05403_),
    .B2(net5454),
    .A2(_05239_),
    .A1(net5453));
 sg13g2_a21oi_1 _19936_ (.A1(_05036_),
    .A2(_05404_),
    .Y(_05405_),
    .B1(net6219));
 sg13g2_nand2_1 _19937_ (.Y(_05406_),
    .A(_05051_),
    .B(net5452));
 sg13g2_nor2_1 _19938_ (.A(_04664_),
    .B(_04805_),
    .Y(_05407_));
 sg13g2_a21oi_1 _19939_ (.A1(_04665_),
    .A2(net5763),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_o21ai_1 _19940_ (.B1(_05408_),
    .Y(_05409_),
    .A1(_04663_),
    .A2(_04797_));
 sg13g2_nor3_1 _19941_ (.A(net5094),
    .B(_05405_),
    .C(_05409_),
    .Y(_05410_));
 sg13g2_nand3_1 _19942_ (.B(_05406_),
    .C(_05410_),
    .A(_05400_),
    .Y(_05411_));
 sg13g2_a21oi_2 _19943_ (.B1(_05411_),
    .Y(_05412_),
    .A2(_05396_),
    .A1(_05394_));
 sg13g2_o21ai_1 _19944_ (.B1(_05393_),
    .Y(_01368_),
    .A1(net5242),
    .A2(_05412_));
 sg13g2_and2_1 _19945_ (.A(_04685_),
    .B(_05394_),
    .X(_05413_));
 sg13g2_xnor2_1 _19946_ (.Y(_05414_),
    .A(_04672_),
    .B(_05413_));
 sg13g2_mux2_1 _19947_ (.A0(\soc_inst.cpu_core.alu.a[23] ),
    .A1(\soc_inst.cpu_core.alu.a[22] ),
    .S(net6258),
    .X(_05415_));
 sg13g2_mux2_1 _19948_ (.A0(_05383_),
    .A1(_05415_),
    .S(net6114),
    .X(_05416_));
 sg13g2_mux2_1 _19949_ (.A0(_05336_),
    .A1(_05416_),
    .S(net6125),
    .X(_05417_));
 sg13g2_a221oi_1 _19950_ (.B2(_04848_),
    .C1(_05082_),
    .B1(_05417_),
    .A1(_05096_),
    .Y(_05418_),
    .A2(_05260_));
 sg13g2_o21ai_1 _19951_ (.B1(_04671_),
    .Y(_05419_),
    .A1(net6287),
    .A2(_04670_));
 sg13g2_o21ai_1 _19952_ (.B1(_05255_),
    .Y(_05420_),
    .A1(_04672_),
    .A2(net5761));
 sg13g2_a221oi_1 _19953_ (.B2(net5767),
    .C1(_05420_),
    .B1(_05419_),
    .A1(_05069_),
    .Y(_05421_),
    .A2(net5452));
 sg13g2_o21ai_1 _19954_ (.B1(_05421_),
    .Y(_05422_),
    .A1(net6218),
    .A2(_05418_));
 sg13g2_a21oi_1 _19955_ (.A1(_04664_),
    .A2(_05398_),
    .Y(_05423_),
    .B1(_04672_));
 sg13g2_nand3_1 _19956_ (.B(_04672_),
    .C(_05398_),
    .A(_04664_),
    .Y(_05424_));
 sg13g2_nor2_1 _19957_ (.A(net5757),
    .B(_05423_),
    .Y(_05425_));
 sg13g2_a221oi_1 _19958_ (.B2(_05425_),
    .C1(_05422_),
    .B1(_05424_),
    .A1(net5772),
    .Y(_05426_),
    .A2(_05414_));
 sg13g2_nand2_1 _19959_ (.Y(_05427_),
    .A(net6394),
    .B(net2964));
 sg13g2_o21ai_1 _19960_ (.B1(_05427_),
    .Y(_01369_),
    .A1(net5241),
    .A2(_05426_));
 sg13g2_nor4_1 _19961_ (.A(_04662_),
    .B(_04666_),
    .C(_04669_),
    .D(_04672_),
    .Y(_05428_));
 sg13g2_o21ai_1 _19962_ (.B1(_05428_),
    .Y(_05429_),
    .A1(_05353_),
    .A2(_05356_));
 sg13g2_o21ai_1 _19963_ (.B1(_04671_),
    .Y(_05430_),
    .A1(_04664_),
    .A2(_04670_));
 sg13g2_nor3_1 _19964_ (.A(_04666_),
    .B(_04672_),
    .C(_05397_),
    .Y(_05431_));
 sg13g2_nor2_1 _19965_ (.A(_05430_),
    .B(_05431_),
    .Y(_05432_));
 sg13g2_nand3_1 _19966_ (.B(_05429_),
    .C(_05432_),
    .A(_04710_),
    .Y(_05433_));
 sg13g2_a21oi_1 _19967_ (.A1(_05429_),
    .A2(_05432_),
    .Y(_05434_),
    .B1(_04710_));
 sg13g2_nor2_1 _19968_ (.A(net5758),
    .B(_05434_),
    .Y(_05435_));
 sg13g2_a221oi_1 _19969_ (.B2(_04707_),
    .C1(_05254_),
    .B1(net5458),
    .A1(_04708_),
    .Y(_05436_),
    .A2(net5460));
 sg13g2_o21ai_1 _19970_ (.B1(_05436_),
    .Y(_05437_),
    .A1(_04710_),
    .A2(net5761));
 sg13g2_and2_1 _19971_ (.A(net5462),
    .B(_05101_),
    .X(_05438_));
 sg13g2_nor2_1 _19972_ (.A(net6135),
    .B(_05097_),
    .Y(_05439_));
 sg13g2_nand2_1 _19973_ (.Y(_05440_),
    .A(net6233),
    .B(_05361_));
 sg13g2_mux2_1 _19974_ (.A0(\soc_inst.cpu_core.alu.a[24] ),
    .A1(\soc_inst.cpu_core.alu.a[23] ),
    .S(net6257),
    .X(_05441_));
 sg13g2_mux2_1 _19975_ (.A0(_05401_),
    .A1(_05441_),
    .S(net6113),
    .X(_05442_));
 sg13g2_a21oi_1 _19976_ (.A1(net6121),
    .A2(_05442_),
    .Y(_05443_),
    .B1(net6225));
 sg13g2_a221oi_1 _19977_ (.B2(_05443_),
    .C1(_04810_),
    .B1(_05440_),
    .A1(net6225),
    .Y(_05444_),
    .A2(_05280_));
 sg13g2_nor4_1 _19978_ (.A(_05437_),
    .B(_05438_),
    .C(_05439_),
    .D(_05444_),
    .Y(_05445_));
 sg13g2_nand2b_1 _19979_ (.Y(_05446_),
    .B(_04710_),
    .A_N(_04699_));
 sg13g2_a21oi_1 _19980_ (.A1(_04699_),
    .A2(_04709_),
    .Y(_05447_),
    .B1(net5770));
 sg13g2_a22oi_1 _19981_ (.Y(_05448_),
    .B1(_05446_),
    .B2(_05447_),
    .A2(_05435_),
    .A1(_05433_));
 sg13g2_a21oi_2 _19982_ (.B1(net5241),
    .Y(_05449_),
    .A2(_05448_),
    .A1(_05445_));
 sg13g2_a21o_1 _19983_ (.A2(net3235),
    .A1(net6360),
    .B1(_05449_),
    .X(_01370_));
 sg13g2_nor3_1 _19984_ (.A(_04707_),
    .B(_04714_),
    .C(_05434_),
    .Y(_05450_));
 sg13g2_o21ai_1 _19985_ (.B1(_04714_),
    .Y(_05451_),
    .A1(_04707_),
    .A2(_05434_));
 sg13g2_nand2_1 _19986_ (.Y(_05452_),
    .A(net5760),
    .B(_05451_));
 sg13g2_nor2_1 _19987_ (.A(_05450_),
    .B(_05452_),
    .Y(_05453_));
 sg13g2_nand2b_1 _19988_ (.Y(_05454_),
    .B(_04715_),
    .A_N(_05446_));
 sg13g2_nand3_1 _19989_ (.B(_04717_),
    .C(_05446_),
    .A(_04714_),
    .Y(_05455_));
 sg13g2_nor2_1 _19990_ (.A(net5770),
    .B(_04718_),
    .Y(_05456_));
 sg13g2_nand3_1 _19991_ (.B(_05455_),
    .C(_05456_),
    .A(_05454_),
    .Y(_05457_));
 sg13g2_nand2_1 _19992_ (.Y(_05458_),
    .A(_05120_),
    .B(net5452));
 sg13g2_a22oi_1 _19993_ (.Y(_05459_),
    .B1(net5458),
    .B2(_04712_),
    .A2(net5460),
    .A1(_04711_));
 sg13g2_a21oi_1 _19994_ (.A1(_04714_),
    .A2(net5763),
    .Y(_05460_),
    .B1(net5094));
 sg13g2_mux2_1 _19995_ (.A0(\soc_inst.cpu_core.alu.a[25] ),
    .A1(\soc_inst.cpu_core.alu.a[24] ),
    .S(net6258),
    .X(_05461_));
 sg13g2_mux2_1 _19996_ (.A0(_05415_),
    .A1(_05461_),
    .S(net6114),
    .X(_05462_));
 sg13g2_mux4_1 _19997_ (.S0(net6125),
    .A0(_05215_),
    .A1(_05298_),
    .A2(_05384_),
    .A3(_05462_),
    .S1(net6132),
    .X(_05463_));
 sg13g2_a22oi_1 _19998_ (.Y(_05464_),
    .B1(_05463_),
    .B2(net5457),
    .A2(_05127_),
    .A1(net6136));
 sg13g2_nand4_1 _19999_ (.B(_05459_),
    .C(_05460_),
    .A(_05458_),
    .Y(_05465_),
    .D(_05464_));
 sg13g2_nor2_1 _20000_ (.A(_05453_),
    .B(_05465_),
    .Y(_05466_));
 sg13g2_a21oi_2 _20001_ (.B1(net5241),
    .Y(_05467_),
    .A2(_05466_),
    .A1(_05457_));
 sg13g2_a21o_1 _20002_ (.A2(net3273),
    .A1(net6354),
    .B1(_05467_),
    .X(_01371_));
 sg13g2_a21oi_1 _20003_ (.A1(_04707_),
    .A2(_04711_),
    .Y(_05468_),
    .B1(_04712_));
 sg13g2_nand3_1 _20004_ (.B(_04713_),
    .C(_05451_),
    .A(_04706_),
    .Y(_05469_));
 sg13g2_a21o_1 _20005_ (.A2(_05451_),
    .A1(_04713_),
    .B1(_04706_),
    .X(_05470_));
 sg13g2_nand3_1 _20006_ (.B(_05469_),
    .C(_05470_),
    .A(net5759),
    .Y(_05471_));
 sg13g2_a21o_1 _20007_ (.A2(_05454_),
    .A1(_04719_),
    .B1(_04705_),
    .X(_05472_));
 sg13g2_nand3_1 _20008_ (.B(_04719_),
    .C(_05454_),
    .A(_04705_),
    .Y(_05473_));
 sg13g2_nand3_1 _20009_ (.B(_05472_),
    .C(_05473_),
    .A(net5772),
    .Y(_05474_));
 sg13g2_nor2_1 _20010_ (.A(net6121),
    .B(_05402_),
    .Y(_05475_));
 sg13g2_mux2_1 _20011_ (.A0(net6267),
    .A1(\soc_inst.cpu_core.alu.a[25] ),
    .S(net6257),
    .X(_05476_));
 sg13g2_mux2_1 _20012_ (.A0(_05441_),
    .A1(_05476_),
    .S(net6113),
    .X(_05477_));
 sg13g2_o21ai_1 _20013_ (.B1(net6134),
    .Y(_05478_),
    .A1(net6233),
    .A2(_05477_));
 sg13g2_nand2_1 _20014_ (.Y(_05479_),
    .A(net6225),
    .B(_05318_));
 sg13g2_o21ai_1 _20015_ (.B1(_05479_),
    .Y(_05480_),
    .A1(_05475_),
    .A2(_05478_));
 sg13g2_o21ai_1 _20016_ (.B1(_04703_),
    .Y(_05481_),
    .A1(net6288),
    .A2(_04704_));
 sg13g2_a221oi_1 _20017_ (.B2(net5767),
    .C1(_05254_),
    .B1(_05481_),
    .A1(_04705_),
    .Y(_05482_),
    .A2(net5763));
 sg13g2_o21ai_1 _20018_ (.B1(_05482_),
    .Y(_05483_),
    .A1(_05145_),
    .A2(_05284_));
 sg13g2_a21oi_1 _20019_ (.A1(net5456),
    .A2(_05480_),
    .Y(_05484_),
    .B1(_05483_));
 sg13g2_or2_1 _20020_ (.X(_05485_),
    .B(_05150_),
    .A(net6218));
 sg13g2_nand4_1 _20021_ (.B(_05474_),
    .C(_05484_),
    .A(_05471_),
    .Y(_05486_),
    .D(_05485_));
 sg13g2_a22oi_1 _20022_ (.Y(_05487_),
    .B1(_04555_),
    .B2(_05486_),
    .A2(net3338),
    .A1(net6426));
 sg13g2_inv_1 _20023_ (.Y(_01372_),
    .A(_05487_));
 sg13g2_a21oi_1 _20024_ (.A1(_04703_),
    .A2(_05470_),
    .Y(_05488_),
    .B1(_04702_));
 sg13g2_nand3_1 _20025_ (.B(_04703_),
    .C(_05470_),
    .A(_04702_),
    .Y(_05489_));
 sg13g2_nor2_1 _20026_ (.A(net5758),
    .B(_05488_),
    .Y(_05490_));
 sg13g2_nand2_1 _20027_ (.Y(_05491_),
    .A(_04721_),
    .B(_05472_));
 sg13g2_xor2_1 _20028_ (.B(_05491_),
    .A(_04702_),
    .X(_05492_));
 sg13g2_a21o_1 _20029_ (.A2(net6258),
    .A1(net6267),
    .B1(_04819_),
    .X(_05493_));
 sg13g2_mux2_1 _20030_ (.A0(_05461_),
    .A1(_05493_),
    .S(net6114),
    .X(_05494_));
 sg13g2_nand2_1 _20031_ (.Y(_05495_),
    .A(net6235),
    .B(_05416_));
 sg13g2_a21oi_1 _20032_ (.A1(net6126),
    .A2(_05494_),
    .Y(_05496_),
    .B1(net6226));
 sg13g2_nor2_1 _20033_ (.A(net6132),
    .B(_05337_),
    .Y(_05497_));
 sg13g2_a21oi_1 _20034_ (.A1(_05495_),
    .A2(_05496_),
    .Y(_05498_),
    .B1(_05497_));
 sg13g2_nand2_1 _20035_ (.Y(_05499_),
    .A(net5456),
    .B(_05498_));
 sg13g2_a221oi_1 _20036_ (.B2(_04701_),
    .C1(net5094),
    .B1(net5458),
    .A1(_04700_),
    .Y(_05500_),
    .A2(net5460));
 sg13g2_o21ai_1 _20037_ (.B1(_05500_),
    .Y(_05501_),
    .A1(_04702_),
    .A2(net5761));
 sg13g2_a221oi_1 _20038_ (.B2(_05164_),
    .C1(_05501_),
    .B1(net5452),
    .A1(net6135),
    .Y(_05502_),
    .A2(_05171_));
 sg13g2_nand2_1 _20039_ (.Y(_05503_),
    .A(_05499_),
    .B(_05502_));
 sg13g2_a221oi_1 _20040_ (.B2(net5773),
    .C1(_05503_),
    .B1(_05492_),
    .A1(_05489_),
    .Y(_05504_),
    .A2(_05490_));
 sg13g2_nand2_1 _20041_ (.Y(_05505_),
    .A(net6395),
    .B(net3204));
 sg13g2_o21ai_1 _20042_ (.B1(_05505_),
    .Y(_01373_),
    .A1(net5241),
    .A2(_05504_));
 sg13g2_or4_1 _20043_ (.A(_04702_),
    .B(_04706_),
    .C(_04710_),
    .D(_04715_),
    .X(_05506_));
 sg13g2_a21oi_1 _20044_ (.A1(_05429_),
    .A2(_05432_),
    .Y(_05507_),
    .B1(_05506_));
 sg13g2_nor2b_1 _20045_ (.A(_04703_),
    .B_N(_04700_),
    .Y(_05508_));
 sg13g2_nor3_1 _20046_ (.A(_04702_),
    .B(_04706_),
    .C(_05468_),
    .Y(_05509_));
 sg13g2_or3_1 _20047_ (.A(_04701_),
    .B(_05508_),
    .C(_05509_),
    .X(_05510_));
 sg13g2_nor2_1 _20048_ (.A(_05507_),
    .B(_05510_),
    .Y(_05511_));
 sg13g2_or2_1 _20049_ (.X(_05512_),
    .B(_05511_),
    .A(_04726_));
 sg13g2_a21oi_1 _20050_ (.A1(_04726_),
    .A2(_05511_),
    .Y(_05513_),
    .B1(net5757));
 sg13g2_nor2_1 _20051_ (.A(_04724_),
    .B(_04726_),
    .Y(_05514_));
 sg13g2_nor2_1 _20052_ (.A(net5770),
    .B(_05514_),
    .Y(_05515_));
 sg13g2_o21ai_1 _20053_ (.B1(net5767),
    .Y(_05516_),
    .A1(\soc_inst.cpu_core.alu.b[28] ),
    .A2(net6264));
 sg13g2_a21oi_1 _20054_ (.A1(net6287),
    .A2(_04725_),
    .Y(_05517_),
    .B1(_05516_));
 sg13g2_o21ai_1 _20055_ (.B1(_05255_),
    .Y(_05518_),
    .A1(_04726_),
    .A2(net5761));
 sg13g2_mux2_1 _20056_ (.A0(net6264),
    .A1(\soc_inst.cpu_core.alu.a[27] ),
    .S(net6257),
    .X(_05519_));
 sg13g2_a22oi_1 _20057_ (.Y(_05520_),
    .B1(_05519_),
    .B2(_04785_),
    .A2(_05476_),
    .A1(_04783_));
 sg13g2_a21oi_1 _20058_ (.A1(net6233),
    .A2(_05442_),
    .Y(_05521_),
    .B1(net6225));
 sg13g2_a221oi_1 _20059_ (.B2(_05521_),
    .C1(_04810_),
    .B1(_05520_),
    .A1(net6225),
    .Y(_05522_),
    .A2(_05363_));
 sg13g2_nor3_1 _20060_ (.A(_05517_),
    .B(_05518_),
    .C(_05522_),
    .Y(_05523_));
 sg13g2_o21ai_1 _20061_ (.B1(_05523_),
    .Y(_05524_),
    .A1(net6218),
    .A2(_05192_));
 sg13g2_a21o_1 _20062_ (.A2(net5452),
    .A1(_05185_),
    .B1(_05524_),
    .X(_05525_));
 sg13g2_a221oi_1 _20063_ (.B2(_04727_),
    .C1(_05525_),
    .B1(_05515_),
    .A1(_05512_),
    .Y(_05526_),
    .A2(_05513_));
 sg13g2_nand2_1 _20064_ (.Y(_05527_),
    .A(net6355),
    .B(net2993));
 sg13g2_o21ai_1 _20065_ (.B1(_05527_),
    .Y(_01374_),
    .A1(net5242),
    .A2(_05526_));
 sg13g2_nand2_1 _20066_ (.Y(_05528_),
    .A(net6367),
    .B(net3095));
 sg13g2_nor2_1 _20067_ (.A(_04559_),
    .B(_04730_),
    .Y(_05529_));
 sg13g2_a21oi_1 _20068_ (.A1(_04559_),
    .A2(_04730_),
    .Y(_05530_),
    .B1(net5771));
 sg13g2_nand2_1 _20069_ (.Y(_05531_),
    .A(_04728_),
    .B(_05530_));
 sg13g2_a21oi_1 _20070_ (.A1(_04727_),
    .A2(_05529_),
    .Y(_05532_),
    .B1(_05531_));
 sg13g2_nand3_1 _20071_ (.B(_04725_),
    .C(_05512_),
    .A(_04559_),
    .Y(_05533_));
 sg13g2_nor2_1 _20072_ (.A(_04559_),
    .B(_04726_),
    .Y(_05534_));
 sg13g2_o21ai_1 _20073_ (.B1(_05534_),
    .Y(_05535_),
    .A1(_05507_),
    .A2(_05510_));
 sg13g2_nor2_1 _20074_ (.A(_04559_),
    .B(_04725_),
    .Y(_05536_));
 sg13g2_nor2_1 _20075_ (.A(net5757),
    .B(_05536_),
    .Y(_05537_));
 sg13g2_and2_1 _20076_ (.A(_05535_),
    .B(_05537_),
    .X(_05538_));
 sg13g2_nor2_1 _20077_ (.A(net6220),
    .B(_05210_),
    .Y(_05539_));
 sg13g2_nor2_1 _20078_ (.A(_04820_),
    .B(_04823_),
    .Y(_05540_));
 sg13g2_o21ai_1 _20079_ (.B1(net6130),
    .Y(_05541_),
    .A1(net5769),
    .A2(_05540_));
 sg13g2_a221oi_1 _20080_ (.B2(_04783_),
    .C1(_05541_),
    .B1(_05493_),
    .A1(net6235),
    .Y(_05542_),
    .A2(_05462_));
 sg13g2_o21ai_1 _20081_ (.B1(net5457),
    .Y(_05543_),
    .A1(net6133),
    .A2(_05385_));
 sg13g2_nor2_1 _20082_ (.A(_05542_),
    .B(_05543_),
    .Y(_05544_));
 sg13g2_nand3_1 _20083_ (.B(net6263),
    .C(net5458),
    .A(\soc_inst.cpu_core.alu.b[29] ),
    .Y(_05545_));
 sg13g2_o21ai_1 _20084_ (.B1(net5460),
    .Y(_05546_),
    .A1(\soc_inst.cpu_core.alu.b[29] ),
    .A2(net6263));
 sg13g2_nor2_1 _20085_ (.A(_04559_),
    .B(net5761),
    .Y(_05547_));
 sg13g2_nand3_1 _20086_ (.B(_05545_),
    .C(_05546_),
    .A(_05255_),
    .Y(_05548_));
 sg13g2_or4_1 _20087_ (.A(_05539_),
    .B(_05544_),
    .C(_05547_),
    .D(_05548_),
    .X(_05549_));
 sg13g2_a221oi_1 _20088_ (.B2(_05538_),
    .C1(_05549_),
    .B1(_05533_),
    .A1(_05218_),
    .Y(_05550_),
    .A2(net5452));
 sg13g2_nor2b_2 _20089_ (.A(_05532_),
    .B_N(_05550_),
    .Y(_05551_));
 sg13g2_o21ai_1 _20090_ (.B1(_05528_),
    .Y(_01375_),
    .A1(net5242),
    .A2(_05551_));
 sg13g2_nand3_1 _20091_ (.B(_04731_),
    .C(_04733_),
    .A(_04728_),
    .Y(_05552_));
 sg13g2_nand3_1 _20092_ (.B(_04735_),
    .C(_05552_),
    .A(net5772),
    .Y(_05553_));
 sg13g2_a21oi_1 _20093_ (.A1(\soc_inst.cpu_core.alu.b[29] ),
    .A2(net6263),
    .Y(_05554_),
    .B1(_05536_));
 sg13g2_a21oi_1 _20094_ (.A1(_05535_),
    .A2(_05554_),
    .Y(_05555_),
    .B1(_04734_));
 sg13g2_nand3_1 _20095_ (.B(_05535_),
    .C(_05554_),
    .A(_04734_),
    .Y(_05556_));
 sg13g2_nor2_1 _20096_ (.A(net5758),
    .B(_05555_),
    .Y(_05557_));
 sg13g2_mux2_1 _20097_ (.A0(\soc_inst.cpu_core.alu.a[30] ),
    .A1(net6263),
    .S(net6257),
    .X(_05558_));
 sg13g2_a22oi_1 _20098_ (.Y(_05559_),
    .B1(_05558_),
    .B2(_04785_),
    .A2(_05519_),
    .A1(_04783_));
 sg13g2_a21oi_1 _20099_ (.A1(net6233),
    .A2(_05477_),
    .Y(_05560_),
    .B1(net6225));
 sg13g2_nor2_1 _20100_ (.A(net6134),
    .B(_05403_),
    .Y(_05561_));
 sg13g2_a21oi_1 _20101_ (.A1(_05559_),
    .A2(_05560_),
    .Y(_05562_),
    .B1(_05561_));
 sg13g2_a22oi_1 _20102_ (.Y(_05563_),
    .B1(_05562_),
    .B2(net5456),
    .A2(_05234_),
    .A1(net6135));
 sg13g2_nand2b_1 _20103_ (.Y(_05564_),
    .B(_05283_),
    .A_N(_05241_));
 sg13g2_o21ai_1 _20104_ (.B1(_04797_),
    .Y(_05565_),
    .A1(_04732_),
    .A2(net5761));
 sg13g2_o21ai_1 _20105_ (.B1(_05565_),
    .Y(_05566_),
    .A1(\soc_inst.cpu_core.alu.b[30] ),
    .A2(\soc_inst.cpu_core.alu.a[30] ));
 sg13g2_a21oi_1 _20106_ (.A1(_04732_),
    .A2(net5458),
    .Y(_05567_),
    .B1(net5094));
 sg13g2_nand4_1 _20107_ (.B(_05564_),
    .C(_05566_),
    .A(_05563_),
    .Y(_05568_),
    .D(_05567_));
 sg13g2_a21oi_1 _20108_ (.A1(_05556_),
    .A2(_05557_),
    .Y(_05569_),
    .B1(_05568_));
 sg13g2_a21oi_1 _20109_ (.A1(_05553_),
    .A2(_05569_),
    .Y(_05570_),
    .B1(net5241));
 sg13g2_a21o_1 _20110_ (.A2(net3329),
    .A1(net6409),
    .B1(_05570_),
    .X(_01376_));
 sg13g2_xnor2_1 _20111_ (.Y(_05571_),
    .A(_04558_),
    .B(_04736_));
 sg13g2_nor3_1 _20112_ (.A(_04558_),
    .B(_04732_),
    .C(_05555_),
    .Y(_05572_));
 sg13g2_o21ai_1 _20113_ (.B1(_04558_),
    .Y(_05573_),
    .A1(_04732_),
    .A2(_05555_));
 sg13g2_nor2_1 _20114_ (.A(net5757),
    .B(_05572_),
    .Y(_05574_));
 sg13g2_a21oi_1 _20115_ (.A1(\soc_inst.cpu_core.alu.a[30] ),
    .A2(net6259),
    .Y(_05575_),
    .B1(net6248));
 sg13g2_a221oi_1 _20116_ (.B2(_04832_),
    .C1(net6235),
    .B1(_05575_),
    .A1(net6247),
    .Y(_05576_),
    .A2(_05540_));
 sg13g2_a21o_1 _20117_ (.A2(_05494_),
    .A1(net6234),
    .B1(_05576_),
    .X(_05577_));
 sg13g2_a221oi_1 _20118_ (.B2(net5454),
    .C1(_05252_),
    .B1(_05577_),
    .A1(net5453),
    .Y(_05578_),
    .A2(_05417_));
 sg13g2_o21ai_1 _20119_ (.B1(net5461),
    .Y(_05579_),
    .A1(\soc_inst.cpu_core.alu.b[31] ),
    .A2(net6261));
 sg13g2_nand3_1 _20120_ (.B(net6261),
    .C(net5459),
    .A(\soc_inst.cpu_core.alu.b[31] ),
    .Y(_05580_));
 sg13g2_a21oi_1 _20121_ (.A1(_04558_),
    .A2(net5764),
    .Y(_05581_),
    .B1(_05075_));
 sg13g2_nand3_1 _20122_ (.B(_05580_),
    .C(_05581_),
    .A(_05579_),
    .Y(_05582_));
 sg13g2_a21oi_1 _20123_ (.A1(_05261_),
    .A2(_05283_),
    .Y(_05583_),
    .B1(_05582_));
 sg13g2_o21ai_1 _20124_ (.B1(_05583_),
    .Y(_05584_),
    .A1(net6218),
    .A2(_05578_));
 sg13g2_a221oi_1 _20125_ (.B2(_05574_),
    .C1(_05584_),
    .B1(_05573_),
    .A1(net5773),
    .Y(_05585_),
    .A2(_05571_));
 sg13g2_nand2_1 _20126_ (.Y(_05586_),
    .A(net6367),
    .B(net1394));
 sg13g2_o21ai_1 _20127_ (.B1(_05586_),
    .Y(_01377_),
    .A1(net5242),
    .A2(_05585_));
 sg13g2_nor3_1 _20128_ (.A(net6376),
    .B(net6306),
    .C(_11403_),
    .Y(_05587_));
 sg13g2_a22oi_1 _20129_ (.Y(_05588_),
    .B1(_11393_),
    .B2(_05587_),
    .A2(net2128),
    .A1(net6370));
 sg13g2_inv_1 _20130_ (.Y(_01378_),
    .A(net2129));
 sg13g2_a21oi_1 _20131_ (.A1(net6413),
    .A2(_08130_),
    .Y(_01379_),
    .B1(_11395_));
 sg13g2_nor2b_2 _20132_ (.A(net6214),
    .B_N(net6216),
    .Y(_05589_));
 sg13g2_nor2b_2 _20133_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .B_N(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .Y(_05590_));
 sg13g2_nand2_1 _20134_ (.Y(_05591_),
    .A(_05589_),
    .B(_05590_));
 sg13g2_nor2_2 _20135_ (.A(_09505_),
    .B(_05591_),
    .Y(_05592_));
 sg13g2_nor2_1 _20136_ (.A(net1949),
    .B(net5444),
    .Y(_05593_));
 sg13g2_a21oi_1 _20137_ (.A1(net4994),
    .A2(net5444),
    .Y(_01380_),
    .B1(_05593_));
 sg13g2_nor2_1 _20138_ (.A(net2311),
    .B(net5444),
    .Y(_05594_));
 sg13g2_a21oi_1 _20139_ (.A1(net4989),
    .A2(net5444),
    .Y(_01381_),
    .B1(_05594_));
 sg13g2_nor2_1 _20140_ (.A(net1575),
    .B(net5444),
    .Y(_05595_));
 sg13g2_a21oi_1 _20141_ (.A1(net4984),
    .A2(net5444),
    .Y(_01382_),
    .B1(_05595_));
 sg13g2_nor2_1 _20142_ (.A(net2308),
    .B(net5442),
    .Y(_05596_));
 sg13g2_a21oi_1 _20143_ (.A1(net4979),
    .A2(net5442),
    .Y(_01383_),
    .B1(_05596_));
 sg13g2_nor2_1 _20144_ (.A(net2184),
    .B(net5450),
    .Y(_05597_));
 sg13g2_a21oi_1 _20145_ (.A1(net4976),
    .A2(net5450),
    .Y(_01384_),
    .B1(_05597_));
 sg13g2_nor2_1 _20146_ (.A(net2240),
    .B(net5450),
    .Y(_05598_));
 sg13g2_a21oi_1 _20147_ (.A1(net4973),
    .A2(net5450),
    .Y(_01385_),
    .B1(_05598_));
 sg13g2_nor2_1 _20148_ (.A(net1379),
    .B(net5445),
    .Y(_05599_));
 sg13g2_a21oi_1 _20149_ (.A1(net4965),
    .A2(net5445),
    .Y(_01386_),
    .B1(_05599_));
 sg13g2_nor2_1 _20150_ (.A(net1157),
    .B(net5447),
    .Y(_05600_));
 sg13g2_a21oi_1 _20151_ (.A1(net4917),
    .A2(net5447),
    .Y(_01387_),
    .B1(_05600_));
 sg13g2_nor2_1 _20152_ (.A(net1221),
    .B(net5444),
    .Y(_05601_));
 sg13g2_a21oi_1 _20153_ (.A1(net4782),
    .A2(net5444),
    .Y(_01388_),
    .B1(_05601_));
 sg13g2_nor2_1 _20154_ (.A(net1609),
    .B(net5450),
    .Y(_05602_));
 sg13g2_a21oi_1 _20155_ (.A1(net4914),
    .A2(net5450),
    .Y(_01389_),
    .B1(_05602_));
 sg13g2_nor2_1 _20156_ (.A(net1884),
    .B(net5449),
    .Y(_05603_));
 sg13g2_a21oi_1 _20157_ (.A1(net4908),
    .A2(net5449),
    .Y(_01390_),
    .B1(_05603_));
 sg13g2_nor2_1 _20158_ (.A(net1275),
    .B(net5445),
    .Y(_05604_));
 sg13g2_a21oi_1 _20159_ (.A1(net4775),
    .A2(net5445),
    .Y(_01391_),
    .B1(_05604_));
 sg13g2_nor2_1 _20160_ (.A(net2376),
    .B(net5448),
    .Y(_05605_));
 sg13g2_a21oi_1 _20161_ (.A1(net4902),
    .A2(net5448),
    .Y(_01392_),
    .B1(_05605_));
 sg13g2_nor2_1 _20162_ (.A(net1555),
    .B(net5448),
    .Y(_05606_));
 sg13g2_a21oi_1 _20163_ (.A1(net4959),
    .A2(net5448),
    .Y(_01393_),
    .B1(_05606_));
 sg13g2_nor2_1 _20164_ (.A(net2290),
    .B(net5442),
    .Y(_05607_));
 sg13g2_a21oi_1 _20165_ (.A1(net4954),
    .A2(net5442),
    .Y(_01394_),
    .B1(_05607_));
 sg13g2_nor2_1 _20166_ (.A(net1782),
    .B(net5448),
    .Y(_05608_));
 sg13g2_a21oi_1 _20167_ (.A1(net4895),
    .A2(net5448),
    .Y(_01395_),
    .B1(_05608_));
 sg13g2_nor2_1 _20168_ (.A(net2107),
    .B(net5447),
    .Y(_05609_));
 sg13g2_a21oi_1 _20169_ (.A1(net4890),
    .A2(net5447),
    .Y(_01396_),
    .B1(_05609_));
 sg13g2_nor2_1 _20170_ (.A(net1527),
    .B(net5443),
    .Y(_05610_));
 sg13g2_a21oi_1 _20171_ (.A1(net4885),
    .A2(net5443),
    .Y(_01397_),
    .B1(_05610_));
 sg13g2_nor2_1 _20172_ (.A(net1601),
    .B(net5448),
    .Y(_05611_));
 sg13g2_a21oi_1 _20173_ (.A1(net4771),
    .A2(net5448),
    .Y(_01398_),
    .B1(_05611_));
 sg13g2_nor2_1 _20174_ (.A(net1847),
    .B(net5447),
    .Y(_05612_));
 sg13g2_a21oi_1 _20175_ (.A1(net4878),
    .A2(net5447),
    .Y(_01399_),
    .B1(_05612_));
 sg13g2_nor2_1 _20176_ (.A(net1589),
    .B(net5449),
    .Y(_05613_));
 sg13g2_a21oi_1 _20177_ (.A1(net4875),
    .A2(net5449),
    .Y(_01400_),
    .B1(_05613_));
 sg13g2_nor2_1 _20178_ (.A(net1898),
    .B(net5450),
    .Y(_05614_));
 sg13g2_a21oi_1 _20179_ (.A1(net4764),
    .A2(net5450),
    .Y(_01401_),
    .B1(_05614_));
 sg13g2_nor2_1 _20180_ (.A(net1781),
    .B(net5443),
    .Y(_05615_));
 sg13g2_a21oi_1 _20181_ (.A1(net4868),
    .A2(net5443),
    .Y(_01402_),
    .B1(_05615_));
 sg13g2_nor2_1 _20182_ (.A(net2082),
    .B(net5449),
    .Y(_05616_));
 sg13g2_a21oi_1 _20183_ (.A1(net4863),
    .A2(net5449),
    .Y(_01403_),
    .B1(_05616_));
 sg13g2_nor2_1 _20184_ (.A(net1495),
    .B(net5443),
    .Y(_05617_));
 sg13g2_a21oi_1 _20185_ (.A1(net4857),
    .A2(net5443),
    .Y(_01404_),
    .B1(_05617_));
 sg13g2_nor2_1 _20186_ (.A(net2119),
    .B(net5442),
    .Y(_05618_));
 sg13g2_a21oi_1 _20187_ (.A1(net4853),
    .A2(net5442),
    .Y(_01405_),
    .B1(_05618_));
 sg13g2_nor2_1 _20188_ (.A(net2165),
    .B(net5447),
    .Y(_05619_));
 sg13g2_a21oi_1 _20189_ (.A1(net4847),
    .A2(net5447),
    .Y(_01406_),
    .B1(_05619_));
 sg13g2_nor2_1 _20190_ (.A(net2123),
    .B(net5442),
    .Y(_05620_));
 sg13g2_a21oi_1 _20191_ (.A1(net4844),
    .A2(net5442),
    .Y(_01407_),
    .B1(_05620_));
 sg13g2_nor2_1 _20192_ (.A(net2285),
    .B(net5443),
    .Y(_05621_));
 sg13g2_a21oi_1 _20193_ (.A1(net4837),
    .A2(net5446),
    .Y(_01408_),
    .B1(_05621_));
 sg13g2_nor2_1 _20194_ (.A(net1736),
    .B(net5445),
    .Y(_05622_));
 sg13g2_a21oi_1 _20195_ (.A1(net4834),
    .A2(net5445),
    .Y(_01409_),
    .B1(_05622_));
 sg13g2_nor2_1 _20196_ (.A(net1780),
    .B(net5451),
    .Y(_05623_));
 sg13g2_a21oi_1 _20197_ (.A1(net4828),
    .A2(net5451),
    .Y(_01410_),
    .B1(_05623_));
 sg13g2_nor2_1 _20198_ (.A(net2071),
    .B(net5449),
    .Y(_05624_));
 sg13g2_a21oi_1 _20199_ (.A1(net4825),
    .A2(net5449),
    .Y(_01411_),
    .B1(_05624_));
 sg13g2_nor2b_2 _20200_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .B_N(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .Y(_05625_));
 sg13g2_nand2_1 _20201_ (.Y(_05626_),
    .A(_05589_),
    .B(_05625_));
 sg13g2_nor2_2 _20202_ (.A(_09505_),
    .B(_05626_),
    .Y(_05627_));
 sg13g2_nor2_1 _20203_ (.A(net1687),
    .B(net5434),
    .Y(_05628_));
 sg13g2_a21oi_1 _20204_ (.A1(net4996),
    .A2(net5434),
    .Y(_01412_),
    .B1(_05628_));
 sg13g2_nor2_1 _20205_ (.A(net1708),
    .B(net5434),
    .Y(_05629_));
 sg13g2_a21oi_1 _20206_ (.A1(net4990),
    .A2(net5434),
    .Y(_01413_),
    .B1(_05629_));
 sg13g2_nor2_1 _20207_ (.A(net1410),
    .B(net5434),
    .Y(_05630_));
 sg13g2_a21oi_1 _20208_ (.A1(net4987),
    .A2(net5434),
    .Y(_01414_),
    .B1(_05630_));
 sg13g2_nor2_1 _20209_ (.A(net1852),
    .B(net5432),
    .Y(_05631_));
 sg13g2_a21oi_1 _20210_ (.A1(net4979),
    .A2(net5432),
    .Y(_01415_),
    .B1(_05631_));
 sg13g2_nor2_1 _20211_ (.A(net2027),
    .B(net5438),
    .Y(_05632_));
 sg13g2_a21oi_1 _20212_ (.A1(net4977),
    .A2(net5438),
    .Y(_01416_),
    .B1(_05632_));
 sg13g2_nor2_1 _20213_ (.A(net2121),
    .B(net5440),
    .Y(_05633_));
 sg13g2_a21oi_1 _20214_ (.A1(net4969),
    .A2(net5440),
    .Y(_01417_),
    .B1(_05633_));
 sg13g2_nor2_1 _20215_ (.A(net1528),
    .B(net5434),
    .Y(_05634_));
 sg13g2_a21oi_1 _20216_ (.A1(net4967),
    .A2(net5434),
    .Y(_01418_),
    .B1(_05634_));
 sg13g2_nor2_1 _20217_ (.A(net1891),
    .B(net5437),
    .Y(_05635_));
 sg13g2_a21oi_1 _20218_ (.A1(net4916),
    .A2(net5437),
    .Y(_01419_),
    .B1(_05635_));
 sg13g2_nor2_1 _20219_ (.A(net1437),
    .B(net5435),
    .Y(_05636_));
 sg13g2_a21oi_1 _20220_ (.A1(_09603_),
    .A2(net5435),
    .Y(_01420_),
    .B1(_05636_));
 sg13g2_nor2_1 _20221_ (.A(net1828),
    .B(net5440),
    .Y(_05637_));
 sg13g2_a21oi_1 _20222_ (.A1(net4913),
    .A2(net5440),
    .Y(_01421_),
    .B1(_05637_));
 sg13g2_nor2_1 _20223_ (.A(net1339),
    .B(net5439),
    .Y(_05638_));
 sg13g2_a21oi_1 _20224_ (.A1(net4905),
    .A2(net5439),
    .Y(_01422_),
    .B1(_05638_));
 sg13g2_nor2_1 _20225_ (.A(net1794),
    .B(net5435),
    .Y(_05639_));
 sg13g2_a21oi_1 _20226_ (.A1(net4776),
    .A2(net5435),
    .Y(_01423_),
    .B1(_05639_));
 sg13g2_nor2_1 _20227_ (.A(net1874),
    .B(net5437),
    .Y(_05640_));
 sg13g2_a21oi_1 _20228_ (.A1(net4901),
    .A2(net5441),
    .Y(_01424_),
    .B1(_05640_));
 sg13g2_nor2_1 _20229_ (.A(net1477),
    .B(net5437),
    .Y(_05641_));
 sg13g2_a21oi_1 _20230_ (.A1(net4961),
    .A2(net5437),
    .Y(_01425_),
    .B1(_05641_));
 sg13g2_nor2_1 _20231_ (.A(net2241),
    .B(net5432),
    .Y(_05642_));
 sg13g2_a21oi_1 _20232_ (.A1(net4957),
    .A2(net5432),
    .Y(_01426_),
    .B1(_05642_));
 sg13g2_nor2_1 _20233_ (.A(net1922),
    .B(net5437),
    .Y(_05643_));
 sg13g2_a21oi_1 _20234_ (.A1(net4895),
    .A2(net5441),
    .Y(_01427_),
    .B1(_05643_));
 sg13g2_nor2_1 _20235_ (.A(net1830),
    .B(net5438),
    .Y(_05644_));
 sg13g2_a21oi_1 _20236_ (.A1(net4889),
    .A2(net5438),
    .Y(_01428_),
    .B1(_05644_));
 sg13g2_nor2_1 _20237_ (.A(net2575),
    .B(net5433),
    .Y(_05645_));
 sg13g2_a21oi_1 _20238_ (.A1(net4884),
    .A2(net5433),
    .Y(_01429_),
    .B1(_05645_));
 sg13g2_nor2_1 _20239_ (.A(net1819),
    .B(net5437),
    .Y(_05646_));
 sg13g2_a21oi_1 _20240_ (.A1(net4771),
    .A2(net5437),
    .Y(_01430_),
    .B1(_05646_));
 sg13g2_nor2_1 _20241_ (.A(net2186),
    .B(net5438),
    .Y(_05647_));
 sg13g2_a21oi_1 _20242_ (.A1(net4879),
    .A2(net5438),
    .Y(_01431_),
    .B1(_05647_));
 sg13g2_nor2_1 _20243_ (.A(net1701),
    .B(net5439),
    .Y(_05648_));
 sg13g2_a21oi_1 _20244_ (.A1(net4875),
    .A2(net5439),
    .Y(_01432_),
    .B1(_05648_));
 sg13g2_nor2_1 _20245_ (.A(net1426),
    .B(net5440),
    .Y(_05649_));
 sg13g2_a21oi_1 _20246_ (.A1(net4763),
    .A2(net5440),
    .Y(_01433_),
    .B1(_05649_));
 sg13g2_nor2_1 _20247_ (.A(net1917),
    .B(net5432),
    .Y(_05650_));
 sg13g2_a21oi_1 _20248_ (.A1(net4871),
    .A2(net5433),
    .Y(_01434_),
    .B1(_05650_));
 sg13g2_nor2_1 _20249_ (.A(net2126),
    .B(net5439),
    .Y(_05651_));
 sg13g2_a21oi_1 _20250_ (.A1(net4863),
    .A2(net5441),
    .Y(_01435_),
    .B1(_05651_));
 sg13g2_nor2_1 _20251_ (.A(net2001),
    .B(net5433),
    .Y(_05652_));
 sg13g2_a21oi_1 _20252_ (.A1(net4860),
    .A2(net5433),
    .Y(_01436_),
    .B1(_05652_));
 sg13g2_nor2_1 _20253_ (.A(net1547),
    .B(net5432),
    .Y(_05653_));
 sg13g2_a21oi_1 _20254_ (.A1(net4854),
    .A2(net5432),
    .Y(_01437_),
    .B1(_05653_));
 sg13g2_nor2_1 _20255_ (.A(net1880),
    .B(net5438),
    .Y(_05654_));
 sg13g2_a21oi_1 _20256_ (.A1(net4848),
    .A2(net5438),
    .Y(_01438_),
    .B1(_05654_));
 sg13g2_nor2_1 _20257_ (.A(net1541),
    .B(net5432),
    .Y(_05655_));
 sg13g2_a21oi_1 _20258_ (.A1(net4842),
    .A2(net5433),
    .Y(_01439_),
    .B1(_05655_));
 sg13g2_nor2_1 _20259_ (.A(net1762),
    .B(net5433),
    .Y(_05656_));
 sg13g2_a21oi_1 _20260_ (.A1(net4837),
    .A2(net5436),
    .Y(_01440_),
    .B1(_05656_));
 sg13g2_nor2_1 _20261_ (.A(net1485),
    .B(net5435),
    .Y(_05657_));
 sg13g2_a21oi_1 _20262_ (.A1(net4832),
    .A2(net5435),
    .Y(_01441_),
    .B1(_05657_));
 sg13g2_nor2_1 _20263_ (.A(net1345),
    .B(net5439),
    .Y(_05658_));
 sg13g2_a21oi_1 _20264_ (.A1(net4829),
    .A2(net5439),
    .Y(_01442_),
    .B1(_05658_));
 sg13g2_nor2_1 _20265_ (.A(net1425),
    .B(net5439),
    .Y(_05659_));
 sg13g2_a21oi_1 _20266_ (.A1(net4823),
    .A2(net5440),
    .Y(_01443_),
    .B1(_05659_));
 sg13g2_nor2_2 _20267_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .Y(_05660_));
 sg13g2_nand3_1 _20268_ (.B(_05589_),
    .C(_05660_),
    .A(net6096),
    .Y(_05661_));
 sg13g2_nand2_1 _20269_ (.Y(_05662_),
    .A(net493),
    .B(net5749));
 sg13g2_o21ai_1 _20270_ (.B1(_05662_),
    .Y(_01444_),
    .A1(net4995),
    .A2(net5749));
 sg13g2_nand2_1 _20271_ (.Y(_05663_),
    .A(net1023),
    .B(net5749));
 sg13g2_o21ai_1 _20272_ (.B1(_05663_),
    .Y(_01445_),
    .A1(net4991),
    .A2(net5749));
 sg13g2_nand2_1 _20273_ (.Y(_05664_),
    .A(net972),
    .B(net5749));
 sg13g2_o21ai_1 _20274_ (.B1(_05664_),
    .Y(_01446_),
    .A1(net4988),
    .A2(net5749));
 sg13g2_nand2_1 _20275_ (.Y(_05665_),
    .A(net599),
    .B(net5747));
 sg13g2_o21ai_1 _20276_ (.B1(_05665_),
    .Y(_01447_),
    .A1(net4983),
    .A2(net5747));
 sg13g2_nand2_1 _20277_ (.Y(_05666_),
    .A(net1050),
    .B(net5753));
 sg13g2_o21ai_1 _20278_ (.B1(_05666_),
    .Y(_01448_),
    .A1(net4975),
    .A2(net5753));
 sg13g2_nand2_1 _20279_ (.Y(_05667_),
    .A(net862),
    .B(net5754));
 sg13g2_o21ai_1 _20280_ (.B1(_05667_),
    .Y(_01449_),
    .A1(net4969),
    .A2(net5754));
 sg13g2_nand2_1 _20281_ (.Y(_05668_),
    .A(net1214),
    .B(net5750));
 sg13g2_o21ai_1 _20282_ (.B1(_05668_),
    .Y(_01450_),
    .A1(net4965),
    .A2(net5750));
 sg13g2_nand2_1 _20283_ (.Y(_05669_),
    .A(net443),
    .B(net5753));
 sg13g2_o21ai_1 _20284_ (.B1(_05669_),
    .Y(_01451_),
    .A1(net4917),
    .A2(net5753));
 sg13g2_nand2_1 _20285_ (.Y(_05670_),
    .A(net1684),
    .B(net5750));
 sg13g2_o21ai_1 _20286_ (.B1(_05670_),
    .Y(_01452_),
    .A1(net4782),
    .A2(net5750));
 sg13g2_nand2_1 _20287_ (.Y(_05671_),
    .A(net459),
    .B(net5754));
 sg13g2_o21ai_1 _20288_ (.B1(_05671_),
    .Y(_01453_),
    .A1(net4911),
    .A2(net5754));
 sg13g2_nand2_1 _20289_ (.Y(_05672_),
    .A(net588),
    .B(net5755));
 sg13g2_o21ai_1 _20290_ (.B1(_05672_),
    .Y(_01454_),
    .A1(net4905),
    .A2(net5755));
 sg13g2_nand2_1 _20291_ (.Y(_05673_),
    .A(net868),
    .B(net5750));
 sg13g2_o21ai_1 _20292_ (.B1(_05673_),
    .Y(_01455_),
    .A1(net4777),
    .A2(net5750));
 sg13g2_nand2_1 _20293_ (.Y(_05674_),
    .A(net861),
    .B(net5752));
 sg13g2_o21ai_1 _20294_ (.B1(_05674_),
    .Y(_01456_),
    .A1(net4899),
    .A2(net5752));
 sg13g2_nand2_1 _20295_ (.Y(_05675_),
    .A(net1611),
    .B(net5752));
 sg13g2_o21ai_1 _20296_ (.B1(_05675_),
    .Y(_01457_),
    .A1(net4960),
    .A2(net5752));
 sg13g2_nand2_1 _20297_ (.Y(_05676_),
    .A(net521),
    .B(net5747));
 sg13g2_o21ai_1 _20298_ (.B1(_05676_),
    .Y(_01458_),
    .A1(net4958),
    .A2(net5747));
 sg13g2_nand2_1 _20299_ (.Y(_05677_),
    .A(net1634),
    .B(net5756));
 sg13g2_o21ai_1 _20300_ (.B1(_05677_),
    .Y(_01459_),
    .A1(net4894),
    .A2(net5756));
 sg13g2_nand2_1 _20301_ (.Y(_05678_),
    .A(net1326),
    .B(net5752));
 sg13g2_o21ai_1 _20302_ (.B1(_05678_),
    .Y(_01460_),
    .A1(net4892),
    .A2(net5752));
 sg13g2_nand2_1 _20303_ (.Y(_05679_),
    .A(net1129),
    .B(net5748));
 sg13g2_o21ai_1 _20304_ (.B1(_05679_),
    .Y(_01461_),
    .A1(net4887),
    .A2(net5748));
 sg13g2_nand2_1 _20305_ (.Y(_05680_),
    .A(net969),
    .B(net5752));
 sg13g2_o21ai_1 _20306_ (.B1(_05680_),
    .Y(_01462_),
    .A1(net4772),
    .A2(net5752));
 sg13g2_nand2_1 _20307_ (.Y(_05681_),
    .A(net968),
    .B(net5753));
 sg13g2_o21ai_1 _20308_ (.B1(_05681_),
    .Y(_01463_),
    .A1(net4882),
    .A2(net5753));
 sg13g2_nand2_1 _20309_ (.Y(_05682_),
    .A(net420),
    .B(net5755));
 sg13g2_o21ai_1 _20310_ (.B1(_05682_),
    .Y(_01464_),
    .A1(net4873),
    .A2(net5755));
 sg13g2_nand2_1 _20311_ (.Y(_05683_),
    .A(net706),
    .B(net5754));
 sg13g2_o21ai_1 _20312_ (.B1(_05683_),
    .Y(_01465_),
    .A1(net4762),
    .A2(net5754));
 sg13g2_nand2_1 _20313_ (.Y(_05684_),
    .A(net879),
    .B(net5747));
 sg13g2_o21ai_1 _20314_ (.B1(_05684_),
    .Y(_01466_),
    .A1(net4868),
    .A2(net5747));
 sg13g2_nand2_1 _20315_ (.Y(_05685_),
    .A(net582),
    .B(net5755));
 sg13g2_o21ai_1 _20316_ (.B1(_05685_),
    .Y(_01467_),
    .A1(net4866),
    .A2(net5755));
 sg13g2_nand2_1 _20317_ (.Y(_05686_),
    .A(net623),
    .B(net5748));
 sg13g2_o21ai_1 _20318_ (.B1(_05686_),
    .Y(_01468_),
    .A1(net4859),
    .A2(net5748));
 sg13g2_nand2_1 _20319_ (.Y(_05687_),
    .A(net714),
    .B(net5747));
 sg13g2_o21ai_1 _20320_ (.B1(_05687_),
    .Y(_01469_),
    .A1(net4855),
    .A2(net5747));
 sg13g2_nand2_1 _20321_ (.Y(_05688_),
    .A(net1047),
    .B(net5753));
 sg13g2_o21ai_1 _20322_ (.B1(_05688_),
    .Y(_01470_),
    .A1(net4847),
    .A2(net5753));
 sg13g2_nand2_1 _20323_ (.Y(_05689_),
    .A(net1552),
    .B(net5748));
 sg13g2_o21ai_1 _20324_ (.B1(_05689_),
    .Y(_01471_),
    .A1(net4845),
    .A2(net5748));
 sg13g2_nand2_1 _20325_ (.Y(_05690_),
    .A(net451),
    .B(net5751));
 sg13g2_o21ai_1 _20326_ (.B1(_05690_),
    .Y(_01472_),
    .A1(net4837),
    .A2(net5748));
 sg13g2_nand2_1 _20327_ (.Y(_05691_),
    .A(net1107),
    .B(net5749));
 sg13g2_o21ai_1 _20328_ (.B1(_05691_),
    .Y(_01473_),
    .A1(net4835),
    .A2(net5749));
 sg13g2_nand2_1 _20329_ (.Y(_05692_),
    .A(net677),
    .B(net5755));
 sg13g2_o21ai_1 _20330_ (.B1(_05692_),
    .Y(_01474_),
    .A1(net4827),
    .A2(net5755));
 sg13g2_nand2_1 _20331_ (.Y(_05693_),
    .A(net540),
    .B(net5754));
 sg13g2_o21ai_1 _20332_ (.B1(_05693_),
    .Y(_01475_),
    .A1(net4826),
    .A2(net5754));
 sg13g2_nor2b_2 _20333_ (.A(net6216),
    .B_N(net6214),
    .Y(_05694_));
 sg13g2_and3_2 _20334_ (.X(_05695_),
    .A(net6096),
    .B(_09507_),
    .C(_05694_));
 sg13g2_nor2_1 _20335_ (.A(net1613),
    .B(net5424),
    .Y(_05696_));
 sg13g2_a21oi_1 _20336_ (.A1(net4995),
    .A2(net5424),
    .Y(_01476_),
    .B1(_05696_));
 sg13g2_nor2_1 _20337_ (.A(net2131),
    .B(net5424),
    .Y(_05697_));
 sg13g2_a21oi_1 _20338_ (.A1(net4990),
    .A2(net5424),
    .Y(_01477_),
    .B1(_05697_));
 sg13g2_nor2_1 _20339_ (.A(net1342),
    .B(net5424),
    .Y(_05698_));
 sg13g2_a21oi_1 _20340_ (.A1(net4987),
    .A2(net5424),
    .Y(_01478_),
    .B1(_05698_));
 sg13g2_nor2_1 _20341_ (.A(net2031),
    .B(net5421),
    .Y(_05699_));
 sg13g2_a21oi_1 _20342_ (.A1(net4981),
    .A2(net5421),
    .Y(_01479_),
    .B1(_05699_));
 sg13g2_nor2_1 _20343_ (.A(net2289),
    .B(net5421),
    .Y(_05700_));
 sg13g2_a21oi_1 _20344_ (.A1(net4978),
    .A2(net5421),
    .Y(_01480_),
    .B1(_05700_));
 sg13g2_nor2_1 _20345_ (.A(net1903),
    .B(net5429),
    .Y(_05701_));
 sg13g2_a21oi_1 _20346_ (.A1(net4970),
    .A2(net5429),
    .Y(_01481_),
    .B1(_05701_));
 sg13g2_nor2_1 _20347_ (.A(net1327),
    .B(net5424),
    .Y(_05702_));
 sg13g2_a21oi_1 _20348_ (.A1(net4966),
    .A2(net5424),
    .Y(_01482_),
    .B1(_05702_));
 sg13g2_nor2_1 _20349_ (.A(net2168),
    .B(net5427),
    .Y(_05703_));
 sg13g2_a21oi_1 _20350_ (.A1(net4918),
    .A2(net5427),
    .Y(_01483_),
    .B1(_05703_));
 sg13g2_nor2_1 _20351_ (.A(net1305),
    .B(net5425),
    .Y(_05704_));
 sg13g2_a21oi_1 _20352_ (.A1(net4779),
    .A2(net5425),
    .Y(_01484_),
    .B1(_05704_));
 sg13g2_nor2_1 _20353_ (.A(net2057),
    .B(net5429),
    .Y(_05705_));
 sg13g2_a21oi_1 _20354_ (.A1(net4913),
    .A2(net5429),
    .Y(_01485_),
    .B1(_05705_));
 sg13g2_nor2_1 _20355_ (.A(net1940),
    .B(net5430),
    .Y(_05706_));
 sg13g2_a21oi_1 _20356_ (.A1(net4907),
    .A2(net5430),
    .Y(_01486_),
    .B1(_05706_));
 sg13g2_nor2_1 _20357_ (.A(net2120),
    .B(net5425),
    .Y(_05707_));
 sg13g2_a21oi_1 _20358_ (.A1(net4776),
    .A2(net5425),
    .Y(_01487_),
    .B1(_05707_));
 sg13g2_nor2_1 _20359_ (.A(net1632),
    .B(net5428),
    .Y(_05708_));
 sg13g2_a21oi_1 _20360_ (.A1(net4901),
    .A2(net5428),
    .Y(_01488_),
    .B1(_05708_));
 sg13g2_nor2_1 _20361_ (.A(net1519),
    .B(net5428),
    .Y(_05709_));
 sg13g2_a21oi_1 _20362_ (.A1(net4962),
    .A2(net5428),
    .Y(_01489_),
    .B1(_05709_));
 sg13g2_nor2_1 _20363_ (.A(net2494),
    .B(net5423),
    .Y(_05710_));
 sg13g2_a21oi_1 _20364_ (.A1(net4957),
    .A2(net5423),
    .Y(_01490_),
    .B1(_05710_));
 sg13g2_nor2_1 _20365_ (.A(net1407),
    .B(net5428),
    .Y(_05711_));
 sg13g2_a21oi_1 _20366_ (.A1(net4894),
    .A2(net5428),
    .Y(_01491_),
    .B1(_05711_));
 sg13g2_nor2_1 _20367_ (.A(net2201),
    .B(net5427),
    .Y(_05712_));
 sg13g2_a21oi_1 _20368_ (.A1(net4891),
    .A2(net5427),
    .Y(_01492_),
    .B1(_05712_));
 sg13g2_nor2_1 _20369_ (.A(net1532),
    .B(net5421),
    .Y(_05713_));
 sg13g2_a21oi_1 _20370_ (.A1(net4887),
    .A2(net5421),
    .Y(_01493_),
    .B1(_05713_));
 sg13g2_nor2_1 _20371_ (.A(net1389),
    .B(net5428),
    .Y(_05714_));
 sg13g2_a21oi_1 _20372_ (.A1(net4772),
    .A2(net5428),
    .Y(_01494_),
    .B1(_05714_));
 sg13g2_nor2_1 _20373_ (.A(net1610),
    .B(net5427),
    .Y(_05715_));
 sg13g2_a21oi_1 _20374_ (.A1(net4881),
    .A2(net5427),
    .Y(_01495_),
    .B1(_05715_));
 sg13g2_nor2_1 _20375_ (.A(net1790),
    .B(net5430),
    .Y(_05716_));
 sg13g2_a21oi_1 _20376_ (.A1(net4874),
    .A2(net5430),
    .Y(_01496_),
    .B1(_05716_));
 sg13g2_nor2_1 _20377_ (.A(net2202),
    .B(net5429),
    .Y(_05717_));
 sg13g2_a21oi_1 _20378_ (.A1(net4766),
    .A2(net5429),
    .Y(_01497_),
    .B1(_05717_));
 sg13g2_nor2_1 _20379_ (.A(net1333),
    .B(net5423),
    .Y(_05718_));
 sg13g2_a21oi_1 _20380_ (.A1(net4867),
    .A2(net5423),
    .Y(_01498_),
    .B1(_05718_));
 sg13g2_nor2_1 _20381_ (.A(net1521),
    .B(net5430),
    .Y(_05719_));
 sg13g2_a21oi_1 _20382_ (.A1(net4862),
    .A2(net5430),
    .Y(_01499_),
    .B1(_05719_));
 sg13g2_nor2_1 _20383_ (.A(net1676),
    .B(net5422),
    .Y(_05720_));
 sg13g2_a21oi_1 _20384_ (.A1(net4860),
    .A2(net5422),
    .Y(_01500_),
    .B1(_05720_));
 sg13g2_nor2_1 _20385_ (.A(net1872),
    .B(net5423),
    .Y(_05721_));
 sg13g2_a21oi_1 _20386_ (.A1(net4854),
    .A2(net5423),
    .Y(_01501_),
    .B1(_05721_));
 sg13g2_nor2_1 _20387_ (.A(net1515),
    .B(net5427),
    .Y(_05722_));
 sg13g2_a21oi_1 _20388_ (.A1(net4850),
    .A2(net5427),
    .Y(_01502_),
    .B1(_05722_));
 sg13g2_nor2_1 _20389_ (.A(net1715),
    .B(net5423),
    .Y(_05723_));
 sg13g2_a21oi_1 _20390_ (.A1(net4844),
    .A2(net5423),
    .Y(_01503_),
    .B1(_05723_));
 sg13g2_nor2_1 _20391_ (.A(net1720),
    .B(net5421),
    .Y(_05724_));
 sg13g2_a21oi_1 _20392_ (.A1(net4839),
    .A2(net5421),
    .Y(_01504_),
    .B1(_05724_));
 sg13g2_nor2_1 _20393_ (.A(net1978),
    .B(net5422),
    .Y(_05725_));
 sg13g2_a21oi_1 _20394_ (.A1(net4833),
    .A2(net5422),
    .Y(_01505_),
    .B1(_05725_));
 sg13g2_nor2_1 _20395_ (.A(net2088),
    .B(net5430),
    .Y(_05726_));
 sg13g2_a21oi_1 _20396_ (.A1(net4829),
    .A2(net5430),
    .Y(_01506_),
    .B1(_05726_));
 sg13g2_nor2_1 _20397_ (.A(net1536),
    .B(net5429),
    .Y(_05727_));
 sg13g2_a21oi_1 _20398_ (.A1(net4823),
    .A2(net5429),
    .Y(_01507_),
    .B1(_05727_));
 sg13g2_nor2_2 _20399_ (.A(net6215),
    .B(net6216),
    .Y(_05728_));
 sg13g2_nor4_1 _20400_ (.A(net6214),
    .B(net6216),
    .C(_09505_),
    .D(_09506_),
    .Y(_05729_));
 sg13g2_nor2_1 _20401_ (.A(net1774),
    .B(net5740),
    .Y(_05730_));
 sg13g2_a21oi_1 _20402_ (.A1(net4994),
    .A2(net5740),
    .Y(_01508_),
    .B1(_05730_));
 sg13g2_nor2_1 _20403_ (.A(net2491),
    .B(net5740),
    .Y(_05731_));
 sg13g2_a21oi_1 _20404_ (.A1(net4991),
    .A2(net5740),
    .Y(_01509_),
    .B1(_05731_));
 sg13g2_nor2_1 _20405_ (.A(net1400),
    .B(net5740),
    .Y(_05732_));
 sg13g2_a21oi_1 _20406_ (.A1(net4987),
    .A2(net5740),
    .Y(_01510_),
    .B1(_05732_));
 sg13g2_nor2_1 _20407_ (.A(net2468),
    .B(net5737),
    .Y(_05733_));
 sg13g2_a21oi_1 _20408_ (.A1(net4979),
    .A2(net5737),
    .Y(_01511_),
    .B1(_05733_));
 sg13g2_nor2_1 _20409_ (.A(net1953),
    .B(net5743),
    .Y(_05734_));
 sg13g2_a21oi_1 _20410_ (.A1(net4975),
    .A2(net5743),
    .Y(_01512_),
    .B1(_05734_));
 sg13g2_nor2_1 _20411_ (.A(net1803),
    .B(net5745),
    .Y(_05735_));
 sg13g2_a21oi_1 _20412_ (.A1(net4970),
    .A2(net5745),
    .Y(_01513_),
    .B1(_05735_));
 sg13g2_nor2_1 _20413_ (.A(net1933),
    .B(net5739),
    .Y(_05736_));
 sg13g2_a21oi_1 _20414_ (.A1(net4966),
    .A2(net5739),
    .Y(_01514_),
    .B1(_05736_));
 sg13g2_nor2_1 _20415_ (.A(net1850),
    .B(net5742),
    .Y(_05737_));
 sg13g2_a21oi_1 _20416_ (.A1(net4916),
    .A2(net5742),
    .Y(_01515_),
    .B1(_05737_));
 sg13g2_nor2_1 _20417_ (.A(net1972),
    .B(net5739),
    .Y(_05738_));
 sg13g2_a21oi_1 _20418_ (.A1(net4780),
    .A2(net5739),
    .Y(_01516_),
    .B1(_05738_));
 sg13g2_nor2_1 _20419_ (.A(net1773),
    .B(net5745),
    .Y(_05739_));
 sg13g2_a21oi_1 _20420_ (.A1(net4911),
    .A2(net5744),
    .Y(_01517_),
    .B1(_05739_));
 sg13g2_nor2_1 _20421_ (.A(net2326),
    .B(net5744),
    .Y(_05740_));
 sg13g2_a21oi_1 _20422_ (.A1(net4909),
    .A2(net5744),
    .Y(_01518_),
    .B1(_05740_));
 sg13g2_nor2_1 _20423_ (.A(net1827),
    .B(net5739),
    .Y(_05741_));
 sg13g2_a21oi_1 _20424_ (.A1(net4777),
    .A2(net5739),
    .Y(_01519_),
    .B1(_05741_));
 sg13g2_nor2_1 _20425_ (.A(net1761),
    .B(net5741),
    .Y(_05742_));
 sg13g2_a21oi_1 _20426_ (.A1(net4899),
    .A2(net5741),
    .Y(_01520_),
    .B1(_05742_));
 sg13g2_nor2_1 _20427_ (.A(net1608),
    .B(net5741),
    .Y(_05743_));
 sg13g2_a21oi_1 _20428_ (.A1(net4959),
    .A2(net5741),
    .Y(_01521_),
    .B1(_05743_));
 sg13g2_nor2_1 _20429_ (.A(net2108),
    .B(net5737),
    .Y(_05744_));
 sg13g2_a21oi_1 _20430_ (.A1(net4954),
    .A2(net5737),
    .Y(_01522_),
    .B1(_05744_));
 sg13g2_nor2_1 _20431_ (.A(net1588),
    .B(net5742),
    .Y(_05745_));
 sg13g2_a21oi_1 _20432_ (.A1(net4897),
    .A2(net5742),
    .Y(_01523_),
    .B1(_05745_));
 sg13g2_nor2_1 _20433_ (.A(net1499),
    .B(net5741),
    .Y(_05746_));
 sg13g2_a21oi_1 _20434_ (.A1(net4893),
    .A2(net5741),
    .Y(_01524_),
    .B1(_05746_));
 sg13g2_nor2_1 _20435_ (.A(net1250),
    .B(net5738),
    .Y(_05747_));
 sg13g2_a21oi_1 _20436_ (.A1(net4884),
    .A2(net5738),
    .Y(_01525_),
    .B1(_05747_));
 sg13g2_nor2_1 _20437_ (.A(net1433),
    .B(net5741),
    .Y(_05748_));
 sg13g2_a21oi_1 _20438_ (.A1(net4772),
    .A2(net5741),
    .Y(_01526_),
    .B1(_05748_));
 sg13g2_nor2_1 _20439_ (.A(net1971),
    .B(net5743),
    .Y(_05749_));
 sg13g2_a21oi_1 _20440_ (.A1(net4878),
    .A2(net5743),
    .Y(_01527_),
    .B1(_05749_));
 sg13g2_nor2_1 _20441_ (.A(net1448),
    .B(net5744),
    .Y(_05750_));
 sg13g2_a21oi_1 _20442_ (.A1(net4876),
    .A2(net5744),
    .Y(_01528_),
    .B1(_05750_));
 sg13g2_nor2_1 _20443_ (.A(net1729),
    .B(net5745),
    .Y(_05751_));
 sg13g2_a21oi_1 _20444_ (.A1(net4764),
    .A2(net5745),
    .Y(_01529_),
    .B1(_05751_));
 sg13g2_nor2_1 _20445_ (.A(net2198),
    .B(net5738),
    .Y(_05752_));
 sg13g2_a21oi_1 _20446_ (.A1(net4868),
    .A2(net5738),
    .Y(_01530_),
    .B1(_05752_));
 sg13g2_nor2_1 _20447_ (.A(net1451),
    .B(net5746),
    .Y(_05753_));
 sg13g2_a21oi_1 _20448_ (.A1(net4865),
    .A2(net5745),
    .Y(_01531_),
    .B1(_05753_));
 sg13g2_nor2_1 _20449_ (.A(net1461),
    .B(net5738),
    .Y(_05754_));
 sg13g2_a21oi_1 _20450_ (.A1(net4858),
    .A2(net5738),
    .Y(_01532_),
    .B1(_05754_));
 sg13g2_nor2_1 _20451_ (.A(net1824),
    .B(net5737),
    .Y(_05755_));
 sg13g2_a21oi_1 _20452_ (.A1(net4852),
    .A2(net5737),
    .Y(_01533_),
    .B1(_05755_));
 sg13g2_nor2_1 _20453_ (.A(net1938),
    .B(net5743),
    .Y(_05756_));
 sg13g2_a21oi_1 _20454_ (.A1(net4849),
    .A2(net5743),
    .Y(_01534_),
    .B1(_05756_));
 sg13g2_nor2_1 _20455_ (.A(net1592),
    .B(net5737),
    .Y(_05757_));
 sg13g2_a21oi_1 _20456_ (.A1(net4844),
    .A2(net5737),
    .Y(_01535_),
    .B1(_05757_));
 sg13g2_nor2_1 _20457_ (.A(net1603),
    .B(net5738),
    .Y(_05758_));
 sg13g2_a21oi_1 _20458_ (.A1(net4837),
    .A2(net5746),
    .Y(_01536_),
    .B1(_05758_));
 sg13g2_nor2_1 _20459_ (.A(net2148),
    .B(net5739),
    .Y(_05759_));
 sg13g2_a21oi_1 _20460_ (.A1(net4833),
    .A2(net5739),
    .Y(_01537_),
    .B1(_05759_));
 sg13g2_nor2_1 _20461_ (.A(net1727),
    .B(net5744),
    .Y(_05760_));
 sg13g2_a21oi_1 _20462_ (.A1(net4828),
    .A2(net5744),
    .Y(_01538_),
    .B1(_05760_));
 sg13g2_nor2_1 _20463_ (.A(net2422),
    .B(net5744),
    .Y(_05761_));
 sg13g2_a21oi_1 _20464_ (.A1(net4822),
    .A2(net5745),
    .Y(_01539_),
    .B1(_05761_));
 sg13g2_nand3_1 _20465_ (.B(_05590_),
    .C(_05728_),
    .A(net6096),
    .Y(_05762_));
 sg13g2_nand2_1 _20466_ (.Y(_05763_),
    .A(net565),
    .B(net5729));
 sg13g2_o21ai_1 _20467_ (.B1(_05763_),
    .Y(_01540_),
    .A1(net4996),
    .A2(net5729));
 sg13g2_nand2_1 _20468_ (.Y(_05764_),
    .A(net1637),
    .B(net5729));
 sg13g2_o21ai_1 _20469_ (.B1(_05764_),
    .Y(_01541_),
    .A1(net4992),
    .A2(net5729));
 sg13g2_nand2_1 _20470_ (.Y(_05765_),
    .A(net634),
    .B(net5729));
 sg13g2_o21ai_1 _20471_ (.B1(_05765_),
    .Y(_01542_),
    .A1(net4986),
    .A2(net5729));
 sg13g2_nand2_1 _20472_ (.Y(_05766_),
    .A(net934),
    .B(net5727));
 sg13g2_o21ai_1 _20473_ (.B1(_05766_),
    .Y(_01543_),
    .A1(net4979),
    .A2(net5727));
 sg13g2_nand2_1 _20474_ (.Y(_05767_),
    .A(net1049),
    .B(net5733));
 sg13g2_o21ai_1 _20475_ (.B1(_05767_),
    .Y(_01544_),
    .A1(net4975),
    .A2(net5733));
 sg13g2_nand2_1 _20476_ (.Y(_05768_),
    .A(net805),
    .B(net5735));
 sg13g2_o21ai_1 _20477_ (.B1(_05768_),
    .Y(_01545_),
    .A1(net4969),
    .A2(net5735));
 sg13g2_nand2_1 _20478_ (.Y(_05769_),
    .A(net811),
    .B(net5730));
 sg13g2_o21ai_1 _20479_ (.B1(_05769_),
    .Y(_01546_),
    .A1(net4968),
    .A2(net5730));
 sg13g2_nand2_1 _20480_ (.Y(_05770_),
    .A(net1328),
    .B(net5732));
 sg13g2_o21ai_1 _20481_ (.B1(_05770_),
    .Y(_01547_),
    .A1(net4917),
    .A2(net5732));
 sg13g2_nand2_1 _20482_ (.Y(_05771_),
    .A(net838),
    .B(net5729));
 sg13g2_o21ai_1 _20483_ (.B1(_05771_),
    .Y(_01548_),
    .A1(net4780),
    .A2(net5730));
 sg13g2_nand2_1 _20484_ (.Y(_05772_),
    .A(net617),
    .B(net5735));
 sg13g2_o21ai_1 _20485_ (.B1(_05772_),
    .Y(_01549_),
    .A1(net4911),
    .A2(net5735));
 sg13g2_nand2_1 _20486_ (.Y(_05773_),
    .A(net624),
    .B(net5734));
 sg13g2_o21ai_1 _20487_ (.B1(_05773_),
    .Y(_01550_),
    .A1(net4905),
    .A2(net5734));
 sg13g2_nand2_1 _20488_ (.Y(_05774_),
    .A(net1201),
    .B(net5730));
 sg13g2_o21ai_1 _20489_ (.B1(_05774_),
    .Y(_01551_),
    .A1(net4776),
    .A2(net5730));
 sg13g2_nand2_1 _20490_ (.Y(_05775_),
    .A(net939),
    .B(net5732));
 sg13g2_o21ai_1 _20491_ (.B1(_05775_),
    .Y(_01552_),
    .A1(net4899),
    .A2(net5736));
 sg13g2_nand2_1 _20492_ (.Y(_05776_),
    .A(net832),
    .B(net5732));
 sg13g2_o21ai_1 _20493_ (.B1(_05776_),
    .Y(_01553_),
    .A1(net4959),
    .A2(net5732));
 sg13g2_nand2_1 _20494_ (.Y(_05777_),
    .A(net1370),
    .B(net5727));
 sg13g2_o21ai_1 _20495_ (.B1(_05777_),
    .Y(_01554_),
    .A1(net4957),
    .A2(net5727));
 sg13g2_nand2_1 _20496_ (.Y(_05778_),
    .A(net606),
    .B(net5732));
 sg13g2_o21ai_1 _20497_ (.B1(_05778_),
    .Y(_01555_),
    .A1(net4898),
    .A2(net5736));
 sg13g2_nand2_1 _20498_ (.Y(_05779_),
    .A(net1080),
    .B(net5733));
 sg13g2_o21ai_1 _20499_ (.B1(_05779_),
    .Y(_01556_),
    .A1(net4889),
    .A2(net5733));
 sg13g2_nand2_1 _20500_ (.Y(_05780_),
    .A(net1171),
    .B(net5728));
 sg13g2_o21ai_1 _20501_ (.B1(_05780_),
    .Y(_01557_),
    .A1(net4885),
    .A2(net5728));
 sg13g2_nand2_1 _20502_ (.Y(_05781_),
    .A(net691),
    .B(net5732));
 sg13g2_o21ai_1 _20503_ (.B1(_05781_),
    .Y(_01558_),
    .A1(net4769),
    .A2(net5732));
 sg13g2_nand2_1 _20504_ (.Y(_05782_),
    .A(net848),
    .B(net5733));
 sg13g2_o21ai_1 _20505_ (.B1(_05782_),
    .Y(_01559_),
    .A1(net4879),
    .A2(net5733));
 sg13g2_nand2_1 _20506_ (.Y(_05783_),
    .A(net686),
    .B(net5734));
 sg13g2_o21ai_1 _20507_ (.B1(_05783_),
    .Y(_01560_),
    .A1(net4872),
    .A2(net5734));
 sg13g2_nand2_1 _20508_ (.Y(_05784_),
    .A(net699),
    .B(net5735));
 sg13g2_o21ai_1 _20509_ (.B1(_05784_),
    .Y(_01561_),
    .A1(net4766),
    .A2(net5735));
 sg13g2_nand2_1 _20510_ (.Y(_05785_),
    .A(net539),
    .B(net5728));
 sg13g2_o21ai_1 _20511_ (.B1(_05785_),
    .Y(_01562_),
    .A1(net4868),
    .A2(net5728));
 sg13g2_nand2_1 _20512_ (.Y(_05786_),
    .A(net740),
    .B(net5736));
 sg13g2_o21ai_1 _20513_ (.B1(_05786_),
    .Y(_01563_),
    .A1(net4865),
    .A2(net5735));
 sg13g2_nand2_1 _20514_ (.Y(_05787_),
    .A(net372),
    .B(net5728));
 sg13g2_o21ai_1 _20515_ (.B1(_05787_),
    .Y(_01564_),
    .A1(net4858),
    .A2(net5728));
 sg13g2_nand2_1 _20516_ (.Y(_05788_),
    .A(net913),
    .B(net5727));
 sg13g2_o21ai_1 _20517_ (.B1(_05788_),
    .Y(_01565_),
    .A1(net4854),
    .A2(net5727));
 sg13g2_nand2_1 _20518_ (.Y(_05789_),
    .A(net755),
    .B(net5733));
 sg13g2_o21ai_1 _20519_ (.B1(_05789_),
    .Y(_01566_),
    .A1(net4848),
    .A2(net5733));
 sg13g2_nand2_1 _20520_ (.Y(_05790_),
    .A(net923),
    .B(net5727));
 sg13g2_o21ai_1 _20521_ (.B1(_05790_),
    .Y(_01567_),
    .A1(net4846),
    .A2(net5727));
 sg13g2_nand2_1 _20522_ (.Y(_05791_),
    .A(net1150),
    .B(net5728));
 sg13g2_o21ai_1 _20523_ (.B1(_05791_),
    .Y(_01568_),
    .A1(net4840),
    .A2(net5731));
 sg13g2_nand2_1 _20524_ (.Y(_05792_),
    .A(net837),
    .B(net5730));
 sg13g2_o21ai_1 _20525_ (.B1(_05792_),
    .Y(_01569_),
    .A1(net4836),
    .A2(net5729));
 sg13g2_nand2_1 _20526_ (.Y(_05793_),
    .A(net1294),
    .B(net5734));
 sg13g2_o21ai_1 _20527_ (.B1(_05793_),
    .Y(_01570_),
    .A1(net4829),
    .A2(net5734));
 sg13g2_nand2_1 _20528_ (.Y(_05794_),
    .A(net920),
    .B(net5734));
 sg13g2_o21ai_1 _20529_ (.B1(_05794_),
    .Y(_01571_),
    .A1(net4823),
    .A2(net5734));
 sg13g2_nand3_1 _20530_ (.B(_05625_),
    .C(_05728_),
    .A(net6096),
    .Y(_05795_));
 sg13g2_nand2_1 _20531_ (.Y(_05796_),
    .A(net954),
    .B(net5718));
 sg13g2_o21ai_1 _20532_ (.B1(_05796_),
    .Y(_01572_),
    .A1(net4994),
    .A2(net5718));
 sg13g2_nand2_1 _20533_ (.Y(_05797_),
    .A(net1257),
    .B(net5718));
 sg13g2_o21ai_1 _20534_ (.B1(_05797_),
    .Y(_01573_),
    .A1(net4989),
    .A2(net5718));
 sg13g2_nand2_1 _20535_ (.Y(_05798_),
    .A(net1239),
    .B(net5718));
 sg13g2_o21ai_1 _20536_ (.B1(_05798_),
    .Y(_01574_),
    .A1(net4984),
    .A2(net5718));
 sg13g2_nand2_1 _20537_ (.Y(_05799_),
    .A(net660),
    .B(net5717));
 sg13g2_o21ai_1 _20538_ (.B1(_05799_),
    .Y(_01575_),
    .A1(net4980),
    .A2(net5716));
 sg13g2_nand2_1 _20539_ (.Y(_05800_),
    .A(net910),
    .B(net5722));
 sg13g2_o21ai_1 _20540_ (.B1(_05800_),
    .Y(_01576_),
    .A1(net4976),
    .A2(net5722));
 sg13g2_nand2_1 _20541_ (.Y(_05801_),
    .A(net959),
    .B(net5722));
 sg13g2_o21ai_1 _20542_ (.B1(_05801_),
    .Y(_01577_),
    .A1(net4971),
    .A2(net5722));
 sg13g2_nand2_1 _20543_ (.Y(_05802_),
    .A(net410),
    .B(net5718));
 sg13g2_o21ai_1 _20544_ (.B1(_05802_),
    .Y(_01578_),
    .A1(net4966),
    .A2(net5718));
 sg13g2_nand2_1 _20545_ (.Y(_05803_),
    .A(net591),
    .B(net5721));
 sg13g2_o21ai_1 _20546_ (.B1(_05803_),
    .Y(_01579_),
    .A1(net4919),
    .A2(net5721));
 sg13g2_nand2_1 _20547_ (.Y(_05804_),
    .A(net1138),
    .B(net5722));
 sg13g2_o21ai_1 _20548_ (.B1(_05804_),
    .Y(_01580_),
    .A1(net4782),
    .A2(net5722));
 sg13g2_nand2_1 _20549_ (.Y(_05805_),
    .A(net831),
    .B(net5723));
 sg13g2_o21ai_1 _20550_ (.B1(_05805_),
    .Y(_01581_),
    .A1(net4911),
    .A2(net5723));
 sg13g2_nand2_1 _20551_ (.Y(_05806_),
    .A(net1038),
    .B(net5725));
 sg13g2_o21ai_1 _20552_ (.B1(_05806_),
    .Y(_01582_),
    .A1(net4905),
    .A2(net5725));
 sg13g2_nand2_1 _20553_ (.Y(_05807_),
    .A(net971),
    .B(net5719));
 sg13g2_o21ai_1 _20554_ (.B1(_05807_),
    .Y(_01583_),
    .A1(net4775),
    .A2(net5719));
 sg13g2_nand2_1 _20555_ (.Y(_05808_),
    .A(net894),
    .B(net5720));
 sg13g2_o21ai_1 _20556_ (.B1(_05808_),
    .Y(_01584_),
    .A1(net4900),
    .A2(net5725));
 sg13g2_nand2_1 _20557_ (.Y(_05809_),
    .A(net1124),
    .B(net5720));
 sg13g2_o21ai_1 _20558_ (.B1(_05809_),
    .Y(_01585_),
    .A1(net4960),
    .A2(net5720));
 sg13g2_nand2_1 _20559_ (.Y(_05810_),
    .A(net779),
    .B(net5716));
 sg13g2_o21ai_1 _20560_ (.B1(_05810_),
    .Y(_01586_),
    .A1(net4954),
    .A2(net5716));
 sg13g2_nand2_1 _20561_ (.Y(_05811_),
    .A(net780),
    .B(net5725));
 sg13g2_o21ai_1 _20562_ (.B1(_05811_),
    .Y(_01587_),
    .A1(net4898),
    .A2(net5725));
 sg13g2_nand2_1 _20563_ (.Y(_05812_),
    .A(net668),
    .B(net5720));
 sg13g2_o21ai_1 _20564_ (.B1(_05812_),
    .Y(_01588_),
    .A1(net4891),
    .A2(net5720));
 sg13g2_nand2_1 _20565_ (.Y(_05813_),
    .A(net629),
    .B(net5717));
 sg13g2_o21ai_1 _20566_ (.B1(_05813_),
    .Y(_01589_),
    .A1(net4885),
    .A2(net5717));
 sg13g2_nand2_1 _20567_ (.Y(_05814_),
    .A(net1113),
    .B(net5720));
 sg13g2_o21ai_1 _20568_ (.B1(_05814_),
    .Y(_01590_),
    .A1(net4768),
    .A2(net5720));
 sg13g2_nand2_1 _20569_ (.Y(_05815_),
    .A(net1059),
    .B(net5721));
 sg13g2_o21ai_1 _20570_ (.B1(_05815_),
    .Y(_01591_),
    .A1(net4879),
    .A2(net5721));
 sg13g2_nand2_1 _20571_ (.Y(_05816_),
    .A(net696),
    .B(net5724));
 sg13g2_o21ai_1 _20572_ (.B1(_05816_),
    .Y(_01592_),
    .A1(net4872),
    .A2(net5724));
 sg13g2_nand2_1 _20573_ (.Y(_05817_),
    .A(net1371),
    .B(net5723));
 sg13g2_o21ai_1 _20574_ (.B1(_05817_),
    .Y(_01593_),
    .A1(net4765),
    .A2(net5723));
 sg13g2_nand2_1 _20575_ (.Y(_05818_),
    .A(net1241),
    .B(net5716));
 sg13g2_o21ai_1 _20576_ (.B1(_05818_),
    .Y(_01594_),
    .A1(net4867),
    .A2(net5716));
 sg13g2_nand2_1 _20577_ (.Y(_05819_),
    .A(net828),
    .B(net5724));
 sg13g2_o21ai_1 _20578_ (.B1(_05819_),
    .Y(_01595_),
    .A1(net4865),
    .A2(net5724));
 sg13g2_nand2_1 _20579_ (.Y(_05820_),
    .A(net753),
    .B(net5717));
 sg13g2_o21ai_1 _20580_ (.B1(_05820_),
    .Y(_01596_),
    .A1(net4857),
    .A2(net5717));
 sg13g2_nand2_1 _20581_ (.Y(_05821_),
    .A(net882),
    .B(net5716));
 sg13g2_o21ai_1 _20582_ (.B1(_05821_),
    .Y(_01597_),
    .A1(net4853),
    .A2(net5716));
 sg13g2_nand2_1 _20583_ (.Y(_05822_),
    .A(net1267),
    .B(net5720));
 sg13g2_o21ai_1 _20584_ (.B1(_05822_),
    .Y(_01598_),
    .A1(net4847),
    .A2(net5721));
 sg13g2_nand2_1 _20585_ (.Y(_05823_),
    .A(net1151),
    .B(net5716));
 sg13g2_o21ai_1 _20586_ (.B1(_05823_),
    .Y(_01599_),
    .A1(net4844),
    .A2(net5717));
 sg13g2_nand2_1 _20587_ (.Y(_05824_),
    .A(net547),
    .B(net5721));
 sg13g2_o21ai_1 _20588_ (.B1(_05824_),
    .Y(_01600_),
    .A1(net4839),
    .A2(net5721));
 sg13g2_nand2_1 _20589_ (.Y(_05825_),
    .A(net585),
    .B(net5719));
 sg13g2_o21ai_1 _20590_ (.B1(_05825_),
    .Y(_01601_),
    .A1(net4832),
    .A2(net5719));
 sg13g2_nand2_1 _20591_ (.Y(_05826_),
    .A(net759),
    .B(net5724));
 sg13g2_o21ai_1 _20592_ (.B1(_05826_),
    .Y(_01602_),
    .A1(net4830),
    .A2(net5724));
 sg13g2_nand2_1 _20593_ (.Y(_05827_),
    .A(net752),
    .B(net5722));
 sg13g2_o21ai_1 _20594_ (.B1(_05827_),
    .Y(_01603_),
    .A1(net4826),
    .A2(net5722));
 sg13g2_nor4_2 _20595_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .C(_09505_),
    .Y(_05828_),
    .D(_09508_));
 sg13g2_nor2_1 _20596_ (.A(net1187),
    .B(net5708),
    .Y(_05829_));
 sg13g2_a21oi_1 _20597_ (.A1(net4995),
    .A2(net5708),
    .Y(_01604_),
    .B1(_05829_));
 sg13g2_nor2_1 _20598_ (.A(net2440),
    .B(net5708),
    .Y(_05830_));
 sg13g2_a21oi_1 _20599_ (.A1(net4990),
    .A2(net5708),
    .Y(_01605_),
    .B1(_05830_));
 sg13g2_nor2_1 _20600_ (.A(net2377),
    .B(net5708),
    .Y(_05831_));
 sg13g2_a21oi_1 _20601_ (.A1(net4984),
    .A2(net5708),
    .Y(_01606_),
    .B1(_05831_));
 sg13g2_nor2_1 _20602_ (.A(net2300),
    .B(net5706),
    .Y(_05832_));
 sg13g2_a21oi_1 _20603_ (.A1(net4980),
    .A2(net5706),
    .Y(_01607_),
    .B1(_05832_));
 sg13g2_nor2_1 _20604_ (.A(net1618),
    .B(net5712),
    .Y(_05833_));
 sg13g2_a21oi_1 _20605_ (.A1(net4975),
    .A2(net5712),
    .Y(_01608_),
    .B1(_05833_));
 sg13g2_nor2_1 _20606_ (.A(net2169),
    .B(net5714),
    .Y(_05834_));
 sg13g2_a21oi_1 _20607_ (.A1(net4969),
    .A2(net5714),
    .Y(_01609_),
    .B1(_05834_));
 sg13g2_nor2_1 _20608_ (.A(net1840),
    .B(net5708),
    .Y(_05835_));
 sg13g2_a21oi_1 _20609_ (.A1(net4967),
    .A2(net5708),
    .Y(_01610_),
    .B1(_05835_));
 sg13g2_nor2_1 _20610_ (.A(net1614),
    .B(net5711),
    .Y(_05836_));
 sg13g2_a21oi_1 _20611_ (.A1(net4916),
    .A2(net5715),
    .Y(_01611_),
    .B1(_05836_));
 sg13g2_nor2_1 _20612_ (.A(net2511),
    .B(net5709),
    .Y(_05837_));
 sg13g2_a21oi_1 _20613_ (.A1(net4782),
    .A2(net5709),
    .Y(_01612_),
    .B1(_05837_));
 sg13g2_nor2_1 _20614_ (.A(net1572),
    .B(net5714),
    .Y(_05838_));
 sg13g2_a21oi_1 _20615_ (.A1(net4915),
    .A2(net5714),
    .Y(_01613_),
    .B1(_05838_));
 sg13g2_nor2_1 _20616_ (.A(net1759),
    .B(net5713),
    .Y(_05839_));
 sg13g2_a21oi_1 _20617_ (.A1(net4907),
    .A2(net5713),
    .Y(_01614_),
    .B1(_05839_));
 sg13g2_nor2_1 _20618_ (.A(net1869),
    .B(net5709),
    .Y(_05840_));
 sg13g2_a21oi_1 _20619_ (.A1(net4775),
    .A2(net5709),
    .Y(_01615_),
    .B1(_05840_));
 sg13g2_nor2_1 _20620_ (.A(net1866),
    .B(net5711),
    .Y(_05841_));
 sg13g2_a21oi_1 _20621_ (.A1(net4900),
    .A2(net5711),
    .Y(_01616_),
    .B1(_05841_));
 sg13g2_nor2_1 _20622_ (.A(net1276),
    .B(net5711),
    .Y(_05842_));
 sg13g2_a21oi_1 _20623_ (.A1(net4961),
    .A2(net5711),
    .Y(_01617_),
    .B1(_05842_));
 sg13g2_nor2_1 _20624_ (.A(net1878),
    .B(net5706),
    .Y(_05843_));
 sg13g2_a21oi_1 _20625_ (.A1(net4954),
    .A2(net5706),
    .Y(_01618_),
    .B1(_05843_));
 sg13g2_nor2_1 _20626_ (.A(net1693),
    .B(net5715),
    .Y(_05844_));
 sg13g2_a21oi_1 _20627_ (.A1(net4896),
    .A2(net5711),
    .Y(_01619_),
    .B1(_05844_));
 sg13g2_nor2_1 _20628_ (.A(net1390),
    .B(net5712),
    .Y(_05845_));
 sg13g2_a21oi_1 _20629_ (.A1(net4892),
    .A2(net5712),
    .Y(_01620_),
    .B1(_05845_));
 sg13g2_nor2_1 _20630_ (.A(net1574),
    .B(net5707),
    .Y(_05846_));
 sg13g2_a21oi_1 _20631_ (.A1(net4886),
    .A2(net5707),
    .Y(_01621_),
    .B1(_05846_));
 sg13g2_nor2_1 _20632_ (.A(net2187),
    .B(net5711),
    .Y(_05847_));
 sg13g2_a21oi_1 _20633_ (.A1(net4769),
    .A2(net5711),
    .Y(_01622_),
    .B1(_05847_));
 sg13g2_nor2_1 _20634_ (.A(net1984),
    .B(net5712),
    .Y(_05848_));
 sg13g2_a21oi_1 _20635_ (.A1(net4881),
    .A2(net5712),
    .Y(_01623_),
    .B1(_05848_));
 sg13g2_nor2_1 _20636_ (.A(net1579),
    .B(net5713),
    .Y(_05849_));
 sg13g2_a21oi_1 _20637_ (.A1(net4874),
    .A2(net5713),
    .Y(_01624_),
    .B1(_05849_));
 sg13g2_nor2_1 _20638_ (.A(net1432),
    .B(net5714),
    .Y(_05850_));
 sg13g2_a21oi_1 _20639_ (.A1(net4764),
    .A2(net5714),
    .Y(_01625_),
    .B1(_05850_));
 sg13g2_nor2_1 _20640_ (.A(net1408),
    .B(net5706),
    .Y(_05851_));
 sg13g2_a21oi_1 _20641_ (.A1(net4869),
    .A2(net5706),
    .Y(_01626_),
    .B1(_05851_));
 sg13g2_nor2_1 _20642_ (.A(net2210),
    .B(net5715),
    .Y(_05852_));
 sg13g2_a21oi_1 _20643_ (.A1(net4863),
    .A2(net5714),
    .Y(_01627_),
    .B1(_05852_));
 sg13g2_nor2_1 _20644_ (.A(net1259),
    .B(net5707),
    .Y(_05853_));
 sg13g2_a21oi_1 _20645_ (.A1(net4860),
    .A2(net5707),
    .Y(_01628_),
    .B1(_05853_));
 sg13g2_nor2_1 _20646_ (.A(net1473),
    .B(net5706),
    .Y(_05854_));
 sg13g2_a21oi_1 _20647_ (.A1(net4855),
    .A2(net5706),
    .Y(_01629_),
    .B1(_05854_));
 sg13g2_nor2_1 _20648_ (.A(net2092),
    .B(net5712),
    .Y(_05855_));
 sg13g2_a21oi_1 _20649_ (.A1(net4849),
    .A2(net5712),
    .Y(_01630_),
    .B1(_05855_));
 sg13g2_nor2_1 _20650_ (.A(net1334),
    .B(net5707),
    .Y(_05856_));
 sg13g2_a21oi_1 _20651_ (.A1(net4844),
    .A2(net5707),
    .Y(_01631_),
    .B1(_05856_));
 sg13g2_nor2_1 _20652_ (.A(net2216),
    .B(net5707),
    .Y(_05857_));
 sg13g2_a21oi_1 _20653_ (.A1(net4837),
    .A2(net5710),
    .Y(_01632_),
    .B1(_05857_));
 sg13g2_nor2_1 _20654_ (.A(net1254),
    .B(net5709),
    .Y(_05858_));
 sg13g2_a21oi_1 _20655_ (.A1(net4833),
    .A2(net5709),
    .Y(_01633_),
    .B1(_05858_));
 sg13g2_nor2_1 _20656_ (.A(net1658),
    .B(net5713),
    .Y(_05859_));
 sg13g2_a21oi_1 _20657_ (.A1(net4830),
    .A2(net5713),
    .Y(_01634_),
    .B1(_05859_));
 sg13g2_nor2_1 _20658_ (.A(net1355),
    .B(net5713),
    .Y(_05860_));
 sg13g2_a21oi_1 _20659_ (.A1(net4822),
    .A2(net5713),
    .Y(_01635_),
    .B1(_05860_));
 sg13g2_nand2_1 _20660_ (.Y(_05861_),
    .A(_05660_),
    .B(_05728_));
 sg13g2_nand3_1 _20661_ (.B(_05660_),
    .C(_05728_),
    .A(net6096),
    .Y(_05862_));
 sg13g2_nand2_1 _20662_ (.Y(_05863_),
    .A(net1008),
    .B(net5697));
 sg13g2_o21ai_1 _20663_ (.B1(_05863_),
    .Y(_01636_),
    .A1(net4998),
    .A2(net5697));
 sg13g2_nand2_1 _20664_ (.Y(_05864_),
    .A(net993),
    .B(net5697));
 sg13g2_o21ai_1 _20665_ (.B1(_05864_),
    .Y(_01637_),
    .A1(net4989),
    .A2(net5697));
 sg13g2_nand2_1 _20666_ (.Y(_05865_),
    .A(net1004),
    .B(net5697));
 sg13g2_o21ai_1 _20667_ (.B1(_05865_),
    .Y(_01638_),
    .A1(net4985),
    .A2(net5697));
 sg13g2_nand2_1 _20668_ (.Y(_05866_),
    .A(net698),
    .B(net5696));
 sg13g2_o21ai_1 _20669_ (.B1(_05866_),
    .Y(_01639_),
    .A1(net4981),
    .A2(net5696));
 sg13g2_nand2_1 _20670_ (.Y(_05867_),
    .A(net526),
    .B(net5700));
 sg13g2_o21ai_1 _20671_ (.B1(_05867_),
    .Y(_01640_),
    .A1(net4977),
    .A2(net5701));
 sg13g2_nand2_1 _20672_ (.Y(_05868_),
    .A(net1176),
    .B(net5704));
 sg13g2_o21ai_1 _20673_ (.B1(_05868_),
    .Y(_01641_),
    .A1(net4971),
    .A2(net5704));
 sg13g2_nand2_1 _20674_ (.Y(_05869_),
    .A(net1095),
    .B(net5704));
 sg13g2_o21ai_1 _20675_ (.B1(_05869_),
    .Y(_01642_),
    .A1(net4966),
    .A2(net5697));
 sg13g2_nand2_1 _20676_ (.Y(_05870_),
    .A(net450),
    .B(net5701));
 sg13g2_o21ai_1 _20677_ (.B1(_05870_),
    .Y(_01643_),
    .A1(net4919),
    .A2(net5701));
 sg13g2_nand2_1 _20678_ (.Y(_05871_),
    .A(net845),
    .B(net5697));
 sg13g2_o21ai_1 _20679_ (.B1(_05871_),
    .Y(_01644_),
    .A1(net4779),
    .A2(net5698));
 sg13g2_nand2_1 _20680_ (.Y(_05872_),
    .A(net840),
    .B(net5704));
 sg13g2_o21ai_1 _20681_ (.B1(_05872_),
    .Y(_01645_),
    .A1(net4911),
    .A2(net5704));
 sg13g2_nand2_1 _20682_ (.Y(_05873_),
    .A(net877),
    .B(net5703));
 sg13g2_o21ai_1 _20683_ (.B1(_05873_),
    .Y(_01646_),
    .A1(net4909),
    .A2(net5703));
 sg13g2_nand2_1 _20684_ (.Y(_05874_),
    .A(net836),
    .B(net5698));
 sg13g2_o21ai_1 _20685_ (.B1(_05874_),
    .Y(_01647_),
    .A1(net4773),
    .A2(net5698));
 sg13g2_nand2_1 _20686_ (.Y(_05875_),
    .A(net984),
    .B(net5701));
 sg13g2_o21ai_1 _20687_ (.B1(_05875_),
    .Y(_01648_),
    .A1(net4899),
    .A2(net5701));
 sg13g2_nand2_1 _20688_ (.Y(_05876_),
    .A(net1211),
    .B(net5702));
 sg13g2_o21ai_1 _20689_ (.B1(_05876_),
    .Y(_01649_),
    .A1(net4963),
    .A2(net5702));
 sg13g2_nand2_1 _20690_ (.Y(_05877_),
    .A(net955),
    .B(net5695));
 sg13g2_o21ai_1 _20691_ (.B1(_05877_),
    .Y(_01650_),
    .A1(net4954),
    .A2(net5695));
 sg13g2_nand2_1 _20692_ (.Y(_05878_),
    .A(net932),
    .B(net5701));
 sg13g2_o21ai_1 _20693_ (.B1(_05878_),
    .Y(_01651_),
    .A1(net4896),
    .A2(net5701));
 sg13g2_nand2_1 _20694_ (.Y(_05879_),
    .A(net1154),
    .B(net5700));
 sg13g2_o21ai_1 _20695_ (.B1(_05879_),
    .Y(_01652_),
    .A1(net4889),
    .A2(net5700));
 sg13g2_nand2_1 _20696_ (.Y(_05880_),
    .A(net460),
    .B(net5696));
 sg13g2_o21ai_1 _20697_ (.B1(_05880_),
    .Y(_01653_),
    .A1(net4885),
    .A2(net5696));
 sg13g2_nand2_1 _20698_ (.Y(_05881_),
    .A(net869),
    .B(net5702));
 sg13g2_o21ai_1 _20699_ (.B1(_05881_),
    .Y(_01654_),
    .A1(net4770),
    .A2(net5702));
 sg13g2_nand2_1 _20700_ (.Y(_05882_),
    .A(net793),
    .B(net5700));
 sg13g2_o21ai_1 _20701_ (.B1(_05882_),
    .Y(_01655_),
    .A1(net4878),
    .A2(net5700));
 sg13g2_nand2_1 _20702_ (.Y(_05883_),
    .A(net411),
    .B(net5703));
 sg13g2_o21ai_1 _20703_ (.B1(_05883_),
    .Y(_01656_),
    .A1(net4873),
    .A2(net5703));
 sg13g2_nand2_1 _20704_ (.Y(_05884_),
    .A(net1517),
    .B(net5704));
 sg13g2_o21ai_1 _20705_ (.B1(_05884_),
    .Y(_01657_),
    .A1(net4762),
    .A2(net5704));
 sg13g2_nand2_1 _20706_ (.Y(_05885_),
    .A(net970),
    .B(net5695));
 sg13g2_o21ai_1 _20707_ (.B1(_05885_),
    .Y(_01658_),
    .A1(net4867),
    .A2(net5695));
 sg13g2_nand2_1 _20708_ (.Y(_05886_),
    .A(net960),
    .B(net5703));
 sg13g2_o21ai_1 _20709_ (.B1(_05886_),
    .Y(_01659_),
    .A1(net4865),
    .A2(net5703));
 sg13g2_nand2_1 _20710_ (.Y(_05887_),
    .A(net801),
    .B(net5696));
 sg13g2_o21ai_1 _20711_ (.B1(_05887_),
    .Y(_01660_),
    .A1(net4859),
    .A2(net5696));
 sg13g2_nand2_1 _20712_ (.Y(_05888_),
    .A(net875),
    .B(net5695));
 sg13g2_o21ai_1 _20713_ (.B1(_05888_),
    .Y(_01661_),
    .A1(net4852),
    .A2(net5695));
 sg13g2_nand2_1 _20714_ (.Y(_05889_),
    .A(net1112),
    .B(net5700));
 sg13g2_o21ai_1 _20715_ (.B1(_05889_),
    .Y(_01662_),
    .A1(net4848),
    .A2(net5700));
 sg13g2_nand2_1 _20716_ (.Y(_05890_),
    .A(net1288),
    .B(net5695));
 sg13g2_o21ai_1 _20717_ (.B1(_05890_),
    .Y(_01663_),
    .A1(net4846),
    .A2(net5695));
 sg13g2_nand2_1 _20718_ (.Y(_05891_),
    .A(net1235),
    .B(net5700));
 sg13g2_o21ai_1 _20719_ (.B1(_05891_),
    .Y(_01664_),
    .A1(net4839),
    .A2(net5696));
 sg13g2_nand2_1 _20720_ (.Y(_05892_),
    .A(net1128),
    .B(net5698));
 sg13g2_o21ai_1 _20721_ (.B1(_05892_),
    .Y(_01665_),
    .A1(net4835),
    .A2(net5698));
 sg13g2_nand2_1 _20722_ (.Y(_05893_),
    .A(net817),
    .B(net5705));
 sg13g2_o21ai_1 _20723_ (.B1(_05893_),
    .Y(_01666_),
    .A1(net4830),
    .A2(net5705));
 sg13g2_nand2_1 _20724_ (.Y(_05894_),
    .A(net961),
    .B(net5703));
 sg13g2_o21ai_1 _20725_ (.B1(_05894_),
    .Y(_01667_),
    .A1(net4824),
    .A2(net5703));
 sg13g2_nor2b_2 _20726_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[4] ),
    .B_N(\soc_inst.cpu_core.mem_reg_we ),
    .Y(_05895_));
 sg13g2_nand2_2 _20727_ (.Y(_05896_),
    .A(_05861_),
    .B(net6070));
 sg13g2_nand4_1 _20728_ (.B(net6216),
    .C(_09507_),
    .A(net6214),
    .Y(_05897_),
    .D(net6071));
 sg13g2_nand2_1 _20729_ (.Y(_05898_),
    .A(net863),
    .B(net5413));
 sg13g2_o21ai_1 _20730_ (.B1(_05898_),
    .Y(_01668_),
    .A1(net4996),
    .A2(net5413));
 sg13g2_nand2_1 _20731_ (.Y(_05899_),
    .A(net982),
    .B(net5413));
 sg13g2_o21ai_1 _20732_ (.B1(_05899_),
    .Y(_01669_),
    .A1(net4992),
    .A2(net5413));
 sg13g2_nand2_1 _20733_ (.Y(_05900_),
    .A(net1011),
    .B(net5413));
 sg13g2_o21ai_1 _20734_ (.B1(_05900_),
    .Y(_01670_),
    .A1(net4986),
    .A2(net5413));
 sg13g2_nand2_1 _20735_ (.Y(_05901_),
    .A(net480),
    .B(net5411));
 sg13g2_o21ai_1 _20736_ (.B1(_05901_),
    .Y(_01671_),
    .A1(net4981),
    .A2(net5411));
 sg13g2_nand2_1 _20737_ (.Y(_05902_),
    .A(net1360),
    .B(net5416));
 sg13g2_o21ai_1 _20738_ (.B1(_05902_),
    .Y(_01672_),
    .A1(net4975),
    .A2(net5416));
 sg13g2_nand2_1 _20739_ (.Y(_05903_),
    .A(net570),
    .B(net5418));
 sg13g2_o21ai_1 _20740_ (.B1(_05903_),
    .Y(_01673_),
    .A1(net4971),
    .A2(net5418));
 sg13g2_nand2_1 _20741_ (.Y(_05904_),
    .A(net947),
    .B(net5414));
 sg13g2_o21ai_1 _20742_ (.B1(_05904_),
    .Y(_01674_),
    .A1(net4964),
    .A2(net5414));
 sg13g2_nand2_1 _20743_ (.Y(_05905_),
    .A(net958),
    .B(net5417));
 sg13g2_o21ai_1 _20744_ (.B1(_05905_),
    .Y(_01675_),
    .A1(net4918),
    .A2(net5417));
 sg13g2_nand2_1 _20745_ (.Y(_05906_),
    .A(net1102),
    .B(net5413));
 sg13g2_o21ai_1 _20746_ (.B1(_05906_),
    .Y(_01676_),
    .A1(net4780),
    .A2(net5413));
 sg13g2_nand2_1 _20747_ (.Y(_05907_),
    .A(net804),
    .B(net5418));
 sg13g2_o21ai_1 _20748_ (.B1(_05907_),
    .Y(_01677_),
    .A1(net4911),
    .A2(net5418));
 sg13g2_nand2_1 _20749_ (.Y(_05908_),
    .A(net646),
    .B(net5419));
 sg13g2_o21ai_1 _20750_ (.B1(_05908_),
    .Y(_01678_),
    .A1(net4908),
    .A2(net5419));
 sg13g2_nand2_1 _20751_ (.Y(_05909_),
    .A(net485),
    .B(net5414));
 sg13g2_o21ai_1 _20752_ (.B1(_05909_),
    .Y(_01679_),
    .A1(net4773),
    .A2(net5414));
 sg13g2_nand2_1 _20753_ (.Y(_05910_),
    .A(net1046),
    .B(net5417));
 sg13g2_o21ai_1 _20754_ (.B1(_05910_),
    .Y(_01680_),
    .A1(net4901),
    .A2(net5417));
 sg13g2_nand2_1 _20755_ (.Y(_05911_),
    .A(net1204),
    .B(net5417));
 sg13g2_o21ai_1 _20756_ (.B1(_05911_),
    .Y(_01681_),
    .A1(net4961),
    .A2(net5420));
 sg13g2_nand2_1 _20757_ (.Y(_05912_),
    .A(net579),
    .B(net5411));
 sg13g2_o21ai_1 _20758_ (.B1(_05912_),
    .Y(_01682_),
    .A1(net4957),
    .A2(net5411));
 sg13g2_nand2_1 _20759_ (.Y(_05913_),
    .A(net610),
    .B(net5417));
 sg13g2_o21ai_1 _20760_ (.B1(_05913_),
    .Y(_01683_),
    .A1(net4895),
    .A2(net5417));
 sg13g2_nand2_1 _20761_ (.Y(_05914_),
    .A(net1258),
    .B(net5416));
 sg13g2_o21ai_1 _20762_ (.B1(_05914_),
    .Y(_01684_),
    .A1(net4889),
    .A2(net5416));
 sg13g2_nand2_1 _20763_ (.Y(_05915_),
    .A(net474),
    .B(net5412));
 sg13g2_o21ai_1 _20764_ (.B1(_05915_),
    .Y(_01685_),
    .A1(net4885),
    .A2(net5412));
 sg13g2_nand2_1 _20765_ (.Y(_05916_),
    .A(net1073),
    .B(net5420));
 sg13g2_o21ai_1 _20766_ (.B1(_05916_),
    .Y(_01686_),
    .A1(net4770),
    .A2(net5420));
 sg13g2_nand2_1 _20767_ (.Y(_05917_),
    .A(net1092),
    .B(net5416));
 sg13g2_o21ai_1 _20768_ (.B1(_05917_),
    .Y(_01687_),
    .A1(net4879),
    .A2(net5416));
 sg13g2_nand2_1 _20769_ (.Y(_05918_),
    .A(net973),
    .B(net5419));
 sg13g2_o21ai_1 _20770_ (.B1(_05918_),
    .Y(_01688_),
    .A1(net4874),
    .A2(net5419));
 sg13g2_nand2_1 _20771_ (.Y(_05919_),
    .A(net362),
    .B(net5418));
 sg13g2_o21ai_1 _20772_ (.B1(_05919_),
    .Y(_01689_),
    .A1(net4765),
    .A2(net5418));
 sg13g2_nand2_1 _20773_ (.Y(_05920_),
    .A(net648),
    .B(net5412));
 sg13g2_o21ai_1 _20774_ (.B1(_05920_),
    .Y(_01690_),
    .A1(net4869),
    .A2(net5412));
 sg13g2_nand2_1 _20775_ (.Y(_05921_),
    .A(net1247),
    .B(net5419));
 sg13g2_o21ai_1 _20776_ (.B1(_05921_),
    .Y(_01691_),
    .A1(net4864),
    .A2(net5419));
 sg13g2_nand2_1 _20777_ (.Y(_05922_),
    .A(net963),
    .B(net5412));
 sg13g2_o21ai_1 _20778_ (.B1(_05922_),
    .Y(_01692_),
    .A1(net4858),
    .A2(net5412));
 sg13g2_nand2_1 _20779_ (.Y(_05923_),
    .A(net967),
    .B(net5411));
 sg13g2_o21ai_1 _20780_ (.B1(_05923_),
    .Y(_01693_),
    .A1(net4855),
    .A2(net5411));
 sg13g2_nand2_1 _20781_ (.Y(_05924_),
    .A(net1651),
    .B(net5416));
 sg13g2_o21ai_1 _20782_ (.B1(_05924_),
    .Y(_01694_),
    .A1(net4848),
    .A2(net5416));
 sg13g2_nand2_1 _20783_ (.Y(_05925_),
    .A(net544),
    .B(net5411));
 sg13g2_o21ai_1 _20784_ (.B1(_05925_),
    .Y(_01695_),
    .A1(net4842),
    .A2(net5411));
 sg13g2_nand2_1 _20785_ (.Y(_05926_),
    .A(net589),
    .B(net5412));
 sg13g2_o21ai_1 _20786_ (.B1(_05926_),
    .Y(_01696_),
    .A1(net4839),
    .A2(net5415));
 sg13g2_nand2_1 _20787_ (.Y(_05927_),
    .A(net538),
    .B(net5414));
 sg13g2_o21ai_1 _20788_ (.B1(_05927_),
    .Y(_01697_),
    .A1(net4833),
    .A2(net5414));
 sg13g2_nand2_1 _20789_ (.Y(_05928_),
    .A(net1012),
    .B(net5419));
 sg13g2_o21ai_1 _20790_ (.B1(_05928_),
    .Y(_01698_),
    .A1(net4830),
    .A2(net5419));
 sg13g2_nand2_1 _20791_ (.Y(_05929_),
    .A(net532),
    .B(net5418));
 sg13g2_o21ai_1 _20792_ (.B1(_05929_),
    .Y(_01699_),
    .A1(net4826),
    .A2(net5418));
 sg13g2_nand3_1 _20793_ (.B(_05660_),
    .C(_05694_),
    .A(net6096),
    .Y(_05930_));
 sg13g2_nand2_1 _20794_ (.Y(_05931_),
    .A(net818),
    .B(net5687));
 sg13g2_o21ai_1 _20795_ (.B1(_05931_),
    .Y(_01700_),
    .A1(net4995),
    .A2(net5687));
 sg13g2_nand2_1 _20796_ (.Y(_05932_),
    .A(net1005),
    .B(net5687));
 sg13g2_o21ai_1 _20797_ (.B1(_05932_),
    .Y(_01701_),
    .A1(net4990),
    .A2(net5687));
 sg13g2_nand2_1 _20798_ (.Y(_05933_),
    .A(net625),
    .B(net5687));
 sg13g2_o21ai_1 _20799_ (.B1(_05933_),
    .Y(_01702_),
    .A1(net4987),
    .A2(net5687));
 sg13g2_nand2_1 _20800_ (.Y(_05934_),
    .A(net900),
    .B(net5685));
 sg13g2_o21ai_1 _20801_ (.B1(_05934_),
    .Y(_01703_),
    .A1(net4979),
    .A2(net5685));
 sg13g2_nand2_1 _20802_ (.Y(_05935_),
    .A(net975),
    .B(net5693));
 sg13g2_o21ai_1 _20803_ (.B1(_05935_),
    .Y(_01704_),
    .A1(net4978),
    .A2(net5686));
 sg13g2_nand2_1 _20804_ (.Y(_05936_),
    .A(net654),
    .B(net5693));
 sg13g2_o21ai_1 _20805_ (.B1(_05936_),
    .Y(_01705_),
    .A1(net4971),
    .A2(net5693));
 sg13g2_nand2_1 _20806_ (.Y(_05937_),
    .A(net846),
    .B(net5687));
 sg13g2_o21ai_1 _20807_ (.B1(_05937_),
    .Y(_01706_),
    .A1(net4968),
    .A2(net5688));
 sg13g2_nand2_1 _20808_ (.Y(_05938_),
    .A(net506),
    .B(net5691));
 sg13g2_o21ai_1 _20809_ (.B1(_05938_),
    .Y(_01707_),
    .A1(net4919),
    .A2(net5691));
 sg13g2_nand2_1 _20810_ (.Y(_05939_),
    .A(net996),
    .B(net5687));
 sg13g2_o21ai_1 _20811_ (.B1(_05939_),
    .Y(_01708_),
    .A1(net4781),
    .A2(net5688));
 sg13g2_nand2_1 _20812_ (.Y(_05940_),
    .A(net682),
    .B(net5692));
 sg13g2_o21ai_1 _20813_ (.B1(_05940_),
    .Y(_01709_),
    .A1(net4913),
    .A2(net5693));
 sg13g2_nand2_1 _20814_ (.Y(_05941_),
    .A(net439),
    .B(net5692));
 sg13g2_o21ai_1 _20815_ (.B1(_05941_),
    .Y(_01710_),
    .A1(net4906),
    .A2(net5692));
 sg13g2_nand2_1 _20816_ (.Y(_05942_),
    .A(net412),
    .B(net5688));
 sg13g2_o21ai_1 _20817_ (.B1(_05942_),
    .Y(_01711_),
    .A1(net4773),
    .A2(net5688));
 sg13g2_nand2_1 _20818_ (.Y(_05943_),
    .A(net600),
    .B(net5690));
 sg13g2_o21ai_1 _20819_ (.B1(_05943_),
    .Y(_01712_),
    .A1(net4904),
    .A2(net5690));
 sg13g2_nand2_1 _20820_ (.Y(_05944_),
    .A(net893),
    .B(net5690));
 sg13g2_o21ai_1 _20821_ (.B1(_05944_),
    .Y(_01713_),
    .A1(net4959),
    .A2(net5690));
 sg13g2_nand2_1 _20822_ (.Y(_05945_),
    .A(net608),
    .B(net5685));
 sg13g2_o21ai_1 _20823_ (.B1(_05945_),
    .Y(_01714_),
    .A1(net4956),
    .A2(net5685));
 sg13g2_nand2_1 _20824_ (.Y(_05946_),
    .A(net1155),
    .B(net5694));
 sg13g2_o21ai_1 _20825_ (.B1(_05946_),
    .Y(_01715_),
    .A1(net4897),
    .A2(net5691));
 sg13g2_nand2_1 _20826_ (.Y(_05947_),
    .A(net631),
    .B(net5690));
 sg13g2_o21ai_1 _20827_ (.B1(_05947_),
    .Y(_01716_),
    .A1(net4891),
    .A2(net5690));
 sg13g2_nand2_1 _20828_ (.Y(_05948_),
    .A(net953),
    .B(net5686));
 sg13g2_o21ai_1 _20829_ (.B1(_05948_),
    .Y(_01717_),
    .A1(net4885),
    .A2(net5686));
 sg13g2_nand2_1 _20830_ (.Y(_05949_),
    .A(net1098),
    .B(net5690));
 sg13g2_o21ai_1 _20831_ (.B1(_05949_),
    .Y(_01718_),
    .A1(net4768),
    .A2(net5690));
 sg13g2_nand2_1 _20832_ (.Y(_05950_),
    .A(net669),
    .B(net5691));
 sg13g2_o21ai_1 _20833_ (.B1(_05950_),
    .Y(_01719_),
    .A1(net4878),
    .A2(net5691));
 sg13g2_nand2_1 _20834_ (.Y(_05951_),
    .A(net1007),
    .B(net5692));
 sg13g2_o21ai_1 _20835_ (.B1(_05951_),
    .Y(_01720_),
    .A1(net4872),
    .A2(net5692));
 sg13g2_nand2_1 _20836_ (.Y(_05952_),
    .A(net933),
    .B(net5693));
 sg13g2_o21ai_1 _20837_ (.B1(_05952_),
    .Y(_01721_),
    .A1(net4764),
    .A2(net5693));
 sg13g2_nand2_1 _20838_ (.Y(_05953_),
    .A(net1213),
    .B(net5686));
 sg13g2_o21ai_1 _20839_ (.B1(_05953_),
    .Y(_01722_),
    .A1(net4871),
    .A2(net5686));
 sg13g2_nand2_1 _20840_ (.Y(_05954_),
    .A(net685),
    .B(net5694));
 sg13g2_o21ai_1 _20841_ (.B1(_05954_),
    .Y(_01723_),
    .A1(net4866),
    .A2(net5693));
 sg13g2_nand2_1 _20842_ (.Y(_05955_),
    .A(net475),
    .B(net5686));
 sg13g2_o21ai_1 _20843_ (.B1(_05955_),
    .Y(_01724_),
    .A1(net4861),
    .A2(net5686));
 sg13g2_nand2_1 _20844_ (.Y(_05956_),
    .A(net653),
    .B(net5685));
 sg13g2_o21ai_1 _20845_ (.B1(_05956_),
    .Y(_01725_),
    .A1(net4852),
    .A2(net5685));
 sg13g2_nand2_1 _20846_ (.Y(_05957_),
    .A(net561),
    .B(net5691));
 sg13g2_o21ai_1 _20847_ (.B1(_05957_),
    .Y(_01726_),
    .A1(net4847),
    .A2(net5691));
 sg13g2_nand2_1 _20848_ (.Y(_05958_),
    .A(net470),
    .B(net5685));
 sg13g2_o21ai_1 _20849_ (.B1(_05958_),
    .Y(_01727_),
    .A1(net4842),
    .A2(net5685));
 sg13g2_nand2_1 _20850_ (.Y(_05959_),
    .A(net1085),
    .B(net5689));
 sg13g2_o21ai_1 _20851_ (.B1(_05959_),
    .Y(_01728_),
    .A1(net4841),
    .A2(net5689));
 sg13g2_nand2_1 _20852_ (.Y(_05960_),
    .A(net743),
    .B(net5688));
 sg13g2_o21ai_1 _20853_ (.B1(_05960_),
    .Y(_01729_),
    .A1(net4832),
    .A2(net5688));
 sg13g2_nand2_1 _20854_ (.Y(_05961_),
    .A(net1164),
    .B(net5692));
 sg13g2_o21ai_1 _20855_ (.B1(_05961_),
    .Y(_01730_),
    .A1(net4829),
    .A2(net5694));
 sg13g2_nand2_1 _20856_ (.Y(_05962_),
    .A(net987),
    .B(net5692));
 sg13g2_o21ai_1 _20857_ (.B1(_05962_),
    .Y(_01731_),
    .A1(net4824),
    .A2(net5692));
 sg13g2_nand4_1 _20858_ (.B(net6216),
    .C(_05590_),
    .A(net6214),
    .Y(_05963_),
    .D(net6071));
 sg13g2_nand2_1 _20859_ (.Y(_05964_),
    .A(net422),
    .B(net5677));
 sg13g2_o21ai_1 _20860_ (.B1(_05964_),
    .Y(_01732_),
    .A1(net4996),
    .A2(net5677));
 sg13g2_nand2_1 _20861_ (.Y(_05965_),
    .A(net1048),
    .B(net5677));
 sg13g2_o21ai_1 _20862_ (.B1(_05965_),
    .Y(_01733_),
    .A1(net4992),
    .A2(net5677));
 sg13g2_nand2_1 _20863_ (.Y(_05966_),
    .A(net533),
    .B(net5677));
 sg13g2_o21ai_1 _20864_ (.B1(_05966_),
    .Y(_01734_),
    .A1(net4986),
    .A2(net5677));
 sg13g2_nand2_1 _20865_ (.Y(_05967_),
    .A(net990),
    .B(net5675));
 sg13g2_o21ai_1 _20866_ (.B1(_05967_),
    .Y(_01735_),
    .A1(net4979),
    .A2(net5675));
 sg13g2_nand2_1 _20867_ (.Y(_05968_),
    .A(net769),
    .B(net5682));
 sg13g2_o21ai_1 _20868_ (.B1(_05968_),
    .Y(_01736_),
    .A1(net4976),
    .A2(net5682));
 sg13g2_nand2_1 _20869_ (.Y(_05969_),
    .A(net700),
    .B(net5682));
 sg13g2_o21ai_1 _20870_ (.B1(_05969_),
    .Y(_01737_),
    .A1(net4970),
    .A2(net5682));
 sg13g2_nand2_1 _20871_ (.Y(_05970_),
    .A(net593),
    .B(net5677));
 sg13g2_o21ai_1 _20872_ (.B1(_05970_),
    .Y(_01738_),
    .A1(net4964),
    .A2(net5677));
 sg13g2_nand2_1 _20873_ (.Y(_05971_),
    .A(net827),
    .B(net5681));
 sg13g2_o21ai_1 _20874_ (.B1(_05971_),
    .Y(_01739_),
    .A1(net4917),
    .A2(net5681));
 sg13g2_nand2_1 _20875_ (.Y(_05972_),
    .A(net1367),
    .B(net5678));
 sg13g2_o21ai_1 _20876_ (.B1(_05972_),
    .Y(_01740_),
    .A1(net4782),
    .A2(net5678));
 sg13g2_nand2_1 _20877_ (.Y(_05973_),
    .A(net447),
    .B(net5682));
 sg13g2_o21ai_1 _20878_ (.B1(_05973_),
    .Y(_01741_),
    .A1(net4912),
    .A2(net5682));
 sg13g2_nand2_1 _20879_ (.Y(_05974_),
    .A(net1278),
    .B(net5684));
 sg13g2_o21ai_1 _20880_ (.B1(_05974_),
    .Y(_01742_),
    .A1(net4907),
    .A2(net5684));
 sg13g2_nand2_1 _20881_ (.Y(_05975_),
    .A(net719),
    .B(net5678));
 sg13g2_o21ai_1 _20882_ (.B1(_05975_),
    .Y(_01743_),
    .A1(net4773),
    .A2(net5678));
 sg13g2_nand2_1 _20883_ (.Y(_05976_),
    .A(net864),
    .B(net5680));
 sg13g2_o21ai_1 _20884_ (.B1(_05976_),
    .Y(_01744_),
    .A1(net4902),
    .A2(net5684));
 sg13g2_nand2_1 _20885_ (.Y(_05977_),
    .A(net1184),
    .B(net5680));
 sg13g2_o21ai_1 _20886_ (.B1(_05977_),
    .Y(_01745_),
    .A1(net4961),
    .A2(net5680));
 sg13g2_nand2_1 _20887_ (.Y(_05978_),
    .A(net1000),
    .B(net5675));
 sg13g2_o21ai_1 _20888_ (.B1(_05978_),
    .Y(_01746_),
    .A1(net4957),
    .A2(net5675));
 sg13g2_nand2_1 _20889_ (.Y(_05979_),
    .A(net614),
    .B(net5680));
 sg13g2_o21ai_1 _20890_ (.B1(_05979_),
    .Y(_01747_),
    .A1(net4895),
    .A2(net5681));
 sg13g2_nand2_1 _20891_ (.Y(_05980_),
    .A(net742),
    .B(net5680));
 sg13g2_o21ai_1 _20892_ (.B1(_05980_),
    .Y(_01748_),
    .A1(net4891),
    .A2(net5680));
 sg13g2_nand2_1 _20893_ (.Y(_05981_),
    .A(net672),
    .B(net5676));
 sg13g2_o21ai_1 _20894_ (.B1(_05981_),
    .Y(_01749_),
    .A1(net4884),
    .A2(net5676));
 sg13g2_nand2_1 _20895_ (.Y(_05982_),
    .A(net637),
    .B(net5680));
 sg13g2_o21ai_1 _20896_ (.B1(_05982_),
    .Y(_01750_),
    .A1(net4770),
    .A2(net5680));
 sg13g2_nand2_1 _20897_ (.Y(_05983_),
    .A(net1530),
    .B(net5681));
 sg13g2_o21ai_1 _20898_ (.B1(_05983_),
    .Y(_01751_),
    .A1(net4879),
    .A2(net5681));
 sg13g2_nand2_1 _20899_ (.Y(_05984_),
    .A(net859),
    .B(net5683));
 sg13g2_o21ai_1 _20900_ (.B1(_05984_),
    .Y(_01752_),
    .A1(net4875),
    .A2(net5683));
 sg13g2_nand2_1 _20901_ (.Y(_05985_),
    .A(net626),
    .B(net5683));
 sg13g2_o21ai_1 _20902_ (.B1(_05985_),
    .Y(_01753_),
    .A1(net4764),
    .A2(net5683));
 sg13g2_nand2_1 _20903_ (.Y(_05986_),
    .A(net657),
    .B(net5675));
 sg13g2_o21ai_1 _20904_ (.B1(_05986_),
    .Y(_01754_),
    .A1(net4870),
    .A2(net5675));
 sg13g2_nand2_1 _20905_ (.Y(_05987_),
    .A(net1175),
    .B(net5683));
 sg13g2_o21ai_1 _20906_ (.B1(_05987_),
    .Y(_01755_),
    .A1(net4863),
    .A2(net5684));
 sg13g2_nand2_1 _20907_ (.Y(_05988_),
    .A(net807),
    .B(net5679));
 sg13g2_o21ai_1 _20908_ (.B1(_05988_),
    .Y(_01756_),
    .A1(net4857),
    .A2(net5676));
 sg13g2_nand2_1 _20909_ (.Y(_05989_),
    .A(net1520),
    .B(net5675));
 sg13g2_o21ai_1 _20910_ (.B1(_05989_),
    .Y(_01757_),
    .A1(net4852),
    .A2(net5675));
 sg13g2_nand2_1 _20911_ (.Y(_05990_),
    .A(net986),
    .B(net5681));
 sg13g2_o21ai_1 _20912_ (.B1(_05990_),
    .Y(_01758_),
    .A1(net4848),
    .A2(net5681));
 sg13g2_nand2_1 _20913_ (.Y(_05991_),
    .A(net649),
    .B(net5676));
 sg13g2_o21ai_1 _20914_ (.B1(_05991_),
    .Y(_01759_),
    .A1(net4842),
    .A2(net5676));
 sg13g2_nand2_1 _20915_ (.Y(_05992_),
    .A(net806),
    .B(net5676));
 sg13g2_o21ai_1 _20916_ (.B1(_05992_),
    .Y(_01760_),
    .A1(net4838),
    .A2(net5676));
 sg13g2_nand2_1 _20917_ (.Y(_05993_),
    .A(net833),
    .B(net5678));
 sg13g2_o21ai_1 _20918_ (.B1(_05993_),
    .Y(_01761_),
    .A1(net4834),
    .A2(net5678));
 sg13g2_nand2_1 _20919_ (.Y(_05994_),
    .A(net711),
    .B(net5683));
 sg13g2_o21ai_1 _20920_ (.B1(_05994_),
    .Y(_01762_),
    .A1(net4827),
    .A2(net5683));
 sg13g2_nand2_1 _20921_ (.Y(_05995_),
    .A(net872),
    .B(net5682));
 sg13g2_o21ai_1 _20922_ (.B1(_05995_),
    .Y(_01763_),
    .A1(net4826),
    .A2(net5682));
 sg13g2_and4_1 _20923_ (.A(net6214),
    .B(net6216),
    .C(net6096),
    .D(_05625_),
    .X(_05996_));
 sg13g2_nor2_1 _20924_ (.A(net2167),
    .B(net5668),
    .Y(_05997_));
 sg13g2_a21oi_1 _20925_ (.A1(net4994),
    .A2(net5668),
    .Y(_01764_),
    .B1(_05997_));
 sg13g2_nor2_1 _20926_ (.A(net1969),
    .B(net5668),
    .Y(_05998_));
 sg13g2_a21oi_1 _20927_ (.A1(net4989),
    .A2(net5668),
    .Y(_01765_),
    .B1(_05998_));
 sg13g2_nor2_1 _20928_ (.A(net2288),
    .B(net5668),
    .Y(_05999_));
 sg13g2_a21oi_1 _20929_ (.A1(net4984),
    .A2(net5668),
    .Y(_01766_),
    .B1(_05999_));
 sg13g2_nor2_1 _20930_ (.A(net1973),
    .B(net5666),
    .Y(_06000_));
 sg13g2_a21oi_1 _20931_ (.A1(net4983),
    .A2(net5666),
    .Y(_01767_),
    .B1(_06000_));
 sg13g2_nor2_1 _20932_ (.A(net1607),
    .B(net5671),
    .Y(_06001_));
 sg13g2_a21oi_1 _20933_ (.A1(net4977),
    .A2(net5671),
    .Y(_01768_),
    .B1(_06001_));
 sg13g2_nor2_1 _20934_ (.A(net2054),
    .B(net5673),
    .Y(_06002_));
 sg13g2_a21oi_1 _20935_ (.A1(net4969),
    .A2(net5673),
    .Y(_01769_),
    .B1(_06002_));
 sg13g2_nor2_1 _20936_ (.A(net1871),
    .B(net5673),
    .Y(_06003_));
 sg13g2_a21oi_1 _20937_ (.A1(net4964),
    .A2(net5673),
    .Y(_01770_),
    .B1(_06003_));
 sg13g2_nor2_1 _20938_ (.A(net1815),
    .B(net5674),
    .Y(_06004_));
 sg13g2_a21oi_1 _20939_ (.A1(net4918),
    .A2(net5674),
    .Y(_01771_),
    .B1(_06004_));
 sg13g2_nor2_1 _20940_ (.A(net1660),
    .B(net5668),
    .Y(_06005_));
 sg13g2_a21oi_1 _20941_ (.A1(net4781),
    .A2(net5668),
    .Y(_01772_),
    .B1(_06005_));
 sg13g2_nor2_1 _20942_ (.A(net2045),
    .B(net5673),
    .Y(_06006_));
 sg13g2_a21oi_1 _20943_ (.A1(net4913),
    .A2(net5673),
    .Y(_01773_),
    .B1(_06006_));
 sg13g2_nor2_1 _20944_ (.A(net1462),
    .B(net5672),
    .Y(_06007_));
 sg13g2_a21oi_1 _20945_ (.A1(net4907),
    .A2(net5672),
    .Y(_01774_),
    .B1(_06007_));
 sg13g2_nor2_1 _20946_ (.A(net1870),
    .B(net5669),
    .Y(_06008_));
 sg13g2_a21oi_1 _20947_ (.A1(net4773),
    .A2(net5669),
    .Y(_01775_),
    .B1(_06008_));
 sg13g2_nor2_1 _20948_ (.A(net2443),
    .B(net5670),
    .Y(_06009_));
 sg13g2_a21oi_1 _20949_ (.A1(net4901),
    .A2(net5670),
    .Y(_01776_),
    .B1(_06009_));
 sg13g2_nor2_1 _20950_ (.A(net1486),
    .B(net5670),
    .Y(_06010_));
 sg13g2_a21oi_1 _20951_ (.A1(net4962),
    .A2(net5670),
    .Y(_01777_),
    .B1(_06010_));
 sg13g2_nor2_1 _20952_ (.A(net2537),
    .B(net5667),
    .Y(_06011_));
 sg13g2_a21oi_1 _20953_ (.A1(net4955),
    .A2(net5667),
    .Y(_01778_),
    .B1(_06011_));
 sg13g2_nor2_1 _20954_ (.A(net1599),
    .B(net5670),
    .Y(_06012_));
 sg13g2_a21oi_1 _20955_ (.A1(net4894),
    .A2(net5670),
    .Y(_01779_),
    .B1(_06012_));
 sg13g2_nor2_1 _20956_ (.A(net1851),
    .B(net5671),
    .Y(_06013_));
 sg13g2_a21oi_1 _20957_ (.A1(net4892),
    .A2(net5671),
    .Y(_01780_),
    .B1(_06013_));
 sg13g2_nor2_1 _20958_ (.A(net1283),
    .B(net5666),
    .Y(_06014_));
 sg13g2_a21oi_1 _20959_ (.A1(net4887),
    .A2(net5666),
    .Y(_01781_),
    .B1(_06014_));
 sg13g2_nor2_1 _20960_ (.A(net1957),
    .B(net5670),
    .Y(_06015_));
 sg13g2_a21oi_1 _20961_ (.A1(net4772),
    .A2(net5670),
    .Y(_01782_),
    .B1(_06015_));
 sg13g2_nor2_1 _20962_ (.A(net1863),
    .B(net5671),
    .Y(_06016_));
 sg13g2_a21oi_1 _20963_ (.A1(net4882),
    .A2(net5671),
    .Y(_01783_),
    .B1(_06016_));
 sg13g2_nor2_1 _20964_ (.A(net1702),
    .B(net5672),
    .Y(_06017_));
 sg13g2_a21oi_1 _20965_ (.A1(net4876),
    .A2(net5672),
    .Y(_01784_),
    .B1(_06017_));
 sg13g2_nor2_1 _20966_ (.A(net2218),
    .B(net5673),
    .Y(_06018_));
 sg13g2_a21oi_1 _20967_ (.A1(net4762),
    .A2(net5673),
    .Y(_01785_),
    .B1(_06018_));
 sg13g2_nor2_1 _20968_ (.A(net1859),
    .B(net5667),
    .Y(_06019_));
 sg13g2_a21oi_1 _20969_ (.A1(net4868),
    .A2(net5667),
    .Y(_01786_),
    .B1(_06019_));
 sg13g2_nor2_1 _20970_ (.A(net1424),
    .B(net5674),
    .Y(_06020_));
 sg13g2_a21oi_1 _20971_ (.A1(net4862),
    .A2(net5674),
    .Y(_01787_),
    .B1(_06020_));
 sg13g2_nor2_1 _20972_ (.A(net1595),
    .B(net5669),
    .Y(_06021_));
 sg13g2_a21oi_1 _20973_ (.A1(net4857),
    .A2(net5669),
    .Y(_01788_),
    .B1(_06021_));
 sg13g2_nor2_1 _20974_ (.A(net1948),
    .B(net5667),
    .Y(_06022_));
 sg13g2_a21oi_1 _20975_ (.A1(net4856),
    .A2(net5667),
    .Y(_01789_),
    .B1(_06022_));
 sg13g2_nor2_1 _20976_ (.A(net2034),
    .B(net5671),
    .Y(_06023_));
 sg13g2_a21oi_1 _20977_ (.A1(net4847),
    .A2(net5671),
    .Y(_01790_),
    .B1(_06023_));
 sg13g2_nor2_1 _20978_ (.A(net1455),
    .B(net5667),
    .Y(_06024_));
 sg13g2_a21oi_1 _20979_ (.A1(net4842),
    .A2(net5667),
    .Y(_01791_),
    .B1(_06024_));
 sg13g2_nor2_1 _20980_ (.A(net1303),
    .B(net5666),
    .Y(_06025_));
 sg13g2_a21oi_1 _20981_ (.A1(net4841),
    .A2(net5666),
    .Y(_01792_),
    .B1(_06025_));
 sg13g2_nor2_1 _20982_ (.A(net2585),
    .B(net5666),
    .Y(_06026_));
 sg13g2_a21oi_1 _20983_ (.A1(net4834),
    .A2(net5666),
    .Y(_01793_),
    .B1(_06026_));
 sg13g2_nor2_1 _20984_ (.A(net1621),
    .B(net5672),
    .Y(_06027_));
 sg13g2_a21oi_1 _20985_ (.A1(net4827),
    .A2(net5672),
    .Y(_01794_),
    .B1(_06027_));
 sg13g2_nor2_1 _20986_ (.A(net2655),
    .B(net5672),
    .Y(_06028_));
 sg13g2_a21oi_1 _20987_ (.A1(net4822),
    .A2(net5672),
    .Y(_01795_),
    .B1(_06028_));
 sg13g2_nand4_1 _20988_ (.B(net6217),
    .C(_05625_),
    .A(net6215),
    .Y(_06029_),
    .D(net6071));
 sg13g2_nand2_1 _20989_ (.Y(_06030_),
    .A(net1045),
    .B(net5658));
 sg13g2_o21ai_1 _20990_ (.B1(_06030_),
    .Y(_01796_),
    .A1(net4994),
    .A2(net5658));
 sg13g2_nand2_1 _20991_ (.Y(_06031_),
    .A(net1256),
    .B(net5658));
 sg13g2_o21ai_1 _20992_ (.B1(_06031_),
    .Y(_01797_),
    .A1(net4990),
    .A2(net5658));
 sg13g2_nand2_1 _20993_ (.Y(_06032_),
    .A(net491),
    .B(net5658));
 sg13g2_o21ai_1 _20994_ (.B1(_06032_),
    .Y(_01798_),
    .A1(net4986),
    .A2(net5658));
 sg13g2_nand2_1 _20995_ (.Y(_06033_),
    .A(net1006),
    .B(net5657));
 sg13g2_o21ai_1 _20996_ (.B1(_06033_),
    .Y(_01799_),
    .A1(net4982),
    .A2(net5657));
 sg13g2_nand2_1 _20997_ (.Y(_06034_),
    .A(net819),
    .B(net5662));
 sg13g2_o21ai_1 _20998_ (.B1(_06034_),
    .Y(_01800_),
    .A1(net4978),
    .A2(net5662));
 sg13g2_nand2_1 _20999_ (.Y(_06035_),
    .A(net809),
    .B(net5664));
 sg13g2_o21ai_1 _21000_ (.B1(_06035_),
    .Y(_01801_),
    .A1(net4971),
    .A2(net5664));
 sg13g2_nand2_1 _21001_ (.Y(_06036_),
    .A(net1127),
    .B(net5664));
 sg13g2_o21ai_1 _21002_ (.B1(_06036_),
    .Y(_01802_),
    .A1(net4965),
    .A2(net5664));
 sg13g2_nand2_1 _21003_ (.Y(_06037_),
    .A(net803),
    .B(net5662));
 sg13g2_o21ai_1 _21004_ (.B1(_06037_),
    .Y(_01803_),
    .A1(net4919),
    .A2(net5662));
 sg13g2_nand2_1 _21005_ (.Y(_06038_),
    .A(net810),
    .B(net5659));
 sg13g2_o21ai_1 _21006_ (.B1(_06038_),
    .Y(_01804_),
    .A1(net4781),
    .A2(net5659));
 sg13g2_nand2_1 _21007_ (.Y(_06039_),
    .A(net697),
    .B(net5665));
 sg13g2_o21ai_1 _21008_ (.B1(_06039_),
    .Y(_01805_),
    .A1(net4911),
    .A2(net5663));
 sg13g2_nand2_1 _21009_ (.Y(_06040_),
    .A(net952),
    .B(net5663));
 sg13g2_o21ai_1 _21010_ (.B1(_06040_),
    .Y(_01806_),
    .A1(net4909),
    .A2(net5663));
 sg13g2_nand2_1 _21011_ (.Y(_06041_),
    .A(net514),
    .B(net5659));
 sg13g2_o21ai_1 _21012_ (.B1(_06041_),
    .Y(_01807_),
    .A1(net4774),
    .A2(net5659));
 sg13g2_nand2_1 _21013_ (.Y(_06042_),
    .A(net1035),
    .B(net5661));
 sg13g2_o21ai_1 _21014_ (.B1(_06042_),
    .Y(_01808_),
    .A1(net4904),
    .A2(net5661));
 sg13g2_nand2_1 _21015_ (.Y(_06043_),
    .A(net1909),
    .B(net5661));
 sg13g2_o21ai_1 _21016_ (.B1(_06043_),
    .Y(_01809_),
    .A1(net4960),
    .A2(net5661));
 sg13g2_nand2_1 _21017_ (.Y(_06044_),
    .A(net598),
    .B(net5656));
 sg13g2_o21ai_1 _21018_ (.B1(_06044_),
    .Y(_01810_),
    .A1(net4956),
    .A2(net5656));
 sg13g2_nand2_1 _21019_ (.Y(_06045_),
    .A(net992),
    .B(net5665));
 sg13g2_o21ai_1 _21020_ (.B1(_06045_),
    .Y(_01811_),
    .A1(net4894),
    .A2(net5665));
 sg13g2_nand2_1 _21021_ (.Y(_06046_),
    .A(net632),
    .B(net5661));
 sg13g2_o21ai_1 _21022_ (.B1(_06046_),
    .Y(_01812_),
    .A1(net4892),
    .A2(net5661));
 sg13g2_nand2_1 _21023_ (.Y(_06047_),
    .A(net676),
    .B(net5657));
 sg13g2_o21ai_1 _21024_ (.B1(_06047_),
    .Y(_01813_),
    .A1(net4887),
    .A2(net5657));
 sg13g2_nand2_1 _21025_ (.Y(_06048_),
    .A(net1109),
    .B(net5661));
 sg13g2_o21ai_1 _21026_ (.B1(_06048_),
    .Y(_01814_),
    .A1(net4772),
    .A2(net5661));
 sg13g2_nand2_1 _21027_ (.Y(_06049_),
    .A(net784),
    .B(net5662));
 sg13g2_o21ai_1 _21028_ (.B1(_06049_),
    .Y(_01815_),
    .A1(net4881),
    .A2(net5662));
 sg13g2_nand2_1 _21029_ (.Y(_06050_),
    .A(net550),
    .B(net5665));
 sg13g2_o21ai_1 _21030_ (.B1(_06050_),
    .Y(_01816_),
    .A1(net4872),
    .A2(net5665));
 sg13g2_nand2_1 _21031_ (.Y(_06051_),
    .A(net768),
    .B(net5664));
 sg13g2_o21ai_1 _21032_ (.B1(_06051_),
    .Y(_01817_),
    .A1(net4763),
    .A2(net5664));
 sg13g2_nand2_1 _21033_ (.Y(_06052_),
    .A(net534),
    .B(net5656));
 sg13g2_o21ai_1 _21034_ (.B1(_06052_),
    .Y(_01818_),
    .A1(net4867),
    .A2(net5656));
 sg13g2_nand2_1 _21035_ (.Y(_06053_),
    .A(net766),
    .B(net5663));
 sg13g2_o21ai_1 _21036_ (.B1(_06053_),
    .Y(_01819_),
    .A1(net4862),
    .A2(net5663));
 sg13g2_nand2_1 _21037_ (.Y(_06054_),
    .A(net940),
    .B(net5657));
 sg13g2_o21ai_1 _21038_ (.B1(_06054_),
    .Y(_01820_),
    .A1(net4857),
    .A2(net5657));
 sg13g2_nand2_1 _21039_ (.Y(_06055_),
    .A(net640),
    .B(net5656));
 sg13g2_o21ai_1 _21040_ (.B1(_06055_),
    .Y(_01821_),
    .A1(net4852),
    .A2(net5656));
 sg13g2_nand2_1 _21041_ (.Y(_06056_),
    .A(net449),
    .B(net5662));
 sg13g2_o21ai_1 _21042_ (.B1(_06056_),
    .Y(_01822_),
    .A1(net4851),
    .A2(net5662));
 sg13g2_nand2_1 _21043_ (.Y(_06057_),
    .A(net499),
    .B(net5656));
 sg13g2_o21ai_1 _21044_ (.B1(_06057_),
    .Y(_01823_),
    .A1(net4842),
    .A2(net5656));
 sg13g2_nand2_1 _21045_ (.Y(_06058_),
    .A(net723),
    .B(net5657));
 sg13g2_o21ai_1 _21046_ (.B1(_06058_),
    .Y(_01824_),
    .A1(net4838),
    .A2(net5657));
 sg13g2_nand2_1 _21047_ (.Y(_06059_),
    .A(net876),
    .B(net5658));
 sg13g2_o21ai_1 _21048_ (.B1(_06059_),
    .Y(_01825_),
    .A1(net4836),
    .A2(net5658));
 sg13g2_nand2_1 _21049_ (.Y(_06060_),
    .A(net1022),
    .B(net5663));
 sg13g2_o21ai_1 _21050_ (.B1(_06060_),
    .Y(_01826_),
    .A1(net4827),
    .A2(net5663));
 sg13g2_nand2_1 _21051_ (.Y(_06061_),
    .A(net387),
    .B(net5663));
 sg13g2_o21ai_1 _21052_ (.B1(_06061_),
    .Y(_01827_),
    .A1(net4826),
    .A2(net5664));
 sg13g2_and4_1 _21053_ (.A(net6214),
    .B(net6216),
    .C(_05660_),
    .D(net6070),
    .X(_06062_));
 sg13g2_nor2_1 _21054_ (.A(net1605),
    .B(net5648),
    .Y(_06063_));
 sg13g2_a21oi_1 _21055_ (.A1(net4998),
    .A2(net5648),
    .Y(_01828_),
    .B1(_06063_));
 sg13g2_nor2_1 _21056_ (.A(net2149),
    .B(net5648),
    .Y(_06064_));
 sg13g2_a21oi_1 _21057_ (.A1(net4989),
    .A2(net5648),
    .Y(_01829_),
    .B1(_06064_));
 sg13g2_nor2_1 _21058_ (.A(net1665),
    .B(net5648),
    .Y(_06065_));
 sg13g2_a21oi_1 _21059_ (.A1(net4985),
    .A2(net5648),
    .Y(_01830_),
    .B1(_06065_));
 sg13g2_nor2_1 _21060_ (.A(net1892),
    .B(net5647),
    .Y(_06066_));
 sg13g2_a21oi_1 _21061_ (.A1(net4983),
    .A2(net5647),
    .Y(_01831_),
    .B1(_06066_));
 sg13g2_nor2_1 _21062_ (.A(net1564),
    .B(net5651),
    .Y(_06067_));
 sg13g2_a21oi_1 _21063_ (.A1(net4976),
    .A2(net5651),
    .Y(_01832_),
    .B1(_06067_));
 sg13g2_nor2_1 _21064_ (.A(net1606),
    .B(net5654),
    .Y(_06068_));
 sg13g2_a21oi_1 _21065_ (.A1(net4971),
    .A2(net5654),
    .Y(_01833_),
    .B1(_06068_));
 sg13g2_nor2_1 _21066_ (.A(net1544),
    .B(net5654),
    .Y(_06069_));
 sg13g2_a21oi_1 _21067_ (.A1(net4967),
    .A2(net5654),
    .Y(_01834_),
    .B1(_06069_));
 sg13g2_nor2_1 _21068_ (.A(net1960),
    .B(net5655),
    .Y(_06070_));
 sg13g2_a21oi_1 _21069_ (.A1(net4919),
    .A2(net5651),
    .Y(_01835_),
    .B1(_06070_));
 sg13g2_nor2_1 _21070_ (.A(net2068),
    .B(net5654),
    .Y(_06071_));
 sg13g2_a21oi_1 _21071_ (.A1(net4779),
    .A2(net5654),
    .Y(_01836_),
    .B1(_06071_));
 sg13g2_nor2_1 _21072_ (.A(net1747),
    .B(net5652),
    .Y(_06072_));
 sg13g2_a21oi_1 _21073_ (.A1(net4911),
    .A2(net5652),
    .Y(_01837_),
    .B1(_06072_));
 sg13g2_nor2_1 _21074_ (.A(net1636),
    .B(net5652),
    .Y(_06073_));
 sg13g2_a21oi_1 _21075_ (.A1(net4905),
    .A2(net5652),
    .Y(_01838_),
    .B1(_06073_));
 sg13g2_nor2_1 _21076_ (.A(net1580),
    .B(net5648),
    .Y(_06074_));
 sg13g2_a21oi_1 _21077_ (.A1(net4775),
    .A2(net5648),
    .Y(_01839_),
    .B1(_06074_));
 sg13g2_nor2_1 _21078_ (.A(net1954),
    .B(net5650),
    .Y(_06075_));
 sg13g2_a21oi_1 _21079_ (.A1(net4904),
    .A2(net5650),
    .Y(_01840_),
    .B1(_06075_));
 sg13g2_nor2_1 _21080_ (.A(net1602),
    .B(net5650),
    .Y(_06076_));
 sg13g2_a21oi_1 _21081_ (.A1(net4959),
    .A2(net5650),
    .Y(_01841_),
    .B1(_06076_));
 sg13g2_nor2_1 _21082_ (.A(net1768),
    .B(net5646),
    .Y(_06077_));
 sg13g2_a21oi_1 _21083_ (.A1(net4954),
    .A2(net5646),
    .Y(_01842_),
    .B1(_06077_));
 sg13g2_nor2_1 _21084_ (.A(net2100),
    .B(net5655),
    .Y(_06078_));
 sg13g2_a21oi_1 _21085_ (.A1(net4894),
    .A2(net5655),
    .Y(_01843_),
    .B1(_06078_));
 sg13g2_nor2_1 _21086_ (.A(net2616),
    .B(net5650),
    .Y(_06079_));
 sg13g2_a21oi_1 _21087_ (.A1(net4889),
    .A2(net5650),
    .Y(_01844_),
    .B1(_06079_));
 sg13g2_nor2_1 _21088_ (.A(net2209),
    .B(net5647),
    .Y(_06080_));
 sg13g2_a21oi_1 _21089_ (.A1(net4885),
    .A2(net5647),
    .Y(_01845_),
    .B1(_06080_));
 sg13g2_nor2_1 _21090_ (.A(net1271),
    .B(net5650),
    .Y(_06081_));
 sg13g2_a21oi_1 _21091_ (.A1(net4769),
    .A2(net5650),
    .Y(_01846_),
    .B1(_06081_));
 sg13g2_nor2_1 _21092_ (.A(net2116),
    .B(net5651),
    .Y(_06082_));
 sg13g2_a21oi_1 _21093_ (.A1(net4880),
    .A2(net5651),
    .Y(_01847_),
    .B1(_06082_));
 sg13g2_nor2_1 _21094_ (.A(net1604),
    .B(net5652),
    .Y(_06083_));
 sg13g2_a21oi_1 _21095_ (.A1(net4873),
    .A2(net5652),
    .Y(_01848_),
    .B1(_06083_));
 sg13g2_nor2_1 _21096_ (.A(net2171),
    .B(net5654),
    .Y(_06084_));
 sg13g2_a21oi_1 _21097_ (.A1(net4762),
    .A2(net5654),
    .Y(_01849_),
    .B1(_06084_));
 sg13g2_nor2_1 _21098_ (.A(net2263),
    .B(net5646),
    .Y(_06085_));
 sg13g2_a21oi_1 _21099_ (.A1(net4868),
    .A2(net5646),
    .Y(_01850_),
    .B1(_06085_));
 sg13g2_nor2_1 _21100_ (.A(net1789),
    .B(net5653),
    .Y(_06086_));
 sg13g2_a21oi_1 _21101_ (.A1(net4866),
    .A2(net5653),
    .Y(_01851_),
    .B1(_06086_));
 sg13g2_nor2_1 _21102_ (.A(net1710),
    .B(net5647),
    .Y(_06087_));
 sg13g2_a21oi_1 _21103_ (.A1(net4859),
    .A2(net5647),
    .Y(_01852_),
    .B1(_06087_));
 sg13g2_nor2_1 _21104_ (.A(net1965),
    .B(net5646),
    .Y(_06088_));
 sg13g2_a21oi_1 _21105_ (.A1(net4853),
    .A2(net5646),
    .Y(_01853_),
    .B1(_06088_));
 sg13g2_nor2_1 _21106_ (.A(net1624),
    .B(net5651),
    .Y(_06089_));
 sg13g2_a21oi_1 _21107_ (.A1(net4850),
    .A2(net5651),
    .Y(_01854_),
    .B1(_06089_));
 sg13g2_nor2_1 _21108_ (.A(net1233),
    .B(net5646),
    .Y(_06090_));
 sg13g2_a21oi_1 _21109_ (.A1(net4843),
    .A2(net5646),
    .Y(_01855_),
    .B1(_06090_));
 sg13g2_nor2_1 _21110_ (.A(net1218),
    .B(net5647),
    .Y(_06091_));
 sg13g2_a21oi_1 _21111_ (.A1(net4837),
    .A2(net5647),
    .Y(_01856_),
    .B1(_06091_));
 sg13g2_nor2_1 _21112_ (.A(net1945),
    .B(net5649),
    .Y(_06092_));
 sg13g2_a21oi_1 _21113_ (.A1(net4834),
    .A2(net5649),
    .Y(_01857_),
    .B1(_06092_));
 sg13g2_nor2_1 _21114_ (.A(net2029),
    .B(net5653),
    .Y(_06093_));
 sg13g2_a21oi_1 _21115_ (.A1(net4829),
    .A2(net5653),
    .Y(_01858_),
    .B1(_06093_));
 sg13g2_nor2_1 _21116_ (.A(net2097),
    .B(net5652),
    .Y(_06094_));
 sg13g2_a21oi_1 _21117_ (.A1(net4822),
    .A2(net5652),
    .Y(_01859_),
    .B1(_06094_));
 sg13g2_nand2_1 _21118_ (.Y(_06095_),
    .A(_05625_),
    .B(_05694_));
 sg13g2_nor2_2 _21119_ (.A(_09505_),
    .B(_06095_),
    .Y(_06096_));
 sg13g2_nor2_1 _21120_ (.A(net1919),
    .B(net5403),
    .Y(_06097_));
 sg13g2_a21oi_1 _21121_ (.A1(net4995),
    .A2(net5403),
    .Y(_01860_),
    .B1(_06097_));
 sg13g2_nor2_1 _21122_ (.A(net1587),
    .B(net5403),
    .Y(_06098_));
 sg13g2_a21oi_1 _21123_ (.A1(net4992),
    .A2(net5403),
    .Y(_01861_),
    .B1(_06098_));
 sg13g2_nor2_1 _21124_ (.A(net1942),
    .B(net5403),
    .Y(_06099_));
 sg13g2_a21oi_1 _21125_ (.A1(net4987),
    .A2(net5403),
    .Y(_01862_),
    .B1(_06099_));
 sg13g2_nor2_1 _21126_ (.A(net2020),
    .B(net5401),
    .Y(_06100_));
 sg13g2_a21oi_1 _21127_ (.A1(net4981),
    .A2(net5401),
    .Y(_01863_),
    .B1(_06100_));
 sg13g2_nor2_1 _21128_ (.A(net2652),
    .B(net5407),
    .Y(_06101_));
 sg13g2_a21oi_1 _21129_ (.A1(net4974),
    .A2(net5402),
    .Y(_01864_),
    .B1(_06101_));
 sg13g2_nor2_1 _21130_ (.A(net1991),
    .B(net5409),
    .Y(_06102_));
 sg13g2_a21oi_1 _21131_ (.A1(net4972),
    .A2(net5409),
    .Y(_01865_),
    .B1(_06102_));
 sg13g2_nor2_1 _21132_ (.A(net1650),
    .B(net5404),
    .Y(_06103_));
 sg13g2_a21oi_1 _21133_ (.A1(net4964),
    .A2(net5404),
    .Y(_01866_),
    .B1(_06103_));
 sg13g2_nor2_1 _21134_ (.A(net1732),
    .B(net5406),
    .Y(_06104_));
 sg13g2_a21oi_1 _21135_ (.A1(net4918),
    .A2(net5406),
    .Y(_01867_),
    .B1(_06104_));
 sg13g2_nor2_1 _21136_ (.A(net2101),
    .B(net5404),
    .Y(_06105_));
 sg13g2_a21oi_1 _21137_ (.A1(net4779),
    .A2(net5404),
    .Y(_01868_),
    .B1(_06105_));
 sg13g2_nor2_1 _21138_ (.A(net1500),
    .B(net5409),
    .Y(_06106_));
 sg13g2_a21oi_1 _21139_ (.A1(net4915),
    .A2(net5409),
    .Y(_01869_),
    .B1(_06106_));
 sg13g2_nor2_1 _21140_ (.A(net1427),
    .B(net5408),
    .Y(_06107_));
 sg13g2_a21oi_1 _21141_ (.A1(net4909),
    .A2(net5408),
    .Y(_01870_),
    .B1(_06107_));
 sg13g2_nor2_1 _21142_ (.A(net1623),
    .B(net5404),
    .Y(_06108_));
 sg13g2_a21oi_1 _21143_ (.A1(net4775),
    .A2(net5404),
    .Y(_01871_),
    .B1(_06108_));
 sg13g2_nor2_1 _21144_ (.A(net1974),
    .B(net5406),
    .Y(_06109_));
 sg13g2_a21oi_1 _21145_ (.A1(net4899),
    .A2(net5406),
    .Y(_01872_),
    .B1(_06109_));
 sg13g2_nor2_1 _21146_ (.A(net1798),
    .B(net5406),
    .Y(_06110_));
 sg13g2_a21oi_1 _21147_ (.A1(net4961),
    .A2(net5406),
    .Y(_01873_),
    .B1(_06110_));
 sg13g2_nor2_1 _21148_ (.A(net1546),
    .B(net5401),
    .Y(_06111_));
 sg13g2_a21oi_1 _21149_ (.A1(net4956),
    .A2(net5401),
    .Y(_01874_),
    .B1(_06111_));
 sg13g2_nor2_1 _21150_ (.A(net1620),
    .B(net5410),
    .Y(_06112_));
 sg13g2_a21oi_1 _21151_ (.A1(net4895),
    .A2(net5410),
    .Y(_01875_),
    .B1(_06112_));
 sg13g2_nor2_1 _21152_ (.A(net1359),
    .B(net5407),
    .Y(_06113_));
 sg13g2_a21oi_1 _21153_ (.A1(net4890),
    .A2(net5407),
    .Y(_01876_),
    .B1(_06113_));
 sg13g2_nor2_1 _21154_ (.A(net2359),
    .B(net5402),
    .Y(_06114_));
 sg13g2_a21oi_1 _21155_ (.A1(net4884),
    .A2(net5402),
    .Y(_01877_),
    .B1(_06114_));
 sg13g2_nor2_1 _21156_ (.A(net1705),
    .B(net5406),
    .Y(_06115_));
 sg13g2_a21oi_1 _21157_ (.A1(net4768),
    .A2(net5406),
    .Y(_01878_),
    .B1(_06115_));
 sg13g2_nor2_1 _21158_ (.A(net1766),
    .B(net5407),
    .Y(_06116_));
 sg13g2_a21oi_1 _21159_ (.A1(net4880),
    .A2(net5407),
    .Y(_01879_),
    .B1(_06116_));
 sg13g2_nor2_1 _21160_ (.A(net1619),
    .B(net5408),
    .Y(_06117_));
 sg13g2_a21oi_1 _21161_ (.A1(net4876),
    .A2(net5410),
    .Y(_01880_),
    .B1(_06117_));
 sg13g2_nor2_1 _21162_ (.A(net1686),
    .B(net5409),
    .Y(_06118_));
 sg13g2_a21oi_1 _21163_ (.A1(net4765),
    .A2(net5409),
    .Y(_01881_),
    .B1(_06118_));
 sg13g2_nor2_1 _21164_ (.A(net1393),
    .B(net5401),
    .Y(_06119_));
 sg13g2_a21oi_1 _21165_ (.A1(net4869),
    .A2(net5402),
    .Y(_01882_),
    .B1(_06119_));
 sg13g2_nor2_1 _21166_ (.A(net1644),
    .B(net5408),
    .Y(_06120_));
 sg13g2_a21oi_1 _21167_ (.A1(net4866),
    .A2(net5408),
    .Y(_01883_),
    .B1(_06120_));
 sg13g2_nor2_1 _21168_ (.A(net2392),
    .B(net5405),
    .Y(_06121_));
 sg13g2_a21oi_1 _21169_ (.A1(net4858),
    .A2(net5405),
    .Y(_01884_),
    .B1(_06121_));
 sg13g2_nor2_1 _21170_ (.A(net2006),
    .B(net5401),
    .Y(_06122_));
 sg13g2_a21oi_1 _21171_ (.A1(net4854),
    .A2(net5401),
    .Y(_01885_),
    .B1(_06122_));
 sg13g2_nor2_1 _21172_ (.A(net1844),
    .B(net5407),
    .Y(_06123_));
 sg13g2_a21oi_1 _21173_ (.A1(net4848),
    .A2(net5407),
    .Y(_01886_),
    .B1(_06123_));
 sg13g2_nor2_1 _21174_ (.A(net1944),
    .B(net5401),
    .Y(_06124_));
 sg13g2_a21oi_1 _21175_ (.A1(net4844),
    .A2(net5402),
    .Y(_01887_),
    .B1(_06124_));
 sg13g2_nor2_1 _21176_ (.A(net1612),
    .B(net5402),
    .Y(_06125_));
 sg13g2_a21oi_1 _21177_ (.A1(net4840),
    .A2(net5402),
    .Y(_01888_),
    .B1(_06125_));
 sg13g2_nor2_1 _21178_ (.A(net2314),
    .B(net5403),
    .Y(_06126_));
 sg13g2_a21oi_1 _21179_ (.A1(net4836),
    .A2(net5403),
    .Y(_01889_),
    .B1(_06126_));
 sg13g2_nor2_1 _21180_ (.A(net1911),
    .B(net5408),
    .Y(_06127_));
 sg13g2_a21oi_1 _21181_ (.A1(net4827),
    .A2(net5408),
    .Y(_01890_),
    .B1(_06127_));
 sg13g2_nor2_1 _21182_ (.A(net1750),
    .B(net5408),
    .Y(_06128_));
 sg13g2_a21oi_1 _21183_ (.A1(net4823),
    .A2(net5409),
    .Y(_01891_),
    .B1(_06128_));
 sg13g2_nand4_1 _21184_ (.B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .C(_05694_),
    .A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .Y(_06129_),
    .D(net6070));
 sg13g2_nand2_1 _21185_ (.Y(_06130_),
    .A(net1029),
    .B(net5636));
 sg13g2_o21ai_1 _21186_ (.B1(_06130_),
    .Y(_01892_),
    .A1(net4998),
    .A2(net5636));
 sg13g2_nand2_1 _21187_ (.Y(_06131_),
    .A(net924),
    .B(net5636));
 sg13g2_o21ai_1 _21188_ (.B1(_06131_),
    .Y(_01893_),
    .A1(net4989),
    .A2(net5636));
 sg13g2_nand2_1 _21189_ (.Y(_06132_),
    .A(net1192),
    .B(net5637));
 sg13g2_o21ai_1 _21190_ (.B1(_06132_),
    .Y(_01894_),
    .A1(net4988),
    .A2(net5637));
 sg13g2_nand2_1 _21191_ (.Y(_06133_),
    .A(net830),
    .B(net5635));
 sg13g2_o21ai_1 _21192_ (.B1(_06133_),
    .Y(_01895_),
    .A1(net4981),
    .A2(net5635));
 sg13g2_nand2_1 _21193_ (.Y(_06134_),
    .A(net847),
    .B(net5639));
 sg13g2_o21ai_1 _21194_ (.B1(_06134_),
    .Y(_01896_),
    .A1(net4974),
    .A2(net5639));
 sg13g2_nand2_1 _21195_ (.Y(_06135_),
    .A(net999),
    .B(net5644));
 sg13g2_o21ai_1 _21196_ (.B1(_06135_),
    .Y(_01897_),
    .A1(net4971),
    .A2(net5644));
 sg13g2_nand2_1 _21197_ (.Y(_06136_),
    .A(net1043),
    .B(net5644));
 sg13g2_o21ai_1 _21198_ (.B1(_06136_),
    .Y(_01898_),
    .A1(net4967),
    .A2(net5644));
 sg13g2_nand2_1 _21199_ (.Y(_06137_),
    .A(net489),
    .B(net5640));
 sg13g2_o21ai_1 _21200_ (.B1(_06137_),
    .Y(_01899_),
    .A1(net4919),
    .A2(net5638));
 sg13g2_nand2_1 _21201_ (.Y(_06138_),
    .A(net659),
    .B(net5644));
 sg13g2_o21ai_1 _21202_ (.B1(_06138_),
    .Y(_01900_),
    .A1(net4780),
    .A2(net5644));
 sg13g2_nand2_1 _21203_ (.Y(_06139_),
    .A(net1079),
    .B(net5642));
 sg13g2_o21ai_1 _21204_ (.B1(_06139_),
    .Y(_01901_),
    .A1(net4914),
    .A2(net5642));
 sg13g2_nand2_1 _21205_ (.Y(_06140_),
    .A(net1234),
    .B(net5642));
 sg13g2_o21ai_1 _21206_ (.B1(_06140_),
    .Y(_01902_),
    .A1(net4906),
    .A2(net5642));
 sg13g2_nand2_1 _21207_ (.Y(_06141_),
    .A(net1325),
    .B(net5636));
 sg13g2_o21ai_1 _21208_ (.B1(_06141_),
    .Y(_01903_),
    .A1(net4773),
    .A2(net5636));
 sg13g2_nand2_1 _21209_ (.Y(_06142_),
    .A(net860),
    .B(net5640));
 sg13g2_o21ai_1 _21210_ (.B1(_06142_),
    .Y(_01904_),
    .A1(net4904),
    .A2(net5640));
 sg13g2_nand2_1 _21211_ (.Y(_06143_),
    .A(net985),
    .B(net5640));
 sg13g2_o21ai_1 _21212_ (.B1(_06143_),
    .Y(_01905_),
    .A1(net4960),
    .A2(net5640));
 sg13g2_nand2_1 _21213_ (.Y(_06144_),
    .A(net1053),
    .B(net5634));
 sg13g2_o21ai_1 _21214_ (.B1(_06144_),
    .Y(_01906_),
    .A1(net4955),
    .A2(net5634));
 sg13g2_nand2_1 _21215_ (.Y(_06145_),
    .A(net509),
    .B(net5641));
 sg13g2_o21ai_1 _21216_ (.B1(_06145_),
    .Y(_01907_),
    .A1(net4898),
    .A2(net5641));
 sg13g2_nand2_1 _21217_ (.Y(_06146_),
    .A(net962),
    .B(net5640));
 sg13g2_o21ai_1 _21218_ (.B1(_06146_),
    .Y(_01908_),
    .A1(net4889),
    .A2(net5638));
 sg13g2_nand2_1 _21219_ (.Y(_06147_),
    .A(net812),
    .B(net5638));
 sg13g2_o21ai_1 _21220_ (.B1(_06147_),
    .Y(_01909_),
    .A1(net4886),
    .A2(net5638));
 sg13g2_nand2_1 _21221_ (.Y(_06148_),
    .A(net835),
    .B(net5640));
 sg13g2_o21ai_1 _21222_ (.B1(_06148_),
    .Y(_01910_),
    .A1(net4769),
    .A2(net5640));
 sg13g2_nand2_1 _21223_ (.Y(_06149_),
    .A(net929),
    .B(net5638));
 sg13g2_o21ai_1 _21224_ (.B1(_06149_),
    .Y(_01911_),
    .A1(net4878),
    .A2(net5638));
 sg13g2_nand2_1 _21225_ (.Y(_06150_),
    .A(net528),
    .B(net5642));
 sg13g2_o21ai_1 _21226_ (.B1(_06150_),
    .Y(_01912_),
    .A1(net4872),
    .A2(net5642));
 sg13g2_nand2_1 _21227_ (.Y(_06151_),
    .A(net1219),
    .B(net5644));
 sg13g2_o21ai_1 _21228_ (.B1(_06151_),
    .Y(_01913_),
    .A1(net4762),
    .A2(net5644));
 sg13g2_nand2_1 _21229_ (.Y(_06152_),
    .A(net434),
    .B(net5634));
 sg13g2_o21ai_1 _21230_ (.B1(_06152_),
    .Y(_01914_),
    .A1(net4867),
    .A2(net5634));
 sg13g2_nand2_1 _21231_ (.Y(_06153_),
    .A(net1173),
    .B(net5643));
 sg13g2_o21ai_1 _21232_ (.B1(_06153_),
    .Y(_01915_),
    .A1(net4866),
    .A2(net5643));
 sg13g2_nand2_1 _21233_ (.Y(_06154_),
    .A(net513),
    .B(net5635));
 sg13g2_o21ai_1 _21234_ (.B1(_06154_),
    .Y(_01916_),
    .A1(net4859),
    .A2(net5635));
 sg13g2_nand2_1 _21235_ (.Y(_06155_),
    .A(net678),
    .B(net5634));
 sg13g2_o21ai_1 _21236_ (.B1(_06155_),
    .Y(_01917_),
    .A1(net4852),
    .A2(net5634));
 sg13g2_nand2_1 _21237_ (.Y(_06156_),
    .A(net471),
    .B(net5639));
 sg13g2_o21ai_1 _21238_ (.B1(_06156_),
    .Y(_01918_),
    .A1(net4850),
    .A2(net5639));
 sg13g2_nand2_1 _21239_ (.Y(_06157_),
    .A(net905),
    .B(net5634));
 sg13g2_o21ai_1 _21240_ (.B1(_06157_),
    .Y(_01919_),
    .A1(net4846),
    .A2(net5634));
 sg13g2_nand2_1 _21241_ (.Y(_06158_),
    .A(net757),
    .B(net5638));
 sg13g2_o21ai_1 _21242_ (.B1(_06158_),
    .Y(_01920_),
    .A1(net4837),
    .A2(net5638));
 sg13g2_nand2_1 _21243_ (.Y(_06159_),
    .A(net490),
    .B(net5636));
 sg13g2_o21ai_1 _21244_ (.B1(_06159_),
    .Y(_01921_),
    .A1(net4835),
    .A2(net5636));
 sg13g2_nand2_1 _21245_ (.Y(_06160_),
    .A(net1074),
    .B(net5643));
 sg13g2_o21ai_1 _21246_ (.B1(_06160_),
    .Y(_01922_),
    .A1(net4829),
    .A2(net5643));
 sg13g2_nand2_1 _21247_ (.Y(_06161_),
    .A(net870),
    .B(net5642));
 sg13g2_o21ai_1 _21248_ (.B1(_06161_),
    .Y(_01923_),
    .A1(net4825),
    .A2(net5642));
 sg13g2_and4_1 _21249_ (.A(net6215),
    .B(net6217),
    .C(_09504_),
    .D(_05590_),
    .X(_06162_));
 sg13g2_nor2_1 _21250_ (.A(net2042),
    .B(net5626),
    .Y(_06163_));
 sg13g2_a21oi_1 _21251_ (.A1(net4994),
    .A2(net5626),
    .Y(_01924_),
    .B1(_06163_));
 sg13g2_nor2_1 _21252_ (.A(net1876),
    .B(net5626),
    .Y(_06164_));
 sg13g2_a21oi_1 _21253_ (.A1(net4991),
    .A2(net5626),
    .Y(_01925_),
    .B1(_06164_));
 sg13g2_nor2_1 _21254_ (.A(net1653),
    .B(net5626),
    .Y(_06165_));
 sg13g2_a21oi_1 _21255_ (.A1(net4986),
    .A2(net5626),
    .Y(_01926_),
    .B1(_06165_));
 sg13g2_nor2_1 _21256_ (.A(net1463),
    .B(net5624),
    .Y(_06166_));
 sg13g2_a21oi_1 _21257_ (.A1(net4980),
    .A2(net5624),
    .Y(_01927_),
    .B1(_06166_));
 sg13g2_nor2_1 _21258_ (.A(net1498),
    .B(net5630),
    .Y(_06167_));
 sg13g2_a21oi_1 _21259_ (.A1(net4974),
    .A2(net5630),
    .Y(_01928_),
    .B1(_06167_));
 sg13g2_nor2_1 _21260_ (.A(net1846),
    .B(net5632),
    .Y(_06168_));
 sg13g2_a21oi_1 _21261_ (.A1(net4972),
    .A2(net5632),
    .Y(_01929_),
    .B1(_06168_));
 sg13g2_nor2_1 _21262_ (.A(net1700),
    .B(net5627),
    .Y(_06169_));
 sg13g2_a21oi_1 _21263_ (.A1(net4964),
    .A2(net5627),
    .Y(_01930_),
    .B1(_06169_));
 sg13g2_nor2_1 _21264_ (.A(net1596),
    .B(net5630),
    .Y(_06170_));
 sg13g2_a21oi_1 _21265_ (.A1(net4917),
    .A2(net5630),
    .Y(_01931_),
    .B1(_06170_));
 sg13g2_nor2_1 _21266_ (.A(net2331),
    .B(net5626),
    .Y(_06171_));
 sg13g2_a21oi_1 _21267_ (.A1(net4780),
    .A2(net5626),
    .Y(_01932_),
    .B1(_06171_));
 sg13g2_nor2_1 _21268_ (.A(net2514),
    .B(net5632),
    .Y(_06172_));
 sg13g2_a21oi_1 _21269_ (.A1(net4913),
    .A2(net5632),
    .Y(_01933_),
    .B1(_06172_));
 sg13g2_nor2_1 _21270_ (.A(net1330),
    .B(net5631),
    .Y(_06173_));
 sg13g2_a21oi_1 _21271_ (.A1(net4908),
    .A2(net5631),
    .Y(_01934_),
    .B1(_06173_));
 sg13g2_nor2_1 _21272_ (.A(net1625),
    .B(net5627),
    .Y(_06174_));
 sg13g2_a21oi_1 _21273_ (.A1(net4773),
    .A2(net5627),
    .Y(_01935_),
    .B1(_06174_));
 sg13g2_nor2_1 _21274_ (.A(net2604),
    .B(net5629),
    .Y(_06175_));
 sg13g2_a21oi_1 _21275_ (.A1(net4901),
    .A2(net5629),
    .Y(_01936_),
    .B1(_06175_));
 sg13g2_nor2_1 _21276_ (.A(net2367),
    .B(net5629),
    .Y(_06176_));
 sg13g2_a21oi_1 _21277_ (.A1(net4961),
    .A2(net5629),
    .Y(_01937_),
    .B1(_06176_));
 sg13g2_nor2_1 _21278_ (.A(net1920),
    .B(net5624),
    .Y(_06177_));
 sg13g2_a21oi_1 _21279_ (.A1(net4956),
    .A2(net5624),
    .Y(_01938_),
    .B1(_06177_));
 sg13g2_nor2_1 _21280_ (.A(net1561),
    .B(net5633),
    .Y(_06178_));
 sg13g2_a21oi_1 _21281_ (.A1(net4895),
    .A2(net5633),
    .Y(_01939_),
    .B1(_06178_));
 sg13g2_nor2_1 _21282_ (.A(net1505),
    .B(net5629),
    .Y(_06179_));
 sg13g2_a21oi_1 _21283_ (.A1(net4893),
    .A2(net5629),
    .Y(_01940_),
    .B1(_06179_));
 sg13g2_nor2_1 _21284_ (.A(net1806),
    .B(net5625),
    .Y(_06180_));
 sg13g2_a21oi_1 _21285_ (.A1(net4887),
    .A2(net5625),
    .Y(_01941_),
    .B1(_06180_));
 sg13g2_nor2_1 _21286_ (.A(net1979),
    .B(net5629),
    .Y(_06181_));
 sg13g2_a21oi_1 _21287_ (.A1(net4770),
    .A2(net5629),
    .Y(_01942_),
    .B1(_06181_));
 sg13g2_nor2_1 _21288_ (.A(net1770),
    .B(net5630),
    .Y(_06182_));
 sg13g2_a21oi_1 _21289_ (.A1(net4881),
    .A2(net5630),
    .Y(_01943_),
    .B1(_06182_));
 sg13g2_nor2_1 _21290_ (.A(net1883),
    .B(net5631),
    .Y(_06183_));
 sg13g2_a21oi_1 _21291_ (.A1(net4874),
    .A2(net5631),
    .Y(_01944_),
    .B1(_06183_));
 sg13g2_nor2_1 _21292_ (.A(net2124),
    .B(net5632),
    .Y(_06184_));
 sg13g2_a21oi_1 _21293_ (.A1(net4762),
    .A2(net5632),
    .Y(_01945_),
    .B1(_06184_));
 sg13g2_nor2_1 _21294_ (.A(net2066),
    .B(net5625),
    .Y(_06185_));
 sg13g2_a21oi_1 _21295_ (.A1(net4868),
    .A2(net5625),
    .Y(_01946_),
    .B1(_06185_));
 sg13g2_nor2_1 _21296_ (.A(net2278),
    .B(net5633),
    .Y(_06186_));
 sg13g2_a21oi_1 _21297_ (.A1(net4862),
    .A2(net5632),
    .Y(_01947_),
    .B1(_06186_));
 sg13g2_nor2_1 _21298_ (.A(net1964),
    .B(net5625),
    .Y(_06187_));
 sg13g2_a21oi_1 _21299_ (.A1(net4860),
    .A2(net5625),
    .Y(_01948_),
    .B1(_06187_));
 sg13g2_nor2_1 _21300_ (.A(net1707),
    .B(net5624),
    .Y(_06188_));
 sg13g2_a21oi_1 _21301_ (.A1(net4853),
    .A2(net5624),
    .Y(_01949_),
    .B1(_06188_));
 sg13g2_nor2_1 _21302_ (.A(net2172),
    .B(net5630),
    .Y(_06189_));
 sg13g2_a21oi_1 _21303_ (.A1(net4850),
    .A2(net5630),
    .Y(_01950_),
    .B1(_06189_));
 sg13g2_nor2_1 _21304_ (.A(net2253),
    .B(net5624),
    .Y(_06190_));
 sg13g2_a21oi_1 _21305_ (.A1(net4843),
    .A2(net5624),
    .Y(_01951_),
    .B1(_06190_));
 sg13g2_nor2_1 _21306_ (.A(net2189),
    .B(net5625),
    .Y(_06191_));
 sg13g2_a21oi_1 _21307_ (.A1(net4837),
    .A2(net5628),
    .Y(_01952_),
    .B1(_06191_));
 sg13g2_nor2_1 _21308_ (.A(net1501),
    .B(net5627),
    .Y(_06192_));
 sg13g2_a21oi_1 _21309_ (.A1(net4832),
    .A2(net5627),
    .Y(_01953_),
    .B1(_06192_));
 sg13g2_nor2_1 _21310_ (.A(net2162),
    .B(net5631),
    .Y(_06193_));
 sg13g2_a21oi_1 _21311_ (.A1(net4829),
    .A2(net5631),
    .Y(_01954_),
    .B1(_06193_));
 sg13g2_nor2_1 _21312_ (.A(net1875),
    .B(net5631),
    .Y(_06194_));
 sg13g2_a21oi_1 _21313_ (.A1(net4824),
    .A2(net5631),
    .Y(_01955_),
    .B1(_06194_));
 sg13g2_nand2_1 _21314_ (.Y(_06195_),
    .A(_05590_),
    .B(_05694_));
 sg13g2_nor2_1 _21315_ (.A(_05896_),
    .B(_06195_),
    .Y(_06196_));
 sg13g2_nor2_1 _21316_ (.A(net1313),
    .B(net5232),
    .Y(_06197_));
 sg13g2_a21oi_1 _21317_ (.A1(net4995),
    .A2(net5232),
    .Y(_01956_),
    .B1(_06197_));
 sg13g2_nor2_1 _21318_ (.A(net2225),
    .B(net5232),
    .Y(_06198_));
 sg13g2_a21oi_1 _21319_ (.A1(net4989),
    .A2(net5232),
    .Y(_01957_),
    .B1(_06198_));
 sg13g2_nor2_1 _21320_ (.A(net1617),
    .B(net5232),
    .Y(_06199_));
 sg13g2_a21oi_1 _21321_ (.A1(net4986),
    .A2(net5232),
    .Y(_01958_),
    .B1(_06199_));
 sg13g2_nor2_1 _21322_ (.A(net2243),
    .B(net5231),
    .Y(_06200_));
 sg13g2_a21oi_1 _21323_ (.A1(net4981),
    .A2(net5231),
    .Y(_01959_),
    .B1(_06200_));
 sg13g2_nor2_1 _21324_ (.A(net1529),
    .B(net5235),
    .Y(_06201_));
 sg13g2_a21oi_1 _21325_ (.A1(net4974),
    .A2(net5235),
    .Y(_01960_),
    .B1(_06201_));
 sg13g2_nor2_1 _21326_ (.A(net1628),
    .B(net5239),
    .Y(_06202_));
 sg13g2_a21oi_1 _21327_ (.A1(net4971),
    .A2(net5239),
    .Y(_01961_),
    .B1(_06202_));
 sg13g2_nor2_1 _21328_ (.A(net2041),
    .B(net5233),
    .Y(_06203_));
 sg13g2_a21oi_1 _21329_ (.A1(net4966),
    .A2(net5233),
    .Y(_01962_),
    .B1(_06203_));
 sg13g2_nor2_1 _21330_ (.A(net1472),
    .B(net5235),
    .Y(_06204_));
 sg13g2_a21oi_1 _21331_ (.A1(net4918),
    .A2(net5235),
    .Y(_01963_),
    .B1(_06204_));
 sg13g2_nor2_1 _21332_ (.A(net1820),
    .B(net5232),
    .Y(_06205_));
 sg13g2_a21oi_1 _21333_ (.A1(net4780),
    .A2(net5232),
    .Y(_01964_),
    .B1(_06205_));
 sg13g2_nor2_1 _21334_ (.A(net2686),
    .B(net5239),
    .Y(_06206_));
 sg13g2_a21oi_1 _21335_ (.A1(net4914),
    .A2(net5239),
    .Y(_01965_),
    .B1(_06206_));
 sg13g2_nor2_1 _21336_ (.A(net1804),
    .B(net5238),
    .Y(_06207_));
 sg13g2_a21oi_1 _21337_ (.A1(net4907),
    .A2(net5238),
    .Y(_01966_),
    .B1(_06207_));
 sg13g2_nor2_1 _21338_ (.A(net2211),
    .B(net5233),
    .Y(_06208_));
 sg13g2_a21oi_1 _21339_ (.A1(net4773),
    .A2(net5233),
    .Y(_01967_),
    .B1(_06208_));
 sg13g2_nor2_1 _21340_ (.A(net1733),
    .B(net5236),
    .Y(_06209_));
 sg13g2_a21oi_1 _21341_ (.A1(net4902),
    .A2(net5236),
    .Y(_01968_),
    .B1(_06209_));
 sg13g2_nor2_1 _21342_ (.A(net2236),
    .B(net5236),
    .Y(_06210_));
 sg13g2_a21oi_1 _21343_ (.A1(net4963),
    .A2(net5236),
    .Y(_01969_),
    .B1(_06210_));
 sg13g2_nor2_1 _21344_ (.A(net1797),
    .B(net5230),
    .Y(_06211_));
 sg13g2_a21oi_1 _21345_ (.A1(net4954),
    .A2(net5230),
    .Y(_01970_),
    .B1(_06211_));
 sg13g2_nor2_1 _21346_ (.A(net1975),
    .B(net5237),
    .Y(_06212_));
 sg13g2_a21oi_1 _21347_ (.A1(net4895),
    .A2(net5237),
    .Y(_01971_),
    .B1(_06212_));
 sg13g2_nor2_1 _21348_ (.A(net1441),
    .B(net5236),
    .Y(_06213_));
 sg13g2_a21oi_1 _21349_ (.A1(net4891),
    .A2(net5236),
    .Y(_01972_),
    .B1(_06213_));
 sg13g2_nor2_1 _21350_ (.A(net2147),
    .B(net5231),
    .Y(_06214_));
 sg13g2_a21oi_1 _21351_ (.A1(net4884),
    .A2(net5231),
    .Y(_01973_),
    .B1(_06214_));
 sg13g2_nor2_1 _21352_ (.A(net2188),
    .B(net5236),
    .Y(_06215_));
 sg13g2_a21oi_1 _21353_ (.A1(net4770),
    .A2(net5236),
    .Y(_01974_),
    .B1(_06215_));
 sg13g2_nor2_1 _21354_ (.A(net1490),
    .B(net5235),
    .Y(_06216_));
 sg13g2_a21oi_1 _21355_ (.A1(net4878),
    .A2(net5235),
    .Y(_01975_),
    .B1(_06216_));
 sg13g2_nor2_1 _21356_ (.A(net1406),
    .B(net5238),
    .Y(_06217_));
 sg13g2_a21oi_1 _21357_ (.A1(net4874),
    .A2(net5238),
    .Y(_01976_),
    .B1(_06217_));
 sg13g2_nor2_1 _21358_ (.A(net1553),
    .B(net5239),
    .Y(_06218_));
 sg13g2_a21oi_1 _21359_ (.A1(net4764),
    .A2(net5239),
    .Y(_01977_),
    .B1(_06218_));
 sg13g2_nor2_1 _21360_ (.A(net1274),
    .B(net5230),
    .Y(_06219_));
 sg13g2_a21oi_1 _21361_ (.A1(net4869),
    .A2(net5230),
    .Y(_01978_),
    .B1(_06219_));
 sg13g2_nor2_1 _21362_ (.A(net1590),
    .B(net5240),
    .Y(_06220_));
 sg13g2_a21oi_1 _21363_ (.A1(net4862),
    .A2(net5239),
    .Y(_01979_),
    .B1(_06220_));
 sg13g2_nor2_1 _21364_ (.A(net2140),
    .B(net5231),
    .Y(_06221_));
 sg13g2_a21oi_1 _21365_ (.A1(net4857),
    .A2(net5231),
    .Y(_01980_),
    .B1(_06221_));
 sg13g2_nor2_1 _21366_ (.A(net1630),
    .B(net5230),
    .Y(_06222_));
 sg13g2_a21oi_1 _21367_ (.A1(net4856),
    .A2(net5230),
    .Y(_01981_),
    .B1(_06222_));
 sg13g2_nor2_1 _21368_ (.A(net2291),
    .B(net5235),
    .Y(_06223_));
 sg13g2_a21oi_1 _21369_ (.A1(net4848),
    .A2(net5235),
    .Y(_01982_),
    .B1(_06223_));
 sg13g2_nor2_1 _21370_ (.A(net1753),
    .B(net5230),
    .Y(_06224_));
 sg13g2_a21oi_1 _21371_ (.A1(net4842),
    .A2(net5230),
    .Y(_01983_),
    .B1(_06224_));
 sg13g2_nor2_1 _21372_ (.A(net2028),
    .B(net5237),
    .Y(_06225_));
 sg13g2_a21oi_1 _21373_ (.A1(net4838),
    .A2(net5237),
    .Y(_01984_),
    .B1(_06225_));
 sg13g2_nor2_1 _21374_ (.A(net1689),
    .B(net5233),
    .Y(_06226_));
 sg13g2_a21oi_1 _21375_ (.A1(net4834),
    .A2(net5233),
    .Y(_01985_),
    .B1(_06226_));
 sg13g2_nor2_1 _21376_ (.A(net1244),
    .B(net5238),
    .Y(_06227_));
 sg13g2_a21oi_1 _21377_ (.A1(net4827),
    .A2(net5238),
    .Y(_01986_),
    .B1(_06227_));
 sg13g2_nor2_1 _21378_ (.A(net1722),
    .B(net5238),
    .Y(_06228_));
 sg13g2_a21oi_1 _21379_ (.A1(net4824),
    .A2(net5238),
    .Y(_01987_),
    .B1(_06228_));
 sg13g2_nor2_1 _21380_ (.A(_05896_),
    .B(_06095_),
    .Y(_06229_));
 sg13g2_nor2_1 _21381_ (.A(net2269),
    .B(net5221),
    .Y(_06230_));
 sg13g2_a21oi_1 _21382_ (.A1(net4996),
    .A2(net5221),
    .Y(_01988_),
    .B1(_06230_));
 sg13g2_nor2_1 _21383_ (.A(net2067),
    .B(net5221),
    .Y(_06231_));
 sg13g2_a21oi_1 _21384_ (.A1(net4991),
    .A2(net5221),
    .Y(_01989_),
    .B1(_06231_));
 sg13g2_nor2_1 _21385_ (.A(net1277),
    .B(net5221),
    .Y(_06232_));
 sg13g2_a21oi_1 _21386_ (.A1(net4987),
    .A2(net5221),
    .Y(_01990_),
    .B1(_06232_));
 sg13g2_nor2_1 _21387_ (.A(net2268),
    .B(net5219),
    .Y(_06233_));
 sg13g2_a21oi_1 _21388_ (.A1(net4979),
    .A2(net5219),
    .Y(_01991_),
    .B1(_06233_));
 sg13g2_nor2_1 _21389_ (.A(net1752),
    .B(net5226),
    .Y(_06234_));
 sg13g2_a21oi_1 _21390_ (.A1(net4975),
    .A2(net5226),
    .Y(_01992_),
    .B1(_06234_));
 sg13g2_nor2_1 _21391_ (.A(net1429),
    .B(net5228),
    .Y(_06235_));
 sg13g2_a21oi_1 _21392_ (.A1(net4970),
    .A2(net5228),
    .Y(_01993_),
    .B1(_06235_));
 sg13g2_nor2_1 _21393_ (.A(net2280),
    .B(net5222),
    .Y(_06236_));
 sg13g2_a21oi_1 _21394_ (.A1(net4967),
    .A2(net5221),
    .Y(_01994_),
    .B1(_06236_));
 sg13g2_nor2_1 _21395_ (.A(net1403),
    .B(net5225),
    .Y(_06237_));
 sg13g2_a21oi_1 _21396_ (.A1(net4916),
    .A2(net5225),
    .Y(_01995_),
    .B1(_06237_));
 sg13g2_nor2_1 _21397_ (.A(net2634),
    .B(net5221),
    .Y(_06238_));
 sg13g2_a21oi_1 _21398_ (.A1(net4782),
    .A2(net5222),
    .Y(_01996_),
    .B1(_06238_));
 sg13g2_nor2_1 _21399_ (.A(net1525),
    .B(net5228),
    .Y(_06239_));
 sg13g2_a21oi_1 _21400_ (.A1(net4912),
    .A2(net5228),
    .Y(_01997_),
    .B1(_06239_));
 sg13g2_nor2_1 _21401_ (.A(net1340),
    .B(net5227),
    .Y(_06240_));
 sg13g2_a21oi_1 _21402_ (.A1(net4905),
    .A2(net5227),
    .Y(_01998_),
    .B1(_06240_));
 sg13g2_nor2_1 _21403_ (.A(net1535),
    .B(net5222),
    .Y(_06241_));
 sg13g2_a21oi_1 _21404_ (.A1(net4774),
    .A2(net5222),
    .Y(_01999_),
    .B1(_06241_));
 sg13g2_nor2_1 _21405_ (.A(net2178),
    .B(net5224),
    .Y(_06242_));
 sg13g2_a21oi_1 _21406_ (.A1(net4900),
    .A2(net5224),
    .Y(_02000_),
    .B1(_06242_));
 sg13g2_nor2_1 _21407_ (.A(net1573),
    .B(net5224),
    .Y(_06243_));
 sg13g2_a21oi_1 _21408_ (.A1(net4963),
    .A2(net5224),
    .Y(_02001_),
    .B1(_06243_));
 sg13g2_nor2_1 _21409_ (.A(net2215),
    .B(net5219),
    .Y(_06244_));
 sg13g2_a21oi_1 _21410_ (.A1(net4956),
    .A2(net5219),
    .Y(_02002_),
    .B1(_06244_));
 sg13g2_nor2_1 _21411_ (.A(net1395),
    .B(net5225),
    .Y(_06245_));
 sg13g2_a21oi_1 _21412_ (.A1(net4896),
    .A2(net5225),
    .Y(_02003_),
    .B1(_06245_));
 sg13g2_nor2_1 _21413_ (.A(net1654),
    .B(net5224),
    .Y(_06246_));
 sg13g2_a21oi_1 _21414_ (.A1(net4891),
    .A2(net5224),
    .Y(_02004_),
    .B1(_06246_));
 sg13g2_nor2_1 _21415_ (.A(net1240),
    .B(net5220),
    .Y(_06247_));
 sg13g2_a21oi_1 _21416_ (.A1(net4884),
    .A2(net5220),
    .Y(_02005_),
    .B1(_06247_));
 sg13g2_nor2_1 _21417_ (.A(net1412),
    .B(net5224),
    .Y(_06248_));
 sg13g2_a21oi_1 _21418_ (.A1(net4770),
    .A2(net5224),
    .Y(_02006_),
    .B1(_06248_));
 sg13g2_nor2_1 _21419_ (.A(net1685),
    .B(net5226),
    .Y(_06249_));
 sg13g2_a21oi_1 _21420_ (.A1(net4879),
    .A2(net5226),
    .Y(_02007_),
    .B1(_06249_));
 sg13g2_nor2_1 _21421_ (.A(net1374),
    .B(net5227),
    .Y(_06250_));
 sg13g2_a21oi_1 _21422_ (.A1(net4872),
    .A2(net5227),
    .Y(_02008_),
    .B1(_06250_));
 sg13g2_nor2_1 _21423_ (.A(net1711),
    .B(net5228),
    .Y(_06251_));
 sg13g2_a21oi_1 _21424_ (.A1(net4765),
    .A2(net5228),
    .Y(_02009_),
    .B1(_06251_));
 sg13g2_nor2_1 _21425_ (.A(net1554),
    .B(net5219),
    .Y(_06252_));
 sg13g2_a21oi_1 _21426_ (.A1(net4870),
    .A2(net5219),
    .Y(_02010_),
    .B1(_06252_));
 sg13g2_nor2_1 _21427_ (.A(net1989),
    .B(net5229),
    .Y(_06253_));
 sg13g2_a21oi_1 _21428_ (.A1(net4864),
    .A2(net5228),
    .Y(_02011_),
    .B1(_06253_));
 sg13g2_nor2_1 _21429_ (.A(net1210),
    .B(net5220),
    .Y(_06254_));
 sg13g2_a21oi_1 _21430_ (.A1(net4857),
    .A2(net5220),
    .Y(_02012_),
    .B1(_06254_));
 sg13g2_nor2_1 _21431_ (.A(net1885),
    .B(net5219),
    .Y(_06255_));
 sg13g2_a21oi_1 _21432_ (.A1(net4854),
    .A2(net5219),
    .Y(_02013_),
    .B1(_06255_));
 sg13g2_nor2_1 _21433_ (.A(net1921),
    .B(net5226),
    .Y(_06256_));
 sg13g2_a21oi_1 _21434_ (.A1(net4849),
    .A2(net5226),
    .Y(_02014_),
    .B1(_06256_));
 sg13g2_nor2_1 _21435_ (.A(net1771),
    .B(net5220),
    .Y(_06257_));
 sg13g2_a21oi_1 _21436_ (.A1(net4845),
    .A2(net5220),
    .Y(_02015_),
    .B1(_06257_));
 sg13g2_nor2_1 _21437_ (.A(net1436),
    .B(net5223),
    .Y(_06258_));
 sg13g2_a21oi_1 _21438_ (.A1(net4838),
    .A2(net5220),
    .Y(_02016_),
    .B1(_06258_));
 sg13g2_nor2_1 _21439_ (.A(net1695),
    .B(net5222),
    .Y(_06259_));
 sg13g2_a21oi_1 _21440_ (.A1(net4834),
    .A2(net5222),
    .Y(_02017_),
    .B1(_06259_));
 sg13g2_nor2_1 _21441_ (.A(net1943),
    .B(net5227),
    .Y(_06260_));
 sg13g2_a21oi_1 _21442_ (.A1(net4831),
    .A2(net5227),
    .Y(_02018_),
    .B1(_06260_));
 sg13g2_nor2_1 _21443_ (.A(net2040),
    .B(net5227),
    .Y(_06261_));
 sg13g2_a21oi_1 _21444_ (.A1(net4822),
    .A2(net5227),
    .Y(_02019_),
    .B1(_06261_));
 sg13g2_nand3_1 _21445_ (.B(_05694_),
    .C(net6070),
    .A(_05660_),
    .Y(_06262_));
 sg13g2_nand2_1 _21446_ (.Y(_06263_),
    .A(net1423),
    .B(net5615));
 sg13g2_o21ai_1 _21447_ (.B1(_06263_),
    .Y(_02020_),
    .A1(net4998),
    .A2(net5615));
 sg13g2_nand2_1 _21448_ (.Y(_06264_),
    .A(net797),
    .B(net5615));
 sg13g2_o21ai_1 _21449_ (.B1(_06264_),
    .Y(_02021_),
    .A1(net4990),
    .A2(net5615));
 sg13g2_nand2_1 _21450_ (.Y(_06265_),
    .A(net1186),
    .B(net5615));
 sg13g2_o21ai_1 _21451_ (.B1(_06265_),
    .Y(_02022_),
    .A1(net4985),
    .A2(net5615));
 sg13g2_nand2_1 _21452_ (.Y(_06266_),
    .A(net636),
    .B(net5614));
 sg13g2_o21ai_1 _21453_ (.B1(_06266_),
    .Y(_02023_),
    .A1(net4983),
    .A2(net5614));
 sg13g2_nand2_1 _21454_ (.Y(_06267_),
    .A(net813),
    .B(net5618));
 sg13g2_o21ai_1 _21455_ (.B1(_06267_),
    .Y(_02024_),
    .A1(net4974),
    .A2(net5618));
 sg13g2_nand2_1 _21456_ (.Y(_06268_),
    .A(net919),
    .B(net5621));
 sg13g2_o21ai_1 _21457_ (.B1(_06268_),
    .Y(_02025_),
    .A1(net4969),
    .A2(net5621));
 sg13g2_nand2_1 _21458_ (.Y(_06269_),
    .A(net1003),
    .B(net5615));
 sg13g2_o21ai_1 _21459_ (.B1(_06269_),
    .Y(_02026_),
    .A1(net4966),
    .A2(net5616));
 sg13g2_nand2_1 _21460_ (.Y(_06270_),
    .A(net467),
    .B(net5620));
 sg13g2_o21ai_1 _21461_ (.B1(_06270_),
    .Y(_02027_),
    .A1(net4916),
    .A2(net5619));
 sg13g2_nand2_1 _21462_ (.Y(_06271_),
    .A(net1130),
    .B(net5621));
 sg13g2_o21ai_1 _21463_ (.B1(_06271_),
    .Y(_02028_),
    .A1(net4782),
    .A2(net5616));
 sg13g2_nand2_1 _21464_ (.Y(_06272_),
    .A(net448),
    .B(net5621));
 sg13g2_o21ai_1 _21465_ (.B1(_06272_),
    .Y(_02029_),
    .A1(net4912),
    .A2(net5621));
 sg13g2_nand2_1 _21466_ (.Y(_06273_),
    .A(net543),
    .B(net5623));
 sg13g2_o21ai_1 _21467_ (.B1(_06273_),
    .Y(_02030_),
    .A1(net4909),
    .A2(net5623));
 sg13g2_nand2_1 _21468_ (.Y(_06274_),
    .A(net707),
    .B(net5616));
 sg13g2_o21ai_1 _21469_ (.B1(_06274_),
    .Y(_02031_),
    .A1(net4775),
    .A2(net5615));
 sg13g2_nand2_1 _21470_ (.Y(_06275_),
    .A(net865),
    .B(net5619));
 sg13g2_o21ai_1 _21471_ (.B1(_06275_),
    .Y(_02032_),
    .A1(net4902),
    .A2(net5619));
 sg13g2_nand2_1 _21472_ (.Y(_06276_),
    .A(net1101),
    .B(net5619));
 sg13g2_o21ai_1 _21473_ (.B1(_06276_),
    .Y(_02033_),
    .A1(net4961),
    .A2(net5619));
 sg13g2_nand2_1 _21474_ (.Y(_06277_),
    .A(net1116),
    .B(net5613));
 sg13g2_o21ai_1 _21475_ (.B1(_06277_),
    .Y(_02034_),
    .A1(net4954),
    .A2(net5613));
 sg13g2_nand2_1 _21476_ (.Y(_06278_),
    .A(net512),
    .B(net5620));
 sg13g2_o21ai_1 _21477_ (.B1(_06278_),
    .Y(_02035_),
    .A1(net4895),
    .A2(net5619));
 sg13g2_nand2_1 _21478_ (.Y(_06279_),
    .A(net652),
    .B(net5618));
 sg13g2_o21ai_1 _21479_ (.B1(_06279_),
    .Y(_02036_),
    .A1(net4889),
    .A2(net5618));
 sg13g2_nand2_1 _21480_ (.Y(_06280_),
    .A(net402),
    .B(net5614));
 sg13g2_o21ai_1 _21481_ (.B1(_06280_),
    .Y(_02037_),
    .A1(net4888),
    .A2(net5614));
 sg13g2_nand2_1 _21482_ (.Y(_06281_),
    .A(net794),
    .B(net5619));
 sg13g2_o21ai_1 _21483_ (.B1(_06281_),
    .Y(_02038_),
    .A1(net4769),
    .A2(net5619));
 sg13g2_nand2_1 _21484_ (.Y(_06282_),
    .A(net1307),
    .B(net5618));
 sg13g2_o21ai_1 _21485_ (.B1(_06282_),
    .Y(_02039_),
    .A1(net4881),
    .A2(net5618));
 sg13g2_nand2_1 _21486_ (.Y(_06283_),
    .A(net1096),
    .B(net5622));
 sg13g2_o21ai_1 _21487_ (.B1(_06283_),
    .Y(_02040_),
    .A1(net4874),
    .A2(net5622));
 sg13g2_nand2_1 _21488_ (.Y(_06284_),
    .A(net754),
    .B(net5621));
 sg13g2_o21ai_1 _21489_ (.B1(_06284_),
    .Y(_02041_),
    .A1(net4765),
    .A2(net5622));
 sg13g2_nand2_1 _21490_ (.Y(_06285_),
    .A(net1296),
    .B(net5613));
 sg13g2_o21ai_1 _21491_ (.B1(_06285_),
    .Y(_02042_),
    .A1(_09734_),
    .A2(net5613));
 sg13g2_nand2_1 _21492_ (.Y(_06286_),
    .A(net1298),
    .B(net5622));
 sg13g2_o21ai_1 _21493_ (.B1(_06286_),
    .Y(_02043_),
    .A1(net4864),
    .A2(net5622));
 sg13g2_nand2_1 _21494_ (.Y(_06287_),
    .A(net609),
    .B(net5614));
 sg13g2_o21ai_1 _21495_ (.B1(_06287_),
    .Y(_02044_),
    .A1(net4860),
    .A2(net5614));
 sg13g2_nand2_1 _21496_ (.Y(_06288_),
    .A(net974),
    .B(net5613));
 sg13g2_o21ai_1 _21497_ (.B1(_06288_),
    .Y(_02045_),
    .A1(net4856),
    .A2(net5613));
 sg13g2_nand2_1 _21498_ (.Y(_06289_),
    .A(net1030),
    .B(net5620));
 sg13g2_o21ai_1 _21499_ (.B1(_06289_),
    .Y(_02046_),
    .A1(net4849),
    .A2(net5620));
 sg13g2_nand2_1 _21500_ (.Y(_06290_),
    .A(net1260),
    .B(net5613));
 sg13g2_o21ai_1 _21501_ (.B1(_06290_),
    .Y(_02047_),
    .A1(net4846),
    .A2(net5613));
 sg13g2_nand2_1 _21502_ (.Y(_06291_),
    .A(net545),
    .B(net5618));
 sg13g2_o21ai_1 _21503_ (.B1(_06291_),
    .Y(_02048_),
    .A1(net4839),
    .A2(net5618));
 sg13g2_nand2_1 _21504_ (.Y(_06292_),
    .A(net546),
    .B(net5616));
 sg13g2_o21ai_1 _21505_ (.B1(_06292_),
    .Y(_02049_),
    .A1(net4833),
    .A2(net5616));
 sg13g2_nand2_1 _21506_ (.Y(_06293_),
    .A(net481),
    .B(net5622));
 sg13g2_o21ai_1 _21507_ (.B1(_06293_),
    .Y(_02050_),
    .A1(_09799_),
    .A2(net5622));
 sg13g2_nand2_1 _21508_ (.Y(_06294_),
    .A(net576),
    .B(net5621));
 sg13g2_o21ai_1 _21509_ (.B1(_06294_),
    .Y(_02051_),
    .A1(net4822),
    .A2(net5621));
 sg13g2_and4_1 _21510_ (.A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .B(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .C(_05589_),
    .D(net6070),
    .X(_06295_));
 sg13g2_nor2_1 _21511_ (.A(net2399),
    .B(net5605),
    .Y(_06296_));
 sg13g2_a21oi_1 _21512_ (.A1(net4998),
    .A2(net5605),
    .Y(_02052_),
    .B1(_06296_));
 sg13g2_nor2_1 _21513_ (.A(net1666),
    .B(net5605),
    .Y(_06297_));
 sg13g2_a21oi_1 _21514_ (.A1(net4989),
    .A2(net5605),
    .Y(_02053_),
    .B1(_06297_));
 sg13g2_nor2_1 _21515_ (.A(net2012),
    .B(net5605),
    .Y(_06298_));
 sg13g2_a21oi_1 _21516_ (.A1(net4984),
    .A2(net5605),
    .Y(_02054_),
    .B1(_06298_));
 sg13g2_nor2_1 _21517_ (.A(net1540),
    .B(net5603),
    .Y(_06299_));
 sg13g2_a21oi_1 _21518_ (.A1(net4983),
    .A2(net5602),
    .Y(_02055_),
    .B1(_06299_));
 sg13g2_nor2_1 _21519_ (.A(net1877),
    .B(net5607),
    .Y(_06300_));
 sg13g2_a21oi_1 _21520_ (.A1(net4975),
    .A2(net5607),
    .Y(_02056_),
    .B1(_06300_));
 sg13g2_nor2_1 _21521_ (.A(net1586),
    .B(net5608),
    .Y(_06301_));
 sg13g2_a21oi_1 _21522_ (.A1(net4970),
    .A2(net5608),
    .Y(_02057_),
    .B1(_06301_));
 sg13g2_nor2_1 _21523_ (.A(net1907),
    .B(net5608),
    .Y(_06302_));
 sg13g2_a21oi_1 _21524_ (.A1(net4967),
    .A2(net5605),
    .Y(_02058_),
    .B1(_06302_));
 sg13g2_nor2_1 _21525_ (.A(net1349),
    .B(net5606),
    .Y(_06303_));
 sg13g2_a21oi_1 _21526_ (.A1(net4916),
    .A2(net5606),
    .Y(_02059_),
    .B1(_06303_));
 sg13g2_nor2_1 _21527_ (.A(net2370),
    .B(net5608),
    .Y(_06304_));
 sg13g2_a21oi_1 _21528_ (.A1(net4779),
    .A2(net5608),
    .Y(_02060_),
    .B1(_06304_));
 sg13g2_nor2_1 _21529_ (.A(net1926),
    .B(net5608),
    .Y(_06305_));
 sg13g2_a21oi_1 _21530_ (.A1(net4913),
    .A2(net5608),
    .Y(_02061_),
    .B1(_06305_));
 sg13g2_nor2_1 _21531_ (.A(net2257),
    .B(net5609),
    .Y(_06306_));
 sg13g2_a21oi_1 _21532_ (.A1(net4907),
    .A2(net5609),
    .Y(_02062_),
    .B1(_06306_));
 sg13g2_nor2_1 _21533_ (.A(net2226),
    .B(net5605),
    .Y(_06307_));
 sg13g2_a21oi_1 _21534_ (.A1(net4776),
    .A2(net5612),
    .Y(_02063_),
    .B1(_06307_));
 sg13g2_nor2_1 _21535_ (.A(net1680),
    .B(net5611),
    .Y(_06308_));
 sg13g2_a21oi_1 _21536_ (.A1(net4901),
    .A2(net5611),
    .Y(_02064_),
    .B1(_06308_));
 sg13g2_nor2_1 _21537_ (.A(net1767),
    .B(net5606),
    .Y(_06309_));
 sg13g2_a21oi_1 _21538_ (.A1(net4962),
    .A2(net5606),
    .Y(_02065_),
    .B1(_06309_));
 sg13g2_nor2_1 _21539_ (.A(net2203),
    .B(net5602),
    .Y(_06310_));
 sg13g2_a21oi_1 _21540_ (.A1(net4955),
    .A2(net5602),
    .Y(_02066_),
    .B1(_06310_));
 sg13g2_nor2_1 _21541_ (.A(net1894),
    .B(net5606),
    .Y(_06311_));
 sg13g2_a21oi_1 _21542_ (.A1(net4894),
    .A2(net5611),
    .Y(_02067_),
    .B1(_06311_));
 sg13g2_nor2_1 _21543_ (.A(net1899),
    .B(net5606),
    .Y(_06312_));
 sg13g2_a21oi_1 _21544_ (.A1(net4892),
    .A2(net5607),
    .Y(_02068_),
    .B1(_06312_));
 sg13g2_nor2_1 _21545_ (.A(net1937),
    .B(net5603),
    .Y(_06313_));
 sg13g2_a21oi_1 _21546_ (.A1(net4888),
    .A2(net5603),
    .Y(_02069_),
    .B1(_06313_));
 sg13g2_nor2_1 _21547_ (.A(net1337),
    .B(net5606),
    .Y(_06314_));
 sg13g2_a21oi_1 _21548_ (.A1(net4768),
    .A2(net5606),
    .Y(_02070_),
    .B1(_06314_));
 sg13g2_nor2_1 _21549_ (.A(net1962),
    .B(net5607),
    .Y(_06315_));
 sg13g2_a21oi_1 _21550_ (.A1(net4882),
    .A2(net5607),
    .Y(_02071_),
    .B1(_06315_));
 sg13g2_nor2_1 _21551_ (.A(net1347),
    .B(net5609),
    .Y(_06316_));
 sg13g2_a21oi_1 _21552_ (.A1(net4875),
    .A2(net5609),
    .Y(_02072_),
    .B1(_06316_));
 sg13g2_nor2_1 _21553_ (.A(net2104),
    .B(net5608),
    .Y(_06317_));
 sg13g2_a21oi_1 _21554_ (.A1(net4766),
    .A2(net5610),
    .Y(_02073_),
    .B1(_06317_));
 sg13g2_nor2_1 _21555_ (.A(net1419),
    .B(net5602),
    .Y(_06318_));
 sg13g2_a21oi_1 _21556_ (.A1(net4869),
    .A2(net5602),
    .Y(_02074_),
    .B1(_06318_));
 sg13g2_nor2_1 _21557_ (.A(net2500),
    .B(net5609),
    .Y(_06319_));
 sg13g2_a21oi_1 _21558_ (.A1(net4864),
    .A2(net5609),
    .Y(_02075_),
    .B1(_06319_));
 sg13g2_nor2_1 _21559_ (.A(net1172),
    .B(net5603),
    .Y(_06320_));
 sg13g2_a21oi_1 _21560_ (.A1(net4860),
    .A2(net5604),
    .Y(_02076_),
    .B1(_06320_));
 sg13g2_nor2_1 _21561_ (.A(net1600),
    .B(net5602),
    .Y(_06321_));
 sg13g2_a21oi_1 _21562_ (.A1(net4856),
    .A2(net5602),
    .Y(_02077_),
    .B1(_06321_));
 sg13g2_nor2_1 _21563_ (.A(net1818),
    .B(net5607),
    .Y(_06322_));
 sg13g2_a21oi_1 _21564_ (.A1(net4847),
    .A2(net5607),
    .Y(_02078_),
    .B1(_06322_));
 sg13g2_nor2_1 _21565_ (.A(net1487),
    .B(net5602),
    .Y(_06323_));
 sg13g2_a21oi_1 _21566_ (.A1(net4846),
    .A2(net5604),
    .Y(_02079_),
    .B1(_06323_));
 sg13g2_nor2_1 _21567_ (.A(net1643),
    .B(net5603),
    .Y(_06324_));
 sg13g2_a21oi_1 _21568_ (.A1(net4839),
    .A2(net5603),
    .Y(_02080_),
    .B1(_06324_));
 sg13g2_nor2_1 _21569_ (.A(net1897),
    .B(net5603),
    .Y(_06325_));
 sg13g2_a21oi_1 _21570_ (.A1(net4833),
    .A2(net5603),
    .Y(_02081_),
    .B1(_06325_));
 sg13g2_nor2_1 _21571_ (.A(net2163),
    .B(net5610),
    .Y(_06326_));
 sg13g2_a21oi_1 _21572_ (.A1(net4830),
    .A2(net5610),
    .Y(_02082_),
    .B1(_06326_));
 sg13g2_nor2_1 _21573_ (.A(net1550),
    .B(net5609),
    .Y(_06327_));
 sg13g2_a21oi_1 _21574_ (.A1(net4822),
    .A2(net5609),
    .Y(_02083_),
    .B1(_06327_));
 sg13g2_nor2_2 _21575_ (.A(_05591_),
    .B(_05896_),
    .Y(_06328_));
 sg13g2_nor2_1 _21576_ (.A(net2026),
    .B(net5211),
    .Y(_06329_));
 sg13g2_a21oi_1 _21577_ (.A1(net4996),
    .A2(net5211),
    .Y(_02084_),
    .B1(_06329_));
 sg13g2_nor2_1 _21578_ (.A(net1506),
    .B(net5211),
    .Y(_06330_));
 sg13g2_a21oi_1 _21579_ (.A1(net4991),
    .A2(net5211),
    .Y(_02085_),
    .B1(_06330_));
 sg13g2_nor2_1 _21580_ (.A(net1814),
    .B(net5211),
    .Y(_06331_));
 sg13g2_a21oi_1 _21581_ (.A1(net4986),
    .A2(net5211),
    .Y(_02086_),
    .B1(_06331_));
 sg13g2_nor2_1 _21582_ (.A(net1524),
    .B(net5209),
    .Y(_06332_));
 sg13g2_a21oi_1 _21583_ (.A1(net4983),
    .A2(net5209),
    .Y(_02087_),
    .B1(_06332_));
 sg13g2_nor2_1 _21584_ (.A(net2395),
    .B(net5210),
    .Y(_06333_));
 sg13g2_a21oi_1 _21585_ (.A1(net4974),
    .A2(net5210),
    .Y(_02088_),
    .B1(_06333_));
 sg13g2_nor2_1 _21586_ (.A(net2404),
    .B(net5217),
    .Y(_06334_));
 sg13g2_a21oi_1 _21587_ (.A1(net4970),
    .A2(net5217),
    .Y(_02089_),
    .B1(_06334_));
 sg13g2_nor2_1 _21588_ (.A(net1706),
    .B(net5211),
    .Y(_06335_));
 sg13g2_a21oi_1 _21589_ (.A1(net4965),
    .A2(net5212),
    .Y(_02090_),
    .B1(_06335_));
 sg13g2_nor2_1 _21590_ (.A(net1629),
    .B(net5215),
    .Y(_06336_));
 sg13g2_a21oi_1 _21591_ (.A1(net4918),
    .A2(net5215),
    .Y(_02091_),
    .B1(_06336_));
 sg13g2_nor2_1 _21592_ (.A(net1409),
    .B(net5211),
    .Y(_06337_));
 sg13g2_a21oi_1 _21593_ (.A1(net4781),
    .A2(net5212),
    .Y(_02092_),
    .B1(_06337_));
 sg13g2_nor2_1 _21594_ (.A(net1475),
    .B(net5217),
    .Y(_06338_));
 sg13g2_a21oi_1 _21595_ (.A1(net4913),
    .A2(net5217),
    .Y(_02093_),
    .B1(_06338_));
 sg13g2_nor2_1 _21596_ (.A(net1584),
    .B(net5216),
    .Y(_06339_));
 sg13g2_a21oi_1 _21597_ (.A1(net4905),
    .A2(net5216),
    .Y(_02094_),
    .B1(_06339_));
 sg13g2_nor2_1 _21598_ (.A(net1735),
    .B(net5212),
    .Y(_06340_));
 sg13g2_a21oi_1 _21599_ (.A1(net4774),
    .A2(net5212),
    .Y(_02095_),
    .B1(_06340_));
 sg13g2_nor2_1 _21600_ (.A(net1682),
    .B(net5218),
    .Y(_06341_));
 sg13g2_a21oi_1 _21601_ (.A1(net4901),
    .A2(net5215),
    .Y(_02096_),
    .B1(_06341_));
 sg13g2_nor2_1 _21602_ (.A(net1663),
    .B(net5214),
    .Y(_06342_));
 sg13g2_a21oi_1 _21603_ (.A1(net4962),
    .A2(net5214),
    .Y(_02097_),
    .B1(_06342_));
 sg13g2_nor2_1 _21604_ (.A(net1661),
    .B(net5209),
    .Y(_06343_));
 sg13g2_a21oi_1 _21605_ (.A1(net4956),
    .A2(net5209),
    .Y(_02098_),
    .B1(_06343_));
 sg13g2_nor2_1 _21606_ (.A(net1755),
    .B(net5214),
    .Y(_06344_));
 sg13g2_a21oi_1 _21607_ (.A1(net4898),
    .A2(net5214),
    .Y(_02099_),
    .B1(_06344_));
 sg13g2_nor2_1 _21608_ (.A(net1422),
    .B(net5214),
    .Y(_06345_));
 sg13g2_a21oi_1 _21609_ (.A1(net4892),
    .A2(net5214),
    .Y(_02100_),
    .B1(_06345_));
 sg13g2_nor2_1 _21610_ (.A(net1681),
    .B(net5210),
    .Y(_06346_));
 sg13g2_a21oi_1 _21611_ (.A1(net4888),
    .A2(net5210),
    .Y(_02101_),
    .B1(_06346_));
 sg13g2_nor2_1 _21612_ (.A(net2155),
    .B(net5214),
    .Y(_06347_));
 sg13g2_a21oi_1 _21613_ (.A1(net4768),
    .A2(net5214),
    .Y(_02102_),
    .B1(_06347_));
 sg13g2_nor2_1 _21614_ (.A(net1763),
    .B(net5215),
    .Y(_06348_));
 sg13g2_a21oi_1 _21615_ (.A1(net4881),
    .A2(net5215),
    .Y(_02103_),
    .B1(_06348_));
 sg13g2_nor2_1 _21616_ (.A(net2000),
    .B(net5216),
    .Y(_06349_));
 sg13g2_a21oi_1 _21617_ (.A1(net4874),
    .A2(net5216),
    .Y(_02104_),
    .B1(_06349_));
 sg13g2_nor2_1 _21618_ (.A(net1585),
    .B(net5217),
    .Y(_06350_));
 sg13g2_a21oi_1 _21619_ (.A1(net4765),
    .A2(net5217),
    .Y(_02105_),
    .B1(_06350_));
 sg13g2_nor2_1 _21620_ (.A(net1793),
    .B(net5209),
    .Y(_06351_));
 sg13g2_a21oi_1 _21621_ (.A1(net4869),
    .A2(net5209),
    .Y(_02106_),
    .B1(_06351_));
 sg13g2_nor2_1 _21622_ (.A(net1699),
    .B(net5216),
    .Y(_06352_));
 sg13g2_a21oi_1 _21623_ (.A1(net4863),
    .A2(net5216),
    .Y(_02107_),
    .B1(_06352_));
 sg13g2_nor2_1 _21624_ (.A(net1578),
    .B(net5210),
    .Y(_06353_));
 sg13g2_a21oi_1 _21625_ (.A1(net4859),
    .A2(net5213),
    .Y(_02108_),
    .B1(_06353_));
 sg13g2_nor2_1 _21626_ (.A(net1659),
    .B(net5209),
    .Y(_06354_));
 sg13g2_a21oi_1 _21627_ (.A1(net4854),
    .A2(net5209),
    .Y(_02109_),
    .B1(_06354_));
 sg13g2_nor2_1 _21628_ (.A(net1626),
    .B(net5215),
    .Y(_06355_));
 sg13g2_a21oi_1 _21629_ (.A1(net4850),
    .A2(net5215),
    .Y(_02110_),
    .B1(_06355_));
 sg13g2_nor2_1 _21630_ (.A(net1713),
    .B(net5210),
    .Y(_06356_));
 sg13g2_a21oi_1 _21631_ (.A1(net4844),
    .A2(net5210),
    .Y(_02111_),
    .B1(_06356_));
 sg13g2_nor2_1 _21632_ (.A(net2450),
    .B(net5213),
    .Y(_06357_));
 sg13g2_a21oi_1 _21633_ (.A1(net4840),
    .A2(net5213),
    .Y(_02112_),
    .B1(_06357_));
 sg13g2_nor2_1 _21634_ (.A(net2320),
    .B(net5212),
    .Y(_06358_));
 sg13g2_a21oi_1 _21635_ (.A1(net4833),
    .A2(net5212),
    .Y(_02113_),
    .B1(_06358_));
 sg13g2_nor2_1 _21636_ (.A(net1300),
    .B(net5218),
    .Y(_06359_));
 sg13g2_a21oi_1 _21637_ (.A1(net4828),
    .A2(net5217),
    .Y(_02114_),
    .B1(_06359_));
 sg13g2_nor2_1 _21638_ (.A(net1635),
    .B(net5216),
    .Y(_06360_));
 sg13g2_a21oi_1 _21639_ (.A1(net4822),
    .A2(net5216),
    .Y(_02115_),
    .B1(_06360_));
 sg13g2_and3_2 _21640_ (.X(_06361_),
    .A(net6096),
    .B(_09507_),
    .C(_05589_));
 sg13g2_nor2_1 _21641_ (.A(net2059),
    .B(net5394),
    .Y(_06362_));
 sg13g2_a21oi_1 _21642_ (.A1(net4996),
    .A2(net5394),
    .Y(_02116_),
    .B1(_06362_));
 sg13g2_nor2_1 _21643_ (.A(net1963),
    .B(net5394),
    .Y(_06363_));
 sg13g2_a21oi_1 _21644_ (.A1(net4992),
    .A2(net5394),
    .Y(_02117_),
    .B1(_06363_));
 sg13g2_nor2_1 _21645_ (.A(net1970),
    .B(net5393),
    .Y(_06364_));
 sg13g2_a21oi_1 _21646_ (.A1(net4988),
    .A2(net5393),
    .Y(_02118_),
    .B1(_06364_));
 sg13g2_nor2_1 _21647_ (.A(net2596),
    .B(net5391),
    .Y(_06365_));
 sg13g2_a21oi_1 _21648_ (.A1(net4981),
    .A2(net5391),
    .Y(_02119_),
    .B1(_06365_));
 sg13g2_nor2_1 _21649_ (.A(net2522),
    .B(net5397),
    .Y(_06366_));
 sg13g2_a21oi_1 _21650_ (.A1(net4976),
    .A2(net5392),
    .Y(_02120_),
    .B1(_06366_));
 sg13g2_nor2_1 _21651_ (.A(net2498),
    .B(net5398),
    .Y(_06367_));
 sg13g2_a21oi_1 _21652_ (.A1(net4969),
    .A2(net5398),
    .Y(_02121_),
    .B1(_06367_));
 sg13g2_nor2_1 _21653_ (.A(net1516),
    .B(net5393),
    .Y(_06368_));
 sg13g2_a21oi_1 _21654_ (.A1(net4966),
    .A2(net5393),
    .Y(_02122_),
    .B1(_06368_));
 sg13g2_nor2_1 _21655_ (.A(net2457),
    .B(net5396),
    .Y(_06369_));
 sg13g2_a21oi_1 _21656_ (.A1(net4917),
    .A2(net5396),
    .Y(_02123_),
    .B1(_06369_));
 sg13g2_nor2_1 _21657_ (.A(net2048),
    .B(net5393),
    .Y(_06370_));
 sg13g2_a21oi_1 _21658_ (.A1(net4781),
    .A2(net5393),
    .Y(_02124_),
    .B1(_06370_));
 sg13g2_nor2_1 _21659_ (.A(net1308),
    .B(net5398),
    .Y(_06371_));
 sg13g2_a21oi_1 _21660_ (.A1(net4915),
    .A2(net5398),
    .Y(_02125_),
    .B1(_06371_));
 sg13g2_nor2_1 _21661_ (.A(net2548),
    .B(net5399),
    .Y(_06372_));
 sg13g2_a21oi_1 _21662_ (.A1(net4907),
    .A2(net5399),
    .Y(_02126_),
    .B1(_06372_));
 sg13g2_nor2_1 _21663_ (.A(net2277),
    .B(net5394),
    .Y(_06373_));
 sg13g2_a21oi_1 _21664_ (.A1(net4775),
    .A2(net5394),
    .Y(_02127_),
    .B1(_06373_));
 sg13g2_nor2_1 _21665_ (.A(net2267),
    .B(net5396),
    .Y(_06374_));
 sg13g2_a21oi_1 _21666_ (.A1(net4901),
    .A2(net5396),
    .Y(_02128_),
    .B1(_06374_));
 sg13g2_nor2_1 _21667_ (.A(net1356),
    .B(net5396),
    .Y(_06375_));
 sg13g2_a21oi_1 _21668_ (.A1(net4961),
    .A2(net5396),
    .Y(_02129_),
    .B1(_06375_));
 sg13g2_nor2_1 _21669_ (.A(net2183),
    .B(net5391),
    .Y(_06376_));
 sg13g2_a21oi_1 _21670_ (.A1(net4957),
    .A2(net5391),
    .Y(_02130_),
    .B1(_06376_));
 sg13g2_nor2_1 _21671_ (.A(net2159),
    .B(net5400),
    .Y(_06377_));
 sg13g2_a21oi_1 _21672_ (.A1(net4897),
    .A2(net5400),
    .Y(_02131_),
    .B1(_06377_));
 sg13g2_nor2_1 _21673_ (.A(net1465),
    .B(net5397),
    .Y(_06378_));
 sg13g2_a21oi_1 _21674_ (.A1(net4893),
    .A2(net5397),
    .Y(_02132_),
    .B1(_06378_));
 sg13g2_nor2_1 _21675_ (.A(net2351),
    .B(net5392),
    .Y(_06379_));
 sg13g2_a21oi_1 _21676_ (.A1(net4886),
    .A2(net5392),
    .Y(_02133_),
    .B1(_06379_));
 sg13g2_nor2_1 _21677_ (.A(net2177),
    .B(net5396),
    .Y(_06380_));
 sg13g2_a21oi_1 _21678_ (.A1(net4768),
    .A2(net5396),
    .Y(_02134_),
    .B1(_06380_));
 sg13g2_nor2_1 _21679_ (.A(net1809),
    .B(net5397),
    .Y(_06381_));
 sg13g2_a21oi_1 _21680_ (.A1(net4878),
    .A2(net5397),
    .Y(_02135_),
    .B1(_06381_));
 sg13g2_nor2_1 _21681_ (.A(net1757),
    .B(net5399),
    .Y(_06382_));
 sg13g2_a21oi_1 _21682_ (.A1(net4877),
    .A2(net5399),
    .Y(_02136_),
    .B1(_06382_));
 sg13g2_nor2_1 _21683_ (.A(net1925),
    .B(net5398),
    .Y(_06383_));
 sg13g2_a21oi_1 _21684_ (.A1(net4765),
    .A2(net5398),
    .Y(_02137_),
    .B1(_06383_));
 sg13g2_nor2_1 _21685_ (.A(net1460),
    .B(net5391),
    .Y(_06384_));
 sg13g2_a21oi_1 _21686_ (.A1(net4868),
    .A2(net5391),
    .Y(_02138_),
    .B1(_06384_));
 sg13g2_nor2_1 _21687_ (.A(net2239),
    .B(net5399),
    .Y(_06385_));
 sg13g2_a21oi_1 _21688_ (.A1(net4863),
    .A2(net5399),
    .Y(_02139_),
    .B1(_06385_));
 sg13g2_nor2_1 _21689_ (.A(net1440),
    .B(net5395),
    .Y(_06386_));
 sg13g2_a21oi_1 _21690_ (.A1(net4857),
    .A2(net5395),
    .Y(_02140_),
    .B1(_06386_));
 sg13g2_nor2_1 _21691_ (.A(net1956),
    .B(net5391),
    .Y(_06387_));
 sg13g2_a21oi_1 _21692_ (.A1(net4854),
    .A2(net5391),
    .Y(_02141_),
    .B1(_06387_));
 sg13g2_nor2_1 _21693_ (.A(net1450),
    .B(net5397),
    .Y(_06388_));
 sg13g2_a21oi_1 _21694_ (.A1(net4850),
    .A2(net5397),
    .Y(_02142_),
    .B1(_06388_));
 sg13g2_nor2_1 _21695_ (.A(net1559),
    .B(net5392),
    .Y(_06389_));
 sg13g2_a21oi_1 _21696_ (.A1(net4843),
    .A2(net5392),
    .Y(_02143_),
    .B1(_06389_));
 sg13g2_nor2_1 _21697_ (.A(net1714),
    .B(net5392),
    .Y(_06390_));
 sg13g2_a21oi_1 _21698_ (.A1(net4838),
    .A2(net5392),
    .Y(_02144_),
    .B1(_06390_));
 sg13g2_nor2_1 _21699_ (.A(net2051),
    .B(net5393),
    .Y(_06391_));
 sg13g2_a21oi_1 _21700_ (.A1(net4832),
    .A2(net5393),
    .Y(_02145_),
    .B1(_06391_));
 sg13g2_nor2_1 _21701_ (.A(net1792),
    .B(net5399),
    .Y(_06392_));
 sg13g2_a21oi_1 _21702_ (.A1(net4830),
    .A2(net5399),
    .Y(_02146_),
    .B1(_06392_));
 sg13g2_nor2_1 _21703_ (.A(net1306),
    .B(net5398),
    .Y(_06393_));
 sg13g2_a21oi_1 _21704_ (.A1(net4823),
    .A2(net5398),
    .Y(_02147_),
    .B1(_06393_));
 sg13g2_nor2_1 _21705_ (.A(_05626_),
    .B(_05896_),
    .Y(_06394_));
 sg13g2_nor2_1 _21706_ (.A(net2004),
    .B(net5201),
    .Y(_06395_));
 sg13g2_a21oi_1 _21707_ (.A1(net4996),
    .A2(net5201),
    .Y(_02148_),
    .B1(_06395_));
 sg13g2_nor2_1 _21708_ (.A(net2019),
    .B(net5201),
    .Y(_06396_));
 sg13g2_a21oi_1 _21709_ (.A1(net4991),
    .A2(net5201),
    .Y(_02149_),
    .B1(_06396_));
 sg13g2_nor2_1 _21710_ (.A(net1523),
    .B(net5201),
    .Y(_06397_));
 sg13g2_a21oi_1 _21711_ (.A1(net4987),
    .A2(net5201),
    .Y(_02150_),
    .B1(_06397_));
 sg13g2_nor2_1 _21712_ (.A(net1754),
    .B(net5198),
    .Y(_06398_));
 sg13g2_a21oi_1 _21713_ (.A1(net4979),
    .A2(net5198),
    .Y(_02151_),
    .B1(_06398_));
 sg13g2_nor2_1 _21714_ (.A(net1955),
    .B(net5204),
    .Y(_06399_));
 sg13g2_a21oi_1 _21715_ (.A1(net4974),
    .A2(net5204),
    .Y(_02152_),
    .B1(_06399_));
 sg13g2_nor2_1 _21716_ (.A(net2197),
    .B(net5205),
    .Y(_06400_));
 sg13g2_a21oi_1 _21717_ (.A1(net4972),
    .A2(net5205),
    .Y(_02153_),
    .B1(_06400_));
 sg13g2_nor2_1 _21718_ (.A(net1344),
    .B(net5202),
    .Y(_06401_));
 sg13g2_a21oi_1 _21719_ (.A1(net4964),
    .A2(net5202),
    .Y(_02154_),
    .B1(_06401_));
 sg13g2_nor2_1 _21720_ (.A(net1435),
    .B(net5203),
    .Y(_06402_));
 sg13g2_a21oi_1 _21721_ (.A1(net4916),
    .A2(net5203),
    .Y(_02155_),
    .B1(_06402_));
 sg13g2_nor2_1 _21722_ (.A(net1551),
    .B(net5202),
    .Y(_06403_));
 sg13g2_a21oi_1 _21723_ (.A1(net4781),
    .A2(net5202),
    .Y(_02156_),
    .B1(_06403_));
 sg13g2_nor2_1 _21724_ (.A(net1997),
    .B(net5205),
    .Y(_06404_));
 sg13g2_a21oi_1 _21725_ (.A1(net4914),
    .A2(net5205),
    .Y(_02157_),
    .B1(_06404_));
 sg13g2_nor2_1 _21726_ (.A(net2132),
    .B(net5206),
    .Y(_06405_));
 sg13g2_a21oi_1 _21727_ (.A1(net4907),
    .A2(net5206),
    .Y(_02158_),
    .B1(_06405_));
 sg13g2_nor2_1 _21728_ (.A(net1990),
    .B(net5202),
    .Y(_06406_));
 sg13g2_a21oi_1 _21729_ (.A1(net4776),
    .A2(net5202),
    .Y(_02159_),
    .B1(_06406_));
 sg13g2_nor2_1 _21730_ (.A(net1788),
    .B(net5203),
    .Y(_06407_));
 sg13g2_a21oi_1 _21731_ (.A1(net4902),
    .A2(net5203),
    .Y(_02160_),
    .B1(_06407_));
 sg13g2_nor2_1 _21732_ (.A(net1633),
    .B(net5203),
    .Y(_06408_));
 sg13g2_a21oi_1 _21733_ (.A1(net4963),
    .A2(net5203),
    .Y(_02161_),
    .B1(_06408_));
 sg13g2_nor2_1 _21734_ (.A(net1691),
    .B(net5198),
    .Y(_06409_));
 sg13g2_a21oi_1 _21735_ (.A1(net4956),
    .A2(net5198),
    .Y(_02162_),
    .B1(_06409_));
 sg13g2_nor2_1 _21736_ (.A(net1507),
    .B(net5207),
    .Y(_06410_));
 sg13g2_a21oi_1 _21737_ (.A1(net4896),
    .A2(net5204),
    .Y(_02163_),
    .B1(_06410_));
 sg13g2_nor2_1 _21738_ (.A(net1243),
    .B(net5204),
    .Y(_06411_));
 sg13g2_a21oi_1 _21739_ (.A1(net4891),
    .A2(net5204),
    .Y(_02164_),
    .B1(_06411_));
 sg13g2_nor2_1 _21740_ (.A(net1531),
    .B(net5200),
    .Y(_06412_));
 sg13g2_a21oi_1 _21741_ (.A1(net4884),
    .A2(net5200),
    .Y(_02165_),
    .B1(_06412_));
 sg13g2_nor2_1 _21742_ (.A(net1728),
    .B(net5203),
    .Y(_06413_));
 sg13g2_a21oi_1 _21743_ (.A1(net4770),
    .A2(net5203),
    .Y(_02166_),
    .B1(_06413_));
 sg13g2_nor2_1 _21744_ (.A(net2222),
    .B(net5200),
    .Y(_06414_));
 sg13g2_a21oi_1 _21745_ (.A1(net4879),
    .A2(net5200),
    .Y(_02167_),
    .B1(_06414_));
 sg13g2_nor2_1 _21746_ (.A(net1476),
    .B(net5206),
    .Y(_06415_));
 sg13g2_a21oi_1 _21747_ (.A1(net4874),
    .A2(net5206),
    .Y(_02168_),
    .B1(_06415_));
 sg13g2_nor2_1 _21748_ (.A(net2091),
    .B(net5205),
    .Y(_06416_));
 sg13g2_a21oi_1 _21749_ (.A1(net4764),
    .A2(net5205),
    .Y(_02169_),
    .B1(_06416_));
 sg13g2_nor2_1 _21750_ (.A(net1352),
    .B(net5198),
    .Y(_06417_));
 sg13g2_a21oi_1 _21751_ (.A1(net4869),
    .A2(net5198),
    .Y(_02170_),
    .B1(_06417_));
 sg13g2_nor2_1 _21752_ (.A(net1647),
    .B(net5206),
    .Y(_06418_));
 sg13g2_a21oi_1 _21753_ (.A1(net4863),
    .A2(net5206),
    .Y(_02171_),
    .B1(_06418_));
 sg13g2_nor2_1 _21754_ (.A(net1721),
    .B(net5199),
    .Y(_06419_));
 sg13g2_a21oi_1 _21755_ (.A1(net4861),
    .A2(net5199),
    .Y(_02172_),
    .B1(_06419_));
 sg13g2_nor2_1 _21756_ (.A(net1502),
    .B(net5198),
    .Y(_06420_));
 sg13g2_a21oi_1 _21757_ (.A1(net4855),
    .A2(net5198),
    .Y(_02173_),
    .B1(_06420_));
 sg13g2_nor2_1 _21758_ (.A(net1675),
    .B(net5204),
    .Y(_06421_));
 sg13g2_a21oi_1 _21759_ (.A1(net4849),
    .A2(net5204),
    .Y(_02174_),
    .B1(_06421_));
 sg13g2_nor2_1 _21760_ (.A(net1474),
    .B(net5199),
    .Y(_06422_));
 sg13g2_a21oi_1 _21761_ (.A1(net4845),
    .A2(net5199),
    .Y(_02175_),
    .B1(_06422_));
 sg13g2_nor2_1 _21762_ (.A(net1185),
    .B(net5200),
    .Y(_06423_));
 sg13g2_a21oi_1 _21763_ (.A1(net4838),
    .A2(net5200),
    .Y(_02176_),
    .B1(_06423_));
 sg13g2_nor2_1 _21764_ (.A(net1431),
    .B(net5201),
    .Y(_06424_));
 sg13g2_a21oi_1 _21765_ (.A1(net4832),
    .A2(net5201),
    .Y(_02177_),
    .B1(_06424_));
 sg13g2_nor2_1 _21766_ (.A(net2170),
    .B(net5206),
    .Y(_06425_));
 sg13g2_a21oi_1 _21767_ (.A1(net4830),
    .A2(net5206),
    .Y(_02178_),
    .B1(_06425_));
 sg13g2_nor2_1 _21768_ (.A(net1690),
    .B(net5205),
    .Y(_06426_));
 sg13g2_a21oi_1 _21769_ (.A1(net4823),
    .A2(net5205),
    .Y(_02179_),
    .B1(_06426_));
 sg13g2_nand3_1 _21770_ (.B(_05660_),
    .C(net6070),
    .A(_05589_),
    .Y(_06427_));
 sg13g2_nand2_1 _21771_ (.Y(_06428_),
    .A(net1168),
    .B(net5594));
 sg13g2_o21ai_1 _21772_ (.B1(_06428_),
    .Y(_02180_),
    .A1(net4994),
    .A2(net5594));
 sg13g2_nand2_1 _21773_ (.Y(_06429_),
    .A(net925),
    .B(net5594));
 sg13g2_o21ai_1 _21774_ (.B1(_06429_),
    .Y(_02181_),
    .A1(net4991),
    .A2(net5594));
 sg13g2_nand2_1 _21775_ (.Y(_06430_),
    .A(net1062),
    .B(net5593));
 sg13g2_o21ai_1 _21776_ (.B1(_06430_),
    .Y(_02182_),
    .A1(net4986),
    .A2(net5594));
 sg13g2_nand2_1 _21777_ (.Y(_06431_),
    .A(net650),
    .B(net5591));
 sg13g2_o21ai_1 _21778_ (.B1(_06431_),
    .Y(_02183_),
    .A1(net4983),
    .A2(net5592));
 sg13g2_nand2_1 _21779_ (.Y(_06432_),
    .A(net1534),
    .B(net5597));
 sg13g2_o21ai_1 _21780_ (.B1(_06432_),
    .Y(_02184_),
    .A1(net4978),
    .A2(net5597));
 sg13g2_nand2_1 _21781_ (.Y(_06433_),
    .A(net1286),
    .B(net5600));
 sg13g2_o21ai_1 _21782_ (.B1(_06433_),
    .Y(_02185_),
    .A1(net4972),
    .A2(net5600));
 sg13g2_nand2_1 _21783_ (.Y(_06434_),
    .A(net911),
    .B(net5600));
 sg13g2_o21ai_1 _21784_ (.B1(_06434_),
    .Y(_02186_),
    .A1(net4968),
    .A2(net5593));
 sg13g2_nand2_1 _21785_ (.Y(_06435_),
    .A(net633),
    .B(net5596));
 sg13g2_o21ai_1 _21786_ (.B1(_06435_),
    .Y(_02187_),
    .A1(net4916),
    .A2(net5596));
 sg13g2_nand2_1 _21787_ (.Y(_06436_),
    .A(net767),
    .B(net5593));
 sg13g2_o21ai_1 _21788_ (.B1(_06436_),
    .Y(_02188_),
    .A1(net4779),
    .A2(net5593));
 sg13g2_nand2_1 _21789_ (.Y(_06437_),
    .A(net1067),
    .B(net5598));
 sg13g2_o21ai_1 _21790_ (.B1(_06437_),
    .Y(_02189_),
    .A1(net4912),
    .A2(net5598));
 sg13g2_nand2_1 _21791_ (.Y(_06438_),
    .A(net890),
    .B(net5598));
 sg13g2_o21ai_1 _21792_ (.B1(_06438_),
    .Y(_02190_),
    .A1(net4905),
    .A2(net5598));
 sg13g2_nand2_1 _21793_ (.Y(_06439_),
    .A(net756),
    .B(net5593));
 sg13g2_o21ai_1 _21794_ (.B1(_06439_),
    .Y(_02191_),
    .A1(net4774),
    .A2(net5593));
 sg13g2_nand2_1 _21795_ (.Y(_06440_),
    .A(net564),
    .B(net5596));
 sg13g2_o21ai_1 _21796_ (.B1(_06440_),
    .Y(_02192_),
    .A1(net4899),
    .A2(net5596));
 sg13g2_nand2_1 _21797_ (.Y(_06441_),
    .A(net1354),
    .B(net5595));
 sg13g2_o21ai_1 _21798_ (.B1(_06441_),
    .Y(_02193_),
    .A1(net4959),
    .A2(net5595));
 sg13g2_nand2_1 _21799_ (.Y(_06442_),
    .A(net1522),
    .B(net5591));
 sg13g2_o21ai_1 _21800_ (.B1(_06442_),
    .Y(_02194_),
    .A1(net4955),
    .A2(net5591));
 sg13g2_nand2_1 _21801_ (.Y(_06443_),
    .A(net607),
    .B(net5596));
 sg13g2_o21ai_1 _21802_ (.B1(_06443_),
    .Y(_02195_),
    .A1(net4896),
    .A2(net5596));
 sg13g2_nand2_1 _21803_ (.Y(_06444_),
    .A(net983),
    .B(net5595));
 sg13g2_o21ai_1 _21804_ (.B1(_06444_),
    .Y(_02196_),
    .A1(net4892),
    .A2(net5595));
 sg13g2_nand2_1 _21805_ (.Y(_06445_),
    .A(net887),
    .B(net5591));
 sg13g2_o21ai_1 _21806_ (.B1(_06445_),
    .Y(_02197_),
    .A1(net4885),
    .A2(net5592));
 sg13g2_nand2_1 _21807_ (.Y(_06446_),
    .A(net1220),
    .B(net5595));
 sg13g2_o21ai_1 _21808_ (.B1(_06446_),
    .Y(_02198_),
    .A1(net4768),
    .A2(net5595));
 sg13g2_nand2_1 _21809_ (.Y(_06447_),
    .A(net1156),
    .B(net5597));
 sg13g2_o21ai_1 _21810_ (.B1(_06447_),
    .Y(_02199_),
    .A1(net4878),
    .A2(net5597));
 sg13g2_nand2_1 _21811_ (.Y(_06448_),
    .A(net914),
    .B(net5599));
 sg13g2_o21ai_1 _21812_ (.B1(_06448_),
    .Y(_02200_),
    .A1(net4872),
    .A2(net5599));
 sg13g2_nand2_1 _21813_ (.Y(_06449_),
    .A(net651),
    .B(net5600));
 sg13g2_o21ai_1 _21814_ (.B1(_06449_),
    .Y(_02201_),
    .A1(net4762),
    .A2(net5600));
 sg13g2_nand2_1 _21815_ (.Y(_06450_),
    .A(net871),
    .B(net5592));
 sg13g2_o21ai_1 _21816_ (.B1(_06450_),
    .Y(_02202_),
    .A1(net4870),
    .A2(net5592));
 sg13g2_nand2_1 _21817_ (.Y(_06451_),
    .A(net751),
    .B(net5598));
 sg13g2_o21ai_1 _21818_ (.B1(_06451_),
    .Y(_02203_),
    .A1(net4862),
    .A2(net5598));
 sg13g2_nand2_1 _21819_ (.Y(_06452_),
    .A(net492),
    .B(net5592));
 sg13g2_o21ai_1 _21820_ (.B1(_06452_),
    .Y(_02204_),
    .A1(net4859),
    .A2(net5592));
 sg13g2_nand2_1 _21821_ (.Y(_06453_),
    .A(net1108),
    .B(net5591));
 sg13g2_o21ai_1 _21822_ (.B1(_06453_),
    .Y(_02205_),
    .A1(net4856),
    .A2(net5591));
 sg13g2_nand2_1 _21823_ (.Y(_06454_),
    .A(net453),
    .B(net5595));
 sg13g2_o21ai_1 _21824_ (.B1(_06454_),
    .Y(_02206_),
    .A1(net4851),
    .A2(net5595));
 sg13g2_nand2_1 _21825_ (.Y(_06455_),
    .A(net1001),
    .B(net5591));
 sg13g2_o21ai_1 _21826_ (.B1(_06455_),
    .Y(_02207_),
    .A1(net4846),
    .A2(net5591));
 sg13g2_nand2_1 _21827_ (.Y(_06456_),
    .A(net1287),
    .B(net5597));
 sg13g2_o21ai_1 _21828_ (.B1(_06456_),
    .Y(_02208_),
    .A1(net4839),
    .A2(net5597));
 sg13g2_nand2_1 _21829_ (.Y(_06457_),
    .A(net720),
    .B(net5593));
 sg13g2_o21ai_1 _21830_ (.B1(_06457_),
    .Y(_02209_),
    .A1(net4832),
    .A2(net5593));
 sg13g2_nand2_1 _21831_ (.Y(_06458_),
    .A(net592),
    .B(net5599));
 sg13g2_o21ai_1 _21832_ (.B1(_06458_),
    .Y(_02210_),
    .A1(net4828),
    .A2(net5599));
 sg13g2_nand2_1 _21833_ (.Y(_06459_),
    .A(net508),
    .B(net5598));
 sg13g2_o21ai_1 _21834_ (.B1(_06459_),
    .Y(_02211_),
    .A1(net4823),
    .A2(net5598));
 sg13g2_and3_2 _21835_ (.X(_06460_),
    .A(_09507_),
    .B(_05728_),
    .C(net6070));
 sg13g2_nor2_1 _21836_ (.A(net1631),
    .B(net5383),
    .Y(_06461_));
 sg13g2_a21oi_1 _21837_ (.A1(net4994),
    .A2(net5383),
    .Y(_02212_),
    .B1(_06461_));
 sg13g2_nor2_1 _21838_ (.A(net1724),
    .B(net5383),
    .Y(_06462_));
 sg13g2_a21oi_1 _21839_ (.A1(net4990),
    .A2(net5383),
    .Y(_02213_),
    .B1(_06462_));
 sg13g2_nor2_1 _21840_ (.A(net1833),
    .B(net5383),
    .Y(_06463_));
 sg13g2_a21oi_1 _21841_ (.A1(net4984),
    .A2(net5383),
    .Y(_02214_),
    .B1(_06463_));
 sg13g2_nor2_1 _21842_ (.A(net1642),
    .B(net5382),
    .Y(_06464_));
 sg13g2_a21oi_1 _21843_ (.A1(net4981),
    .A2(net5382),
    .Y(_02215_),
    .B1(_06464_));
 sg13g2_nor2_1 _21844_ (.A(net2330),
    .B(net5389),
    .Y(_06465_));
 sg13g2_a21oi_1 _21845_ (.A1(net4976),
    .A2(net5389),
    .Y(_02216_),
    .B1(_06465_));
 sg13g2_nor2_1 _21846_ (.A(net1212),
    .B(net5389),
    .Y(_06466_));
 sg13g2_a21oi_1 _21847_ (.A1(net4970),
    .A2(net5389),
    .Y(_02217_),
    .B1(_06466_));
 sg13g2_nor2_1 _21848_ (.A(net1791),
    .B(net5383),
    .Y(_06467_));
 sg13g2_a21oi_1 _21849_ (.A1(net4965),
    .A2(net5383),
    .Y(_02218_),
    .B1(_06467_));
 sg13g2_nor2_1 _21850_ (.A(net1810),
    .B(net5386),
    .Y(_06468_));
 sg13g2_a21oi_1 _21851_ (.A1(net4917),
    .A2(net5386),
    .Y(_02219_),
    .B1(_06468_));
 sg13g2_nor2_1 _21852_ (.A(net1464),
    .B(net5384),
    .Y(_06469_));
 sg13g2_a21oi_1 _21853_ (.A1(net4779),
    .A2(net5384),
    .Y(_02220_),
    .B1(_06469_));
 sg13g2_nor2_1 _21854_ (.A(net1324),
    .B(net5390),
    .Y(_06470_));
 sg13g2_a21oi_1 _21855_ (.A1(net4912),
    .A2(net5390),
    .Y(_02221_),
    .B1(_06470_));
 sg13g2_nor2_1 _21856_ (.A(net1683),
    .B(net5388),
    .Y(_06471_));
 sg13g2_a21oi_1 _21857_ (.A1(net4908),
    .A2(net5388),
    .Y(_02222_),
    .B1(_06471_));
 sg13g2_nor2_1 _21858_ (.A(net1581),
    .B(net5384),
    .Y(_06472_));
 sg13g2_a21oi_1 _21859_ (.A1(net4777),
    .A2(net5384),
    .Y(_02223_),
    .B1(_06472_));
 sg13g2_nor2_1 _21860_ (.A(net2070),
    .B(net5387),
    .Y(_06473_));
 sg13g2_a21oi_1 _21861_ (.A1(net4899),
    .A2(net5387),
    .Y(_02224_),
    .B1(_06473_));
 sg13g2_nor2_1 _21862_ (.A(net1914),
    .B(net5387),
    .Y(_06474_));
 sg13g2_a21oi_1 _21863_ (.A1(net4963),
    .A2(net5387),
    .Y(_02225_),
    .B1(_06474_));
 sg13g2_nor2_1 _21864_ (.A(net1741),
    .B(net5381),
    .Y(_06475_));
 sg13g2_a21oi_1 _21865_ (.A1(net4956),
    .A2(net5381),
    .Y(_02226_),
    .B1(_06475_));
 sg13g2_nor2_1 _21866_ (.A(net1692),
    .B(net5387),
    .Y(_06476_));
 sg13g2_a21oi_1 _21867_ (.A1(net4896),
    .A2(net5387),
    .Y(_02227_),
    .B1(_06476_));
 sg13g2_nor2_1 _21868_ (.A(net1449),
    .B(net5386),
    .Y(_06477_));
 sg13g2_a21oi_1 _21869_ (.A1(net4889),
    .A2(net5386),
    .Y(_02228_),
    .B1(_06477_));
 sg13g2_nor2_1 _21870_ (.A(net1895),
    .B(net5382),
    .Y(_06478_));
 sg13g2_a21oi_1 _21871_ (.A1(net4886),
    .A2(net5382),
    .Y(_02229_),
    .B1(_06478_));
 sg13g2_nor2_1 _21872_ (.A(net1879),
    .B(net5387),
    .Y(_06479_));
 sg13g2_a21oi_1 _21873_ (.A1(net4770),
    .A2(net5387),
    .Y(_02230_),
    .B1(_06479_));
 sg13g2_nor2_1 _21874_ (.A(net2214),
    .B(net5386),
    .Y(_06480_));
 sg13g2_a21oi_1 _21875_ (.A1(net4880),
    .A2(net5386),
    .Y(_02231_),
    .B1(_06480_));
 sg13g2_nor2_1 _21876_ (.A(net2081),
    .B(net5388),
    .Y(_06481_));
 sg13g2_a21oi_1 _21877_ (.A1(net4876),
    .A2(net5388),
    .Y(_02232_),
    .B1(_06481_));
 sg13g2_nor2_1 _21878_ (.A(net1459),
    .B(net5389),
    .Y(_06482_));
 sg13g2_a21oi_1 _21879_ (.A1(net4763),
    .A2(net5389),
    .Y(_02233_),
    .B1(_06482_));
 sg13g2_nor2_1 _21880_ (.A(net2242),
    .B(net5381),
    .Y(_06483_));
 sg13g2_a21oi_1 _21881_ (.A1(net4867),
    .A2(net5381),
    .Y(_02234_),
    .B1(_06483_));
 sg13g2_nor2_1 _21882_ (.A(net1295),
    .B(net5388),
    .Y(_06484_));
 sg13g2_a21oi_1 _21883_ (.A1(net4862),
    .A2(net5388),
    .Y(_02235_),
    .B1(_06484_));
 sg13g2_nor2_1 _21884_ (.A(net1571),
    .B(net5382),
    .Y(_06485_));
 sg13g2_a21oi_1 _21885_ (.A1(net4860),
    .A2(net5382),
    .Y(_02236_),
    .B1(_06485_));
 sg13g2_nor2_1 _21886_ (.A(net1421),
    .B(net5381),
    .Y(_06486_));
 sg13g2_a21oi_1 _21887_ (.A1(net4852),
    .A2(net5381),
    .Y(_02237_),
    .B1(_06486_));
 sg13g2_nor2_1 _21888_ (.A(net1236),
    .B(net5386),
    .Y(_06487_));
 sg13g2_a21oi_1 _21889_ (.A1(net4849),
    .A2(net5386),
    .Y(_02238_),
    .B1(_06487_));
 sg13g2_nor2_1 _21890_ (.A(net1918),
    .B(net5381),
    .Y(_06488_));
 sg13g2_a21oi_1 _21891_ (.A1(net4842),
    .A2(net5381),
    .Y(_02239_),
    .B1(_06488_));
 sg13g2_nor2_1 _21892_ (.A(net2152),
    .B(net5382),
    .Y(_06489_));
 sg13g2_a21oi_1 _21893_ (.A1(net4838),
    .A2(net5382),
    .Y(_02240_),
    .B1(_06489_));
 sg13g2_nor2_1 _21894_ (.A(net1597),
    .B(net5384),
    .Y(_06490_));
 sg13g2_a21oi_1 _21895_ (.A1(net4832),
    .A2(net5384),
    .Y(_02241_),
    .B1(_06490_));
 sg13g2_nor2_1 _21896_ (.A(net1667),
    .B(net5388),
    .Y(_06491_));
 sg13g2_a21oi_1 _21897_ (.A1(net4827),
    .A2(net5388),
    .Y(_02242_),
    .B1(_06491_));
 sg13g2_nor2_1 _21898_ (.A(net1657),
    .B(net5389),
    .Y(_06492_));
 sg13g2_a21oi_1 _21899_ (.A1(net4826),
    .A2(net5389),
    .Y(_02243_),
    .B1(_06492_));
 sg13g2_nor2_2 _21900_ (.A(_09505_),
    .B(_06195_),
    .Y(_06493_));
 sg13g2_nor2_1 _21901_ (.A(net1717),
    .B(net5373),
    .Y(_06494_));
 sg13g2_a21oi_1 _21902_ (.A1(net4995),
    .A2(net5373),
    .Y(_02244_),
    .B1(_06494_));
 sg13g2_nor2_1 _21903_ (.A(net2217),
    .B(net5373),
    .Y(_06495_));
 sg13g2_a21oi_1 _21904_ (.A1(net4991),
    .A2(net5373),
    .Y(_02245_),
    .B1(_06495_));
 sg13g2_nor2_1 _21905_ (.A(net2305),
    .B(net5373),
    .Y(_06496_));
 sg13g2_a21oi_1 _21906_ (.A1(net4984),
    .A2(net5373),
    .Y(_02246_),
    .B1(_06496_));
 sg13g2_nor2_1 _21907_ (.A(net2069),
    .B(net5371),
    .Y(_06497_));
 sg13g2_a21oi_1 _21908_ (.A1(net4980),
    .A2(net5371),
    .Y(_02247_),
    .B1(_06497_));
 sg13g2_nor2_1 _21909_ (.A(net1873),
    .B(net5372),
    .Y(_06498_));
 sg13g2_a21oi_1 _21910_ (.A1(net4978),
    .A2(net5372),
    .Y(_02248_),
    .B1(_06498_));
 sg13g2_nor2_1 _21911_ (.A(net2127),
    .B(net5379),
    .Y(_06499_));
 sg13g2_a21oi_1 _21912_ (.A1(net4972),
    .A2(net5379),
    .Y(_02249_),
    .B1(_06499_));
 sg13g2_nor2_1 _21913_ (.A(net1537),
    .B(net5373),
    .Y(_06500_));
 sg13g2_a21oi_1 _21914_ (.A1(net4966),
    .A2(net5374),
    .Y(_02250_),
    .B1(_06500_));
 sg13g2_nor2_1 _21915_ (.A(net1322),
    .B(net5376),
    .Y(_06501_));
 sg13g2_a21oi_1 _21916_ (.A1(net4919),
    .A2(net5376),
    .Y(_02251_),
    .B1(_06501_));
 sg13g2_nor2_1 _21917_ (.A(net1821),
    .B(net5373),
    .Y(_06502_));
 sg13g2_a21oi_1 _21918_ (.A1(net4781),
    .A2(net5374),
    .Y(_02252_),
    .B1(_06502_));
 sg13g2_nor2_1 _21919_ (.A(net1932),
    .B(net5379),
    .Y(_06503_));
 sg13g2_a21oi_1 _21920_ (.A1(net4914),
    .A2(net5379),
    .Y(_02253_),
    .B1(_06503_));
 sg13g2_nor2_1 _21921_ (.A(net2139),
    .B(net5378),
    .Y(_06504_));
 sg13g2_a21oi_1 _21922_ (.A1(net4906),
    .A2(net5378),
    .Y(_02254_),
    .B1(_06504_));
 sg13g2_nor2_1 _21923_ (.A(net2614),
    .B(net5374),
    .Y(_06505_));
 sg13g2_a21oi_1 _21924_ (.A1(net4775),
    .A2(net5374),
    .Y(_02255_),
    .B1(_06505_));
 sg13g2_nor2_1 _21925_ (.A(net1674),
    .B(net5376),
    .Y(_06506_));
 sg13g2_a21oi_1 _21926_ (.A1(net4899),
    .A2(net5376),
    .Y(_02256_),
    .B1(_06506_));
 sg13g2_nor2_1 _21927_ (.A(net1543),
    .B(net5376),
    .Y(_06507_));
 sg13g2_a21oi_1 _21928_ (.A1(net4959),
    .A2(net5376),
    .Y(_02257_),
    .B1(_06507_));
 sg13g2_nor2_1 _21929_ (.A(net1900),
    .B(net5371),
    .Y(_06508_));
 sg13g2_a21oi_1 _21930_ (.A1(net4958),
    .A2(net5371),
    .Y(_02258_),
    .B1(_06508_));
 sg13g2_nor2_1 _21931_ (.A(net2164),
    .B(net5380),
    .Y(_06509_));
 sg13g2_a21oi_1 _21932_ (.A1(net4894),
    .A2(net5377),
    .Y(_02259_),
    .B1(_06509_));
 sg13g2_nor2_1 _21933_ (.A(net1896),
    .B(net5377),
    .Y(_06510_));
 sg13g2_a21oi_1 _21934_ (.A1(net4890),
    .A2(net5377),
    .Y(_02260_),
    .B1(_06510_));
 sg13g2_nor2_1 _21935_ (.A(net2270),
    .B(net5372),
    .Y(_06511_));
 sg13g2_a21oi_1 _21936_ (.A1(net4887),
    .A2(net5372),
    .Y(_02261_),
    .B1(_06511_));
 sg13g2_nor2_1 _21937_ (.A(net1908),
    .B(net5376),
    .Y(_06512_));
 sg13g2_a21oi_1 _21938_ (.A1(net4772),
    .A2(net5376),
    .Y(_02262_),
    .B1(_06512_));
 sg13g2_nor2_1 _21939_ (.A(net1725),
    .B(net5377),
    .Y(_06513_));
 sg13g2_a21oi_1 _21940_ (.A1(net4882),
    .A2(net5377),
    .Y(_02263_),
    .B1(_06513_));
 sg13g2_nor2_1 _21941_ (.A(net1284),
    .B(net5378),
    .Y(_06514_));
 sg13g2_a21oi_1 _21942_ (.A1(net4872),
    .A2(net5378),
    .Y(_02264_),
    .B1(_06514_));
 sg13g2_nor2_1 _21943_ (.A(net2294),
    .B(net5379),
    .Y(_06515_));
 sg13g2_a21oi_1 _21944_ (.A1(net4764),
    .A2(net5379),
    .Y(_02265_),
    .B1(_06515_));
 sg13g2_nor2_1 _21945_ (.A(net2421),
    .B(net5371),
    .Y(_06516_));
 sg13g2_a21oi_1 _21946_ (.A1(net4869),
    .A2(net5371),
    .Y(_02266_),
    .B1(_06516_));
 sg13g2_nor2_1 _21947_ (.A(net2032),
    .B(net5378),
    .Y(_06517_));
 sg13g2_a21oi_1 _21948_ (.A1(net4865),
    .A2(net5378),
    .Y(_02267_),
    .B1(_06517_));
 sg13g2_nor2_1 _21949_ (.A(net1315),
    .B(net5372),
    .Y(_06518_));
 sg13g2_a21oi_1 _21950_ (.A1(net4859),
    .A2(net5375),
    .Y(_02268_),
    .B1(_06518_));
 sg13g2_nor2_1 _21951_ (.A(net1941),
    .B(net5371),
    .Y(_06519_));
 sg13g2_a21oi_1 _21952_ (.A1(net4854),
    .A2(net5371),
    .Y(_02269_),
    .B1(_06519_));
 sg13g2_nor2_1 _21953_ (.A(net1510),
    .B(net5377),
    .Y(_06520_));
 sg13g2_a21oi_1 _21954_ (.A1(net4847),
    .A2(net5377),
    .Y(_02270_),
    .B1(_06520_));
 sg13g2_nor2_1 _21955_ (.A(net1511),
    .B(net5372),
    .Y(_06521_));
 sg13g2_a21oi_1 _21956_ (.A1(net4843),
    .A2(net5372),
    .Y(_02271_),
    .B1(_06521_));
 sg13g2_nor2_1 _21957_ (.A(net2007),
    .B(net5375),
    .Y(_06522_));
 sg13g2_a21oi_1 _21958_ (.A1(net4838),
    .A2(net5375),
    .Y(_02272_),
    .B1(_06522_));
 sg13g2_nor2_1 _21959_ (.A(net1817),
    .B(net5374),
    .Y(_06523_));
 sg13g2_a21oi_1 _21960_ (.A1(net4834),
    .A2(net5374),
    .Y(_02273_),
    .B1(_06523_));
 sg13g2_nor2_1 _21961_ (.A(net1834),
    .B(net5379),
    .Y(_06524_));
 sg13g2_a21oi_1 _21962_ (.A1(net4830),
    .A2(net5380),
    .Y(_02274_),
    .B1(_06524_));
 sg13g2_nor2_1 _21963_ (.A(net2321),
    .B(net5378),
    .Y(_06525_));
 sg13g2_a21oi_1 _21964_ (.A1(net4824),
    .A2(net5378),
    .Y(_02275_),
    .B1(_06525_));
 sg13g2_nand3_1 _21965_ (.B(_05728_),
    .C(net6071),
    .A(_05590_),
    .Y(_06526_));
 sg13g2_nand2_1 _21966_ (.Y(_06527_),
    .A(net744),
    .B(net5583));
 sg13g2_o21ai_1 _21967_ (.B1(_06527_),
    .Y(_02276_),
    .A1(net4995),
    .A2(net5583));
 sg13g2_nand2_1 _21968_ (.Y(_06528_),
    .A(net679),
    .B(net5583));
 sg13g2_o21ai_1 _21969_ (.B1(_06528_),
    .Y(_02277_),
    .A1(net4992),
    .A2(net5583));
 sg13g2_nand2_1 _21970_ (.Y(_06529_),
    .A(net966),
    .B(net5582));
 sg13g2_o21ai_1 _21971_ (.B1(_06529_),
    .Y(_02278_),
    .A1(net4987),
    .A2(net5582));
 sg13g2_nand2_1 _21972_ (.Y(_06530_),
    .A(net452),
    .B(net5580));
 sg13g2_o21ai_1 _21973_ (.B1(_06530_),
    .Y(_02279_),
    .A1(net4980),
    .A2(net5580));
 sg13g2_nand2_1 _21974_ (.Y(_06531_),
    .A(net731),
    .B(net5584));
 sg13g2_o21ai_1 _21975_ (.B1(_06531_),
    .Y(_02280_),
    .A1(net4974),
    .A2(net5584));
 sg13g2_nand2_1 _21976_ (.Y(_06532_),
    .A(net1253),
    .B(net5589));
 sg13g2_o21ai_1 _21977_ (.B1(_06532_),
    .Y(_02281_),
    .A1(net4969),
    .A2(net5589));
 sg13g2_nand2_1 _21978_ (.Y(_06533_),
    .A(net692),
    .B(net5582));
 sg13g2_o21ai_1 _21979_ (.B1(_06533_),
    .Y(_02282_),
    .A1(net4964),
    .A2(net5582));
 sg13g2_nand2_1 _21980_ (.Y(_06534_),
    .A(net461),
    .B(net5584));
 sg13g2_o21ai_1 _21981_ (.B1(_06534_),
    .Y(_02283_),
    .A1(net4918),
    .A2(net5584));
 sg13g2_nand2_1 _21982_ (.Y(_06535_),
    .A(net454),
    .B(net5582));
 sg13g2_o21ai_1 _21983_ (.B1(_06535_),
    .Y(_02284_),
    .A1(net4781),
    .A2(net5582));
 sg13g2_nand2_1 _21984_ (.Y(_06536_),
    .A(net622),
    .B(net5587));
 sg13g2_o21ai_1 _21985_ (.B1(_06536_),
    .Y(_02285_),
    .A1(net4913),
    .A2(net5587));
 sg13g2_nand2_1 _21986_ (.Y(_06537_),
    .A(net527),
    .B(net5587));
 sg13g2_o21ai_1 _21987_ (.B1(_06537_),
    .Y(_02286_),
    .A1(net4909),
    .A2(net5587));
 sg13g2_nand2_1 _21988_ (.Y(_06538_),
    .A(net781),
    .B(net5583));
 sg13g2_o21ai_1 _21989_ (.B1(_06538_),
    .Y(_02287_),
    .A1(net4777),
    .A2(net5583));
 sg13g2_nand2_1 _21990_ (.Y(_06539_),
    .A(net393),
    .B(net5585));
 sg13g2_o21ai_1 _21991_ (.B1(_06539_),
    .Y(_02288_),
    .A1(net4904),
    .A2(net5585));
 sg13g2_nand2_1 _21992_ (.Y(_06540_),
    .A(net790),
    .B(net5585));
 sg13g2_o21ai_1 _21993_ (.B1(_06540_),
    .Y(_02289_),
    .A1(net4959),
    .A2(net5585));
 sg13g2_nand2_1 _21994_ (.Y(_06541_),
    .A(net930),
    .B(net5580));
 sg13g2_o21ai_1 _21995_ (.B1(_06541_),
    .Y(_02290_),
    .A1(net4957),
    .A2(net5580));
 sg13g2_nand2_1 _21996_ (.Y(_06542_),
    .A(net560),
    .B(net5586));
 sg13g2_o21ai_1 _21997_ (.B1(_06542_),
    .Y(_02291_),
    .A1(net4894),
    .A2(net5586));
 sg13g2_nand2_1 _21998_ (.Y(_06543_),
    .A(net951),
    .B(net5585));
 sg13g2_o21ai_1 _21999_ (.B1(_06543_),
    .Y(_02292_),
    .A1(net4891),
    .A2(net5585));
 sg13g2_nand2_1 _22000_ (.Y(_06544_),
    .A(net1131),
    .B(net5581));
 sg13g2_o21ai_1 _22001_ (.B1(_06544_),
    .Y(_02293_),
    .A1(net4884),
    .A2(net5581));
 sg13g2_nand2_1 _22002_ (.Y(_06545_),
    .A(net758),
    .B(net5585));
 sg13g2_o21ai_1 _22003_ (.B1(_06545_),
    .Y(_02294_),
    .A1(net4768),
    .A2(net5585));
 sg13g2_nand2_1 _22004_ (.Y(_06546_),
    .A(net849),
    .B(net5584));
 sg13g2_o21ai_1 _22005_ (.B1(_06546_),
    .Y(_02295_),
    .A1(net4879),
    .A2(net5584));
 sg13g2_nand2_1 _22006_ (.Y(_06547_),
    .A(net618),
    .B(net5587));
 sg13g2_o21ai_1 _22007_ (.B1(_06547_),
    .Y(_02296_),
    .A1(net4876),
    .A2(net5587));
 sg13g2_nand2_1 _22008_ (.Y(_06548_),
    .A(net895),
    .B(net5589));
 sg13g2_o21ai_1 _22009_ (.B1(_06548_),
    .Y(_02297_),
    .A1(net4763),
    .A2(net5589));
 sg13g2_nand2_1 _22010_ (.Y(_06549_),
    .A(net433),
    .B(net5581));
 sg13g2_o21ai_1 _22011_ (.B1(_06549_),
    .Y(_02298_),
    .A1(net4870),
    .A2(net5581));
 sg13g2_nand2_1 _22012_ (.Y(_06550_),
    .A(net834),
    .B(net5588));
 sg13g2_o21ai_1 _22013_ (.B1(_06550_),
    .Y(_02299_),
    .A1(net4862),
    .A2(net5588));
 sg13g2_nand2_1 _22014_ (.Y(_06551_),
    .A(net531),
    .B(net5581));
 sg13g2_o21ai_1 _22015_ (.B1(_06551_),
    .Y(_02300_),
    .A1(net4859),
    .A2(net5581));
 sg13g2_nand2_1 _22016_ (.Y(_06552_),
    .A(net1037),
    .B(net5580));
 sg13g2_o21ai_1 _22017_ (.B1(_06552_),
    .Y(_02301_),
    .A1(net4855),
    .A2(net5580));
 sg13g2_nand2_1 _22018_ (.Y(_06553_),
    .A(net647),
    .B(net5584));
 sg13g2_o21ai_1 _22019_ (.B1(_06553_),
    .Y(_02302_),
    .A1(net4849),
    .A2(net5584));
 sg13g2_nand2_1 _22020_ (.Y(_06554_),
    .A(net435),
    .B(net5580));
 sg13g2_o21ai_1 _22021_ (.B1(_06554_),
    .Y(_02303_),
    .A1(net4845),
    .A2(net5580));
 sg13g2_nand2_1 _22022_ (.Y(_06555_),
    .A(net1002),
    .B(net5586));
 sg13g2_o21ai_1 _22023_ (.B1(_06555_),
    .Y(_02304_),
    .A1(net4840),
    .A2(net5586));
 sg13g2_nand2_1 _22024_ (.Y(_06556_),
    .A(net1285),
    .B(net5582));
 sg13g2_o21ai_1 _22025_ (.B1(_06556_),
    .Y(_02305_),
    .A1(net4835),
    .A2(net5582));
 sg13g2_nand2_1 _22026_ (.Y(_06557_),
    .A(net658),
    .B(net5588));
 sg13g2_o21ai_1 _22027_ (.B1(_06557_),
    .Y(_02306_),
    .A1(net4827),
    .A2(net5588));
 sg13g2_nand2_1 _22028_ (.Y(_06558_),
    .A(net1242),
    .B(net5587));
 sg13g2_o21ai_1 _22029_ (.B1(_06558_),
    .Y(_02307_),
    .A1(net4823),
    .A2(net5587));
 sg13g2_nand3_1 _22030_ (.B(_05728_),
    .C(net6070),
    .A(_05625_),
    .Y(_06559_));
 sg13g2_nand2_1 _22031_ (.Y(_06560_),
    .A(net1209),
    .B(net5576));
 sg13g2_o21ai_1 _22032_ (.B1(_06560_),
    .Y(_02308_),
    .A1(net4998),
    .A2(net5576));
 sg13g2_nand2_1 _22033_ (.Y(_06561_),
    .A(net1139),
    .B(net5576));
 sg13g2_o21ai_1 _22034_ (.B1(_06561_),
    .Y(_02309_),
    .A1(_09533_),
    .A2(net5576));
 sg13g2_nand2_1 _22035_ (.Y(_06562_),
    .A(net507),
    .B(net5573));
 sg13g2_o21ai_1 _22036_ (.B1(_06562_),
    .Y(_02310_),
    .A1(net4985),
    .A2(net5573));
 sg13g2_nand2_1 _22037_ (.Y(_06563_),
    .A(net1142),
    .B(net5577));
 sg13g2_o21ai_1 _22038_ (.B1(_06563_),
    .Y(_02311_),
    .A1(_09551_),
    .A2(net5577));
 sg13g2_nand2_1 _22039_ (.Y(_06564_),
    .A(net444),
    .B(net5577));
 sg13g2_o21ai_1 _22040_ (.B1(_06564_),
    .Y(_02312_),
    .A1(_09560_),
    .A2(net5577));
 sg13g2_nand2_1 _22041_ (.Y(_06565_),
    .A(net1044),
    .B(net5574));
 sg13g2_o21ai_1 _22042_ (.B1(_06565_),
    .Y(_02313_),
    .A1(_09569_),
    .A2(net5574));
 sg13g2_nand2_1 _22043_ (.Y(_06566_),
    .A(net1094),
    .B(net5576));
 sg13g2_o21ai_1 _22044_ (.B1(_06566_),
    .Y(_02314_),
    .A1(_09578_),
    .A2(net5576));
 sg13g2_nand2_1 _22045_ (.Y(_06567_),
    .A(net798),
    .B(net5571));
 sg13g2_o21ai_1 _22046_ (.B1(_06567_),
    .Y(_02315_),
    .A1(_09589_),
    .A2(net5571));
 sg13g2_nand2_1 _22047_ (.Y(_06568_),
    .A(net488),
    .B(net5574));
 sg13g2_o21ai_1 _22048_ (.B1(_06568_),
    .Y(_02316_),
    .A1(_09603_),
    .A2(net5574));
 sg13g2_nand2_1 _22049_ (.Y(_06569_),
    .A(net673),
    .B(net5574));
 sg13g2_o21ai_1 _22050_ (.B1(_06569_),
    .Y(_02317_),
    .A1(_09612_),
    .A2(net5573));
 sg13g2_nand2_1 _22051_ (.Y(_06570_),
    .A(net684),
    .B(net5573));
 sg13g2_o21ai_1 _22052_ (.B1(_06570_),
    .Y(_02318_),
    .A1(net4910),
    .A2(net5573));
 sg13g2_nand2_1 _22053_ (.Y(_06571_),
    .A(net991),
    .B(net5575));
 sg13g2_o21ai_1 _22054_ (.B1(_06571_),
    .Y(_02319_),
    .A1(net4778),
    .A2(net5575));
 sg13g2_nand2_1 _22055_ (.Y(_06572_),
    .A(net479),
    .B(net5571));
 sg13g2_o21ai_1 _22056_ (.B1(_06572_),
    .Y(_02320_),
    .A1(_09641_),
    .A2(net5572));
 sg13g2_nand2_1 _22057_ (.Y(_06573_),
    .A(net808),
    .B(net5569));
 sg13g2_o21ai_1 _22058_ (.B1(_06573_),
    .Y(_02321_),
    .A1(_09650_),
    .A2(net5569));
 sg13g2_nand2_1 _22059_ (.Y(_06574_),
    .A(net839),
    .B(net5569));
 sg13g2_o21ai_1 _22060_ (.B1(_06574_),
    .Y(_02322_),
    .A1(_09659_),
    .A2(net5569));
 sg13g2_nand2_1 _22061_ (.Y(_06575_),
    .A(net641),
    .B(net5570));
 sg13g2_o21ai_1 _22062_ (.B1(_06575_),
    .Y(_02323_),
    .A1(_09669_),
    .A2(net5570));
 sg13g2_nand2_1 _22063_ (.Y(_06576_),
    .A(net1734),
    .B(net5569));
 sg13g2_o21ai_1 _22064_ (.B1(_06576_),
    .Y(_02324_),
    .A1(_09680_),
    .A2(net5569));
 sg13g2_nand2_1 _22065_ (.Y(_06577_),
    .A(net1196),
    .B(net5571));
 sg13g2_o21ai_1 _22066_ (.B1(_06577_),
    .Y(_02325_),
    .A1(_09689_),
    .A2(net5571));
 sg13g2_nand2_1 _22067_ (.Y(_06578_),
    .A(net1036),
    .B(net5569));
 sg13g2_o21ai_1 _22068_ (.B1(_06578_),
    .Y(_02326_),
    .A1(_09698_),
    .A2(net5569));
 sg13g2_nand2_1 _22069_ (.Y(_06579_),
    .A(net392),
    .B(net5577));
 sg13g2_o21ai_1 _22070_ (.B1(_06579_),
    .Y(_02327_),
    .A1(net4881),
    .A2(net5578));
 sg13g2_nand2_1 _22071_ (.Y(_06580_),
    .A(net2735),
    .B(net5578));
 sg13g2_o21ai_1 _22072_ (.B1(_06580_),
    .Y(_02328_),
    .A1(net4877),
    .A2(net5578));
 sg13g2_nand2_1 _22073_ (.Y(_06581_),
    .A(net878),
    .B(net5578));
 sg13g2_o21ai_1 _22074_ (.B1(_06581_),
    .Y(_02329_),
    .A1(net4762),
    .A2(net5578));
 sg13g2_nand2_1 _22075_ (.Y(_06582_),
    .A(net635),
    .B(net5572));
 sg13g2_o21ai_1 _22076_ (.B1(_06582_),
    .Y(_02330_),
    .A1(net4867),
    .A2(net5572));
 sg13g2_nand2_1 _22077_ (.Y(_06583_),
    .A(net390),
    .B(net5578));
 sg13g2_o21ai_1 _22078_ (.B1(_06583_),
    .Y(_02331_),
    .A1(_09743_),
    .A2(net5579));
 sg13g2_nand2_1 _22079_ (.Y(_06584_),
    .A(net1304),
    .B(net5571));
 sg13g2_o21ai_1 _22080_ (.B1(_06584_),
    .Y(_02332_),
    .A1(net4861),
    .A2(net5571));
 sg13g2_nand2_1 _22081_ (.Y(_06585_),
    .A(net1097),
    .B(net5570));
 sg13g2_o21ai_1 _22082_ (.B1(_06585_),
    .Y(_02333_),
    .A1(net4856),
    .A2(net5570));
 sg13g2_nand2_1 _22083_ (.Y(_06586_),
    .A(net912),
    .B(net5577));
 sg13g2_o21ai_1 _22084_ (.B1(_06586_),
    .Y(_02334_),
    .A1(net4849),
    .A2(net5578));
 sg13g2_nand2_1 _22085_ (.Y(_06587_),
    .A(net829),
    .B(net5571));
 sg13g2_o21ai_1 _22086_ (.B1(_06587_),
    .Y(_02335_),
    .A1(net4846),
    .A2(net5572));
 sg13g2_nand2_1 _22087_ (.Y(_06588_),
    .A(net484),
    .B(net5577));
 sg13g2_o21ai_1 _22088_ (.B1(_06588_),
    .Y(_02336_),
    .A1(net4841),
    .A2(net5577));
 sg13g2_nand2_1 _22089_ (.Y(_06589_),
    .A(net741),
    .B(net5573));
 sg13g2_o21ai_1 _22090_ (.B1(_06589_),
    .Y(_02337_),
    .A1(net4836),
    .A2(net5574));
 sg13g2_nand2_1 _22091_ (.Y(_06590_),
    .A(net816),
    .B(net5579));
 sg13g2_o21ai_1 _22092_ (.B1(_06590_),
    .Y(_02338_),
    .A1(_09799_),
    .A2(net5579));
 sg13g2_nand2_1 _22093_ (.Y(_06591_),
    .A(net555),
    .B(net5573));
 sg13g2_o21ai_1 _22094_ (.B1(_06591_),
    .Y(_02339_),
    .A1(_09807_),
    .A2(net5573));
 sg13g2_nand3_1 _22095_ (.B(_09043_),
    .C(_09514_),
    .A(_09024_),
    .Y(_06592_));
 sg13g2_nand2_2 _22096_ (.Y(_06593_),
    .A(_09893_),
    .B(_10267_));
 sg13g2_a21oi_1 _22097_ (.A1(net2827),
    .A2(_06593_),
    .Y(_06594_),
    .B1(_11137_));
 sg13g2_nor2b_1 _22098_ (.A(_11139_),
    .B_N(_06593_),
    .Y(_06595_));
 sg13g2_nor3_1 _22099_ (.A(_06592_),
    .B(_06594_),
    .C(_06595_),
    .Y(_06596_));
 sg13g2_a21o_1 _22100_ (.A2(_06592_),
    .A1(net2827),
    .B1(_06596_),
    .X(_02340_));
 sg13g2_a21oi_1 _22101_ (.A1(net2502),
    .A2(_06593_),
    .Y(_06597_),
    .B1(_11147_));
 sg13g2_nor2b_1 _22102_ (.A(_11149_),
    .B_N(_06593_),
    .Y(_06598_));
 sg13g2_nor3_1 _22103_ (.A(_06592_),
    .B(_06597_),
    .C(_06598_),
    .Y(_06599_));
 sg13g2_a21o_1 _22104_ (.A2(_06592_),
    .A1(net2502),
    .B1(_06599_),
    .X(_02341_));
 sg13g2_nand2_1 _22105_ (.Y(_06600_),
    .A(\soc_inst.cpu_core.id_imm[0] ),
    .B(\soc_inst.cpu_core.id_pc[0] ));
 sg13g2_xor2_1 _22106_ (.B(\soc_inst.cpu_core.id_pc[0] ),
    .A(\soc_inst.cpu_core.id_imm[0] ),
    .X(_06601_));
 sg13g2_nand2_2 _22107_ (.Y(_06602_),
    .A(_08056_),
    .B(\soc_inst.cpu_core.id_rs1_data[31] ));
 sg13g2_nor2_1 _22108_ (.A(_08056_),
    .B(\soc_inst.cpu_core.id_rs1_data[31] ),
    .Y(_06603_));
 sg13g2_o21ai_1 _22109_ (.B1(_06602_),
    .Y(_06604_),
    .A1(\soc_inst.cpu_core.id_rs1_data[24] ),
    .A2(_08067_));
 sg13g2_nand2b_1 _22110_ (.Y(_06605_),
    .B(\soc_inst.cpu_core.id_rs1_data[28] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[28] ));
 sg13g2_o21ai_1 _22111_ (.B1(_06605_),
    .Y(_06606_),
    .A1(_08059_),
    .A2(\soc_inst.cpu_core.id_rs2_data[29] ));
 sg13g2_nand2_1 _22112_ (.Y(_06607_),
    .A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .B(_08067_));
 sg13g2_o21ai_1 _22113_ (.B1(_06607_),
    .Y(_06608_),
    .A1(_08065_),
    .A2(\soc_inst.cpu_core.id_rs2_data[25] ));
 sg13g2_a22oi_1 _22114_ (.Y(_06609_),
    .B1(\soc_inst.cpu_core.id_rs1_data[26] ),
    .B2(_08064_),
    .A2(_08062_),
    .A1(\soc_inst.cpu_core.id_rs1_data[27] ));
 sg13g2_nand2b_1 _22115_ (.Y(_06610_),
    .B(\soc_inst.cpu_core.id_rs1_data[30] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[30] ));
 sg13g2_nand2b_1 _22116_ (.Y(_06611_),
    .B(_06610_),
    .A_N(_06603_));
 sg13g2_a221oi_1 _22117_ (.B2(\soc_inst.cpu_core.id_rs2_data[29] ),
    .C1(_06611_),
    .B1(_08059_),
    .A1(_08058_),
    .Y(_06612_),
    .A2(\soc_inst.cpu_core.id_rs2_data[30] ));
 sg13g2_nand2_1 _22118_ (.Y(_06613_),
    .A(_08065_),
    .B(\soc_inst.cpu_core.id_rs2_data[25] ));
 sg13g2_o21ai_1 _22119_ (.B1(_06613_),
    .Y(_06614_),
    .A1(\soc_inst.cpu_core.id_rs1_data[26] ),
    .A2(_08064_));
 sg13g2_a22oi_1 _22120_ (.Y(_06615_),
    .B1(_08061_),
    .B2(\soc_inst.cpu_core.id_rs2_data[27] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[28] ),
    .A1(_08060_));
 sg13g2_nor4_1 _22121_ (.A(_06604_),
    .B(_06606_),
    .C(_06608_),
    .D(_06614_),
    .Y(_06616_));
 sg13g2_nand4_1 _22122_ (.B(_06612_),
    .C(_06615_),
    .A(_06609_),
    .Y(_06617_),
    .D(_06616_));
 sg13g2_a22oi_1 _22123_ (.Y(_06618_),
    .B1(\soc_inst.cpu_core.id_rs1_data[22] ),
    .B2(_08071_),
    .A2(_08069_),
    .A1(\soc_inst.cpu_core.id_rs1_data[23] ));
 sg13g2_o21ai_1 _22124_ (.B1(_06618_),
    .Y(_06619_),
    .A1(\soc_inst.cpu_core.id_rs1_data[21] ),
    .A2(_08072_));
 sg13g2_a221oi_1 _22125_ (.B2(\soc_inst.cpu_core.id_rs2_data[22] ),
    .C1(_06619_),
    .B1(_08070_),
    .A1(_08068_),
    .Y(_06620_),
    .A2(\soc_inst.cpu_core.id_rs2_data[23] ));
 sg13g2_nand2_1 _22126_ (.Y(_06621_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(_08072_));
 sg13g2_o21ai_1 _22127_ (.B1(_06621_),
    .Y(_06622_),
    .A1(_08073_),
    .A2(\soc_inst.cpu_core.id_rs2_data[20] ));
 sg13g2_a221oi_1 _22128_ (.B2(\soc_inst.cpu_core.id_rs2_data[17] ),
    .C1(_06622_),
    .B1(_08078_),
    .A1(_08076_),
    .Y(_06623_),
    .A2(\soc_inst.cpu_core.id_rs2_data[18] ));
 sg13g2_nand2_1 _22129_ (.Y(_06624_),
    .A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B(_08075_));
 sg13g2_o21ai_1 _22130_ (.B1(_06624_),
    .Y(_06625_),
    .A1(_08076_),
    .A2(\soc_inst.cpu_core.id_rs2_data[18] ));
 sg13g2_a22oi_1 _22131_ (.Y(_06626_),
    .B1(_08074_),
    .B2(\soc_inst.cpu_core.id_rs2_data[19] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[20] ),
    .A1(_08073_));
 sg13g2_nor2b_1 _22132_ (.A(_06625_),
    .B_N(_06626_),
    .Y(_06627_));
 sg13g2_nand3_1 _22133_ (.B(_06623_),
    .C(_06627_),
    .A(_06620_),
    .Y(_06628_));
 sg13g2_a22oi_1 _22134_ (.Y(_06629_),
    .B1(\soc_inst.cpu_core.id_rs1_data[16] ),
    .B2(_08081_),
    .A2(_08079_),
    .A1(\soc_inst.cpu_core.id_rs1_data[17] ));
 sg13g2_o21ai_1 _22135_ (.B1(_06629_),
    .Y(_06630_),
    .A1(\soc_inst.cpu_core.id_rs1_data[16] ),
    .A2(_08081_));
 sg13g2_or2_1 _22136_ (.X(_06631_),
    .B(_06630_),
    .A(_06628_));
 sg13g2_a22oi_1 _22137_ (.Y(_06632_),
    .B1(_08047_),
    .B2(\soc_inst.cpu_core.id_rs2_data[12] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[13] ),
    .A1(_08045_));
 sg13g2_inv_1 _22138_ (.Y(_06633_),
    .A(_06632_));
 sg13g2_a22oi_1 _22139_ (.Y(_06634_),
    .B1(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B2(_08046_),
    .A2(_08044_),
    .A1(\soc_inst.cpu_core.id_rs1_data[14] ));
 sg13g2_a22oi_1 _22140_ (.Y(_06635_),
    .B1(_08043_),
    .B2(\soc_inst.cpu_core.id_rs2_data[14] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[15] ),
    .A1(_08041_));
 sg13g2_nand3_1 _22141_ (.B(_06634_),
    .C(_06635_),
    .A(_06632_),
    .Y(_06636_));
 sg13g2_nand2b_1 _22142_ (.Y(_06637_),
    .B(\soc_inst.cpu_core.id_rs1_data[8] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[8] ));
 sg13g2_nand2_1 _22143_ (.Y(_06638_),
    .A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .B(_08051_));
 sg13g2_nand2b_1 _22144_ (.Y(_06639_),
    .B(\soc_inst.cpu_core.id_rs1_data[9] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[9] ));
 sg13g2_nand3_1 _22145_ (.B(_06638_),
    .C(_06639_),
    .A(_06637_),
    .Y(_06640_));
 sg13g2_nand2b_1 _22146_ (.Y(_06641_),
    .B(\soc_inst.cpu_core.id_rs2_data[9] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[9] ));
 sg13g2_nand2b_1 _22147_ (.Y(_06642_),
    .B(\soc_inst.cpu_core.id_rs2_data[10] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[10] ));
 sg13g2_nand2b_1 _22148_ (.Y(_06643_),
    .B(\soc_inst.cpu_core.id_rs1_data[11] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[11] ));
 sg13g2_nand3_1 _22149_ (.B(_06642_),
    .C(_06643_),
    .A(_06641_),
    .Y(_06644_));
 sg13g2_a22oi_1 _22150_ (.Y(_06645_),
    .B1(_08054_),
    .B2(\soc_inst.cpu_core.id_rs2_data[8] ),
    .A2(_08042_),
    .A1(\soc_inst.cpu_core.id_rs1_data[15] ));
 sg13g2_nand2_1 _22151_ (.Y(_06646_),
    .A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .B(_08048_));
 sg13g2_nand2_1 _22152_ (.Y(_06647_),
    .A(_08049_),
    .B(\soc_inst.cpu_core.id_rs2_data[11] ));
 sg13g2_nand3_1 _22153_ (.B(_06646_),
    .C(_06647_),
    .A(_06645_),
    .Y(_06648_));
 sg13g2_nor4_1 _22154_ (.A(_06636_),
    .B(_06640_),
    .C(_06644_),
    .D(_06648_),
    .Y(_06649_));
 sg13g2_a22oi_1 _22155_ (.Y(_06650_),
    .B1(\soc_inst.cpu_core.id_rs1_data[6] ),
    .B2(_08036_),
    .A2(_08034_),
    .A1(\soc_inst.cpu_core.id_rs1_data[7] ));
 sg13g2_a21oi_1 _22156_ (.A1(_08033_),
    .A2(\soc_inst.cpu_core.id_rs2_data[7] ),
    .Y(_06651_),
    .B1(_06650_));
 sg13g2_a22oi_1 _22157_ (.Y(_06652_),
    .B1(_08035_),
    .B2(\soc_inst.cpu_core.id_rs2_data[6] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[7] ),
    .A1(_08033_));
 sg13g2_nand2_1 _22158_ (.Y(_06653_),
    .A(_06650_),
    .B(_06652_));
 sg13g2_nand2_1 _22159_ (.Y(_06654_),
    .A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .B(_08038_));
 sg13g2_nand2_1 _22160_ (.Y(_06655_),
    .A(_08037_),
    .B(\soc_inst.cpu_core.id_rs2_data[5] ));
 sg13g2_o21ai_1 _22161_ (.B1(_06655_),
    .Y(_06656_),
    .A1(\soc_inst.cpu_core.id_rs1_data[4] ),
    .A2(_08040_));
 sg13g2_nand2b_1 _22162_ (.Y(_06657_),
    .B(\soc_inst.cpu_core.id_rs1_data[2] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[2] ));
 sg13g2_nand2b_1 _22163_ (.Y(_06658_),
    .B(\soc_inst.cpu_core.id_rs1_data[3] ),
    .A_N(\soc_inst.cpu_core.id_rs2_data[3] ));
 sg13g2_nand2_1 _22164_ (.Y(_06659_),
    .A(_06657_),
    .B(_06658_));
 sg13g2_nand2b_1 _22165_ (.Y(_06660_),
    .B(\soc_inst.cpu_core.id_rs2_data[2] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[2] ));
 sg13g2_nand2b_1 _22166_ (.Y(_06661_),
    .B(\soc_inst.cpu_core.id_rs2_data[3] ),
    .A_N(\soc_inst.cpu_core.id_rs1_data[3] ));
 sg13g2_and4_1 _22167_ (.A(_06657_),
    .B(_06658_),
    .C(_06660_),
    .D(_06661_),
    .X(_06662_));
 sg13g2_a22oi_1 _22168_ (.Y(_06663_),
    .B1(_08030_),
    .B2(\soc_inst.cpu_core.id_rs2_data[1] ),
    .A2(\soc_inst.cpu_core.id_rs2_data[0] ),
    .A1(_08029_));
 sg13g2_nand2_1 _22169_ (.Y(_06664_),
    .A(_06662_),
    .B(_06663_));
 sg13g2_nor2b_1 _22170_ (.A(\soc_inst.cpu_core.id_rs2_data[1] ),
    .B_N(\soc_inst.cpu_core.id_rs1_data[1] ),
    .Y(_06665_));
 sg13g2_nor2_1 _22171_ (.A(_08039_),
    .B(\soc_inst.cpu_core.id_rs2_data[4] ),
    .Y(_06666_));
 sg13g2_a221oi_1 _22172_ (.B2(_06665_),
    .C1(_06666_),
    .B1(_06662_),
    .A1(_06659_),
    .Y(_06667_),
    .A2(_06661_));
 sg13g2_a21o_1 _22173_ (.A2(_06667_),
    .A1(_06664_),
    .B1(_06656_),
    .X(_06668_));
 sg13g2_a21oi_1 _22174_ (.A1(_06654_),
    .A2(_06668_),
    .Y(_06669_),
    .B1(_06653_));
 sg13g2_o21ai_1 _22175_ (.B1(_06649_),
    .Y(_06670_),
    .A1(_06651_),
    .A2(_06669_));
 sg13g2_and2_1 _22176_ (.A(_06637_),
    .B(_06639_),
    .X(_06671_));
 sg13g2_o21ai_1 _22177_ (.B1(_06638_),
    .Y(_06672_),
    .A1(_06644_),
    .A2(_06671_));
 sg13g2_nand2_1 _22178_ (.Y(_06673_),
    .A(_06643_),
    .B(_06646_));
 sg13g2_a21oi_1 _22179_ (.A1(_06647_),
    .A2(_06672_),
    .Y(_06674_),
    .B1(_06673_));
 sg13g2_o21ai_1 _22180_ (.B1(_06634_),
    .Y(_06675_),
    .A1(_06633_),
    .A2(_06674_));
 sg13g2_a22oi_1 _22181_ (.Y(_06676_),
    .B1(_06635_),
    .B2(_06675_),
    .A2(_08042_),
    .A1(\soc_inst.cpu_core.id_rs1_data[15] ));
 sg13g2_a21oi_1 _22182_ (.A1(_06670_),
    .A2(_06676_),
    .Y(_06677_),
    .B1(_06631_));
 sg13g2_a21oi_1 _22183_ (.A1(_08068_),
    .A2(\soc_inst.cpu_core.id_rs2_data[23] ),
    .Y(_06678_),
    .B1(_06618_));
 sg13g2_a21oi_1 _22184_ (.A1(_06625_),
    .A2(_06626_),
    .Y(_06679_),
    .B1(_06622_));
 sg13g2_nor2b_1 _22185_ (.A(_06679_),
    .B_N(_06620_),
    .Y(_06680_));
 sg13g2_nor2_1 _22186_ (.A(_06628_),
    .B(_06629_),
    .Y(_06681_));
 sg13g2_nor4_1 _22187_ (.A(_06677_),
    .B(_06678_),
    .C(_06680_),
    .D(_06681_),
    .Y(_06682_));
 sg13g2_nand3b_1 _22188_ (.B(_06615_),
    .C(_06608_),
    .Y(_06683_),
    .A_N(_06614_));
 sg13g2_nand2b_1 _22189_ (.Y(_06684_),
    .B(_06615_),
    .A_N(_06609_));
 sg13g2_nand3b_1 _22190_ (.B(_06683_),
    .C(_06684_),
    .Y(_06685_),
    .A_N(_06606_));
 sg13g2_o21ai_1 _22191_ (.B1(_06602_),
    .Y(_06686_),
    .A1(_06603_),
    .A2(_06610_));
 sg13g2_a21oi_1 _22192_ (.A1(_06612_),
    .A2(_06685_),
    .Y(_06687_),
    .B1(_06686_));
 sg13g2_o21ai_1 _22193_ (.B1(_06687_),
    .Y(_06688_),
    .A1(_06617_),
    .A2(_06682_));
 sg13g2_a21oi_2 _22194_ (.B1(_06603_),
    .Y(_06689_),
    .A2(_06688_),
    .A1(_06602_));
 sg13g2_nor2b_1 _22195_ (.A(\soc_inst.cpu_core.id_funct3[0] ),
    .B_N(\soc_inst.cpu_core.id_funct3[2] ),
    .Y(_06690_));
 sg13g2_nand2_1 _22196_ (.Y(_06691_),
    .A(\soc_inst.cpu_core.id_funct3[2] ),
    .B(\soc_inst.cpu_core.id_funct3[0] ));
 sg13g2_nand3b_1 _22197_ (.B(_06689_),
    .C(_06690_),
    .Y(_06692_),
    .A_N(\soc_inst.cpu_core.id_funct3[1] ));
 sg13g2_or3_1 _22198_ (.A(\soc_inst.cpu_core.id_funct3[1] ),
    .B(_06689_),
    .C(_06691_),
    .X(_06693_));
 sg13g2_o21ai_1 _22199_ (.B1(\soc_inst.cpu_core.id_funct3[1] ),
    .Y(_06694_),
    .A1(_06688_),
    .A2(_06690_));
 sg13g2_a21o_1 _22200_ (.A2(_06691_),
    .A1(_06688_),
    .B1(_06694_),
    .X(_06695_));
 sg13g2_nand3_1 _22201_ (.B(_06693_),
    .C(_06695_),
    .A(_06692_),
    .Y(_06696_));
 sg13g2_nor2b_1 _22202_ (.A(_06601_),
    .B_N(_06696_),
    .Y(_06697_));
 sg13g2_nand2_2 _22203_ (.Y(_06698_),
    .A(\soc_inst.cpu_core.id_funct3[0] ),
    .B(_11397_));
 sg13g2_o21ai_1 _22204_ (.B1(_06698_),
    .Y(_06699_),
    .A1(\soc_inst.cpu_core.id_pc[0] ),
    .A2(_06696_));
 sg13g2_o21ai_1 _22205_ (.B1(_06654_),
    .Y(_06700_),
    .A1(_08029_),
    .A2(\soc_inst.cpu_core.id_rs2_data[0] ));
 sg13g2_or4_1 _22206_ (.A(_06656_),
    .B(_06665_),
    .C(_06666_),
    .D(_06700_),
    .X(_06701_));
 sg13g2_nor4_1 _22207_ (.A(_06617_),
    .B(_06653_),
    .C(_06664_),
    .D(_06701_),
    .Y(_06702_));
 sg13g2_nand3b_1 _22208_ (.B(_06649_),
    .C(_06702_),
    .Y(_06703_),
    .A_N(_06631_));
 sg13g2_nor2b_2 _22209_ (.A(_06698_),
    .B_N(_06703_),
    .Y(_06704_));
 sg13g2_nor2_1 _22210_ (.A(_06698_),
    .B(_06703_),
    .Y(_06705_));
 sg13g2_a22oi_1 _22211_ (.Y(_06706_),
    .B1(_06705_),
    .B2(\soc_inst.cpu_core.id_pc[0] ),
    .A2(_06704_),
    .A1(_06601_));
 sg13g2_o21ai_1 _22212_ (.B1(_06706_),
    .Y(_06707_),
    .A1(_06697_),
    .A2(_06699_));
 sg13g2_and2_1 _22213_ (.A(_11398_),
    .B(_06703_),
    .X(_06708_));
 sg13g2_and4_1 _22214_ (.A(_00257_),
    .B(\soc_inst.cpu_core.id_instr[5] ),
    .C(net6306),
    .D(_11393_),
    .X(_06709_));
 sg13g2_nand4_1 _22215_ (.B(\soc_inst.cpu_core.id_instr[5] ),
    .C(net6306),
    .A(_00257_),
    .Y(_06710_),
    .D(_11393_));
 sg13g2_nor2_2 _22216_ (.A(_11399_),
    .B(_06703_),
    .Y(_06711_));
 sg13g2_a21oi_1 _22217_ (.A1(\soc_inst.cpu_core.id_pc[0] ),
    .A2(_06708_),
    .Y(_06712_),
    .B1(net5369));
 sg13g2_a22oi_1 _22218_ (.Y(_06713_),
    .B1(_06711_),
    .B2(_06601_),
    .A2(_06707_),
    .A1(_11399_));
 sg13g2_nand2_1 _22219_ (.Y(_06714_),
    .A(net5517),
    .B(_06601_));
 sg13g2_a221oi_1 _22220_ (.B2(net5370),
    .C1(net6369),
    .B1(_06714_),
    .A1(_06712_),
    .Y(_06715_),
    .A2(_06713_));
 sg13g2_a21o_1 _22221_ (.A2(net6366),
    .A1(net2434),
    .B1(_06715_),
    .X(_02342_));
 sg13g2_nor2_1 _22222_ (.A(_06696_),
    .B(_06704_),
    .Y(_06716_));
 sg13g2_nand2_1 _22223_ (.Y(_06717_),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xnor2_1 _22224_ (.Y(_06718_),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xor2_1 _22225_ (.B(_06718_),
    .A(_06600_),
    .X(_06719_));
 sg13g2_nand2_1 _22226_ (.Y(_06720_),
    .A(_08083_),
    .B(\soc_inst.cpu_core.id_is_compressed ));
 sg13g2_xor2_1 _22227_ (.B(\soc_inst.cpu_core.id_is_compressed ),
    .A(\soc_inst.cpu_core.id_pc[1] ),
    .X(_06721_));
 sg13g2_nor3_1 _22228_ (.A(_06696_),
    .B(_06704_),
    .C(_06721_),
    .Y(_06722_));
 sg13g2_o21ai_1 _22229_ (.B1(_11399_),
    .Y(_06723_),
    .A1(_06716_),
    .A2(_06719_));
 sg13g2_a221oi_1 _22230_ (.B2(_06708_),
    .C1(net5370),
    .B1(_06721_),
    .A1(_06711_),
    .Y(_06724_),
    .A2(_06719_));
 sg13g2_o21ai_1 _22231_ (.B1(_06724_),
    .Y(_06725_),
    .A1(_06722_),
    .A2(_06723_));
 sg13g2_nand2_1 _22232_ (.Y(_06726_),
    .A(\soc_inst.cpu_core.id_rs1_data[0] ),
    .B(\soc_inst.cpu_core.id_imm[0] ));
 sg13g2_nand2_1 _22233_ (.Y(_06727_),
    .A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xnor2_1 _22234_ (.Y(_06728_),
    .A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .B(\soc_inst.cpu_core.id_imm[1] ));
 sg13g2_xor2_1 _22235_ (.B(_06728_),
    .A(_06726_),
    .X(_06729_));
 sg13g2_a221oi_1 _22236_ (.B2(net6002),
    .C1(_06709_),
    .B1(_06729_),
    .A1(net5517),
    .Y(_06730_),
    .A2(_06719_));
 sg13g2_nor2_1 _22237_ (.A(net6369),
    .B(_06730_),
    .Y(_06731_));
 sg13g2_a22oi_1 _22238_ (.Y(_06732_),
    .B1(_06725_),
    .B2(_06731_),
    .A2(net3012),
    .A1(net6371));
 sg13g2_inv_1 _22239_ (.Y(_02343_),
    .A(_06732_));
 sg13g2_nand2_1 _22240_ (.Y(_06733_),
    .A(net6369),
    .B(net1784));
 sg13g2_nand2_1 _22241_ (.Y(_06734_),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .B(_06720_));
 sg13g2_xnor2_1 _22242_ (.Y(_06735_),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .B(_06720_));
 sg13g2_nor3_2 _22243_ (.A(_06696_),
    .B(_06704_),
    .C(_06711_),
    .Y(_06736_));
 sg13g2_and2_1 _22244_ (.A(_06709_),
    .B(_06736_),
    .X(_06737_));
 sg13g2_nand2_2 _22245_ (.Y(_06738_),
    .A(_06709_),
    .B(_06736_));
 sg13g2_and2_1 _22246_ (.A(\soc_inst.cpu_core.id_pc[2] ),
    .B(\soc_inst.cpu_core.id_imm[2] ),
    .X(_06739_));
 sg13g2_xor2_1 _22247_ (.B(\soc_inst.cpu_core.id_imm[2] ),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .X(_06740_));
 sg13g2_o21ai_1 _22248_ (.B1(_06717_),
    .Y(_06741_),
    .A1(_06600_),
    .A2(_06718_));
 sg13g2_xor2_1 _22249_ (.B(_06741_),
    .A(_06740_),
    .X(_06742_));
 sg13g2_and2_1 _22250_ (.A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .B(\soc_inst.cpu_core.id_imm[2] ),
    .X(_06743_));
 sg13g2_xor2_1 _22251_ (.B(\soc_inst.cpu_core.id_imm[2] ),
    .A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .X(_06744_));
 sg13g2_o21ai_1 _22252_ (.B1(_06727_),
    .Y(_06745_),
    .A1(_06726_),
    .A2(_06728_));
 sg13g2_nand2_1 _22253_ (.Y(_06746_),
    .A(_06744_),
    .B(_06745_));
 sg13g2_o21ai_1 _22254_ (.B1(net6002),
    .Y(_06747_),
    .A1(_06744_),
    .A2(_06745_));
 sg13g2_inv_1 _22255_ (.Y(_06748_),
    .A(_06747_));
 sg13g2_a22oi_1 _22256_ (.Y(_06749_),
    .B1(_06746_),
    .B2(_06748_),
    .A2(_06742_),
    .A1(net5517));
 sg13g2_nor2_2 _22257_ (.A(net5369),
    .B(_06736_),
    .Y(_06750_));
 sg13g2_nand2b_2 _22258_ (.Y(_06751_),
    .B(_06709_),
    .A_N(_06736_));
 sg13g2_a22oi_1 _22259_ (.Y(_06752_),
    .B1(_06749_),
    .B2(net5370),
    .A2(net4716),
    .A1(_06735_));
 sg13g2_o21ai_1 _22260_ (.B1(_06752_),
    .Y(_06753_),
    .A1(_06742_),
    .A2(_06751_));
 sg13g2_o21ai_1 _22261_ (.B1(_06733_),
    .Y(_02344_),
    .A1(net6370),
    .A2(_06753_));
 sg13g2_xnor2_1 _22262_ (.Y(_06754_),
    .A(\soc_inst.cpu_core.id_pc[3] ),
    .B(_06734_));
 sg13g2_nand2_1 _22263_ (.Y(_06755_),
    .A(\soc_inst.cpu_core.id_pc[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_xnor2_1 _22264_ (.Y(_06756_),
    .A(\soc_inst.cpu_core.id_pc[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_a21oi_1 _22265_ (.A1(_06740_),
    .A2(_06741_),
    .Y(_06757_),
    .B1(_06739_));
 sg13g2_xor2_1 _22266_ (.B(_06757_),
    .A(_06756_),
    .X(_06758_));
 sg13g2_nor2_1 _22267_ (.A(_06751_),
    .B(_06758_),
    .Y(_06759_));
 sg13g2_nand2_1 _22268_ (.Y(_06760_),
    .A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_xnor2_1 _22269_ (.Y(_06761_),
    .A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .B(\soc_inst.cpu_core.id_imm[3] ));
 sg13g2_a21oi_1 _22270_ (.A1(_06744_),
    .A2(_06745_),
    .Y(_06762_),
    .B1(_06743_));
 sg13g2_nor2_1 _22271_ (.A(_06761_),
    .B(_06762_),
    .Y(_06763_));
 sg13g2_a21o_1 _22272_ (.A2(_06762_),
    .A1(_06761_),
    .B1(net5999),
    .X(_06764_));
 sg13g2_a21oi_1 _22273_ (.A1(net5517),
    .A2(_06758_),
    .Y(_06765_),
    .B1(_06709_));
 sg13g2_o21ai_1 _22274_ (.B1(_06765_),
    .Y(_06766_),
    .A1(_06763_),
    .A2(_06764_));
 sg13g2_o21ai_1 _22275_ (.B1(_06766_),
    .Y(_06767_),
    .A1(_06738_),
    .A2(_06754_));
 sg13g2_nor3_1 _22276_ (.A(net6406),
    .B(_06759_),
    .C(_06767_),
    .Y(_06768_));
 sg13g2_a21o_1 _22277_ (.A2(net2914),
    .A1(net6411),
    .B1(_06768_),
    .X(_02345_));
 sg13g2_nor2_1 _22278_ (.A(_08087_),
    .B(_08088_),
    .Y(_06769_));
 sg13g2_xor2_1 _22279_ (.B(\soc_inst.cpu_core.id_imm[4] ),
    .A(\soc_inst.cpu_core.id_pc[4] ),
    .X(_06770_));
 sg13g2_o21ai_1 _22280_ (.B1(_06755_),
    .Y(_06771_),
    .A1(_06756_),
    .A2(_06757_));
 sg13g2_xor2_1 _22281_ (.B(_06771_),
    .A(_06770_),
    .X(_06772_));
 sg13g2_nor2_1 _22282_ (.A(_06751_),
    .B(_06772_),
    .Y(_06773_));
 sg13g2_nand4_1 _22283_ (.B(\soc_inst.cpu_core.id_pc[3] ),
    .C(\soc_inst.cpu_core.id_pc[4] ),
    .A(\soc_inst.cpu_core.id_pc[2] ),
    .Y(_06774_),
    .D(_06720_));
 sg13g2_o21ai_1 _22284_ (.B1(_08087_),
    .Y(_06775_),
    .A1(_08085_),
    .A2(_06734_));
 sg13g2_a21oi_1 _22285_ (.A1(_06774_),
    .A2(_06775_),
    .Y(_06776_),
    .B1(_06738_));
 sg13g2_nor2_1 _22286_ (.A(_08039_),
    .B(_08088_),
    .Y(_06777_));
 sg13g2_xor2_1 _22287_ (.B(\soc_inst.cpu_core.id_imm[4] ),
    .A(\soc_inst.cpu_core.id_rs1_data[4] ),
    .X(_06778_));
 sg13g2_o21ai_1 _22288_ (.B1(_06760_),
    .Y(_06779_),
    .A1(_06761_),
    .A2(_06762_));
 sg13g2_nand2_1 _22289_ (.Y(_06780_),
    .A(_06778_),
    .B(_06779_));
 sg13g2_nor2_1 _22290_ (.A(_06778_),
    .B(_06779_),
    .Y(_06781_));
 sg13g2_nor2_1 _22291_ (.A(net5999),
    .B(_06781_),
    .Y(_06782_));
 sg13g2_a221oi_1 _22292_ (.B2(_06782_),
    .C1(_06709_),
    .B1(_06780_),
    .A1(net5517),
    .Y(_06783_),
    .A2(_06772_));
 sg13g2_nor4_1 _22293_ (.A(net6407),
    .B(_06773_),
    .C(_06776_),
    .D(_06783_),
    .Y(_06784_));
 sg13g2_a21o_1 _22294_ (.A2(net2876),
    .A1(net6411),
    .B1(_06784_),
    .X(_02346_));
 sg13g2_nor2_1 _22295_ (.A(_08089_),
    .B(_06774_),
    .Y(_06785_));
 sg13g2_xnor2_1 _22296_ (.Y(_06786_),
    .A(_08089_),
    .B(_06774_));
 sg13g2_a21oi_1 _22297_ (.A1(_06770_),
    .A2(_06771_),
    .Y(_06787_),
    .B1(_06769_));
 sg13g2_nor2_1 _22298_ (.A(\soc_inst.cpu_core.id_pc[5] ),
    .B(\soc_inst.cpu_core.id_imm[5] ),
    .Y(_06788_));
 sg13g2_xor2_1 _22299_ (.B(\soc_inst.cpu_core.id_imm[5] ),
    .A(\soc_inst.cpu_core.id_pc[5] ),
    .X(_06789_));
 sg13g2_xnor2_1 _22300_ (.Y(_06790_),
    .A(_06787_),
    .B(_06789_));
 sg13g2_a21oi_1 _22301_ (.A1(_06778_),
    .A2(_06779_),
    .Y(_06791_),
    .B1(_06777_));
 sg13g2_nor2_1 _22302_ (.A(_08037_),
    .B(_08090_),
    .Y(_06792_));
 sg13g2_nor2_2 _22303_ (.A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .B(\soc_inst.cpu_core.id_imm[5] ),
    .Y(_06793_));
 sg13g2_nor3_1 _22304_ (.A(_06791_),
    .B(_06792_),
    .C(_06793_),
    .Y(_06794_));
 sg13g2_o21ai_1 _22305_ (.B1(_06791_),
    .Y(_06795_),
    .A1(_06792_),
    .A2(_06793_));
 sg13g2_nor2_1 _22306_ (.A(net5999),
    .B(_06794_),
    .Y(_06796_));
 sg13g2_a22oi_1 _22307_ (.Y(_06797_),
    .B1(_06795_),
    .B2(_06796_),
    .A2(_06790_),
    .A1(_11408_));
 sg13g2_a21oi_1 _22308_ (.A1(net5369),
    .A2(_06797_),
    .Y(_06798_),
    .B1(net6414));
 sg13g2_o21ai_1 _22309_ (.B1(_06798_),
    .Y(_06799_),
    .A1(_06751_),
    .A2(_06790_));
 sg13g2_a21oi_1 _22310_ (.A1(net4716),
    .A2(_06786_),
    .Y(_06800_),
    .B1(_06799_));
 sg13g2_a21o_1 _22311_ (.A2(net3073),
    .A1(net6411),
    .B1(_06800_),
    .X(_02347_));
 sg13g2_xnor2_1 _22312_ (.Y(_06801_),
    .A(\soc_inst.cpu_core.id_pc[6] ),
    .B(\soc_inst.cpu_core.id_imm[6] ));
 sg13g2_a221oi_1 _22313_ (.B2(_06771_),
    .C1(_06769_),
    .B1(_06770_),
    .A1(\soc_inst.cpu_core.id_pc[5] ),
    .Y(_06802_),
    .A2(\soc_inst.cpu_core.id_imm[5] ));
 sg13g2_nor3_1 _22314_ (.A(_06788_),
    .B(_06801_),
    .C(_06802_),
    .Y(_06803_));
 sg13g2_o21ai_1 _22315_ (.B1(_06801_),
    .Y(_06804_),
    .A1(_06788_),
    .A2(_06802_));
 sg13g2_nor2b_1 _22316_ (.A(_06803_),
    .B_N(_06804_),
    .Y(_06805_));
 sg13g2_nor2_1 _22317_ (.A(_06751_),
    .B(_06805_),
    .Y(_06806_));
 sg13g2_nor2_1 _22318_ (.A(_08035_),
    .B(_08092_),
    .Y(_06807_));
 sg13g2_xnor2_1 _22319_ (.Y(_06808_),
    .A(\soc_inst.cpu_core.id_rs1_data[6] ),
    .B(\soc_inst.cpu_core.id_imm[6] ));
 sg13g2_a221oi_1 _22320_ (.B2(_06779_),
    .C1(_06777_),
    .B1(_06778_),
    .A1(\soc_inst.cpu_core.id_rs1_data[5] ),
    .Y(_06809_),
    .A2(\soc_inst.cpu_core.id_imm[5] ));
 sg13g2_nor3_1 _22321_ (.A(_06793_),
    .B(_06808_),
    .C(_06809_),
    .Y(_06810_));
 sg13g2_o21ai_1 _22322_ (.B1(_06808_),
    .Y(_06811_),
    .A1(_06793_),
    .A2(_06809_));
 sg13g2_nor2_1 _22323_ (.A(net5999),
    .B(_06810_),
    .Y(_06812_));
 sg13g2_a22oi_1 _22324_ (.Y(_06813_),
    .B1(_06811_),
    .B2(_06812_),
    .A2(_06805_),
    .A1(_11408_));
 sg13g2_nor3_1 _22325_ (.A(_08089_),
    .B(_08091_),
    .C(_06774_),
    .Y(_06814_));
 sg13g2_xnor2_1 _22326_ (.Y(_06815_),
    .A(\soc_inst.cpu_core.id_pc[6] ),
    .B(_06785_));
 sg13g2_a221oi_1 _22327_ (.B2(net4716),
    .C1(_06806_),
    .B1(_06815_),
    .A1(net5369),
    .Y(_06816_),
    .A2(_06813_));
 sg13g2_mux2_1 _22328_ (.A0(net3036),
    .A1(_06816_),
    .S(net6156),
    .X(_02348_));
 sg13g2_nor2_2 _22329_ (.A(net5517),
    .B(_06750_),
    .Y(_06817_));
 sg13g2_nand2_2 _22330_ (.Y(_06818_),
    .A(_11409_),
    .B(_06751_));
 sg13g2_a21oi_1 _22331_ (.A1(\soc_inst.cpu_core.id_pc[6] ),
    .A2(\soc_inst.cpu_core.id_imm[6] ),
    .Y(_06819_),
    .B1(_06803_));
 sg13g2_nand2_1 _22332_ (.Y(_06820_),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .B(\soc_inst.cpu_core.id_imm[7] ));
 sg13g2_nor2_1 _22333_ (.A(\soc_inst.cpu_core.id_pc[7] ),
    .B(\soc_inst.cpu_core.id_imm[7] ),
    .Y(_06821_));
 sg13g2_xor2_1 _22334_ (.B(\soc_inst.cpu_core.id_imm[7] ),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .X(_06822_));
 sg13g2_xnor2_1 _22335_ (.Y(_06823_),
    .A(_06819_),
    .B(_06822_));
 sg13g2_nand2_1 _22336_ (.Y(_06824_),
    .A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .B(\soc_inst.cpu_core.id_imm[7] ));
 sg13g2_xor2_1 _22337_ (.B(\soc_inst.cpu_core.id_imm[7] ),
    .A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .X(_06825_));
 sg13g2_o21ai_1 _22338_ (.B1(_06825_),
    .Y(_06826_),
    .A1(_06807_),
    .A2(_06810_));
 sg13g2_nor3_1 _22339_ (.A(_06807_),
    .B(_06810_),
    .C(_06825_),
    .Y(_06827_));
 sg13g2_nor2_1 _22340_ (.A(net5999),
    .B(_06827_),
    .Y(_06828_));
 sg13g2_a21oi_1 _22341_ (.A1(_06826_),
    .A2(_06828_),
    .Y(_06829_),
    .B1(net6407));
 sg13g2_xnor2_1 _22342_ (.Y(_06830_),
    .A(_08093_),
    .B(_06814_));
 sg13g2_a22oi_1 _22343_ (.Y(_06831_),
    .B1(_06830_),
    .B2(net4716),
    .A2(_06823_),
    .A1(_06818_));
 sg13g2_a22oi_1 _22344_ (.Y(_02349_),
    .B1(_06829_),
    .B2(_06831_),
    .A2(_08119_),
    .A1(net6406));
 sg13g2_nand3_1 _22345_ (.B(\soc_inst.cpu_core.id_pc[8] ),
    .C(_06814_),
    .A(\soc_inst.cpu_core.id_pc[7] ),
    .Y(_06832_));
 sg13g2_a21o_1 _22346_ (.A2(_06814_),
    .A1(\soc_inst.cpu_core.id_pc[7] ),
    .B1(\soc_inst.cpu_core.id_pc[8] ),
    .X(_06833_));
 sg13g2_nand2_1 _22347_ (.Y(_06834_),
    .A(_06832_),
    .B(_06833_));
 sg13g2_nand2_1 _22348_ (.Y(_06835_),
    .A(\soc_inst.cpu_core.id_pc[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_xnor2_1 _22349_ (.Y(_06836_),
    .A(\soc_inst.cpu_core.id_pc[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_a21oi_1 _22350_ (.A1(_06819_),
    .A2(_06820_),
    .Y(_06837_),
    .B1(_06821_));
 sg13g2_inv_1 _22351_ (.Y(_06838_),
    .A(_06837_));
 sg13g2_xnor2_1 _22352_ (.Y(_06839_),
    .A(_06836_),
    .B(_06837_));
 sg13g2_xnor2_1 _22353_ (.Y(_06840_),
    .A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .B(\soc_inst.cpu_core.id_imm[8] ));
 sg13g2_a21oi_1 _22354_ (.A1(_06824_),
    .A2(_06826_),
    .Y(_06841_),
    .B1(_06840_));
 sg13g2_nand3_1 _22355_ (.B(_06826_),
    .C(_06840_),
    .A(_06824_),
    .Y(_06842_));
 sg13g2_nor2_1 _22356_ (.A(net5999),
    .B(_06841_),
    .Y(_06843_));
 sg13g2_a22oi_1 _22357_ (.Y(_06844_),
    .B1(_06842_),
    .B2(_06843_),
    .A2(_06839_),
    .A1(_11408_));
 sg13g2_o21ai_1 _22358_ (.B1(net6155),
    .Y(_06845_),
    .A1(_06751_),
    .A2(_06839_));
 sg13g2_a221oi_1 _22359_ (.B2(net5369),
    .C1(_06845_),
    .B1(_06844_),
    .A1(net4716),
    .Y(_06846_),
    .A2(_06834_));
 sg13g2_a21o_1 _22360_ (.A2(net2839),
    .A1(net6404),
    .B1(_06846_),
    .X(_02350_));
 sg13g2_xor2_1 _22361_ (.B(\soc_inst.cpu_core.id_imm[9] ),
    .A(\soc_inst.cpu_core.id_pc[9] ),
    .X(_06847_));
 sg13g2_o21ai_1 _22362_ (.B1(_06835_),
    .Y(_06848_),
    .A1(_06836_),
    .A2(_06838_));
 sg13g2_xnor2_1 _22363_ (.Y(_06849_),
    .A(_06847_),
    .B(_06848_));
 sg13g2_or2_1 _22364_ (.X(_06850_),
    .B(_06832_),
    .A(_08097_));
 sg13g2_xnor2_1 _22365_ (.Y(_06851_),
    .A(_08097_),
    .B(_06832_));
 sg13g2_xnor2_1 _22366_ (.Y(_06852_),
    .A(\soc_inst.cpu_core.id_rs1_data[9] ),
    .B(\soc_inst.cpu_core.id_imm[9] ));
 sg13g2_inv_1 _22367_ (.Y(_06853_),
    .A(_06852_));
 sg13g2_a21oi_1 _22368_ (.A1(\soc_inst.cpu_core.id_rs1_data[8] ),
    .A2(\soc_inst.cpu_core.id_imm[8] ),
    .Y(_06854_),
    .B1(_06841_));
 sg13g2_nand3_1 _22369_ (.B(\soc_inst.cpu_core.id_imm[8] ),
    .C(_06853_),
    .A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .Y(_06855_));
 sg13g2_o21ai_1 _22370_ (.B1(net6002),
    .Y(_06856_),
    .A1(_06852_),
    .A2(_06854_));
 sg13g2_a21oi_1 _22371_ (.A1(_06852_),
    .A2(_06854_),
    .Y(_06857_),
    .B1(_06856_));
 sg13g2_o21ai_1 _22372_ (.B1(net5369),
    .Y(_06858_),
    .A1(_11409_),
    .A2(_06849_));
 sg13g2_o21ai_1 _22373_ (.B1(net6155),
    .Y(_06859_),
    .A1(_06857_),
    .A2(_06858_));
 sg13g2_a221oi_1 _22374_ (.B2(net4716),
    .C1(_06859_),
    .B1(_06851_),
    .A1(_06750_),
    .Y(_06860_),
    .A2(_06849_));
 sg13g2_a21o_1 _22375_ (.A2(net2780),
    .A1(net6404),
    .B1(_06860_),
    .X(_02351_));
 sg13g2_nand2_1 _22376_ (.Y(_06861_),
    .A(\soc_inst.cpu_core.id_pc[10] ),
    .B(\soc_inst.cpu_core.id_imm[10] ));
 sg13g2_xor2_1 _22377_ (.B(\soc_inst.cpu_core.id_imm[10] ),
    .A(\soc_inst.cpu_core.id_pc[10] ),
    .X(_06862_));
 sg13g2_inv_1 _22378_ (.Y(_06863_),
    .A(_06862_));
 sg13g2_a21oi_1 _22379_ (.A1(_08097_),
    .A2(_08098_),
    .Y(_06864_),
    .B1(_06835_));
 sg13g2_nor2b_1 _22380_ (.A(_06836_),
    .B_N(_06847_),
    .Y(_06865_));
 sg13g2_a221oi_1 _22381_ (.B2(_06865_),
    .C1(_06864_),
    .B1(_06837_),
    .A1(\soc_inst.cpu_core.id_pc[9] ),
    .Y(_06866_),
    .A2(\soc_inst.cpu_core.id_imm[9] ));
 sg13g2_xnor2_1 _22382_ (.Y(_06867_),
    .A(_06862_),
    .B(_06866_));
 sg13g2_or2_1 _22383_ (.X(_06868_),
    .B(_06850_),
    .A(_08099_));
 sg13g2_xnor2_1 _22384_ (.Y(_06869_),
    .A(\soc_inst.cpu_core.id_pc[10] ),
    .B(_06850_));
 sg13g2_mux2_1 _22385_ (.A0(_06869_),
    .A1(_06867_),
    .S(_06696_),
    .X(_06870_));
 sg13g2_nand2_1 _22386_ (.Y(_06871_),
    .A(_06698_),
    .B(_06870_));
 sg13g2_a22oi_1 _22387_ (.Y(_06872_),
    .B1(_06869_),
    .B2(_06705_),
    .A2(_06867_),
    .A1(_06704_));
 sg13g2_nand2_1 _22388_ (.Y(_06873_),
    .A(_06871_),
    .B(_06872_));
 sg13g2_a21oi_1 _22389_ (.A1(_06708_),
    .A2(_06869_),
    .Y(_06874_),
    .B1(net5369));
 sg13g2_a22oi_1 _22390_ (.Y(_06875_),
    .B1(_06873_),
    .B2(_11399_),
    .A2(_06867_),
    .A1(_06711_));
 sg13g2_nand2_1 _22391_ (.Y(_06876_),
    .A(_08050_),
    .B(_08100_));
 sg13g2_nand2_1 _22392_ (.Y(_06877_),
    .A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .B(\soc_inst.cpu_core.id_imm[10] ));
 sg13g2_nand2_1 _22393_ (.Y(_06878_),
    .A(_06876_),
    .B(_06877_));
 sg13g2_o21ai_1 _22394_ (.B1(_06855_),
    .Y(_06879_),
    .A1(_08052_),
    .A2(_08098_));
 sg13g2_a21oi_1 _22395_ (.A1(_06841_),
    .A2(_06853_),
    .Y(_06880_),
    .B1(_06879_));
 sg13g2_or2_1 _22396_ (.X(_06881_),
    .B(_06880_),
    .A(_06878_));
 sg13g2_a21oi_1 _22397_ (.A1(_06878_),
    .A2(_06880_),
    .Y(_06882_),
    .B1(net5999));
 sg13g2_a22oi_1 _22398_ (.Y(_06883_),
    .B1(_06881_),
    .B2(_06882_),
    .A2(_06867_),
    .A1(net5517));
 sg13g2_a221oi_1 _22399_ (.B2(net5369),
    .C1(net6367),
    .B1(_06883_),
    .A1(_06874_),
    .Y(_06884_),
    .A2(_06875_));
 sg13g2_a21o_1 _22400_ (.A2(net2721),
    .A1(net6368),
    .B1(_06884_),
    .X(_02352_));
 sg13g2_nand2_1 _22401_ (.Y(_06885_),
    .A(net6404),
    .B(net1513));
 sg13g2_nand2_1 _22402_ (.Y(_06886_),
    .A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .B(\soc_inst.cpu_core.id_imm[11] ));
 sg13g2_xnor2_1 _22403_ (.Y(_06887_),
    .A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .B(\soc_inst.cpu_core.id_imm[11] ));
 sg13g2_a21o_1 _22404_ (.A2(_06881_),
    .A1(_06877_),
    .B1(_06887_),
    .X(_06888_));
 sg13g2_nand3_1 _22405_ (.B(_06881_),
    .C(_06887_),
    .A(_06877_),
    .Y(_06889_));
 sg13g2_xor2_1 _22406_ (.B(\soc_inst.cpu_core.id_imm[11] ),
    .A(\soc_inst.cpu_core.id_pc[11] ),
    .X(_06890_));
 sg13g2_o21ai_1 _22407_ (.B1(_06861_),
    .Y(_06891_),
    .A1(_06863_),
    .A2(_06866_));
 sg13g2_xnor2_1 _22408_ (.Y(_06892_),
    .A(_06890_),
    .B(_06891_));
 sg13g2_nand3_1 _22409_ (.B(_06888_),
    .C(_06889_),
    .A(net6002),
    .Y(_06893_));
 sg13g2_o21ai_1 _22410_ (.B1(_06893_),
    .Y(_06894_),
    .A1(_11409_),
    .A2(_06892_));
 sg13g2_nor2_2 _22411_ (.A(_08101_),
    .B(_06868_),
    .Y(_06895_));
 sg13g2_xnor2_1 _22412_ (.Y(_06896_),
    .A(_08101_),
    .B(_06868_));
 sg13g2_a22oi_1 _22413_ (.Y(_06897_),
    .B1(_06896_),
    .B2(_06737_),
    .A2(_06892_),
    .A1(_06750_));
 sg13g2_o21ai_1 _22414_ (.B1(_06897_),
    .Y(_06898_),
    .A1(_06709_),
    .A2(_06894_));
 sg13g2_o21ai_1 _22415_ (.B1(_06885_),
    .Y(_02353_),
    .A1(net6404),
    .A2(_06898_));
 sg13g2_nand2_1 _22416_ (.Y(_06899_),
    .A(net6356),
    .B(net2741));
 sg13g2_xnor2_1 _22417_ (.Y(_06900_),
    .A(\soc_inst.cpu_core.id_pc[12] ),
    .B(\soc_inst.cpu_core.id_imm[12] ));
 sg13g2_a21oi_1 _22418_ (.A1(_08101_),
    .A2(_08102_),
    .Y(_06901_),
    .B1(_06861_));
 sg13g2_a21oi_1 _22419_ (.A1(\soc_inst.cpu_core.id_pc[11] ),
    .A2(\soc_inst.cpu_core.id_imm[11] ),
    .Y(_06902_),
    .B1(_06901_));
 sg13g2_nand2_1 _22420_ (.Y(_06903_),
    .A(_06862_),
    .B(_06890_));
 sg13g2_o21ai_1 _22421_ (.B1(_06902_),
    .Y(_06904_),
    .A1(_06866_),
    .A2(_06903_));
 sg13g2_nor2b_1 _22422_ (.A(_06900_),
    .B_N(_06904_),
    .Y(_06905_));
 sg13g2_xnor2_1 _22423_ (.Y(_06906_),
    .A(_06900_),
    .B(_06904_));
 sg13g2_nor2b_1 _22424_ (.A(_06876_),
    .B_N(_06886_),
    .Y(_06907_));
 sg13g2_and2_1 _22425_ (.A(_06877_),
    .B(_06886_),
    .X(_06908_));
 sg13g2_a221oi_1 _22426_ (.B2(_06908_),
    .C1(_06907_),
    .B1(_06880_),
    .A1(_08049_),
    .Y(_06909_),
    .A2(_08102_));
 sg13g2_nand2_1 _22427_ (.Y(_06910_),
    .A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .B(\soc_inst.cpu_core.id_imm[12] ));
 sg13g2_xor2_1 _22428_ (.B(\soc_inst.cpu_core.id_imm[12] ),
    .A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .X(_06911_));
 sg13g2_inv_1 _22429_ (.Y(_06912_),
    .A(_06911_));
 sg13g2_and2_1 _22430_ (.A(_06909_),
    .B(_06911_),
    .X(_06913_));
 sg13g2_o21ai_1 _22431_ (.B1(net6001),
    .Y(_06914_),
    .A1(_06909_),
    .A2(_06911_));
 sg13g2_o21ai_1 _22432_ (.B1(net5370),
    .Y(_06915_),
    .A1(_06913_),
    .A2(_06914_));
 sg13g2_a21oi_1 _22433_ (.A1(net5517),
    .A2(_06906_),
    .Y(_06916_),
    .B1(_06915_));
 sg13g2_xnor2_1 _22434_ (.Y(_06917_),
    .A(\soc_inst.cpu_core.id_pc[12] ),
    .B(_06895_));
 sg13g2_a21oi_1 _22435_ (.A1(_06737_),
    .A2(_06917_),
    .Y(_06918_),
    .B1(net6355));
 sg13g2_o21ai_1 _22436_ (.B1(_06918_),
    .Y(_06919_),
    .A1(_06751_),
    .A2(_06906_));
 sg13g2_o21ai_1 _22437_ (.B1(_06899_),
    .Y(_02354_),
    .A1(_06916_),
    .A2(_06919_));
 sg13g2_nand3_1 _22438_ (.B(\soc_inst.cpu_core.id_pc[13] ),
    .C(_06895_),
    .A(\soc_inst.cpu_core.id_pc[12] ),
    .Y(_06920_));
 sg13g2_a21o_1 _22439_ (.A2(_06895_),
    .A1(\soc_inst.cpu_core.id_pc[12] ),
    .B1(\soc_inst.cpu_core.id_pc[13] ),
    .X(_06921_));
 sg13g2_nand2_1 _22440_ (.Y(_06922_),
    .A(_06920_),
    .B(_06921_));
 sg13g2_nand2_1 _22441_ (.Y(_06923_),
    .A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ));
 sg13g2_xnor2_1 _22442_ (.Y(_06924_),
    .A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ));
 sg13g2_a21oi_1 _22443_ (.A1(\soc_inst.cpu_core.id_rs1_data[12] ),
    .A2(\soc_inst.cpu_core.id_imm[12] ),
    .Y(_06925_),
    .B1(_06913_));
 sg13g2_nor2_1 _22444_ (.A(_06912_),
    .B(_06924_),
    .Y(_06926_));
 sg13g2_a21oi_1 _22445_ (.A1(_06924_),
    .A2(_06925_),
    .Y(_06927_),
    .B1(net5998));
 sg13g2_o21ai_1 _22446_ (.B1(_06927_),
    .Y(_06928_),
    .A1(_06924_),
    .A2(_06925_));
 sg13g2_o21ai_1 _22447_ (.B1(_06928_),
    .Y(_06929_),
    .A1(_06738_),
    .A2(_06922_));
 sg13g2_nor2_1 _22448_ (.A(net6355),
    .B(_06929_),
    .Y(_06930_));
 sg13g2_or2_1 _22449_ (.X(_06931_),
    .B(\soc_inst.cpu_core.id_imm[13] ),
    .A(\soc_inst.cpu_core.id_pc[13] ));
 sg13g2_nand2_1 _22450_ (.Y(_06932_),
    .A(\soc_inst.cpu_core.id_pc[13] ),
    .B(\soc_inst.cpu_core.id_imm[13] ));
 sg13g2_nand2_1 _22451_ (.Y(_06933_),
    .A(_06931_),
    .B(_06932_));
 sg13g2_a21oi_1 _22452_ (.A1(\soc_inst.cpu_core.id_pc[12] ),
    .A2(\soc_inst.cpu_core.id_imm[12] ),
    .Y(_06934_),
    .B1(_06905_));
 sg13g2_o21ai_1 _22453_ (.B1(net4713),
    .Y(_06935_),
    .A1(_06933_),
    .A2(_06934_));
 sg13g2_a21o_1 _22454_ (.A2(_06934_),
    .A1(_06933_),
    .B1(_06935_),
    .X(_06936_));
 sg13g2_a22oi_1 _22455_ (.Y(_02355_),
    .B1(_06930_),
    .B2(_06936_),
    .A2(_08120_),
    .A1(net6354));
 sg13g2_nor2_1 _22456_ (.A(\soc_inst.cpu_core.id_pc[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ),
    .Y(_06937_));
 sg13g2_and2_1 _22457_ (.A(\soc_inst.cpu_core.id_pc[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ),
    .X(_06938_));
 sg13g2_nand2_1 _22458_ (.Y(_06939_),
    .A(\soc_inst.cpu_core.id_pc[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ));
 sg13g2_nor2_1 _22459_ (.A(_06937_),
    .B(_06938_),
    .Y(_06940_));
 sg13g2_o21ai_1 _22460_ (.B1(_06932_),
    .Y(_06941_),
    .A1(_08103_),
    .A2(_08104_));
 sg13g2_o21ai_1 _22461_ (.B1(_06931_),
    .Y(_06942_),
    .A1(_06905_),
    .A2(_06941_));
 sg13g2_xnor2_1 _22462_ (.Y(_06943_),
    .A(_06940_),
    .B(_06942_));
 sg13g2_nand2_1 _22463_ (.Y(_06944_),
    .A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ));
 sg13g2_xnor2_1 _22464_ (.Y(_06945_),
    .A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .B(\soc_inst.cpu_core.id_imm[14] ));
 sg13g2_o21ai_1 _22465_ (.B1(_06923_),
    .Y(_06946_),
    .A1(_06910_),
    .A2(_06924_));
 sg13g2_a21oi_1 _22466_ (.A1(_06909_),
    .A2(_06926_),
    .Y(_06947_),
    .B1(_06946_));
 sg13g2_nand2_1 _22467_ (.Y(_06948_),
    .A(_06945_),
    .B(_06947_));
 sg13g2_nor2_1 _22468_ (.A(_06945_),
    .B(_06947_),
    .Y(_06949_));
 sg13g2_nor2_1 _22469_ (.A(net5998),
    .B(_06949_),
    .Y(_06950_));
 sg13g2_or2_1 _22470_ (.X(_06951_),
    .B(_06920_),
    .A(_08106_));
 sg13g2_xnor2_1 _22471_ (.Y(_06952_),
    .A(\soc_inst.cpu_core.id_pc[14] ),
    .B(_06920_));
 sg13g2_a22oi_1 _22472_ (.Y(_06953_),
    .B1(_06952_),
    .B2(net4716),
    .A2(_06950_),
    .A1(_06948_));
 sg13g2_a21oi_1 _22473_ (.A1(net4713),
    .A2(_06943_),
    .Y(_06954_),
    .B1(net6353));
 sg13g2_a22oi_1 _22474_ (.Y(_02356_),
    .B1(_06953_),
    .B2(_06954_),
    .A2(_08121_),
    .A1(net6352));
 sg13g2_xnor2_1 _22475_ (.Y(_06955_),
    .A(\soc_inst.cpu_core.id_pc[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_o21ai_1 _22476_ (.B1(_06939_),
    .Y(_06956_),
    .A1(_06937_),
    .A2(_06942_));
 sg13g2_nand2_1 _22477_ (.Y(_06957_),
    .A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_nor2_1 _22478_ (.A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ),
    .Y(_06958_));
 sg13g2_xnor2_1 _22479_ (.Y(_06959_),
    .A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .B(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_a21oi_1 _22480_ (.A1(\soc_inst.cpu_core.id_rs1_data[14] ),
    .A2(\soc_inst.cpu_core.id_imm[14] ),
    .Y(_06960_),
    .B1(_06949_));
 sg13g2_nor2_1 _22481_ (.A(_08107_),
    .B(_06951_),
    .Y(_06961_));
 sg13g2_nand2_1 _22482_ (.Y(_06962_),
    .A(_08107_),
    .B(_06951_));
 sg13g2_nand3b_1 _22483_ (.B(_06962_),
    .C(net4715),
    .Y(_06963_),
    .A_N(_06961_));
 sg13g2_xor2_1 _22484_ (.B(_06956_),
    .A(_06955_),
    .X(_06964_));
 sg13g2_nor2_1 _22485_ (.A(_06817_),
    .B(_06964_),
    .Y(_06965_));
 sg13g2_o21ai_1 _22486_ (.B1(net6001),
    .Y(_06966_),
    .A1(_06959_),
    .A2(_06960_));
 sg13g2_a21oi_1 _22487_ (.A1(_06959_),
    .A2(_06960_),
    .Y(_06967_),
    .B1(_06966_));
 sg13g2_nor3_1 _22488_ (.A(net6352),
    .B(_06965_),
    .C(_06967_),
    .Y(_06968_));
 sg13g2_a22oi_1 _22489_ (.Y(_02357_),
    .B1(_06963_),
    .B2(_06968_),
    .A2(_08122_),
    .A1(net6344));
 sg13g2_nor2_1 _22490_ (.A(net6143),
    .B(net2005),
    .Y(_06969_));
 sg13g2_nor2_1 _22491_ (.A(_06945_),
    .B(_06959_),
    .Y(_06970_));
 sg13g2_and2_1 _22492_ (.A(_06926_),
    .B(_06970_),
    .X(_06971_));
 sg13g2_o21ai_1 _22493_ (.B1(_06957_),
    .Y(_06972_),
    .A1(_06944_),
    .A2(_06958_));
 sg13g2_a221oi_1 _22494_ (.B2(_06909_),
    .C1(_06972_),
    .B1(_06971_),
    .A1(_06946_),
    .Y(_06973_),
    .A2(_06970_));
 sg13g2_xor2_1 _22495_ (.B(\soc_inst.cpu_core.id_imm[16] ),
    .A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .X(_06974_));
 sg13g2_nor2b_1 _22496_ (.A(_06973_),
    .B_N(_06974_),
    .Y(_06975_));
 sg13g2_nand2b_1 _22497_ (.Y(_06976_),
    .B(_06974_),
    .A_N(_06973_));
 sg13g2_nor2b_1 _22498_ (.A(_06974_),
    .B_N(_06973_),
    .Y(_06977_));
 sg13g2_nor2_1 _22499_ (.A(net5998),
    .B(_06977_),
    .Y(_06978_));
 sg13g2_nor3_1 _22500_ (.A(_06937_),
    .B(_06938_),
    .C(_06955_),
    .Y(_06979_));
 sg13g2_inv_1 _22501_ (.Y(_06980_),
    .A(_06979_));
 sg13g2_nor3_1 _22502_ (.A(_06900_),
    .B(_06933_),
    .C(_06980_),
    .Y(_06981_));
 sg13g2_o21ai_1 _22503_ (.B1(_06938_),
    .Y(_06982_),
    .A1(\soc_inst.cpu_core.id_pc[15] ),
    .A2(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_nand3_1 _22504_ (.B(_06941_),
    .C(_06979_),
    .A(_06931_),
    .Y(_06983_));
 sg13g2_nand2_1 _22505_ (.Y(_06984_),
    .A(_06982_),
    .B(_06983_));
 sg13g2_a221oi_1 _22506_ (.B2(_06981_),
    .C1(_06984_),
    .B1(_06904_),
    .A1(\soc_inst.cpu_core.id_pc[15] ),
    .Y(_06985_),
    .A2(\soc_inst.cpu_core.id_imm[15] ));
 sg13g2_nand2_1 _22507_ (.Y(_06986_),
    .A(\soc_inst.cpu_core.id_pc[16] ),
    .B(\soc_inst.cpu_core.id_imm[16] ));
 sg13g2_xnor2_1 _22508_ (.Y(_06987_),
    .A(\soc_inst.cpu_core.id_pc[16] ),
    .B(\soc_inst.cpu_core.id_imm[16] ));
 sg13g2_xnor2_1 _22509_ (.Y(_06988_),
    .A(_08108_),
    .B(_06961_));
 sg13g2_o21ai_1 _22510_ (.B1(net4713),
    .Y(_06989_),
    .A1(_06985_),
    .A2(_06987_));
 sg13g2_a21oi_1 _22511_ (.A1(_06985_),
    .A2(_06987_),
    .Y(_06990_),
    .B1(_06989_));
 sg13g2_a221oi_1 _22512_ (.B2(net4715),
    .C1(_06990_),
    .B1(_06988_),
    .A1(_06976_),
    .Y(_06991_),
    .A2(_06978_));
 sg13g2_a21oi_1 _22513_ (.A1(net6143),
    .A2(_06991_),
    .Y(_02358_),
    .B1(_06969_));
 sg13g2_nand2_1 _22514_ (.Y(_06992_),
    .A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ));
 sg13g2_xor2_1 _22515_ (.B(\soc_inst.cpu_core.id_imm[17] ),
    .A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .X(_06993_));
 sg13g2_a21oi_1 _22516_ (.A1(\soc_inst.cpu_core.id_rs1_data[16] ),
    .A2(\soc_inst.cpu_core.id_imm[16] ),
    .Y(_06994_),
    .B1(_06993_));
 sg13g2_nand2b_1 _22517_ (.Y(_06995_),
    .B(_06994_),
    .A_N(_06975_));
 sg13g2_nand2_1 _22518_ (.Y(_06996_),
    .A(_06974_),
    .B(_06993_));
 sg13g2_nand2_1 _22519_ (.Y(_06997_),
    .A(_06975_),
    .B(_06993_));
 sg13g2_nand3_1 _22520_ (.B(\soc_inst.cpu_core.id_imm[16] ),
    .C(_06993_),
    .A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .Y(_06998_));
 sg13g2_and4_1 _22521_ (.A(net6000),
    .B(_06995_),
    .C(_06997_),
    .D(_06998_),
    .X(_06999_));
 sg13g2_nor4_2 _22522_ (.A(_08107_),
    .B(_08108_),
    .C(_08109_),
    .Y(_07000_),
    .D(_06951_));
 sg13g2_a21oi_1 _22523_ (.A1(\soc_inst.cpu_core.id_pc[16] ),
    .A2(_06961_),
    .Y(_07001_),
    .B1(\soc_inst.cpu_core.id_pc[17] ));
 sg13g2_nor3_1 _22524_ (.A(_06738_),
    .B(_07000_),
    .C(_07001_),
    .Y(_07002_));
 sg13g2_nor2_1 _22525_ (.A(\soc_inst.cpu_core.id_pc[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ),
    .Y(_07003_));
 sg13g2_xnor2_1 _22526_ (.Y(_07004_),
    .A(\soc_inst.cpu_core.id_pc[17] ),
    .B(\soc_inst.cpu_core.id_imm[17] ));
 sg13g2_o21ai_1 _22527_ (.B1(_06986_),
    .Y(_07005_),
    .A1(_06985_),
    .A2(_06987_));
 sg13g2_xnor2_1 _22528_ (.Y(_07006_),
    .A(_07004_),
    .B(_07005_));
 sg13g2_nand2_1 _22529_ (.Y(_07007_),
    .A(net4713),
    .B(_07006_));
 sg13g2_nor3_1 _22530_ (.A(net6345),
    .B(_06999_),
    .C(_07002_),
    .Y(_07008_));
 sg13g2_a22oi_1 _22531_ (.Y(_02359_),
    .B1(_07007_),
    .B2(_07008_),
    .A2(_08123_),
    .A1(net6345));
 sg13g2_or2_1 _22532_ (.X(_07009_),
    .B(\soc_inst.cpu_core.id_imm[18] ),
    .A(\soc_inst.cpu_core.id_pc[18] ));
 sg13g2_nand2_1 _22533_ (.Y(_07010_),
    .A(\soc_inst.cpu_core.id_pc[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_inv_1 _22534_ (.Y(_07011_),
    .A(_07010_));
 sg13g2_nand2_1 _22535_ (.Y(_07012_),
    .A(_07009_),
    .B(_07010_));
 sg13g2_a22oi_1 _22536_ (.Y(_07013_),
    .B1(\soc_inst.cpu_core.id_pc[17] ),
    .B2(\soc_inst.cpu_core.id_imm[17] ),
    .A2(\soc_inst.cpu_core.id_imm[16] ),
    .A1(\soc_inst.cpu_core.id_pc[16] ));
 sg13g2_o21ai_1 _22537_ (.B1(_07013_),
    .Y(_07014_),
    .A1(_06985_),
    .A2(_06987_));
 sg13g2_nor2b_1 _22538_ (.A(_07003_),
    .B_N(_07014_),
    .Y(_07015_));
 sg13g2_xnor2_1 _22539_ (.Y(_07016_),
    .A(_07012_),
    .B(_07015_));
 sg13g2_xnor2_1 _22540_ (.Y(_07017_),
    .A(_08110_),
    .B(_07000_));
 sg13g2_a221oi_1 _22541_ (.B2(net4715),
    .C1(net6345),
    .B1(_07017_),
    .A1(net4713),
    .Y(_07018_),
    .A2(_07016_));
 sg13g2_nand2_1 _22542_ (.Y(_07019_),
    .A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_xnor2_1 _22543_ (.Y(_07020_),
    .A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .B(\soc_inst.cpu_core.id_imm[18] ));
 sg13g2_and2_1 _22544_ (.A(_06992_),
    .B(_06998_),
    .X(_07021_));
 sg13g2_a21o_1 _22545_ (.A2(_07021_),
    .A1(_06997_),
    .B1(_07020_),
    .X(_07022_));
 sg13g2_nand3_1 _22546_ (.B(_07020_),
    .C(_07021_),
    .A(_06997_),
    .Y(_07023_));
 sg13g2_nand3_1 _22547_ (.B(_07022_),
    .C(_07023_),
    .A(net6000),
    .Y(_07024_));
 sg13g2_a22oi_1 _22548_ (.Y(_02360_),
    .B1(_07018_),
    .B2(_07024_),
    .A2(_08124_),
    .A1(net6381));
 sg13g2_nor2_1 _22549_ (.A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ),
    .Y(_07025_));
 sg13g2_xnor2_1 _22550_ (.Y(_07026_),
    .A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ));
 sg13g2_nand3_1 _22551_ (.B(_07022_),
    .C(_07026_),
    .A(_07019_),
    .Y(_07027_));
 sg13g2_a21o_1 _22552_ (.A2(_07022_),
    .A1(_07019_),
    .B1(_07026_),
    .X(_07028_));
 sg13g2_nand3_1 _22553_ (.B(_07027_),
    .C(_07028_),
    .A(net6000),
    .Y(_07029_));
 sg13g2_nand2_1 _22554_ (.Y(_07030_),
    .A(\soc_inst.cpu_core.id_pc[19] ),
    .B(\soc_inst.cpu_core.id_imm[19] ));
 sg13g2_or2_1 _22555_ (.X(_07031_),
    .B(\soc_inst.cpu_core.id_imm[19] ),
    .A(\soc_inst.cpu_core.id_pc[19] ));
 sg13g2_nand2_1 _22556_ (.Y(_07032_),
    .A(_07030_),
    .B(_07031_));
 sg13g2_a21oi_1 _22557_ (.A1(_07009_),
    .A2(_07015_),
    .Y(_07033_),
    .B1(_07011_));
 sg13g2_xor2_1 _22558_ (.B(_07033_),
    .A(_07032_),
    .X(_07034_));
 sg13g2_nand3_1 _22559_ (.B(\soc_inst.cpu_core.id_pc[19] ),
    .C(_07000_),
    .A(\soc_inst.cpu_core.id_pc[18] ),
    .Y(_07035_));
 sg13g2_a21o_1 _22560_ (.A2(_07000_),
    .A1(\soc_inst.cpu_core.id_pc[18] ),
    .B1(\soc_inst.cpu_core.id_pc[19] ),
    .X(_07036_));
 sg13g2_and2_1 _22561_ (.A(_07035_),
    .B(_07036_),
    .X(_07037_));
 sg13g2_a221oi_1 _22562_ (.B2(net4715),
    .C1(net6381),
    .B1(_07037_),
    .A1(net4713),
    .Y(_07038_),
    .A2(_07034_));
 sg13g2_a22oi_1 _22563_ (.Y(_02361_),
    .B1(_07029_),
    .B2(_07038_),
    .A2(_08125_),
    .A1(net6381));
 sg13g2_or2_1 _22564_ (.X(_07039_),
    .B(_07032_),
    .A(_07012_));
 sg13g2_or3_1 _22565_ (.A(_06987_),
    .B(_07004_),
    .C(_07039_),
    .X(_07040_));
 sg13g2_nand2_1 _22566_ (.Y(_07041_),
    .A(_07010_),
    .B(_07030_));
 sg13g2_nor3_1 _22567_ (.A(_07003_),
    .B(_07013_),
    .C(_07039_),
    .Y(_07042_));
 sg13g2_a21oi_1 _22568_ (.A1(_07031_),
    .A2(_07041_),
    .Y(_07043_),
    .B1(_07042_));
 sg13g2_o21ai_1 _22569_ (.B1(_07043_),
    .Y(_07044_),
    .A1(_06985_),
    .A2(_07040_));
 sg13g2_xnor2_1 _22570_ (.Y(_07045_),
    .A(\soc_inst.cpu_core.id_pc[20] ),
    .B(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_xnor2_1 _22571_ (.Y(_07046_),
    .A(_07044_),
    .B(_07045_));
 sg13g2_nor2_1 _22572_ (.A(_08112_),
    .B(_07035_),
    .Y(_07047_));
 sg13g2_xnor2_1 _22573_ (.Y(_07048_),
    .A(\soc_inst.cpu_core.id_pc[20] ),
    .B(_07035_));
 sg13g2_a221oi_1 _22574_ (.B2(net4715),
    .C1(net6383),
    .B1(_07048_),
    .A1(net4714),
    .Y(_07049_),
    .A2(_07046_));
 sg13g2_nand2_1 _22575_ (.Y(_07050_),
    .A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .B(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_xor2_1 _22576_ (.B(\soc_inst.cpu_core.id_imm[20] ),
    .A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .X(_07051_));
 sg13g2_inv_1 _22577_ (.Y(_07052_),
    .A(_07051_));
 sg13g2_or2_1 _22578_ (.X(_07053_),
    .B(_07026_),
    .A(_07020_));
 sg13g2_nor3_1 _22579_ (.A(_06973_),
    .B(_06996_),
    .C(_07053_),
    .Y(_07054_));
 sg13g2_or2_1 _22580_ (.X(_07055_),
    .B(_07025_),
    .A(_07019_));
 sg13g2_inv_1 _22581_ (.Y(_07056_),
    .A(_07055_));
 sg13g2_a21oi_1 _22582_ (.A1(\soc_inst.cpu_core.id_rs1_data[19] ),
    .A2(\soc_inst.cpu_core.id_imm[19] ),
    .Y(_07057_),
    .B1(_07056_));
 sg13g2_o21ai_1 _22583_ (.B1(_07057_),
    .Y(_07058_),
    .A1(_07021_),
    .A2(_07053_));
 sg13g2_or3_1 _22584_ (.A(_07051_),
    .B(_07054_),
    .C(_07058_),
    .X(_07059_));
 sg13g2_o21ai_1 _22585_ (.B1(_07051_),
    .Y(_07060_),
    .A1(_07054_),
    .A2(_07058_));
 sg13g2_nand3_1 _22586_ (.B(_07059_),
    .C(_07060_),
    .A(net6000),
    .Y(_07061_));
 sg13g2_a22oi_1 _22587_ (.Y(_02362_),
    .B1(_07049_),
    .B2(_07061_),
    .A2(_08126_),
    .A1(net6382));
 sg13g2_nand2_1 _22588_ (.Y(_07062_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_nor2_1 _22589_ (.A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ),
    .Y(_07063_));
 sg13g2_xnor2_1 _22590_ (.Y(_07064_),
    .A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_nand3_1 _22591_ (.B(_07060_),
    .C(_07064_),
    .A(_07050_),
    .Y(_07065_));
 sg13g2_a21o_1 _22592_ (.A2(_07060_),
    .A1(_07050_),
    .B1(_07064_),
    .X(_07066_));
 sg13g2_and2_1 _22593_ (.A(net6000),
    .B(_07065_),
    .X(_07067_));
 sg13g2_xnor2_1 _22594_ (.Y(_07068_),
    .A(\soc_inst.cpu_core.id_pc[21] ),
    .B(\soc_inst.cpu_core.id_imm[21] ));
 sg13g2_a21o_1 _22595_ (.A2(\soc_inst.cpu_core.id_imm[20] ),
    .A1(\soc_inst.cpu_core.id_pc[20] ),
    .B1(_07044_),
    .X(_07069_));
 sg13g2_o21ai_1 _22596_ (.B1(_07069_),
    .Y(_07070_),
    .A1(\soc_inst.cpu_core.id_pc[20] ),
    .A2(\soc_inst.cpu_core.id_imm[20] ));
 sg13g2_xor2_1 _22597_ (.B(_07070_),
    .A(_07068_),
    .X(_07071_));
 sg13g2_nand2_1 _22598_ (.Y(_07072_),
    .A(net4714),
    .B(_07071_));
 sg13g2_nor3_1 _22599_ (.A(_08112_),
    .B(_08113_),
    .C(_07035_),
    .Y(_07073_));
 sg13g2_xnor2_1 _22600_ (.Y(_07074_),
    .A(_08113_),
    .B(_07047_));
 sg13g2_a221oi_1 _22601_ (.B2(net4715),
    .C1(net6382),
    .B1(_07074_),
    .A1(_07066_),
    .Y(_07075_),
    .A2(_07067_));
 sg13g2_a22oi_1 _22602_ (.Y(_02363_),
    .B1(_07072_),
    .B2(_07075_),
    .A2(_08127_),
    .A1(net6383));
 sg13g2_and2_1 _22603_ (.A(net3403),
    .B(\soc_inst.cpu_core.id_imm[22] ),
    .X(_07076_));
 sg13g2_xnor2_1 _22604_ (.Y(_07077_),
    .A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ));
 sg13g2_nand3_1 _22605_ (.B(_07066_),
    .C(_07077_),
    .A(_07062_),
    .Y(_07078_));
 sg13g2_a21oi_1 _22606_ (.A1(_07062_),
    .A2(_07066_),
    .Y(_07079_),
    .B1(_07077_));
 sg13g2_nor2_1 _22607_ (.A(net5998),
    .B(_07079_),
    .Y(_07080_));
 sg13g2_nor2_1 _22608_ (.A(\soc_inst.cpu_core.id_pc[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ),
    .Y(_07081_));
 sg13g2_nand2_1 _22609_ (.Y(_07082_),
    .A(\soc_inst.cpu_core.id_pc[22] ),
    .B(\soc_inst.cpu_core.id_imm[22] ));
 sg13g2_nor2b_1 _22610_ (.A(_07081_),
    .B_N(_07082_),
    .Y(_07083_));
 sg13g2_a22oi_1 _22611_ (.Y(_07084_),
    .B1(\soc_inst.cpu_core.id_pc[21] ),
    .B2(\soc_inst.cpu_core.id_imm[21] ),
    .A2(\soc_inst.cpu_core.id_imm[20] ),
    .A1(\soc_inst.cpu_core.id_pc[20] ));
 sg13g2_nor2_1 _22612_ (.A(_07045_),
    .B(_07068_),
    .Y(_07085_));
 sg13g2_a21oi_1 _22613_ (.A1(_08113_),
    .A2(_08114_),
    .Y(_07086_),
    .B1(_07084_));
 sg13g2_a21oi_1 _22614_ (.A1(_07044_),
    .A2(_07085_),
    .Y(_07087_),
    .B1(_07086_));
 sg13g2_nand2_1 _22615_ (.Y(_07088_),
    .A(\soc_inst.cpu_core.id_pc[22] ),
    .B(_07073_));
 sg13g2_xnor2_1 _22616_ (.Y(_07089_),
    .A(_08115_),
    .B(_07073_));
 sg13g2_xnor2_1 _22617_ (.Y(_07090_),
    .A(_07083_),
    .B(_07087_));
 sg13g2_nand2_1 _22618_ (.Y(_07091_),
    .A(net4713),
    .B(_07090_));
 sg13g2_a221oi_1 _22619_ (.B2(net4715),
    .C1(net6382),
    .B1(_07089_),
    .A1(_07078_),
    .Y(_07092_),
    .A2(_07080_));
 sg13g2_a22oi_1 _22620_ (.Y(_02364_),
    .B1(_07091_),
    .B2(_07092_),
    .A2(_08128_),
    .A1(net6382));
 sg13g2_xor2_1 _22621_ (.B(\soc_inst.cpu_core.id_imm[23] ),
    .A(\soc_inst.cpu_core.id_rs1_data[23] ),
    .X(_07093_));
 sg13g2_o21ai_1 _22622_ (.B1(_07093_),
    .Y(_07094_),
    .A1(_07076_),
    .A2(_07079_));
 sg13g2_or3_1 _22623_ (.A(_07076_),
    .B(_07079_),
    .C(_07093_),
    .X(_07095_));
 sg13g2_nand3_1 _22624_ (.B(net3404),
    .C(_07095_),
    .A(net6000),
    .Y(_07096_));
 sg13g2_nor2_1 _22625_ (.A(\soc_inst.cpu_core.id_pc[23] ),
    .B(\soc_inst.cpu_core.id_imm[23] ),
    .Y(_07097_));
 sg13g2_nand2_1 _22626_ (.Y(_07098_),
    .A(\soc_inst.cpu_core.id_pc[23] ),
    .B(\soc_inst.cpu_core.id_imm[23] ));
 sg13g2_nor2b_2 _22627_ (.A(_07097_),
    .B_N(_07098_),
    .Y(_07099_));
 sg13g2_o21ai_1 _22628_ (.B1(_07082_),
    .Y(_07100_),
    .A1(_07081_),
    .A2(_07087_));
 sg13g2_nor2_1 _22629_ (.A(_08116_),
    .B(_07088_),
    .Y(_07101_));
 sg13g2_xnor2_1 _22630_ (.Y(_07102_),
    .A(_08116_),
    .B(_07088_));
 sg13g2_nor2_1 _22631_ (.A(net5370),
    .B(_07102_),
    .Y(_07103_));
 sg13g2_o21ai_1 _22632_ (.B1(_06817_),
    .Y(_07104_),
    .A1(net5370),
    .A2(_07102_));
 sg13g2_xor2_1 _22633_ (.B(_07100_),
    .A(_07099_),
    .X(_07105_));
 sg13g2_a221oi_1 _22634_ (.B2(_07105_),
    .C1(net6382),
    .B1(_07104_),
    .A1(_06736_),
    .Y(_07106_),
    .A2(_07103_));
 sg13g2_a22oi_1 _22635_ (.Y(_02365_),
    .B1(_07096_),
    .B2(_07106_),
    .A2(_08129_),
    .A1(net6382));
 sg13g2_nand2_1 _22636_ (.Y(_07107_),
    .A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .B(\soc_inst.cpu_core.id_imm[24] ));
 sg13g2_xnor2_1 _22637_ (.Y(_07108_),
    .A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .B(\soc_inst.cpu_core.id_imm[24] ));
 sg13g2_inv_1 _22638_ (.Y(_07109_),
    .A(_07108_));
 sg13g2_nand2b_1 _22639_ (.Y(_07110_),
    .B(_07093_),
    .A_N(_07077_));
 sg13g2_nor2_1 _22640_ (.A(_07052_),
    .B(_07064_),
    .Y(_07111_));
 sg13g2_nand2b_1 _22641_ (.Y(_07112_),
    .B(_07111_),
    .A_N(_07110_));
 sg13g2_o21ai_1 _22642_ (.B1(_07076_),
    .Y(_07113_),
    .A1(\soc_inst.cpu_core.id_rs1_data[23] ),
    .A2(\soc_inst.cpu_core.id_imm[23] ));
 sg13g2_o21ai_1 _22643_ (.B1(_07062_),
    .Y(_07114_),
    .A1(_07050_),
    .A2(_07063_));
 sg13g2_nor4_1 _22644_ (.A(_06973_),
    .B(_06996_),
    .C(_07053_),
    .D(_07112_),
    .Y(_07115_));
 sg13g2_a21oi_1 _22645_ (.A1(_07058_),
    .A2(_07111_),
    .Y(_07116_),
    .B1(_07114_));
 sg13g2_nor2_1 _22646_ (.A(_07110_),
    .B(_07116_),
    .Y(_07117_));
 sg13g2_a21oi_1 _22647_ (.A1(\soc_inst.cpu_core.id_rs1_data[23] ),
    .A2(\soc_inst.cpu_core.id_imm[23] ),
    .Y(_07118_),
    .B1(_07117_));
 sg13g2_nand2_1 _22648_ (.Y(_07119_),
    .A(_07113_),
    .B(_07118_));
 sg13g2_o21ai_1 _22649_ (.B1(_07109_),
    .Y(_07120_),
    .A1(_07115_),
    .A2(_07119_));
 sg13g2_or3_1 _22650_ (.A(_07109_),
    .B(_07115_),
    .C(_07119_),
    .X(_07121_));
 sg13g2_nand3_1 _22651_ (.B(_07120_),
    .C(_07121_),
    .A(net6001),
    .Y(_07122_));
 sg13g2_and3_1 _22652_ (.X(_07123_),
    .A(_07083_),
    .B(_07085_),
    .C(_07099_));
 sg13g2_o21ai_1 _22653_ (.B1(_07098_),
    .Y(_07124_),
    .A1(_07082_),
    .A2(_07097_));
 sg13g2_nand3_1 _22654_ (.B(_07086_),
    .C(_07099_),
    .A(_07083_),
    .Y(_07125_));
 sg13g2_nand2b_1 _22655_ (.Y(_07126_),
    .B(_07125_),
    .A_N(_07124_));
 sg13g2_a21o_2 _22656_ (.A2(_07123_),
    .A1(_07044_),
    .B1(_07126_),
    .X(_07127_));
 sg13g2_xor2_1 _22657_ (.B(_07127_),
    .A(\soc_inst.cpu_core.id_imm[24] ),
    .X(_07128_));
 sg13g2_a221oi_1 _22658_ (.B2(net4714),
    .C1(net6383),
    .B1(_07128_),
    .A1(net4715),
    .Y(_07129_),
    .A2(_07101_));
 sg13g2_a22oi_1 _22659_ (.Y(_02366_),
    .B1(_07122_),
    .B2(_07129_),
    .A2(_08178_),
    .A1(net6384));
 sg13g2_nor2_1 _22660_ (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B(\soc_inst.cpu_core.id_imm[25] ),
    .Y(_07130_));
 sg13g2_and2_1 _22661_ (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B(\soc_inst.cpu_core.id_imm[25] ),
    .X(_07131_));
 sg13g2_nand2_1 _22662_ (.Y(_07132_),
    .A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .B(\soc_inst.cpu_core.id_imm[25] ));
 sg13g2_nand2b_1 _22663_ (.Y(_07133_),
    .B(_07132_),
    .A_N(_07130_));
 sg13g2_a21oi_1 _22664_ (.A1(_07107_),
    .A2(_07120_),
    .Y(_07134_),
    .B1(_07133_));
 sg13g2_nand3_1 _22665_ (.B(_07120_),
    .C(_07133_),
    .A(_07107_),
    .Y(_07135_));
 sg13g2_nor2_1 _22666_ (.A(net5998),
    .B(_07134_),
    .Y(_07136_));
 sg13g2_a21oi_1 _22667_ (.A1(\soc_inst.cpu_core.id_imm[24] ),
    .A2(_07127_),
    .Y(_07137_),
    .B1(\soc_inst.cpu_core.id_imm[25] ));
 sg13g2_and3_2 _22668_ (.X(_07138_),
    .A(\soc_inst.cpu_core.id_imm[24] ),
    .B(\soc_inst.cpu_core.id_imm[25] ),
    .C(_07127_));
 sg13g2_or3_1 _22669_ (.A(_06817_),
    .B(_07137_),
    .C(_07138_),
    .X(_07139_));
 sg13g2_a21oi_1 _22670_ (.A1(_07135_),
    .A2(_07136_),
    .Y(_07140_),
    .B1(net6383));
 sg13g2_a22oi_1 _22671_ (.Y(_02367_),
    .B1(_07139_),
    .B2(_07140_),
    .A2(_08180_),
    .A1(net6384));
 sg13g2_nor2_1 _22672_ (.A(net6147),
    .B(net2303),
    .Y(_07141_));
 sg13g2_nand2_1 _22673_ (.Y(_07142_),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .B(\soc_inst.cpu_core.id_imm[26] ));
 sg13g2_xor2_1 _22674_ (.B(\soc_inst.cpu_core.id_imm[26] ),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .X(_07143_));
 sg13g2_xnor2_1 _22675_ (.Y(_07144_),
    .A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .B(\soc_inst.cpu_core.id_imm[26] ));
 sg13g2_nor3_1 _22676_ (.A(_07131_),
    .B(_07134_),
    .C(_07143_),
    .Y(_07145_));
 sg13g2_o21ai_1 _22677_ (.B1(_07143_),
    .Y(_07146_),
    .A1(_07131_),
    .A2(_07134_));
 sg13g2_and2_1 _22678_ (.A(\soc_inst.cpu_core.id_imm[26] ),
    .B(_07138_),
    .X(_07147_));
 sg13g2_xor2_1 _22679_ (.B(_07138_),
    .A(\soc_inst.cpu_core.id_imm[26] ),
    .X(_07148_));
 sg13g2_nor2_1 _22680_ (.A(net5998),
    .B(_07145_),
    .Y(_07149_));
 sg13g2_a22oi_1 _22681_ (.Y(_07150_),
    .B1(_07149_),
    .B2(_07146_),
    .A2(_07148_),
    .A1(net4713));
 sg13g2_a21oi_1 _22682_ (.A1(net6147),
    .A2(_07150_),
    .Y(_02368_),
    .B1(_07141_));
 sg13g2_xnor2_1 _22683_ (.Y(_07151_),
    .A(\soc_inst.cpu_core.id_rs1_data[27] ),
    .B(\soc_inst.cpu_core.id_imm[27] ));
 sg13g2_nand2_1 _22684_ (.Y(_07152_),
    .A(_07142_),
    .B(_07146_));
 sg13g2_xor2_1 _22685_ (.B(_07152_),
    .A(_07151_),
    .X(_07153_));
 sg13g2_a21oi_1 _22686_ (.A1(\soc_inst.cpu_core.id_imm[27] ),
    .A2(_07147_),
    .Y(_07154_),
    .B1(_06817_));
 sg13g2_o21ai_1 _22687_ (.B1(_07154_),
    .Y(_07155_),
    .A1(\soc_inst.cpu_core.id_imm[27] ),
    .A2(_07147_));
 sg13g2_o21ai_1 _22688_ (.B1(_07155_),
    .Y(_07156_),
    .A1(net5998),
    .A2(_07153_));
 sg13g2_mux2_1 _22689_ (.A0(net3093),
    .A1(_07156_),
    .S(net6150),
    .X(_02369_));
 sg13g2_nor2_1 _22690_ (.A(_07144_),
    .B(_07151_),
    .Y(_07157_));
 sg13g2_nand2b_1 _22691_ (.Y(_07158_),
    .B(_07157_),
    .A_N(_07133_));
 sg13g2_o21ai_1 _22692_ (.B1(_07132_),
    .Y(_07159_),
    .A1(_07107_),
    .A2(_07130_));
 sg13g2_a21oi_1 _22693_ (.A1(_08061_),
    .A2(_08117_),
    .Y(_07160_),
    .B1(_07142_));
 sg13g2_a221oi_1 _22694_ (.B2(_07159_),
    .C1(_07160_),
    .B1(_07157_),
    .A1(\soc_inst.cpu_core.id_rs1_data[27] ),
    .Y(_07161_),
    .A2(\soc_inst.cpu_core.id_imm[27] ));
 sg13g2_o21ai_1 _22695_ (.B1(_07161_),
    .Y(_07162_),
    .A1(_07120_),
    .A2(_07158_));
 sg13g2_xor2_1 _22696_ (.B(\soc_inst.cpu_core.id_imm[28] ),
    .A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .X(_07163_));
 sg13g2_or2_1 _22697_ (.X(_07164_),
    .B(_07163_),
    .A(_07162_));
 sg13g2_nand2_1 _22698_ (.Y(_07165_),
    .A(_07162_),
    .B(_07163_));
 sg13g2_nand3_1 _22699_ (.B(_07164_),
    .C(_07165_),
    .A(net6000),
    .Y(_07166_));
 sg13g2_a21oi_1 _22700_ (.A1(\soc_inst.cpu_core.id_imm[27] ),
    .A2(_07147_),
    .Y(_07167_),
    .B1(\soc_inst.cpu_core.id_imm[28] ));
 sg13g2_and4_1 _22701_ (.A(\soc_inst.cpu_core.id_imm[26] ),
    .B(\soc_inst.cpu_core.id_imm[27] ),
    .C(\soc_inst.cpu_core.id_imm[28] ),
    .D(_07138_),
    .X(_07168_));
 sg13g2_nor3_1 _22702_ (.A(_06817_),
    .B(_07167_),
    .C(_07168_),
    .Y(_07169_));
 sg13g2_nor2_1 _22703_ (.A(net6385),
    .B(_07169_),
    .Y(_07170_));
 sg13g2_a22oi_1 _22704_ (.Y(_02370_),
    .B1(_07166_),
    .B2(_07170_),
    .A2(_08181_),
    .A1(net6386));
 sg13g2_a21oi_1 _22705_ (.A1(\soc_inst.cpu_core.id_imm[29] ),
    .A2(_07168_),
    .Y(_07171_),
    .B1(_06817_));
 sg13g2_o21ai_1 _22706_ (.B1(_07171_),
    .Y(_07172_),
    .A1(\soc_inst.cpu_core.id_imm[29] ),
    .A2(_07168_));
 sg13g2_xor2_1 _22707_ (.B(\soc_inst.cpu_core.id_imm[29] ),
    .A(\soc_inst.cpu_core.id_rs1_data[29] ),
    .X(_07173_));
 sg13g2_a21oi_1 _22708_ (.A1(\soc_inst.cpu_core.id_rs1_data[28] ),
    .A2(\soc_inst.cpu_core.id_imm[28] ),
    .Y(_07174_),
    .B1(_07173_));
 sg13g2_and2_1 _22709_ (.A(_07163_),
    .B(_07173_),
    .X(_07175_));
 sg13g2_nand2_1 _22710_ (.Y(_07176_),
    .A(_07162_),
    .B(_07175_));
 sg13g2_nand3_1 _22711_ (.B(\soc_inst.cpu_core.id_imm[28] ),
    .C(_07173_),
    .A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .Y(_07177_));
 sg13g2_inv_1 _22712_ (.Y(_07178_),
    .A(_07177_));
 sg13g2_a21oi_1 _22713_ (.A1(_07165_),
    .A2(_07174_),
    .Y(_07179_),
    .B1(_07178_));
 sg13g2_and2_1 _22714_ (.A(net6000),
    .B(_07179_),
    .X(_07180_));
 sg13g2_a21oi_1 _22715_ (.A1(_07176_),
    .A2(_07180_),
    .Y(_07181_),
    .B1(net6387));
 sg13g2_a22oi_1 _22716_ (.Y(_02371_),
    .B1(_07172_),
    .B2(_07181_),
    .A2(_08182_),
    .A1(net6387));
 sg13g2_a221oi_1 _22717_ (.B2(_07175_),
    .C1(_07178_),
    .B1(_07162_),
    .A1(\soc_inst.cpu_core.id_rs1_data[29] ),
    .Y(_07182_),
    .A2(\soc_inst.cpu_core.id_imm[29] ));
 sg13g2_nand2_1 _22718_ (.Y(_07183_),
    .A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .B(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_xnor2_1 _22719_ (.Y(_07184_),
    .A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .B(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_a21oi_1 _22720_ (.A1(_07182_),
    .A2(_07184_),
    .Y(_07185_),
    .B1(net5998));
 sg13g2_o21ai_1 _22721_ (.B1(_07185_),
    .Y(_07186_),
    .A1(_07182_),
    .A2(_07184_));
 sg13g2_a21oi_1 _22722_ (.A1(\soc_inst.cpu_core.id_imm[29] ),
    .A2(_07168_),
    .Y(_07187_),
    .B1(\soc_inst.cpu_core.id_imm[30] ));
 sg13g2_nand3_1 _22723_ (.B(\soc_inst.cpu_core.id_imm[30] ),
    .C(_07168_),
    .A(\soc_inst.cpu_core.id_imm[29] ),
    .Y(_07188_));
 sg13g2_nor2_1 _22724_ (.A(_06817_),
    .B(_07187_),
    .Y(_07189_));
 sg13g2_a21oi_1 _22725_ (.A1(_07188_),
    .A2(_07189_),
    .Y(_07190_),
    .B1(net6393));
 sg13g2_a22oi_1 _22726_ (.Y(_02372_),
    .B1(_07186_),
    .B2(_07190_),
    .A2(_08183_),
    .A1(net6393));
 sg13g2_o21ai_1 _22727_ (.B1(_07183_),
    .Y(_07191_),
    .A1(_07182_),
    .A2(_07184_));
 sg13g2_xnor2_1 _22728_ (.Y(_07192_),
    .A(\soc_inst.cpu_core.id_rs1_data[31] ),
    .B(\soc_inst.cpu_core.id_imm[31] ));
 sg13g2_xnor2_1 _22729_ (.Y(_07193_),
    .A(_07191_),
    .B(_07192_));
 sg13g2_xnor2_1 _22730_ (.Y(_07194_),
    .A(\soc_inst.cpu_core.id_imm[31] ),
    .B(_07188_));
 sg13g2_a221oi_1 _22731_ (.B2(net4714),
    .C1(net6393),
    .B1(_07194_),
    .A1(net6001),
    .Y(_07195_),
    .A2(_07193_));
 sg13g2_a21oi_1 _22732_ (.A1(net6394),
    .A2(_08185_),
    .Y(_02373_),
    .B1(_07195_));
 sg13g2_nor3_2 _22733_ (.A(_11022_),
    .B(_11329_),
    .C(net3345),
    .Y(_07196_));
 sg13g2_a21oi_1 _22734_ (.A1(net6501),
    .A2(_08414_),
    .Y(_07197_),
    .B1(_11338_));
 sg13g2_nor2_1 _22735_ (.A(net6483),
    .B(net6202),
    .Y(_07198_));
 sg13g2_nor3_1 _22736_ (.A(_11340_),
    .B(_07197_),
    .C(_07198_),
    .Y(_07199_));
 sg13g2_mux2_1 _22737_ (.A0(net6202),
    .A1(_07199_),
    .S(_07196_),
    .X(_02374_));
 sg13g2_nand2_1 _22738_ (.Y(_07200_),
    .A(_11339_),
    .B(_11342_));
 sg13g2_a21oi_1 _22739_ (.A1(_11340_),
    .A2(_07196_),
    .Y(_07201_),
    .B1(net6201));
 sg13g2_a21oi_1 _22740_ (.A1(_07196_),
    .A2(_07200_),
    .Y(_02375_),
    .B1(_07201_));
 sg13g2_nand2_2 _22741_ (.Y(_07202_),
    .A(_09029_),
    .B(_09513_));
 sg13g2_inv_1 _22742_ (.Y(_07203_),
    .A(_07202_));
 sg13g2_nand2_2 _22743_ (.Y(_07204_),
    .A(_09042_),
    .B(_09513_));
 sg13g2_and3_2 _22744_ (.X(_07205_),
    .A(_09042_),
    .B(net5146),
    .C(_09513_));
 sg13g2_a21o_1 _22745_ (.A2(net4928),
    .A1(net4944),
    .B1(_07205_),
    .X(_07206_));
 sg13g2_a21oi_1 _22746_ (.A1(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .A2(net6100),
    .Y(_07207_),
    .B1(net5047));
 sg13g2_nor2_1 _22747_ (.A(net6213),
    .B(net5071),
    .Y(_07208_));
 sg13g2_nor2_1 _22748_ (.A(\soc_inst.cpu_core.ex_branch_target[5] ),
    .B(net5159),
    .Y(_07209_));
 sg13g2_nor2_1 _22749_ (.A(\soc_inst.cpu_core.ex_alu_result[5] ),
    .B(net5167),
    .Y(_07210_));
 sg13g2_nor4_1 _22750_ (.A(_07207_),
    .B(_07208_),
    .C(_07209_),
    .D(_07210_),
    .Y(_07211_));
 sg13g2_a21oi_1 _22751_ (.A1(net2312),
    .A2(_09894_),
    .Y(_07212_),
    .B1(\soc_inst.cpu_core.mem_rs1_data[5] ));
 sg13g2_a21oi_1 _22752_ (.A1(net5148),
    .A2(net5527),
    .Y(_07213_),
    .B1(_09895_));
 sg13g2_nor2_1 _22753_ (.A(_07212_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_mux2_1 _22754_ (.A0(_07214_),
    .A1(_07211_),
    .S(net4929),
    .X(_07215_));
 sg13g2_a21o_1 _22755_ (.A2(net4748),
    .A1(net2312),
    .B1(_07215_),
    .X(_02376_));
 sg13g2_a22oi_1 _22756_ (.Y(_07216_),
    .B1(net5163),
    .B2(\soc_inst.cpu_core.ex_branch_target[6] ),
    .A2(net5076),
    .A1(\soc_inst.cpu_core.ex_instr[6] ));
 sg13g2_nor2_1 _22757_ (.A(\soc_inst.cpu_core.ex_alu_result[6] ),
    .B(net5166),
    .Y(_07217_));
 sg13g2_a21oi_1 _22758_ (.A1(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .A2(net6100),
    .Y(_07218_),
    .B1(_08950_));
 sg13g2_nor4_1 _22759_ (.A(net5076),
    .B(net5163),
    .C(_07217_),
    .D(_07218_),
    .Y(_07219_));
 sg13g2_a21oi_1 _22760_ (.A1(net1202),
    .A2(net4949),
    .Y(_07220_),
    .B1(_07219_));
 sg13g2_a221oi_1 _22761_ (.B2(net1202),
    .C1(net4785),
    .B1(_09901_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .Y(_07221_),
    .A2(net5326));
 sg13g2_and3_1 _22762_ (.X(_07222_),
    .A(net4784),
    .B(_07216_),
    .C(_07220_));
 sg13g2_nand2_1 _22763_ (.Y(_07223_),
    .A(net1202),
    .B(_07205_));
 sg13g2_o21ai_1 _22764_ (.B1(_07223_),
    .Y(_02377_),
    .A1(_07221_),
    .A2(_07222_));
 sg13g2_a21oi_1 _22765_ (.A1(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .A2(net6100),
    .Y(_07224_),
    .B1(net5048));
 sg13g2_a221oi_1 _22766_ (.B2(_08119_),
    .C1(_07224_),
    .B1(_08964_),
    .A1(_08165_),
    .Y(_07225_),
    .A2(net5169));
 sg13g2_o21ai_1 _22767_ (.B1(_07225_),
    .Y(_07226_),
    .A1(\soc_inst.cpu_core.ex_instr[7] ),
    .A2(net5072));
 sg13g2_a221oi_1 _22768_ (.B2(net2264),
    .C1(net4929),
    .B1(_11139_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .Y(_07227_),
    .A2(net5326));
 sg13g2_a221oi_1 _22769_ (.B2(net4784),
    .C1(_07227_),
    .B1(_07226_),
    .A1(net5148),
    .Y(_07228_),
    .A2(_07203_));
 sg13g2_a21o_1 _22770_ (.A2(net4749),
    .A1(net2264),
    .B1(_07228_),
    .X(_02378_));
 sg13g2_a21oi_1 _22771_ (.A1(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .A2(net6101),
    .Y(_07229_),
    .B1(net5048));
 sg13g2_nor2_1 _22772_ (.A(\soc_inst.cpu_core.ex_instr[8] ),
    .B(net5072),
    .Y(_07230_));
 sg13g2_nor2_1 _22773_ (.A(\soc_inst.cpu_core.ex_branch_target[8] ),
    .B(net5158),
    .Y(_07231_));
 sg13g2_nor2_1 _22774_ (.A(\soc_inst.cpu_core.ex_alu_result[8] ),
    .B(net5166),
    .Y(_07232_));
 sg13g2_nor4_1 _22775_ (.A(_07229_),
    .B(_07230_),
    .C(_07231_),
    .D(_07232_),
    .Y(_07233_));
 sg13g2_a21oi_1 _22776_ (.A1(net2786),
    .A2(net4951),
    .Y(_07234_),
    .B1(_07233_));
 sg13g2_a221oi_1 _22777_ (.B2(net2786),
    .C1(net4930),
    .B1(_09905_),
    .A1(net1413),
    .Y(_07235_),
    .A2(_09899_));
 sg13g2_a21oi_1 _22778_ (.A1(net4784),
    .A2(_07234_),
    .Y(_07236_),
    .B1(_07235_));
 sg13g2_a21o_1 _22779_ (.A2(_07205_),
    .A1(net2786),
    .B1(_07236_),
    .X(_02379_));
 sg13g2_nand2b_1 _22780_ (.Y(_07237_),
    .B(_08145_),
    .A_N(net5048));
 sg13g2_nor2_1 _22781_ (.A(\soc_inst.cpu_core.ex_instr[9] ),
    .B(net5071),
    .Y(_07238_));
 sg13g2_nor2_1 _22782_ (.A(\soc_inst.cpu_core.ex_alu_result[9] ),
    .B(net5166),
    .Y(_07239_));
 sg13g2_nor2_1 _22783_ (.A(\soc_inst.cpu_core.ex_branch_target[9] ),
    .B(net5158),
    .Y(_07240_));
 sg13g2_nor4_1 _22784_ (.A(_09137_),
    .B(_07238_),
    .C(_07239_),
    .D(_07240_),
    .Y(_07241_));
 sg13g2_a22oi_1 _22785_ (.Y(_07242_),
    .B1(_07237_),
    .B2(_07241_),
    .A2(net4950),
    .A1(net2396));
 sg13g2_a221oi_1 _22786_ (.B2(net2396),
    .C1(net4930),
    .B1(_09909_),
    .A1(net1456),
    .Y(_07243_),
    .A2(net5326));
 sg13g2_a21oi_1 _22787_ (.A1(net4784),
    .A2(_07242_),
    .Y(_07244_),
    .B1(_07243_));
 sg13g2_a21o_1 _22788_ (.A2(_07205_),
    .A1(net2396),
    .B1(_07244_),
    .X(_02380_));
 sg13g2_a21oi_1 _22789_ (.A1(net1401),
    .A2(net6101),
    .Y(_07245_),
    .B1(net5047));
 sg13g2_nor2_1 _22790_ (.A(\soc_inst.cpu_core.ex_instr[10] ),
    .B(net5072),
    .Y(_07246_));
 sg13g2_nor2_1 _22791_ (.A(\soc_inst.cpu_core.ex_branch_target[10] ),
    .B(net5158),
    .Y(_07247_));
 sg13g2_nor2_1 _22792_ (.A(\soc_inst.cpu_core.ex_alu_result[10] ),
    .B(net5166),
    .Y(_07248_));
 sg13g2_nor4_1 _22793_ (.A(_07245_),
    .B(_07246_),
    .C(_07247_),
    .D(_07248_),
    .Y(_07249_));
 sg13g2_nand2_1 _22794_ (.Y(_07250_),
    .A(net4929),
    .B(_07249_));
 sg13g2_a22oi_1 _22795_ (.Y(_07251_),
    .B1(_09915_),
    .B2(net5534),
    .A2(_09913_),
    .A1(net2261));
 sg13g2_o21ai_1 _22796_ (.B1(_07250_),
    .Y(_07252_),
    .A1(net4929),
    .A2(_07251_));
 sg13g2_a21o_1 _22797_ (.A2(net4748),
    .A1(net2261),
    .B1(_07252_),
    .X(_02381_));
 sg13g2_a21oi_1 _22798_ (.A1(net3409),
    .A2(net6101),
    .Y(_07253_),
    .B1(net5047));
 sg13g2_nor2_1 _22799_ (.A(\soc_inst.cpu_core.ex_instr[11] ),
    .B(net5072),
    .Y(_07254_));
 sg13g2_nor2_1 _22800_ (.A(\soc_inst.cpu_core.ex_branch_target[11] ),
    .B(net5158),
    .Y(_07255_));
 sg13g2_nor2_1 _22801_ (.A(\soc_inst.cpu_core.ex_alu_result[11] ),
    .B(net5167),
    .Y(_07256_));
 sg13g2_nor4_2 _22802_ (.A(_07253_),
    .B(_07254_),
    .C(_07255_),
    .Y(_07257_),
    .D(_07256_));
 sg13g2_a21oi_1 _22803_ (.A1(net2252),
    .A2(net4948),
    .Y(_07258_),
    .B1(_07257_));
 sg13g2_a221oi_1 _22804_ (.B2(net2252),
    .C1(net4929),
    .B1(_11149_),
    .A1(net1582),
    .Y(_07259_),
    .A2(net5326));
 sg13g2_a21oi_1 _22805_ (.A1(net4785),
    .A2(_07258_),
    .Y(_07260_),
    .B1(_07259_));
 sg13g2_a21o_1 _22806_ (.A2(_07205_),
    .A1(net2252),
    .B1(_07260_),
    .X(_02382_));
 sg13g2_a21oi_1 _22807_ (.A1(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .A2(net6101),
    .Y(_07261_),
    .B1(net5047));
 sg13g2_nor2_1 _22808_ (.A(\soc_inst.cpu_core.ex_funct3[0] ),
    .B(net5072),
    .Y(_07262_));
 sg13g2_nor2_1 _22809_ (.A(\soc_inst.cpu_core.ex_branch_target[12] ),
    .B(net5158),
    .Y(_07263_));
 sg13g2_nor2_1 _22810_ (.A(\soc_inst.cpu_core.ex_alu_result[12] ),
    .B(net5165),
    .Y(_07264_));
 sg13g2_nor4_1 _22811_ (.A(_07261_),
    .B(_07262_),
    .C(_07263_),
    .D(_07264_),
    .Y(_07265_));
 sg13g2_a21oi_1 _22812_ (.A1(net2458),
    .A2(net4948),
    .Y(_07266_),
    .B1(_07265_));
 sg13g2_a221oi_1 _22813_ (.B2(net2458),
    .C1(net4929),
    .B1(_11153_),
    .A1(net1299),
    .Y(_07267_),
    .A2(net5326));
 sg13g2_a21oi_1 _22814_ (.A1(net4784),
    .A2(_07266_),
    .Y(_07268_),
    .B1(_07267_));
 sg13g2_a21o_1 _22815_ (.A2(_07205_),
    .A1(net2458),
    .B1(_07268_),
    .X(_02383_));
 sg13g2_a21oi_1 _22816_ (.A1(net1867),
    .A2(net6099),
    .Y(_07269_),
    .B1(net5046));
 sg13g2_nor2_1 _22817_ (.A(\soc_inst.cpu_core.ex_funct3[1] ),
    .B(net5071),
    .Y(_07270_));
 sg13g2_nor2_1 _22818_ (.A(net2446),
    .B(net5159),
    .Y(_07271_));
 sg13g2_nor2_1 _22819_ (.A(\soc_inst.cpu_core.ex_alu_result[13] ),
    .B(net5165),
    .Y(_07272_));
 sg13g2_nor4_1 _22820_ (.A(_07269_),
    .B(_07270_),
    .C(_07271_),
    .D(_07272_),
    .Y(_07273_));
 sg13g2_nor2_1 _22821_ (.A(net3252),
    .B(net1452),
    .Y(_07274_));
 sg13g2_a21oi_1 _22822_ (.A1(net1452),
    .A2(net5525),
    .Y(_07275_),
    .B1(_11157_));
 sg13g2_nor3_1 _22823_ (.A(net4928),
    .B(_07274_),
    .C(_07275_),
    .Y(_07276_));
 sg13g2_a221oi_1 _22824_ (.B2(net4928),
    .C1(_07276_),
    .B1(_07273_),
    .A1(net3252),
    .Y(_07277_),
    .A2(net4747));
 sg13g2_inv_1 _22825_ (.Y(_02384_),
    .A(net3253));
 sg13g2_a21o_1 _22826_ (.A2(net6102),
    .A1(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .B1(net5045),
    .X(_07278_));
 sg13g2_o21ai_1 _22827_ (.B1(_07278_),
    .Y(_07279_),
    .A1(\soc_inst.cpu_core.ex_alu_result[14] ),
    .A2(net5164));
 sg13g2_a221oi_1 _22828_ (.B2(_08121_),
    .C1(_07279_),
    .B1(net5160),
    .A1(_07869_),
    .Y(_07280_),
    .A2(net5074));
 sg13g2_nor2_1 _22829_ (.A(net3232),
    .B(net1378),
    .Y(_07281_));
 sg13g2_a21oi_1 _22830_ (.A1(net1378),
    .A2(net5525),
    .Y(_07282_),
    .B1(_11161_));
 sg13g2_nor3_1 _22831_ (.A(net4927),
    .B(_07281_),
    .C(_07282_),
    .Y(_07283_));
 sg13g2_a221oi_1 _22832_ (.B2(net4926),
    .C1(_07283_),
    .B1(_07280_),
    .A1(net3232),
    .Y(_07284_),
    .A2(net4748));
 sg13g2_inv_1 _22833_ (.Y(_02385_),
    .A(net3233));
 sg13g2_a21o_1 _22834_ (.A2(net6099),
    .A1(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .B1(net5045),
    .X(_07285_));
 sg13g2_o21ai_1 _22835_ (.B1(_07285_),
    .Y(_07286_),
    .A1(\soc_inst.cpu_core.ex_alu_result[15] ),
    .A2(net5164));
 sg13g2_a221oi_1 _22836_ (.B2(_08122_),
    .C1(_07286_),
    .B1(net5160),
    .A1(_08173_),
    .Y(_07287_),
    .A2(net5074));
 sg13g2_nor2_1 _22837_ (.A(net3238),
    .B(net2221),
    .Y(_07288_));
 sg13g2_a21oi_1 _22838_ (.A1(net2221),
    .A2(net5525),
    .Y(_07289_),
    .B1(_11165_));
 sg13g2_nor3_1 _22839_ (.A(net4925),
    .B(_07288_),
    .C(_07289_),
    .Y(_07290_));
 sg13g2_a221oi_1 _22840_ (.B2(net4927),
    .C1(_07290_),
    .B1(_07287_),
    .A1(net3238),
    .Y(_07291_),
    .A2(net4747));
 sg13g2_inv_1 _22841_ (.Y(_02386_),
    .A(net3239));
 sg13g2_a21oi_1 _22842_ (.A1(net2231),
    .A2(net6099),
    .Y(_07292_),
    .B1(net5045));
 sg13g2_nor2_1 _22843_ (.A(\soc_inst.cpu_core.ex_instr[16] ),
    .B(net5071),
    .Y(_07293_));
 sg13g2_nor2_1 _22844_ (.A(net2005),
    .B(net5159),
    .Y(_07294_));
 sg13g2_nor2_1 _22845_ (.A(net2299),
    .B(net5164),
    .Y(_07295_));
 sg13g2_nor4_1 _22846_ (.A(_07292_),
    .B(_07293_),
    .C(_07294_),
    .D(_07295_),
    .Y(_07296_));
 sg13g2_nor2_1 _22847_ (.A(net3224),
    .B(net1787),
    .Y(_07297_));
 sg13g2_a21oi_1 _22848_ (.A1(net1787),
    .A2(net5526),
    .Y(_07298_),
    .B1(_11169_));
 sg13g2_nor3_1 _22849_ (.A(net4926),
    .B(_07297_),
    .C(_07298_),
    .Y(_07299_));
 sg13g2_a221oi_1 _22850_ (.B2(net4927),
    .C1(_07299_),
    .B1(_07296_),
    .A1(net3224),
    .Y(_07300_),
    .A2(net4747));
 sg13g2_inv_1 _22851_ (.Y(_02387_),
    .A(_07300_));
 sg13g2_a21o_1 _22852_ (.A2(net6102),
    .A1(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .B1(net5045),
    .X(_07301_));
 sg13g2_o21ai_1 _22853_ (.B1(_07301_),
    .Y(_07302_),
    .A1(\soc_inst.cpu_core.ex_alu_result[17] ),
    .A2(net5164));
 sg13g2_a221oi_1 _22854_ (.B2(_08123_),
    .C1(_07302_),
    .B1(net5160),
    .A1(_08175_),
    .Y(_07303_),
    .A2(net5074));
 sg13g2_nor2_1 _22855_ (.A(net3268),
    .B(net1716),
    .Y(_07304_));
 sg13g2_a21oi_1 _22856_ (.A1(net1716),
    .A2(net5526),
    .Y(_07305_),
    .B1(_11173_));
 sg13g2_nor3_1 _22857_ (.A(net4926),
    .B(_07304_),
    .C(_07305_),
    .Y(_07306_));
 sg13g2_a221oi_1 _22858_ (.B2(net4926),
    .C1(_07306_),
    .B1(_07303_),
    .A1(net3268),
    .Y(_07307_),
    .A2(net4747));
 sg13g2_inv_1 _22859_ (.Y(_02388_),
    .A(net3269));
 sg13g2_nand2b_2 _22860_ (.Y(_07308_),
    .B(_08154_),
    .A_N(net5045));
 sg13g2_nor2_1 _22861_ (.A(\soc_inst.cpu_core.ex_branch_target[18] ),
    .B(net5159),
    .Y(_07309_));
 sg13g2_nor3_1 _22862_ (.A(\soc_inst.cpu_core.ex_instr[18] ),
    .B(net5073),
    .C(net5162),
    .Y(_07310_));
 sg13g2_nor2_1 _22863_ (.A(\soc_inst.cpu_core.ex_alu_result[18] ),
    .B(net5168),
    .Y(_07311_));
 sg13g2_nor4_1 _22864_ (.A(_09137_),
    .B(_07309_),
    .C(_07310_),
    .D(_07311_),
    .Y(_07312_));
 sg13g2_or2_1 _22865_ (.X(_07313_),
    .B(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A(net771));
 sg13g2_a21oi_1 _22866_ (.A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .A2(net5525),
    .Y(_07314_),
    .B1(_11177_));
 sg13g2_a221oi_1 _22867_ (.B2(_07312_),
    .C1(_09143_),
    .B1(_07308_),
    .A1(net771),
    .Y(_07315_),
    .A2(net4946));
 sg13g2_a221oi_1 _22868_ (.B2(_07313_),
    .C1(net4784),
    .B1(_11177_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .Y(_07316_),
    .A2(net5525));
 sg13g2_nand2_1 _22869_ (.Y(_07317_),
    .A(net771),
    .B(_07205_));
 sg13g2_o21ai_1 _22870_ (.B1(_07317_),
    .Y(_02389_),
    .A1(_07315_),
    .A2(_07316_));
 sg13g2_a21oi_1 _22871_ (.A1(net1764),
    .A2(net6102),
    .Y(_07318_),
    .B1(net5045));
 sg13g2_nor2_1 _22872_ (.A(\soc_inst.cpu_core.ex_instr[19] ),
    .B(net5073),
    .Y(_07319_));
 sg13g2_nor2_1 _22873_ (.A(\soc_inst.cpu_core.ex_alu_result[19] ),
    .B(net5164),
    .Y(_07320_));
 sg13g2_nor2_1 _22874_ (.A(net2441),
    .B(net5159),
    .Y(_07321_));
 sg13g2_nor4_1 _22875_ (.A(_07318_),
    .B(_07319_),
    .C(_07320_),
    .D(_07321_),
    .Y(_07322_));
 sg13g2_nor2_1 _22876_ (.A(net3300),
    .B(net1772),
    .Y(_07323_));
 sg13g2_a21oi_1 _22877_ (.A1(net1772),
    .A2(net5526),
    .Y(_07324_),
    .B1(_11181_));
 sg13g2_nor3_1 _22878_ (.A(net4926),
    .B(_07323_),
    .C(_07324_),
    .Y(_07325_));
 sg13g2_a221oi_1 _22879_ (.B2(net4926),
    .C1(_07325_),
    .B1(_07322_),
    .A1(net3300),
    .Y(_07326_),
    .A2(net4747));
 sg13g2_inv_1 _22880_ (.Y(_02390_),
    .A(net3301));
 sg13g2_a21o_1 _22881_ (.A2(net6099),
    .A1(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .B1(net5046),
    .X(_07327_));
 sg13g2_o21ai_1 _22882_ (.B1(_07327_),
    .Y(_07328_),
    .A1(\soc_inst.cpu_core.ex_alu_result[20] ),
    .A2(net5165));
 sg13g2_a221oi_1 _22883_ (.B2(_08126_),
    .C1(_07328_),
    .B1(net5160),
    .A1(_08176_),
    .Y(_07329_),
    .A2(net5074));
 sg13g2_nor2_1 _22884_ (.A(net3278),
    .B(net2260),
    .Y(_07330_));
 sg13g2_a21oi_1 _22885_ (.A1(net2260),
    .A2(net5526),
    .Y(_07331_),
    .B1(_11185_));
 sg13g2_nor3_1 _22886_ (.A(net4927),
    .B(_07330_),
    .C(_07331_),
    .Y(_07332_));
 sg13g2_a221oi_1 _22887_ (.B2(net4926),
    .C1(_07332_),
    .B1(_07329_),
    .A1(net3278),
    .Y(_07333_),
    .A2(net4747));
 sg13g2_inv_1 _22888_ (.Y(_02391_),
    .A(_07333_));
 sg13g2_a21oi_1 _22889_ (.A1(net1801),
    .A2(net6099),
    .Y(_07334_),
    .B1(net5046));
 sg13g2_nor2_1 _22890_ (.A(net2487),
    .B(net5073),
    .Y(_07335_));
 sg13g2_nor2_1 _22891_ (.A(net2754),
    .B(net5159),
    .Y(_07336_));
 sg13g2_nor2_1 _22892_ (.A(net2879),
    .B(net5164),
    .Y(_07337_));
 sg13g2_nor4_1 _22893_ (.A(_07334_),
    .B(_07335_),
    .C(_07336_),
    .D(_07337_),
    .Y(_07338_));
 sg13g2_nor2_1 _22894_ (.A(net3223),
    .B(net2445),
    .Y(_07339_));
 sg13g2_a21oi_1 _22895_ (.A1(net2445),
    .A2(net5525),
    .Y(_07340_),
    .B1(_11189_));
 sg13g2_nor3_1 _22896_ (.A(net4925),
    .B(_07339_),
    .C(_07340_),
    .Y(_07341_));
 sg13g2_a221oi_1 _22897_ (.B2(net4925),
    .C1(_07341_),
    .B1(_07338_),
    .A1(net3223),
    .Y(_07342_),
    .A2(net4747));
 sg13g2_inv_1 _22898_ (.Y(_02392_),
    .A(_07342_));
 sg13g2_a21o_1 _22899_ (.A2(net6099),
    .A1(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .B1(net5045),
    .X(_07343_));
 sg13g2_o21ai_1 _22900_ (.B1(_07343_),
    .Y(_07344_),
    .A1(\soc_inst.cpu_core.ex_alu_result[22] ),
    .A2(net5164));
 sg13g2_a221oi_1 _22901_ (.B2(_08128_),
    .C1(_07344_),
    .B1(net5160),
    .A1(_08177_),
    .Y(_07345_),
    .A2(net5074));
 sg13g2_nor2_1 _22902_ (.A(net3117),
    .B(net2337),
    .Y(_07346_));
 sg13g2_a21oi_1 _22903_ (.A1(net2337),
    .A2(net5525),
    .Y(_07347_),
    .B1(_11193_));
 sg13g2_nor3_1 _22904_ (.A(net4925),
    .B(_07346_),
    .C(_07347_),
    .Y(_07348_));
 sg13g2_a221oi_1 _22905_ (.B2(net4925),
    .C1(_07348_),
    .B1(_07345_),
    .A1(net3117),
    .Y(_07349_),
    .A2(net4746));
 sg13g2_inv_1 _22906_ (.Y(_02393_),
    .A(_07349_));
 sg13g2_a21oi_1 _22907_ (.A1(net1668),
    .A2(net6099),
    .Y(_07350_),
    .B1(net5045));
 sg13g2_nor2_1 _22908_ (.A(net2715),
    .B(net5073),
    .Y(_07351_));
 sg13g2_nor2_1 _22909_ (.A(net2238),
    .B(net5159),
    .Y(_07352_));
 sg13g2_nor2_1 _22910_ (.A(net2964),
    .B(net5164),
    .Y(_07353_));
 sg13g2_nor4_1 _22911_ (.A(_07350_),
    .B(_07351_),
    .C(_07352_),
    .D(_07353_),
    .Y(_07354_));
 sg13g2_nor2_1 _22912_ (.A(net3167),
    .B(net2599),
    .Y(_07355_));
 sg13g2_a21oi_1 _22913_ (.A1(net2599),
    .A2(net5525),
    .Y(_07356_),
    .B1(_11197_));
 sg13g2_nor3_1 _22914_ (.A(net4925),
    .B(_07355_),
    .C(_07356_),
    .Y(_07357_));
 sg13g2_a221oi_1 _22915_ (.B2(net4926),
    .C1(_07357_),
    .B1(_07354_),
    .A1(net3167),
    .Y(_07358_),
    .A2(net4747));
 sg13g2_inv_1 _22916_ (.Y(_02394_),
    .A(net3168));
 sg13g2_a221oi_1 _22917_ (.B2(\soc_inst.cpu_core.ex_instr[24] ),
    .C1(net5163),
    .B1(net5076),
    .A1(\soc_inst.cpu_core.ex_alu_result[24] ),
    .Y(_07359_),
    .A2(_08950_));
 sg13g2_a21oi_2 _22918_ (.B1(_07359_),
    .Y(_07360_),
    .A2(net5162),
    .A1(_08178_));
 sg13g2_o21ai_1 _22919_ (.B1(net3193),
    .Y(_07361_),
    .A1(net6025),
    .A2(_11202_));
 sg13g2_nand2_1 _22920_ (.Y(_07362_),
    .A(net5531),
    .B(_11200_));
 sg13g2_a21oi_1 _22921_ (.A1(_07361_),
    .A2(_07362_),
    .Y(_07363_),
    .B1(net4925));
 sg13g2_a221oi_1 _22922_ (.B2(net4925),
    .C1(_07363_),
    .B1(_07360_),
    .A1(net3193),
    .Y(_07364_),
    .A2(net4746));
 sg13g2_inv_1 _22923_ (.Y(_02395_),
    .A(net3194));
 sg13g2_a22oi_1 _22924_ (.Y(_07365_),
    .B1(net5161),
    .B2(net2681),
    .A2(net5169),
    .A1(\soc_inst.cpu_core.ex_alu_result[25] ));
 sg13g2_o21ai_1 _22925_ (.B1(_07365_),
    .Y(_07366_),
    .A1(_08179_),
    .A2(net5073));
 sg13g2_nand2_1 _22926_ (.Y(_07367_),
    .A(net4928),
    .B(_07366_));
 sg13g2_nand3_1 _22927_ (.B(net5145),
    .C(_11207_),
    .A(net3107),
    .Y(_07368_));
 sg13g2_a21oi_1 _22928_ (.A1(net3107),
    .A2(net6026),
    .Y(_07369_),
    .B1(_11205_));
 sg13g2_nand2_2 _22929_ (.Y(_07370_),
    .A(net5145),
    .B(net5326));
 sg13g2_o21ai_1 _22930_ (.B1(_07368_),
    .Y(_07371_),
    .A1(_07369_),
    .A2(_07370_));
 sg13g2_a22oi_1 _22931_ (.Y(_07372_),
    .B1(_07371_),
    .B2(_09037_),
    .A2(net4749),
    .A1(net3107));
 sg13g2_nand2_1 _22932_ (.Y(_02396_),
    .A(_07367_),
    .B(_07372_));
 sg13g2_nand2_1 _22933_ (.Y(_07373_),
    .A(\soc_inst.cpu_core.ex_alu_result[26] ),
    .B(net5169));
 sg13g2_a22oi_1 _22934_ (.Y(_07374_),
    .B1(net5160),
    .B2(\soc_inst.cpu_core.ex_branch_target[26] ),
    .A2(net5074),
    .A1(\soc_inst.cpu_core.ex_funct7[1] ));
 sg13g2_a21oi_2 _22935_ (.B1(_09143_),
    .Y(_07375_),
    .A2(_07374_),
    .A1(_07373_));
 sg13g2_nand3_1 _22936_ (.B(net5142),
    .C(_11212_),
    .A(net3198),
    .Y(_07376_));
 sg13g2_a21oi_1 _22937_ (.A1(net3198),
    .A2(net6026),
    .Y(_07377_),
    .B1(_11210_));
 sg13g2_o21ai_1 _22938_ (.B1(_07376_),
    .Y(_07378_),
    .A1(_07370_),
    .A2(_07377_));
 sg13g2_a221oi_1 _22939_ (.B2(net4936),
    .C1(_07375_),
    .B1(_07378_),
    .A1(net3198),
    .Y(_07379_),
    .A2(net4746));
 sg13g2_inv_1 _22940_ (.Y(_02397_),
    .A(net3199));
 sg13g2_nand2_1 _22941_ (.Y(_07380_),
    .A(\soc_inst.cpu_core.ex_alu_result[27] ),
    .B(net5169));
 sg13g2_a22oi_1 _22942_ (.Y(_07381_),
    .B1(net5160),
    .B2(\soc_inst.cpu_core.ex_branch_target[27] ),
    .A2(net5075),
    .A1(\soc_inst.cpu_core.ex_funct7[2] ));
 sg13g2_a21oi_1 _22943_ (.A1(_07380_),
    .A2(_07381_),
    .Y(_07382_),
    .B1(_09143_));
 sg13g2_nand3_1 _22944_ (.B(net5145),
    .C(_11217_),
    .A(net3227),
    .Y(_07383_));
 sg13g2_a21oi_1 _22945_ (.A1(net3227),
    .A2(net6026),
    .Y(_07384_),
    .B1(_11215_));
 sg13g2_o21ai_1 _22946_ (.B1(_07383_),
    .Y(_07385_),
    .A1(_07370_),
    .A2(_07384_));
 sg13g2_a221oi_1 _22947_ (.B2(net4936),
    .C1(_07382_),
    .B1(_07385_),
    .A1(net3227),
    .Y(_07386_),
    .A2(net4746));
 sg13g2_inv_1 _22948_ (.Y(_02398_),
    .A(net3228));
 sg13g2_nand2_1 _22949_ (.Y(_07387_),
    .A(net2993),
    .B(net5169));
 sg13g2_a22oi_1 _22950_ (.Y(_07388_),
    .B1(net5162),
    .B2(\soc_inst.cpu_core.ex_branch_target[28] ),
    .A2(net5075),
    .A1(\soc_inst.cpu_core.ex_funct7[3] ));
 sg13g2_a21oi_2 _22951_ (.B1(_09143_),
    .Y(_07389_),
    .A2(_07388_),
    .A1(_07387_));
 sg13g2_nand3_1 _22952_ (.B(net5144),
    .C(_11222_),
    .A(net3118),
    .Y(_07390_));
 sg13g2_a21oi_1 _22953_ (.A1(net3118),
    .A2(net6026),
    .Y(_07391_),
    .B1(_11220_));
 sg13g2_o21ai_1 _22954_ (.B1(_07390_),
    .Y(_07392_),
    .A1(_07370_),
    .A2(_07391_));
 sg13g2_a221oi_1 _22955_ (.B2(net4936),
    .C1(_07389_),
    .B1(_07392_),
    .A1(net3118),
    .Y(_07393_),
    .A2(net4746));
 sg13g2_inv_1 _22956_ (.Y(_02399_),
    .A(_07393_));
 sg13g2_nand2_1 _22957_ (.Y(_07394_),
    .A(net3095),
    .B(net5169));
 sg13g2_a22oi_1 _22958_ (.Y(_07395_),
    .B1(net5160),
    .B2(\soc_inst.cpu_core.ex_branch_target[29] ),
    .A2(net5074),
    .A1(\soc_inst.cpu_core.ex_funct7[4] ));
 sg13g2_a21oi_2 _22959_ (.B1(_09143_),
    .Y(_07396_),
    .A2(_07395_),
    .A1(_07394_));
 sg13g2_nand3_1 _22960_ (.B(net5143),
    .C(_11227_),
    .A(net3153),
    .Y(_07397_));
 sg13g2_a21oi_1 _22961_ (.A1(net3153),
    .A2(net6026),
    .Y(_07398_),
    .B1(_11225_));
 sg13g2_o21ai_1 _22962_ (.B1(_07397_),
    .Y(_07399_),
    .A1(_07370_),
    .A2(_07398_));
 sg13g2_a221oi_1 _22963_ (.B2(net4936),
    .C1(_07396_),
    .B1(_07399_),
    .A1(net3153),
    .Y(_07400_),
    .A2(net4746));
 sg13g2_inv_1 _22964_ (.Y(_02400_),
    .A(net3154));
 sg13g2_nand2_1 _22965_ (.Y(_07401_),
    .A(\soc_inst.cpu_core.ex_alu_result[30] ),
    .B(net5169));
 sg13g2_a22oi_1 _22966_ (.Y(_07402_),
    .B1(net5161),
    .B2(\soc_inst.cpu_core.ex_branch_target[30] ),
    .A2(net5074),
    .A1(\soc_inst.cpu_core.ex_funct7[5] ));
 sg13g2_a21oi_2 _22967_ (.B1(_09143_),
    .Y(_07403_),
    .A2(_07402_),
    .A1(_07401_));
 sg13g2_nand3_1 _22968_ (.B(net5144),
    .C(_11232_),
    .A(net3108),
    .Y(_07404_));
 sg13g2_a21oi_1 _22969_ (.A1(net3108),
    .A2(net6026),
    .Y(_07405_),
    .B1(_11230_));
 sg13g2_o21ai_1 _22970_ (.B1(_07404_),
    .Y(_07406_),
    .A1(_07370_),
    .A2(_07405_));
 sg13g2_a221oi_1 _22971_ (.B2(net4936),
    .C1(_07403_),
    .B1(_07406_),
    .A1(net3108),
    .Y(_07407_),
    .A2(net4746));
 sg13g2_inv_1 _22972_ (.Y(_02401_),
    .A(net3109));
 sg13g2_a22oi_1 _22973_ (.Y(_07408_),
    .B1(net5161),
    .B2(\soc_inst.cpu_core.ex_branch_target[31] ),
    .A2(net5075),
    .A1(\soc_inst.cpu_core.ex_funct7[6] ));
 sg13g2_o21ai_1 _22974_ (.B1(_07408_),
    .Y(_07409_),
    .A1(_08184_),
    .A2(net5168));
 sg13g2_or2_1 _22975_ (.X(_07410_),
    .B(net1398),
    .A(net3067));
 sg13g2_a22oi_1 _22976_ (.Y(_07411_),
    .B1(_11235_),
    .B2(_07410_),
    .A2(net5527),
    .A1(net1398));
 sg13g2_a22oi_1 _22977_ (.Y(_07412_),
    .B1(_07409_),
    .B2(net4784),
    .A2(net4746),
    .A1(net3067));
 sg13g2_o21ai_1 _22978_ (.B1(_07412_),
    .Y(_02402_),
    .A1(net4784),
    .A2(_07411_));
 sg13g2_a21oi_1 _22979_ (.A1(_09898_),
    .A2(net4759),
    .Y(_07413_),
    .B1(net776));
 sg13g2_nor2_1 _22980_ (.A(_09513_),
    .B(_09923_),
    .Y(_07414_));
 sg13g2_a21oi_1 _22981_ (.A1(_11132_),
    .A2(net4744),
    .Y(_02403_),
    .B1(net777));
 sg13g2_a21oi_1 _22982_ (.A1(_09903_),
    .A2(net4758),
    .Y(_07415_),
    .B1(net715));
 sg13g2_a21oi_1 _22983_ (.A1(_11136_),
    .A2(net4744),
    .Y(_02404_),
    .B1(net716));
 sg13g2_a21oi_1 _22984_ (.A1(net4758),
    .A2(_11137_),
    .Y(_07416_),
    .B1(net1193));
 sg13g2_a21oi_1 _22985_ (.A1(_11140_),
    .A2(net4744),
    .Y(_02405_),
    .B1(net1194));
 sg13g2_a21oi_1 _22986_ (.A1(_09907_),
    .A2(net4759),
    .Y(_07417_),
    .B1(net500));
 sg13g2_a21oi_1 _22987_ (.A1(_11142_),
    .A2(net4745),
    .Y(_02406_),
    .B1(net501));
 sg13g2_a21oi_1 _22988_ (.A1(_09911_),
    .A2(net4759),
    .Y(_07418_),
    .B1(net1068));
 sg13g2_a21oi_1 _22989_ (.A1(_11144_),
    .A2(net4745),
    .Y(_02407_),
    .B1(net1069));
 sg13g2_a21oi_1 _22990_ (.A1(_09915_),
    .A2(net4759),
    .Y(_07419_),
    .B1(net1056));
 sg13g2_a21oi_1 _22991_ (.A1(_11146_),
    .A2(net4745),
    .Y(_02408_),
    .B1(net1057));
 sg13g2_a21oi_1 _22992_ (.A1(net4758),
    .A2(_11147_),
    .Y(_07420_),
    .B1(net535));
 sg13g2_a21oi_1 _22993_ (.A1(_11150_),
    .A2(net4745),
    .Y(_02409_),
    .B1(net536));
 sg13g2_a21oi_1 _22994_ (.A1(net4755),
    .A2(_11151_),
    .Y(_07421_),
    .B1(net693));
 sg13g2_a21oi_1 _22995_ (.A1(_11154_),
    .A2(net4744),
    .Y(_02410_),
    .B1(net694));
 sg13g2_a21oi_1 _22996_ (.A1(net4755),
    .A2(_11155_),
    .Y(_07422_),
    .B1(net708));
 sg13g2_a21oi_1 _22997_ (.A1(_11158_),
    .A2(net4743),
    .Y(_02411_),
    .B1(net709));
 sg13g2_a21oi_1 _22998_ (.A1(net4756),
    .A2(_11159_),
    .Y(_07423_),
    .B1(net516));
 sg13g2_a21oi_1 _22999_ (.A1(_11162_),
    .A2(net4744),
    .Y(_02412_),
    .B1(net517));
 sg13g2_a21oi_1 _23000_ (.A1(net4755),
    .A2(_11163_),
    .Y(_07424_),
    .B1(net503));
 sg13g2_a21oi_1 _23001_ (.A1(_11166_),
    .A2(net4743),
    .Y(_02413_),
    .B1(net504));
 sg13g2_a21oi_1 _23002_ (.A1(net4755),
    .A2(_11167_),
    .Y(_07425_),
    .B1(net1143));
 sg13g2_a21oi_1 _23003_ (.A1(_11170_),
    .A2(net4743),
    .Y(_02414_),
    .B1(net1144));
 sg13g2_a21oi_1 _23004_ (.A1(net4756),
    .A2(_11171_),
    .Y(_07426_),
    .B1(net1024));
 sg13g2_a21oi_1 _23005_ (.A1(_11174_),
    .A2(net4744),
    .Y(_02415_),
    .B1(net1025));
 sg13g2_a21oi_1 _23006_ (.A1(net4756),
    .A2(_11175_),
    .Y(_07427_),
    .B1(net464));
 sg13g2_a21oi_1 _23007_ (.A1(_11178_),
    .A2(net4744),
    .Y(_02416_),
    .B1(net465));
 sg13g2_a21oi_1 _23008_ (.A1(net4756),
    .A2(_11179_),
    .Y(_07428_),
    .B1(net611));
 sg13g2_a21oi_1 _23009_ (.A1(_11182_),
    .A2(net4743),
    .Y(_02417_),
    .B1(net612));
 sg13g2_a21oi_1 _23010_ (.A1(net4755),
    .A2(_11183_),
    .Y(_07429_),
    .B1(net344));
 sg13g2_a21oi_1 _23011_ (.A1(_11186_),
    .A2(net4743),
    .Y(_02418_),
    .B1(net345));
 sg13g2_a21oi_1 _23012_ (.A1(net4755),
    .A2(_11187_),
    .Y(_07430_),
    .B1(net842));
 sg13g2_a21oi_1 _23013_ (.A1(_11190_),
    .A2(net4743),
    .Y(_02419_),
    .B1(net843));
 sg13g2_a21oi_1 _23014_ (.A1(net4755),
    .A2(_11191_),
    .Y(_07431_),
    .B1(net1181));
 sg13g2_a21oi_1 _23015_ (.A1(_11194_),
    .A2(net4743),
    .Y(_02420_),
    .B1(net1182));
 sg13g2_a21oi_1 _23016_ (.A1(net4755),
    .A2(_11195_),
    .Y(_07432_),
    .B1(net948));
 sg13g2_a21oi_1 _23017_ (.A1(_11198_),
    .A2(net4743),
    .Y(_02421_),
    .B1(net949));
 sg13g2_nor2_2 _23018_ (.A(_09058_),
    .B(_07204_),
    .Y(_07433_));
 sg13g2_o21ai_1 _23019_ (.B1(_09061_),
    .Y(_07434_),
    .A1(_09058_),
    .A2(_07202_));
 sg13g2_nor3_1 _23020_ (.A(_07871_),
    .B(_08089_),
    .C(net4999),
    .Y(_07435_));
 sg13g2_a21oi_1 _23021_ (.A1(net1268),
    .A2(net4999),
    .Y(_07436_),
    .B1(_07435_));
 sg13g2_a221oi_1 _23022_ (.B2(net1664),
    .C1(net4790),
    .B1(net5326),
    .A1(net2256),
    .Y(_07437_),
    .A2(_09895_));
 sg13g2_a21oi_1 _23023_ (.A1(net4790),
    .A2(_07436_),
    .Y(_07438_),
    .B1(_07437_));
 sg13g2_a21o_1 _23024_ (.A2(net4718),
    .A1(net2256),
    .B1(_07438_),
    .X(_02422_));
 sg13g2_nand3_1 _23025_ (.B(_08091_),
    .C(net5002),
    .A(net6480),
    .Y(_07439_));
 sg13g2_o21ai_1 _23026_ (.B1(_07439_),
    .Y(_07440_),
    .A1(net1384),
    .A2(net5002));
 sg13g2_nor2_1 _23027_ (.A(_09059_),
    .B(_07440_),
    .Y(_07441_));
 sg13g2_nand2_1 _23028_ (.Y(_07442_),
    .A(net1420),
    .B(_09901_));
 sg13g2_a21oi_1 _23029_ (.A1(_09904_),
    .A2(_07442_),
    .Y(_07443_),
    .B1(net4789));
 sg13g2_nor3_1 _23030_ (.A(net4742),
    .B(_07441_),
    .C(_07443_),
    .Y(_07444_));
 sg13g2_a21oi_1 _23031_ (.A1(_08004_),
    .A2(net4718),
    .Y(_02423_),
    .B1(_07444_));
 sg13g2_nand3_1 _23032_ (.B(_08093_),
    .C(net5007),
    .A(net6480),
    .Y(_07445_));
 sg13g2_o21ai_1 _23033_ (.B1(_07445_),
    .Y(_07446_),
    .A1(net1697),
    .A2(net5007));
 sg13g2_nor2_1 _23034_ (.A(net4761),
    .B(_07446_),
    .Y(_07447_));
 sg13g2_nor3_1 _23035_ (.A(_08005_),
    .B(net2390),
    .C(net6019),
    .Y(_07448_));
 sg13g2_nor2_1 _23036_ (.A(net5326),
    .B(_07448_),
    .Y(_07449_));
 sg13g2_a21oi_1 _23037_ (.A1(net2706),
    .A2(_11139_),
    .Y(_07450_),
    .B1(_11137_));
 sg13g2_nor3_1 _23038_ (.A(net4789),
    .B(_07449_),
    .C(_07450_),
    .Y(_07451_));
 sg13g2_nor3_1 _23039_ (.A(net4742),
    .B(_07447_),
    .C(_07451_),
    .Y(_07452_));
 sg13g2_a21oi_1 _23040_ (.A1(_08005_),
    .A2(net4718),
    .Y(_02424_),
    .B1(_07452_));
 sg13g2_nand3_1 _23041_ (.B(_08095_),
    .C(net5007),
    .A(net6480),
    .Y(_07453_));
 sg13g2_o21ai_1 _23042_ (.B1(_07453_),
    .Y(_07454_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .A2(net5006));
 sg13g2_nor2_1 _23043_ (.A(_09059_),
    .B(_07454_),
    .Y(_07455_));
 sg13g2_nand2_1 _23044_ (.Y(_07456_),
    .A(net1261),
    .B(_09905_));
 sg13g2_a21oi_1 _23045_ (.A1(_09908_),
    .A2(_07456_),
    .Y(_07457_),
    .B1(net4790));
 sg13g2_nor3_1 _23046_ (.A(net4742),
    .B(_07455_),
    .C(_07457_),
    .Y(_07458_));
 sg13g2_a21oi_1 _23047_ (.A1(_08006_),
    .A2(net4718),
    .Y(_02425_),
    .B1(_07458_));
 sg13g2_nand3_1 _23048_ (.B(_08097_),
    .C(net5002),
    .A(net6480),
    .Y(_07459_));
 sg13g2_o21ai_1 _23049_ (.B1(_07459_),
    .Y(_07460_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .A2(net5002));
 sg13g2_nor2_1 _23050_ (.A(net4761),
    .B(_07460_),
    .Y(_07461_));
 sg13g2_nand2_1 _23051_ (.Y(_07462_),
    .A(net1292),
    .B(_09909_));
 sg13g2_a21oi_1 _23052_ (.A1(_09912_),
    .A2(_07462_),
    .Y(_07463_),
    .B1(net4790));
 sg13g2_nor3_1 _23053_ (.A(net4742),
    .B(_07461_),
    .C(_07463_),
    .Y(_07464_));
 sg13g2_a21oi_1 _23054_ (.A1(_08007_),
    .A2(_07434_),
    .Y(_02426_),
    .B1(_07464_));
 sg13g2_nand3_1 _23055_ (.B(_08099_),
    .C(net5006),
    .A(net6481),
    .Y(_07465_));
 sg13g2_o21ai_1 _23056_ (.B1(_07465_),
    .Y(_07466_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .A2(net5006));
 sg13g2_nor2_1 _23057_ (.A(net4761),
    .B(_07466_),
    .Y(_07467_));
 sg13g2_nand2_1 _23058_ (.Y(_07468_),
    .A(net1216),
    .B(_09913_));
 sg13g2_a21oi_1 _23059_ (.A1(_09916_),
    .A2(_07468_),
    .Y(_07469_),
    .B1(net4790));
 sg13g2_nor3_1 _23060_ (.A(_07433_),
    .B(_07467_),
    .C(_07469_),
    .Y(_07470_));
 sg13g2_a21oi_1 _23061_ (.A1(_08008_),
    .A2(_07434_),
    .Y(_02427_),
    .B1(_07470_));
 sg13g2_a21oi_1 _23062_ (.A1(net6480),
    .A2(_08101_),
    .Y(_07471_),
    .B1(net5000));
 sg13g2_a21oi_1 _23063_ (.A1(net2292),
    .A2(net5000),
    .Y(_07472_),
    .B1(_07471_));
 sg13g2_a21oi_1 _23064_ (.A1(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .A2(net5527),
    .Y(_07473_),
    .B1(_11149_));
 sg13g2_nor2_1 _23065_ (.A(net3225),
    .B(net1582),
    .Y(_07474_));
 sg13g2_o21ai_1 _23066_ (.B1(net4761),
    .Y(_07475_),
    .A1(_07473_),
    .A2(_07474_));
 sg13g2_nor2_1 _23067_ (.A(net3225),
    .B(net4942),
    .Y(_07476_));
 sg13g2_o21ai_1 _23068_ (.B1(net4790),
    .Y(_07477_),
    .A1(_07472_),
    .A2(_07476_));
 sg13g2_and2_1 _23069_ (.A(net3225),
    .B(_07433_),
    .X(_07478_));
 sg13g2_a21o_1 _23070_ (.A2(_07477_),
    .A1(_07475_),
    .B1(_07478_),
    .X(_02428_));
 sg13g2_nand3_1 _23071_ (.B(_08103_),
    .C(net5006),
    .A(net6481),
    .Y(_07479_));
 sg13g2_o21ai_1 _23072_ (.B1(_07479_),
    .Y(_07480_),
    .A1(net1453),
    .A2(net5006));
 sg13g2_nor2_1 _23073_ (.A(net4761),
    .B(_07480_),
    .Y(_07481_));
 sg13g2_a21oi_1 _23074_ (.A1(net1299),
    .A2(net5527),
    .Y(_07482_),
    .B1(_11153_));
 sg13g2_nor2_1 _23075_ (.A(net2077),
    .B(net1299),
    .Y(_07483_));
 sg13g2_nor3_1 _23076_ (.A(net4788),
    .B(_07482_),
    .C(_07483_),
    .Y(_07484_));
 sg13g2_nor3_1 _23077_ (.A(_07433_),
    .B(_07481_),
    .C(_07484_),
    .Y(_07485_));
 sg13g2_a21oi_1 _23078_ (.A1(_08009_),
    .A2(_07434_),
    .Y(_02429_),
    .B1(_07485_));
 sg13g2_nand3_1 _23079_ (.B(_08105_),
    .C(net5002),
    .A(net6479),
    .Y(_07486_));
 sg13g2_o21ai_1 _23080_ (.B1(_07486_),
    .Y(_07487_),
    .A1(net1867),
    .A2(net5002));
 sg13g2_nand2b_1 _23081_ (.Y(_07488_),
    .B(net4791),
    .A_N(_07487_));
 sg13g2_a21oi_1 _23082_ (.A1(net5531),
    .A2(_11155_),
    .Y(_07489_),
    .B1(net2346));
 sg13g2_nor3_1 _23083_ (.A(net4788),
    .B(_07275_),
    .C(_07489_),
    .Y(_07490_));
 sg13g2_nor2_1 _23084_ (.A(net4741),
    .B(_07490_),
    .Y(_07491_));
 sg13g2_a22oi_1 _23085_ (.Y(_02430_),
    .B1(_07488_),
    .B2(_07491_),
    .A2(net4718),
    .A1(_08011_));
 sg13g2_nand3_1 _23086_ (.B(_08106_),
    .C(net5005),
    .A(net6478),
    .Y(_07492_));
 sg13g2_o21ai_1 _23087_ (.B1(_07492_),
    .Y(_07493_),
    .A1(net1382),
    .A2(net5004));
 sg13g2_nand2b_1 _23088_ (.Y(_07494_),
    .B(net4786),
    .A_N(_07493_));
 sg13g2_a21oi_1 _23089_ (.A1(net5532),
    .A2(_11159_),
    .Y(_07495_),
    .B1(net2510));
 sg13g2_nor3_1 _23090_ (.A(net4788),
    .B(_07282_),
    .C(_07495_),
    .Y(_07496_));
 sg13g2_nor2_1 _23091_ (.A(net4741),
    .B(_07496_),
    .Y(_07497_));
 sg13g2_a22oi_1 _23092_ (.Y(_02431_),
    .B1(_07494_),
    .B2(_07497_),
    .A2(net4718),
    .A1(_08013_));
 sg13g2_nand3_1 _23093_ (.B(_08107_),
    .C(net5003),
    .A(net6478),
    .Y(_07498_));
 sg13g2_o21ai_1 _23094_ (.B1(_07498_),
    .Y(_07499_),
    .A1(net1822),
    .A2(net5001));
 sg13g2_nand2b_1 _23095_ (.Y(_07500_),
    .B(net4787),
    .A_N(_07499_));
 sg13g2_a21oi_1 _23096_ (.A1(net5531),
    .A2(_11163_),
    .Y(_07501_),
    .B1(net2449));
 sg13g2_nor3_1 _23097_ (.A(net4788),
    .B(_07289_),
    .C(_07501_),
    .Y(_07502_));
 sg13g2_nor2_1 _23098_ (.A(net4741),
    .B(_07502_),
    .Y(_07503_));
 sg13g2_a22oi_1 _23099_ (.Y(_02432_),
    .B1(_07500_),
    .B2(_07503_),
    .A2(net4717),
    .A1(_08015_));
 sg13g2_nand3_1 _23100_ (.B(_08108_),
    .C(net5003),
    .A(net6478),
    .Y(_07504_));
 sg13g2_o21ai_1 _23101_ (.B1(_07504_),
    .Y(_07505_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .A2(net5004));
 sg13g2_nand2b_1 _23102_ (.Y(_07506_),
    .B(net4786),
    .A_N(_07505_));
 sg13g2_a21oi_1 _23103_ (.A1(net5531),
    .A2(_11167_),
    .Y(_07507_),
    .B1(net2114));
 sg13g2_nor3_1 _23104_ (.A(net4786),
    .B(_07298_),
    .C(_07507_),
    .Y(_07508_));
 sg13g2_nor2_1 _23105_ (.A(net4741),
    .B(_07508_),
    .Y(_07509_));
 sg13g2_a22oi_1 _23106_ (.Y(_02433_),
    .B1(_07506_),
    .B2(_07509_),
    .A2(net4717),
    .A1(_08016_));
 sg13g2_nand3_1 _23107_ (.B(_08109_),
    .C(net5005),
    .A(net6478),
    .Y(_07510_));
 sg13g2_o21ai_1 _23108_ (.B1(_07510_),
    .Y(_07511_),
    .A1(net1778),
    .A2(net5004));
 sg13g2_nand2b_1 _23109_ (.Y(_07512_),
    .B(net4786),
    .A_N(_07511_));
 sg13g2_a21oi_1 _23110_ (.A1(net5532),
    .A2(_11171_),
    .Y(_07513_),
    .B1(net1966));
 sg13g2_nor3_1 _23111_ (.A(net4787),
    .B(_07305_),
    .C(_07513_),
    .Y(_07514_));
 sg13g2_nor2_1 _23112_ (.A(net4742),
    .B(_07514_),
    .Y(_07515_));
 sg13g2_a22oi_1 _23113_ (.Y(_02434_),
    .B1(_07512_),
    .B2(_07515_),
    .A2(net4717),
    .A1(_08017_));
 sg13g2_nand3_1 _23114_ (.B(_08110_),
    .C(net5003),
    .A(net6479),
    .Y(_07516_));
 sg13g2_o21ai_1 _23115_ (.B1(_07516_),
    .Y(_07517_),
    .A1(\soc_inst.cpu_core.ex_exception_pc[18] ),
    .A2(net5003));
 sg13g2_nor2_1 _23116_ (.A(net4761),
    .B(_07517_),
    .Y(_07518_));
 sg13g2_a21oi_1 _23117_ (.A1(net5532),
    .A2(_11175_),
    .Y(_07519_),
    .B1(net2534));
 sg13g2_nor3_1 _23118_ (.A(net4788),
    .B(_07314_),
    .C(_07519_),
    .Y(_07520_));
 sg13g2_nor3_1 _23119_ (.A(net4741),
    .B(_07518_),
    .C(_07520_),
    .Y(_07521_));
 sg13g2_a21oi_1 _23120_ (.A1(_08018_),
    .A2(net4717),
    .Y(_02435_),
    .B1(_07521_));
 sg13g2_nand3_1 _23121_ (.B(_08111_),
    .C(net5003),
    .A(net6478),
    .Y(_07522_));
 sg13g2_o21ai_1 _23122_ (.B1(_07522_),
    .Y(_07523_),
    .A1(net1764),
    .A2(net5003));
 sg13g2_nand2b_1 _23123_ (.Y(_07524_),
    .B(net4786),
    .A_N(_07523_));
 sg13g2_a21oi_1 _23124_ (.A1(net5531),
    .A2(_11179_),
    .Y(_07525_),
    .B1(net2796));
 sg13g2_nor3_1 _23125_ (.A(net4786),
    .B(_07324_),
    .C(_07525_),
    .Y(_07526_));
 sg13g2_nor2_1 _23126_ (.A(net4742),
    .B(_07526_),
    .Y(_07527_));
 sg13g2_a22oi_1 _23127_ (.Y(_02436_),
    .B1(_07524_),
    .B2(_07527_),
    .A2(net4717),
    .A1(_08019_));
 sg13g2_nand3_1 _23128_ (.B(_08112_),
    .C(net5003),
    .A(net6478),
    .Y(_07528_));
 sg13g2_o21ai_1 _23129_ (.B1(_07528_),
    .Y(_07529_),
    .A1(net1562),
    .A2(net5001));
 sg13g2_nor2_1 _23130_ (.A(net4761),
    .B(_07529_),
    .Y(_07530_));
 sg13g2_a21oi_1 _23131_ (.A1(net5532),
    .A2(_11183_),
    .Y(_07531_),
    .B1(net1576));
 sg13g2_nor3_1 _23132_ (.A(net4786),
    .B(_07331_),
    .C(_07531_),
    .Y(_07532_));
 sg13g2_nor3_1 _23133_ (.A(net4742),
    .B(_07530_),
    .C(_07532_),
    .Y(_07533_));
 sg13g2_a21oi_1 _23134_ (.A1(_08020_),
    .A2(net4718),
    .Y(_02437_),
    .B1(_07533_));
 sg13g2_nand3_1 _23135_ (.B(_08113_),
    .C(net5001),
    .A(net6479),
    .Y(_07534_));
 sg13g2_o21ai_1 _23136_ (.B1(_07534_),
    .Y(_07535_),
    .A1(net1801),
    .A2(net5001));
 sg13g2_nand2b_1 _23137_ (.Y(_07536_),
    .B(net4787),
    .A_N(_07535_));
 sg13g2_a21oi_1 _23138_ (.A1(net5531),
    .A2(_11187_),
    .Y(_07537_),
    .B1(net2586));
 sg13g2_nor3_1 _23139_ (.A(net4788),
    .B(_07340_),
    .C(_07537_),
    .Y(_07538_));
 sg13g2_nor2_1 _23140_ (.A(net4741),
    .B(_07538_),
    .Y(_07539_));
 sg13g2_a22oi_1 _23141_ (.Y(_02438_),
    .B1(_07536_),
    .B2(_07539_),
    .A2(net4717),
    .A1(_08021_));
 sg13g2_nand3_1 _23142_ (.B(_08115_),
    .C(net5005),
    .A(net6478),
    .Y(_07540_));
 sg13g2_o21ai_1 _23143_ (.B1(_07540_),
    .Y(_07541_),
    .A1(net1853),
    .A2(net5003));
 sg13g2_nor2_1 _23144_ (.A(net4761),
    .B(_07541_),
    .Y(_07542_));
 sg13g2_a21oi_1 _23145_ (.A1(net5531),
    .A2(_11191_),
    .Y(_07543_),
    .B1(net2133));
 sg13g2_nor3_1 _23146_ (.A(net4788),
    .B(_07347_),
    .C(_07543_),
    .Y(_07544_));
 sg13g2_nor3_1 _23147_ (.A(net4741),
    .B(_07542_),
    .C(_07544_),
    .Y(_07545_));
 sg13g2_a21oi_1 _23148_ (.A1(_08023_),
    .A2(net4717),
    .Y(_02439_),
    .B1(_07545_));
 sg13g2_nand3_1 _23149_ (.B(_08116_),
    .C(net5001),
    .A(net6479),
    .Y(_07546_));
 sg13g2_o21ai_1 _23150_ (.B1(_07546_),
    .Y(_07547_),
    .A1(net1668),
    .A2(net5001));
 sg13g2_nand2b_1 _23151_ (.Y(_07548_),
    .B(net4786),
    .A_N(_07547_));
 sg13g2_a21oi_1 _23152_ (.A1(net5531),
    .A2(_11195_),
    .Y(_07549_),
    .B1(net2460));
 sg13g2_nor3_1 _23153_ (.A(net4788),
    .B(_07356_),
    .C(_07549_),
    .Y(_07550_));
 sg13g2_nor2_1 _23154_ (.A(net4741),
    .B(_07550_),
    .Y(_07551_));
 sg13g2_a22oi_1 _23155_ (.Y(_02440_),
    .B1(_07548_),
    .B2(_07551_),
    .A2(net4717),
    .A1(_08025_));
 sg13g2_o21ai_1 _23156_ (.B1(net5001),
    .Y(_07552_),
    .A1(\soc_inst.cpu_core.id_int_is_interrupt ),
    .A2(net3070));
 sg13g2_nand2_1 _23157_ (.Y(_07553_),
    .A(net4934),
    .B(_07552_));
 sg13g2_o21ai_1 _23158_ (.B1(net6025),
    .Y(_07554_),
    .A1(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .A2(_09117_));
 sg13g2_o21ai_1 _23159_ (.B1(_09117_),
    .Y(_07555_),
    .A1(net6304),
    .A2(_09513_));
 sg13g2_nand3_1 _23160_ (.B(net5341),
    .C(net5527),
    .A(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .Y(_07556_));
 sg13g2_nand2_1 _23161_ (.Y(_07557_),
    .A(net3070),
    .B(_11235_));
 sg13g2_nand4_1 _23162_ (.B(_07555_),
    .C(_07556_),
    .A(_07554_),
    .Y(_07558_),
    .D(_07557_));
 sg13g2_o21ai_1 _23163_ (.B1(_07553_),
    .Y(_07559_),
    .A1(_09044_),
    .A2(_07558_));
 sg13g2_o21ai_1 _23164_ (.B1(_07559_),
    .Y(_02441_),
    .A1(_09802_),
    .A2(_07202_));
 sg13g2_nand2_1 _23165_ (.Y(_07560_),
    .A(_08908_),
    .B(_09426_));
 sg13g2_nand2_1 _23166_ (.Y(_07561_),
    .A(net1105),
    .B(_07560_));
 sg13g2_o21ai_1 _23167_ (.B1(_07561_),
    .Y(_02442_),
    .A1(_07785_),
    .A2(_07560_));
 sg13g2_a22oi_1 _23168_ (.Y(_07562_),
    .B1(_11139_),
    .B2(net2626),
    .A2(_11137_),
    .A1(net5533));
 sg13g2_nand2_1 _23169_ (.Y(_07563_),
    .A(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .B(net4939));
 sg13g2_o21ai_1 _23170_ (.B1(net4945),
    .Y(_07564_),
    .A1(net6472),
    .A2(net2626));
 sg13g2_nand3b_1 _23171_ (.B(_07563_),
    .C(_07564_),
    .Y(_07565_),
    .A_N(net4792));
 sg13g2_nand3_1 _23172_ (.B(_09043_),
    .C(_07562_),
    .A(net5156),
    .Y(_07566_));
 sg13g2_nor2_1 _23173_ (.A(_09023_),
    .B(_07204_),
    .Y(_07567_));
 sg13g2_a22oi_1 _23174_ (.Y(_07568_),
    .B1(_07567_),
    .B2(net2626),
    .A2(_07566_),
    .A1(_07565_));
 sg13g2_inv_1 _23175_ (.Y(_02443_),
    .A(net2627));
 sg13g2_o21ai_1 _23176_ (.B1(net4738),
    .Y(_07569_),
    .A1(net2792),
    .A2(net6472));
 sg13g2_nor2_1 _23177_ (.A(_07790_),
    .B(_11147_),
    .Y(_07570_));
 sg13g2_o21ai_1 _23178_ (.B1(net4792),
    .Y(_07571_),
    .A1(_07473_),
    .A2(_07570_));
 sg13g2_nor3_1 _23179_ (.A(net2792),
    .B(_09023_),
    .C(_07202_),
    .Y(_07572_));
 sg13g2_a21oi_1 _23180_ (.A1(_07569_),
    .A2(_07571_),
    .Y(_02444_),
    .B1(_07572_));
 sg13g2_o21ai_1 _23181_ (.B1(net4738),
    .Y(_07573_),
    .A1(net2771),
    .A2(net6472));
 sg13g2_nor2_1 _23182_ (.A(_07789_),
    .B(_11151_),
    .Y(_07574_));
 sg13g2_o21ai_1 _23183_ (.B1(net4792),
    .Y(_07575_),
    .A1(_07482_),
    .A2(_07574_));
 sg13g2_nor3_1 _23184_ (.A(net2771),
    .B(_09023_),
    .C(_07202_),
    .Y(_07576_));
 sg13g2_a21oi_1 _23185_ (.A1(_07573_),
    .A2(_07575_),
    .Y(_02445_),
    .B1(_07576_));
 sg13g2_nor2b_1 _23186_ (.A(\soc_inst.gpio_inst.gpio_sync2[6] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[6] ),
    .Y(_07577_));
 sg13g2_a21oi_1 _23187_ (.A1(net86),
    .A2(_07577_),
    .Y(_07578_),
    .B1(net703));
 sg13g2_a21oi_1 _23188_ (.A1(net6457),
    .A2(_09440_),
    .Y(_02446_),
    .B1(net704));
 sg13g2_nor2b_1 _23189_ (.A(\soc_inst.gpio_inst.gpio_sync2[5] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[5] ),
    .Y(_07579_));
 sg13g2_a21oi_1 _23190_ (.A1(net84),
    .A2(_07579_),
    .Y(_07580_),
    .B1(net407));
 sg13g2_a21oi_1 _23191_ (.A1(net6460),
    .A2(_09440_),
    .Y(_02447_),
    .B1(net408));
 sg13g2_nor2b_1 _23192_ (.A(\soc_inst.gpio_inst.gpio_sync2[4] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[4] ),
    .Y(_07581_));
 sg13g2_a21oi_1 _23193_ (.A1(net87),
    .A2(_07581_),
    .Y(_07582_),
    .B1(\soc_inst.gpio_inst.int_pend_reg[4] ));
 sg13g2_a21oi_1 _23194_ (.A1(net245),
    .A2(_09440_),
    .Y(_02448_),
    .B1(_07582_));
 sg13g2_nor2b_1 _23195_ (.A(\soc_inst.gpio_inst.gpio_sync2[3] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[3] ),
    .Y(_07583_));
 sg13g2_a21oi_1 _23196_ (.A1(net88),
    .A2(_07583_),
    .Y(_07584_),
    .B1(\soc_inst.gpio_inst.int_pend_reg[3] ));
 sg13g2_a21oi_1 _23197_ (.A1(net212),
    .A2(_09440_),
    .Y(_02449_),
    .B1(_07584_));
 sg13g2_nor2b_1 _23198_ (.A(\soc_inst.gpio_inst.gpio_sync2[2] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[2] ),
    .Y(_07585_));
 sg13g2_a21oi_1 _23199_ (.A1(net83),
    .A2(_07585_),
    .Y(_07586_),
    .B1(net428));
 sg13g2_a21oi_1 _23200_ (.A1(net6467),
    .A2(_09440_),
    .Y(_02450_),
    .B1(net429));
 sg13g2_nor2b_1 _23201_ (.A(\soc_inst.gpio_inst.gpio_sync2[1] ),
    .B_N(\soc_inst.gpio_inst.int_en_reg[1] ),
    .Y(_07587_));
 sg13g2_a21oi_1 _23202_ (.A1(net81),
    .A2(_07587_),
    .Y(_07588_),
    .B1(net290));
 sg13g2_a21oi_1 _23203_ (.A1(net6469),
    .A2(_09440_),
    .Y(_02451_),
    .B1(net291));
 sg13g2_nor2_1 _23204_ (.A(net6406),
    .B(net2809),
    .Y(_07589_));
 sg13g2_a21oi_1 _23205_ (.A1(net6369),
    .A2(_08082_),
    .Y(_02452_),
    .B1(_07589_));
 sg13g2_nor2_1 _23206_ (.A(net6414),
    .B(net2093),
    .Y(_07590_));
 sg13g2_a21oi_1 _23207_ (.A1(net6414),
    .A2(_08083_),
    .Y(_02453_),
    .B1(_07590_));
 sg13g2_nor2_1 _23208_ (.A(net6413),
    .B(net1316),
    .Y(_07591_));
 sg13g2_a21oi_1 _23209_ (.A1(net6413),
    .A2(_08084_),
    .Y(_02454_),
    .B1(_07591_));
 sg13g2_nor2_1 _23210_ (.A(net6406),
    .B(net2324),
    .Y(_07592_));
 sg13g2_a21oi_1 _23211_ (.A1(net6406),
    .A2(_08085_),
    .Y(_02455_),
    .B1(_07592_));
 sg13g2_nor2_1 _23212_ (.A(net6414),
    .B(net2046),
    .Y(_07593_));
 sg13g2_a21oi_1 _23213_ (.A1(net6414),
    .A2(_08087_),
    .Y(_02456_),
    .B1(_07593_));
 sg13g2_nor2_1 _23214_ (.A(net6414),
    .B(net1748),
    .Y(_07594_));
 sg13g2_a21oi_1 _23215_ (.A1(net6414),
    .A2(_08089_),
    .Y(_02457_),
    .B1(_07594_));
 sg13g2_nor2_1 _23216_ (.A(net6407),
    .B(net1946),
    .Y(_07595_));
 sg13g2_a21oi_1 _23217_ (.A1(net6407),
    .A2(_08091_),
    .Y(_02458_),
    .B1(_07595_));
 sg13g2_nor2_1 _23218_ (.A(net6407),
    .B(net2271),
    .Y(_07596_));
 sg13g2_a21oi_1 _23219_ (.A1(net6408),
    .A2(_08093_),
    .Y(_02459_),
    .B1(_07596_));
 sg13g2_nor2_1 _23220_ (.A(net6405),
    .B(net2258),
    .Y(_07597_));
 sg13g2_a21oi_1 _23221_ (.A1(net6405),
    .A2(_08095_),
    .Y(_02460_),
    .B1(_07597_));
 sg13g2_a21o_1 _23222_ (.A2(net3056),
    .A1(net6404),
    .B1(_04358_),
    .X(_02461_));
 sg13g2_a21o_1 _23223_ (.A2(net3106),
    .A1(net6409),
    .B1(_04360_),
    .X(_02462_));
 sg13g2_a21o_1 _23224_ (.A2(net3075),
    .A1(net6404),
    .B1(_04362_),
    .X(_02463_));
 sg13g2_a21o_1 _23225_ (.A2(net3221),
    .A1(net6391),
    .B1(_04364_),
    .X(_02464_));
 sg13g2_a21o_1 _23226_ (.A2(net2928),
    .A1(net6390),
    .B1(_04366_),
    .X(_02465_));
 sg13g2_a21o_1 _23227_ (.A2(net3146),
    .A1(net6388),
    .B1(_04368_),
    .X(_02466_));
 sg13g2_a21o_1 _23228_ (.A2(net3184),
    .A1(net6390),
    .B1(_04370_),
    .X(_02467_));
 sg13g2_a21o_1 _23229_ (.A2(net3305),
    .A1(net6386),
    .B1(_04372_),
    .X(_02468_));
 sg13g2_a21o_1 _23230_ (.A2(net3137),
    .A1(net6381),
    .B1(_04374_),
    .X(_02469_));
 sg13g2_a21o_1 _23231_ (.A2(net3008),
    .A1(net6381),
    .B1(_04376_),
    .X(_02470_));
 sg13g2_a21o_1 _23232_ (.A2(net3053),
    .A1(net6381),
    .B1(_04378_),
    .X(_02471_));
 sg13g2_a21o_1 _23233_ (.A2(net3314),
    .A1(net6399),
    .B1(_04380_),
    .X(_02472_));
 sg13g2_nor2_1 _23234_ (.A(net6383),
    .B(net2078),
    .Y(_07598_));
 sg13g2_a21oi_1 _23235_ (.A1(net6383),
    .A2(_08113_),
    .Y(_02473_),
    .B1(_07598_));
 sg13g2_a21o_1 _23236_ (.A2(net3176),
    .A1(net6399),
    .B1(_04385_),
    .X(_02474_));
 sg13g2_nor2_1 _23237_ (.A(net6383),
    .B(\soc_inst.cpu_core.if_pc[23] ),
    .Y(_07599_));
 sg13g2_a21oi_1 _23238_ (.A1(net6382),
    .A2(_08116_),
    .Y(_02475_),
    .B1(_07599_));
 sg13g2_nand4_1 _23239_ (.B(\soc_inst.core_mem_addr[13] ),
    .C(_08230_),
    .A(net6205),
    .Y(_07600_),
    .D(_08793_));
 sg13g2_nor2_2 _23240_ (.A(_08672_),
    .B(_07600_),
    .Y(_07601_));
 sg13g2_nor2_1 _23241_ (.A(net2037),
    .B(net5092),
    .Y(_07602_));
 sg13g2_a21oi_1 _23242_ (.A1(net6471),
    .A2(net5092),
    .Y(_02476_),
    .B1(_07602_));
 sg13g2_nor2_1 _23243_ (.A(net1703),
    .B(net5093),
    .Y(_07603_));
 sg13g2_a21oi_1 _23244_ (.A1(net6469),
    .A2(net5093),
    .Y(_02477_),
    .B1(_07603_));
 sg13g2_nor2_1 _23245_ (.A(net2670),
    .B(net5093),
    .Y(_07604_));
 sg13g2_a21oi_1 _23246_ (.A1(net6466),
    .A2(net5093),
    .Y(_02478_),
    .B1(_07604_));
 sg13g2_nor2_1 _23247_ (.A(net2235),
    .B(net5093),
    .Y(_07605_));
 sg13g2_a21oi_1 _23248_ (.A1(net6464),
    .A2(_07601_),
    .Y(_02479_),
    .B1(_07605_));
 sg13g2_nor2_1 _23249_ (.A(net2309),
    .B(net5092),
    .Y(_07606_));
 sg13g2_a21oi_1 _23250_ (.A1(net6462),
    .A2(net5092),
    .Y(_02480_),
    .B1(_07606_));
 sg13g2_nor2_1 _23251_ (.A(net2021),
    .B(net5092),
    .Y(_07607_));
 sg13g2_a21oi_1 _23252_ (.A1(net6459),
    .A2(net5092),
    .Y(_02481_),
    .B1(_07607_));
 sg13g2_nor2_1 _23253_ (.A(net2080),
    .B(net5092),
    .Y(_07608_));
 sg13g2_a21oi_1 _23254_ (.A1(net6458),
    .A2(net5092),
    .Y(_02482_),
    .B1(_07608_));
 sg13g2_nor2_1 _23255_ (.A(net1641),
    .B(net5093),
    .Y(_07609_));
 sg13g2_a21oi_1 _23256_ (.A1(net6456),
    .A2(net5093),
    .Y(_02483_),
    .B1(_07609_));
 sg13g2_nor2_1 _23257_ (.A(net2506),
    .B(net5090),
    .Y(_07610_));
 sg13g2_a21oi_1 _23258_ (.A1(net6454),
    .A2(net5089),
    .Y(_02484_),
    .B1(_07610_));
 sg13g2_nor2_1 _23259_ (.A(net2363),
    .B(net5089),
    .Y(_07611_));
 sg13g2_a21oi_1 _23260_ (.A1(net6453),
    .A2(net5089),
    .Y(_02485_),
    .B1(_07611_));
 sg13g2_nor2_1 _23261_ (.A(net2592),
    .B(net5089),
    .Y(_07612_));
 sg13g2_a21oi_1 _23262_ (.A1(net1533),
    .A2(net5089),
    .Y(_02486_),
    .B1(_07612_));
 sg13g2_nor2_1 _23263_ (.A(net2373),
    .B(net5091),
    .Y(_07613_));
 sg13g2_a21oi_1 _23264_ (.A1(\soc_inst.core_mem_wdata[11] ),
    .A2(net5091),
    .Y(_02487_),
    .B1(_07613_));
 sg13g2_nor2_1 _23265_ (.A(_00279_),
    .B(net5091),
    .Y(_07614_));
 sg13g2_a21oi_1 _23266_ (.A1(net1825),
    .A2(net5090),
    .Y(_02488_),
    .B1(_07614_));
 sg13g2_nor2_1 _23267_ (.A(net2540),
    .B(net5089),
    .Y(_07615_));
 sg13g2_a21oi_1 _23268_ (.A1(net1321),
    .A2(net5090),
    .Y(_02489_),
    .B1(_07615_));
 sg13g2_nor2_1 _23269_ (.A(net2413),
    .B(net5089),
    .Y(_07616_));
 sg13g2_a21oi_1 _23270_ (.A1(net1503),
    .A2(net5090),
    .Y(_02490_),
    .B1(_07616_));
 sg13g2_nor2_1 _23271_ (.A(net2683),
    .B(net5089),
    .Y(_07617_));
 sg13g2_a21oi_1 _23272_ (.A1(\soc_inst.core_mem_wdata[15] ),
    .A2(net5090),
    .Y(_02491_),
    .B1(_07617_));
 sg13g2_nand2_2 _23273_ (.Y(_07618_),
    .A(_11311_),
    .B(_11313_));
 sg13g2_nand2_2 _23274_ (.Y(_07619_),
    .A(net6003),
    .B(_07618_));
 sg13g2_and2_1 _23275_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ),
    .B(net6003),
    .X(_07620_));
 sg13g2_a21oi_1 _23276_ (.A1(net1648),
    .A2(_11290_),
    .Y(_07621_),
    .B1(_07620_));
 sg13g2_o21ai_1 _23277_ (.B1(net6549),
    .Y(_07622_),
    .A1(net2386),
    .A2(net5054));
 sg13g2_a21oi_1 _23278_ (.A1(net5054),
    .A2(_07621_),
    .Y(_02492_),
    .B1(_07622_));
 sg13g2_and2_1 _23279_ (.A(net2194),
    .B(net6003),
    .X(_07623_));
 sg13g2_a21oi_1 _23280_ (.A1(net172),
    .A2(_11290_),
    .Y(_07624_),
    .B1(_07623_));
 sg13g2_o21ai_1 _23281_ (.B1(net6547),
    .Y(_07625_),
    .A1(net2512),
    .A2(net5054));
 sg13g2_a21oi_1 _23282_ (.A1(net5054),
    .A2(_07624_),
    .Y(_02493_),
    .B1(_07625_));
 sg13g2_and2_1 _23283_ (.A(net1994),
    .B(net6003),
    .X(_07626_));
 sg13g2_a21oi_1 _23284_ (.A1(net1388),
    .A2(_11290_),
    .Y(_07627_),
    .B1(_07626_));
 sg13g2_o21ai_1 _23285_ (.B1(net6547),
    .Y(_07628_),
    .A1(net2194),
    .A2(net5054));
 sg13g2_a21oi_1 _23286_ (.A1(net5054),
    .A2(_07627_),
    .Y(_02494_),
    .B1(_07628_));
 sg13g2_and2_1 _23287_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .B(net6003),
    .X(_07629_));
 sg13g2_a21oi_1 _23288_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ),
    .A2(_11290_),
    .Y(_07630_),
    .B1(_07629_));
 sg13g2_o21ai_1 _23289_ (.B1(net6547),
    .Y(_07631_),
    .A1(net1994),
    .A2(net5054));
 sg13g2_a21oi_1 _23290_ (.A1(_07619_),
    .A2(_07630_),
    .Y(_02495_),
    .B1(_07631_));
 sg13g2_and2_1 _23291_ (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ),
    .B(net6003),
    .X(_07632_));
 sg13g2_a21oi_1 _23292_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .A2(_11290_),
    .Y(_07633_),
    .B1(_07632_));
 sg13g2_o21ai_1 _23293_ (.B1(net6547),
    .Y(_07634_),
    .A1(net2015),
    .A2(_07619_));
 sg13g2_a21oi_1 _23294_ (.A1(_07619_),
    .A2(_07633_),
    .Y(_02496_),
    .B1(_07634_));
 sg13g2_a22oi_1 _23295_ (.Y(_07635_),
    .B1(_07618_),
    .B2(_07632_),
    .A2(_11290_),
    .A1(net1712));
 sg13g2_and2_1 _23296_ (.A(net2969),
    .B(net6003),
    .X(_07636_));
 sg13g2_nand2_1 _23297_ (.Y(_07637_),
    .A(net5054),
    .B(_07636_));
 sg13g2_a21oi_1 _23298_ (.A1(_07635_),
    .A2(_07637_),
    .Y(_02497_),
    .B1(_07884_));
 sg13g2_nand2_1 _23299_ (.Y(_07638_),
    .A(net3302),
    .B(_11291_));
 sg13g2_a22oi_1 _23300_ (.Y(_07639_),
    .B1(_07618_),
    .B2(_07636_),
    .A2(_11290_),
    .A1(net1696));
 sg13g2_o21ai_1 _23301_ (.B1(_07639_),
    .Y(_07640_),
    .A1(_07618_),
    .A2(net3303));
 sg13g2_and2_1 _23302_ (.A(net6549),
    .B(_07640_),
    .X(_02498_));
 sg13g2_mux2_1 _23303_ (.A0(net799),
    .A1(net6468),
    .S(_09301_),
    .X(_02499_));
 sg13g2_nor2_1 _23304_ (.A(net6050),
    .B(_07600_),
    .Y(_07641_));
 sg13g2_nor2_1 _23305_ (.A(net2160),
    .B(net5079),
    .Y(_07642_));
 sg13g2_a21oi_1 _23306_ (.A1(net6471),
    .A2(net5079),
    .Y(_02500_),
    .B1(_07642_));
 sg13g2_nor2_1 _23307_ (.A(net2110),
    .B(net5080),
    .Y(_07643_));
 sg13g2_a21oi_1 _23308_ (.A1(net6469),
    .A2(net5079),
    .Y(_02501_),
    .B1(_07643_));
 sg13g2_nor2_1 _23309_ (.A(net2002),
    .B(net5080),
    .Y(_07644_));
 sg13g2_a21oi_1 _23310_ (.A1(net6466),
    .A2(net5080),
    .Y(_02502_),
    .B1(_07644_));
 sg13g2_nor2_1 _23311_ (.A(net2284),
    .B(net5079),
    .Y(_07645_));
 sg13g2_a21oi_1 _23312_ (.A1(net6464),
    .A2(net5080),
    .Y(_02503_),
    .B1(_07645_));
 sg13g2_nor2_1 _23313_ (.A(net2279),
    .B(net5079),
    .Y(_07646_));
 sg13g2_a21oi_1 _23314_ (.A1(net6462),
    .A2(net5079),
    .Y(_02504_),
    .B1(_07646_));
 sg13g2_nor2_1 _23315_ (.A(net2193),
    .B(net5079),
    .Y(_07647_));
 sg13g2_a21oi_1 _23316_ (.A1(net6459),
    .A2(net5079),
    .Y(_02505_),
    .B1(_07647_));
 sg13g2_nor2_1 _23317_ (.A(net1758),
    .B(net5080),
    .Y(_07648_));
 sg13g2_a21oi_1 _23318_ (.A1(net6458),
    .A2(net5081),
    .Y(_02506_),
    .B1(_07648_));
 sg13g2_nor2_1 _23319_ (.A(net1319),
    .B(net5081),
    .Y(_07649_));
 sg13g2_a21oi_1 _23320_ (.A1(net6456),
    .A2(net5081),
    .Y(_02507_),
    .B1(_07649_));
 sg13g2_nor2_1 _23321_ (.A(net2553),
    .B(net5077),
    .Y(_07650_));
 sg13g2_a21oi_1 _23322_ (.A1(net6454),
    .A2(net5078),
    .Y(_02508_),
    .B1(_07650_));
 sg13g2_nor2_1 _23323_ (.A(_00292_),
    .B(net5077),
    .Y(_07651_));
 sg13g2_a21oi_1 _23324_ (.A1(net219),
    .A2(net5078),
    .Y(_02509_),
    .B1(_07651_));
 sg13g2_nor2_1 _23325_ (.A(net2362),
    .B(net5077),
    .Y(_07652_));
 sg13g2_a21oi_1 _23326_ (.A1(net1533),
    .A2(net5077),
    .Y(_02510_),
    .B1(_07652_));
 sg13g2_nor2_1 _23327_ (.A(net2227),
    .B(net5077),
    .Y(_07653_));
 sg13g2_a21oi_1 _23328_ (.A1(\soc_inst.core_mem_wdata[11] ),
    .A2(net5077),
    .Y(_02511_),
    .B1(_07653_));
 sg13g2_nor2_1 _23329_ (.A(net1996),
    .B(net5078),
    .Y(_07654_));
 sg13g2_a21oi_1 _23330_ (.A1(net1825),
    .A2(net5078),
    .Y(_02512_),
    .B1(_07654_));
 sg13g2_nor2_1 _23331_ (.A(net2310),
    .B(net5078),
    .Y(_07655_));
 sg13g2_a21oi_1 _23332_ (.A1(net1321),
    .A2(net5077),
    .Y(_02513_),
    .B1(_07655_));
 sg13g2_nor2_1 _23333_ (.A(net1457),
    .B(net5078),
    .Y(_07656_));
 sg13g2_a21oi_1 _23334_ (.A1(\soc_inst.core_mem_wdata[14] ),
    .A2(net5088),
    .Y(_02514_),
    .B1(_07656_));
 sg13g2_nor2_1 _23335_ (.A(net1855),
    .B(net5078),
    .Y(_07657_));
 sg13g2_a21oi_1 _23336_ (.A1(\soc_inst.core_mem_wdata[15] ),
    .A2(net5077),
    .Y(_02515_),
    .B1(_07657_));
 sg13g2_nor2_1 _23337_ (.A(_00299_),
    .B(net5084),
    .Y(_07658_));
 sg13g2_a21oi_1 _23338_ (.A1(net225),
    .A2(net5084),
    .Y(_02516_),
    .B1(_07658_));
 sg13g2_nor2_1 _23339_ (.A(_00300_),
    .B(net5082),
    .Y(_07659_));
 sg13g2_a21oi_1 _23340_ (.A1(net160),
    .A2(net5084),
    .Y(_02517_),
    .B1(_07659_));
 sg13g2_nor2_1 _23341_ (.A(_00301_),
    .B(net5082),
    .Y(_07660_));
 sg13g2_a21oi_1 _23342_ (.A1(net1272),
    .A2(net5082),
    .Y(_02518_),
    .B1(_07660_));
 sg13g2_nor2_1 _23343_ (.A(_00302_),
    .B(net5082),
    .Y(_07661_));
 sg13g2_a21oi_1 _23344_ (.A1(net295),
    .A2(net5083),
    .Y(_02519_),
    .B1(_07661_));
 sg13g2_nor2_1 _23345_ (.A(_00303_),
    .B(net5082),
    .Y(_07662_));
 sg13g2_a21oi_1 _23346_ (.A1(net548),
    .A2(net5082),
    .Y(_02520_),
    .B1(_07662_));
 sg13g2_nor2_1 _23347_ (.A(_00304_),
    .B(net5083),
    .Y(_07663_));
 sg13g2_a21oi_1 _23348_ (.A1(net571),
    .A2(net5083),
    .Y(_02521_),
    .B1(_07663_));
 sg13g2_nor2_1 _23349_ (.A(_00305_),
    .B(net5083),
    .Y(_07664_));
 sg13g2_a21oi_1 _23350_ (.A1(net1311),
    .A2(net5083),
    .Y(_02522_),
    .B1(_07664_));
 sg13g2_nor2_1 _23351_ (.A(net1931),
    .B(net5082),
    .Y(_07665_));
 sg13g2_a21oi_1 _23352_ (.A1(net1329),
    .A2(net5082),
    .Y(_02523_),
    .B1(_07665_));
 sg13g2_nor2_1 _23353_ (.A(_00307_),
    .B(net5085),
    .Y(_07666_));
 sg13g2_a21oi_1 _23354_ (.A1(net268),
    .A2(net5085),
    .Y(_02524_),
    .B1(_07666_));
 sg13g2_nor2_1 _23355_ (.A(_00308_),
    .B(net5085),
    .Y(_07667_));
 sg13g2_a21oi_1 _23356_ (.A1(net233),
    .A2(net5085),
    .Y(_02525_),
    .B1(_07667_));
 sg13g2_nor2_1 _23357_ (.A(_00309_),
    .B(net5086),
    .Y(_07668_));
 sg13g2_a21oi_1 _23358_ (.A1(net1016),
    .A2(net5086),
    .Y(_02526_),
    .B1(_07668_));
 sg13g2_nor2_1 _23359_ (.A(_00310_),
    .B(net5086),
    .Y(_07669_));
 sg13g2_a21oi_1 _23360_ (.A1(net712),
    .A2(net5084),
    .Y(_02527_),
    .B1(_07669_));
 sg13g2_nor2_1 _23361_ (.A(_00311_),
    .B(net5087),
    .Y(_07670_));
 sg13g2_a21oi_1 _23362_ (.A1(net369),
    .A2(net5087),
    .Y(_02528_),
    .B1(_07670_));
 sg13g2_nor2_1 _23363_ (.A(_00312_),
    .B(net5087),
    .Y(_07671_));
 sg13g2_a21oi_1 _23364_ (.A1(net313),
    .A2(net5087),
    .Y(_02529_),
    .B1(_07671_));
 sg13g2_nor2_1 _23365_ (.A(_00313_),
    .B(net5085),
    .Y(_07672_));
 sg13g2_a21oi_1 _23366_ (.A1(net734),
    .A2(net5085),
    .Y(_02530_),
    .B1(_07672_));
 sg13g2_nor2_1 _23367_ (.A(_00314_),
    .B(net5085),
    .Y(_07673_));
 sg13g2_a21oi_1 _23368_ (.A1(net854),
    .A2(net5085),
    .Y(_02531_),
    .B1(_07673_));
 sg13g2_nand3_1 _23369_ (.B(_09308_),
    .C(_09426_),
    .A(net6204),
    .Y(_07674_));
 sg13g2_mux2_1 _23370_ (.A0(net6470),
    .A1(net1648),
    .S(net5053),
    .X(_02532_));
 sg13g2_nand2_1 _23371_ (.Y(_07675_),
    .A(net172),
    .B(net5053));
 sg13g2_o21ai_1 _23372_ (.B1(_07675_),
    .Y(_02533_),
    .A1(_07784_),
    .A2(_07674_));
 sg13g2_mux2_1 _23373_ (.A0(net6465),
    .A1(net1388),
    .S(net5053),
    .X(_02534_));
 sg13g2_mux2_1 _23374_ (.A0(net6463),
    .A1(net2112),
    .S(net5053),
    .X(_02535_));
 sg13g2_mux2_1 _23375_ (.A0(net6461),
    .A1(net2329),
    .S(net5053),
    .X(_02536_));
 sg13g2_mux2_1 _23376_ (.A0(net6459),
    .A1(net1712),
    .S(net5053),
    .X(_02537_));
 sg13g2_mux2_1 _23377_ (.A0(net6457),
    .A1(net1696),
    .S(net5053),
    .X(_02538_));
 sg13g2_mux2_1 _23378_ (.A0(net6455),
    .A1(net494),
    .S(net5053),
    .X(_02539_));
 sg13g2_nand2_1 _23379_ (.Y(_07676_),
    .A(net494),
    .B(_11290_));
 sg13g2_a21oi_1 _23380_ (.A1(_07638_),
    .A2(net495),
    .Y(_02540_),
    .B1(_07884_));
 sg13g2_and2_1 _23381_ (.A(net6487),
    .B(_11311_),
    .X(_07677_));
 sg13g2_nor2_1 _23382_ (.A(net2406),
    .B(_07677_),
    .Y(_07678_));
 sg13g2_nand4_1 _23383_ (.B(_07782_),
    .C(_07799_),
    .A(net2746),
    .Y(_07679_),
    .D(_11287_));
 sg13g2_nand3_1 _23384_ (.B(net6549),
    .C(_07679_),
    .A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ),
    .Y(_07680_));
 sg13g2_and2_1 _23385_ (.A(net2406),
    .B(_07677_),
    .X(_07681_));
 sg13g2_nor3_1 _23386_ (.A(net2407),
    .B(_07680_),
    .C(_07681_),
    .Y(_02541_));
 sg13g2_nor2_1 _23387_ (.A(net1860),
    .B(_07681_),
    .Y(_07682_));
 sg13g2_and2_1 _23388_ (.A(net1860),
    .B(_07681_),
    .X(_07683_));
 sg13g2_nor3_1 _23389_ (.A(_07680_),
    .B(net1861),
    .C(_07683_),
    .Y(_02542_));
 sg13g2_nand2_1 _23390_ (.Y(_07684_),
    .A(net2432),
    .B(_07683_));
 sg13g2_xnor2_1 _23391_ (.Y(_07685_),
    .A(net2432),
    .B(_07683_));
 sg13g2_nor2_1 _23392_ (.A(_07680_),
    .B(_07685_),
    .Y(_02543_));
 sg13g2_xor2_1 _23393_ (.B(_07684_),
    .A(net2746),
    .X(_07686_));
 sg13g2_nor2_1 _23394_ (.A(_07680_),
    .B(_07686_),
    .Y(_02544_));
 sg13g2_nor3_1 _23395_ (.A(net3308),
    .B(net2919),
    .C(net6487),
    .Y(_07687_));
 sg13g2_nor2b_1 _23396_ (.A(_10274_),
    .B_N(net3308),
    .Y(_07688_));
 sg13g2_nor3_1 _23397_ (.A(net5108),
    .B(_07687_),
    .C(_07688_),
    .Y(_02545_));
 sg13g2_and2_1 _23398_ (.A(net2254),
    .B(_07688_),
    .X(_07689_));
 sg13g2_nor2_1 _23399_ (.A(net2254),
    .B(_07688_),
    .Y(_07690_));
 sg13g2_nor3_1 _23400_ (.A(net5108),
    .B(_07689_),
    .C(net2255),
    .Y(_02546_));
 sg13g2_and2_1 _23401_ (.A(net2340),
    .B(_07689_),
    .X(_07691_));
 sg13g2_nor2_1 _23402_ (.A(net2340),
    .B(_07689_),
    .Y(_07692_));
 sg13g2_nor3_1 _23403_ (.A(net5107),
    .B(_07691_),
    .C(net2341),
    .Y(_02547_));
 sg13g2_and2_1 _23404_ (.A(net2714),
    .B(_07691_),
    .X(_07693_));
 sg13g2_nor2_1 _23405_ (.A(net2714),
    .B(_07691_),
    .Y(_07694_));
 sg13g2_nor3_1 _23406_ (.A(net5107),
    .B(_07693_),
    .C(_07694_),
    .Y(_02548_));
 sg13g2_and2_1 _23407_ (.A(net2508),
    .B(_07693_),
    .X(_07695_));
 sg13g2_nor2_1 _23408_ (.A(net2508),
    .B(_07693_),
    .Y(_07696_));
 sg13g2_nor3_1 _23409_ (.A(net5107),
    .B(_07695_),
    .C(net2509),
    .Y(_02549_));
 sg13g2_xnor2_1 _23410_ (.Y(_07697_),
    .A(net2725),
    .B(_07695_));
 sg13g2_nor2_1 _23411_ (.A(net5107),
    .B(_07697_),
    .Y(_02550_));
 sg13g2_a21oi_1 _23412_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .A2(_07695_),
    .Y(_07698_),
    .B1(net1469));
 sg13g2_and3_1 _23413_ (.X(_07699_),
    .A(net1469),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .C(_07695_));
 sg13g2_nor3_1 _23414_ (.A(net5107),
    .B(net1470),
    .C(_07699_),
    .Y(_02551_));
 sg13g2_nor2_1 _23415_ (.A(net2675),
    .B(_07699_),
    .Y(_07700_));
 sg13g2_and2_1 _23416_ (.A(net2675),
    .B(_07699_),
    .X(_07701_));
 sg13g2_nor3_1 _23417_ (.A(net5107),
    .B(net2676),
    .C(_07701_),
    .Y(_02552_));
 sg13g2_nor2_1 _23418_ (.A(net2495),
    .B(_07701_),
    .Y(_07702_));
 sg13g2_and2_1 _23419_ (.A(net2495),
    .B(_07701_),
    .X(_07703_));
 sg13g2_nor3_1 _23420_ (.A(net5107),
    .B(net2496),
    .C(_07703_),
    .Y(_02553_));
 sg13g2_a21oi_1 _23421_ (.A1(net2963),
    .A2(_07703_),
    .Y(_07704_),
    .B1(net5107));
 sg13g2_o21ai_1 _23422_ (.B1(_07704_),
    .Y(_07705_),
    .A1(net2963),
    .A2(_07703_));
 sg13g2_inv_1 _23423_ (.Y(_02554_),
    .A(_07705_));
 sg13g2_and3_1 _23424_ (.X(_07706_),
    .A(net6204),
    .B(_09308_),
    .C(_10275_));
 sg13g2_nor2_1 _23425_ (.A(net2708),
    .B(net5052),
    .Y(_07707_));
 sg13g2_a21oi_1 _23426_ (.A1(_07785_),
    .A2(net5052),
    .Y(_02555_),
    .B1(_07707_));
 sg13g2_nor2_1 _23427_ (.A(net3124),
    .B(net5050),
    .Y(_07708_));
 sg13g2_a21oi_1 _23428_ (.A1(_07784_),
    .A2(net5050),
    .Y(_02556_),
    .B1(_07708_));
 sg13g2_nor2_1 _23429_ (.A(net3220),
    .B(net5051),
    .Y(_07709_));
 sg13g2_a21oi_1 _23430_ (.A1(net6465),
    .A2(net5050),
    .Y(_02557_),
    .B1(_07709_));
 sg13g2_nor2_1 _23431_ (.A(net3304),
    .B(net5051),
    .Y(_07710_));
 sg13g2_a21oi_1 _23432_ (.A1(net6463),
    .A2(net5050),
    .Y(_02558_),
    .B1(_07710_));
 sg13g2_mux2_1 _23433_ (.A0(net3331),
    .A1(net6461),
    .S(net5051),
    .X(_02559_));
 sg13g2_nor2_1 _23434_ (.A(net3295),
    .B(net5050),
    .Y(_07711_));
 sg13g2_a21oi_1 _23435_ (.A1(net6459),
    .A2(net5050),
    .Y(_02560_),
    .B1(_07711_));
 sg13g2_mux2_1 _23436_ (.A0(net2753),
    .A1(net6457),
    .S(net5050),
    .X(_02561_));
 sg13g2_mux2_1 _23437_ (.A0(net3337),
    .A1(net6455),
    .S(net5050),
    .X(_02562_));
 sg13g2_mux2_1 _23438_ (.A0(net3306),
    .A1(net6454),
    .S(net5052),
    .X(_02563_));
 sg13g2_nor2_1 _23439_ (.A(net2997),
    .B(net5052),
    .Y(_07712_));
 sg13g2_a21oi_1 _23440_ (.A1(net6453),
    .A2(net5052),
    .Y(_02564_),
    .B1(_07712_));
 sg13g2_nor2b_1 _23441_ (.A(net2386),
    .B_N(_11313_),
    .Y(_07713_));
 sg13g2_o21ai_1 _23442_ (.B1(net6549),
    .Y(_02565_),
    .A1(_11295_),
    .A2(_07713_));
 sg13g2_o21ai_1 _23443_ (.B1(net6550),
    .Y(_07714_),
    .A1(net6176),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ));
 sg13g2_a21oi_1 _23444_ (.A1(_07776_),
    .A2(net6176),
    .Y(_02566_),
    .B1(_07714_));
 sg13g2_o21ai_1 _23445_ (.B1(net6550),
    .Y(_07715_),
    .A1(net6176),
    .A2(net1655));
 sg13g2_a21oi_1 _23446_ (.A1(_07775_),
    .A2(net6176),
    .Y(_02567_),
    .B1(_07715_));
 sg13g2_o21ai_1 _23447_ (.B1(net6550),
    .Y(_07716_),
    .A1(net6176),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ));
 sg13g2_a21oi_1 _23448_ (.A1(_07774_),
    .A2(net6176),
    .Y(_02568_),
    .B1(_07716_));
 sg13g2_o21ai_1 _23449_ (.B1(net6551),
    .Y(_07717_),
    .A1(net6176),
    .A2(net1992));
 sg13g2_a21oi_1 _23450_ (.A1(_07773_),
    .A2(net6178),
    .Y(_02569_),
    .B1(_07717_));
 sg13g2_o21ai_1 _23451_ (.B1(net6552),
    .Y(_07718_),
    .A1(net6177),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ));
 sg13g2_a21oi_1 _23452_ (.A1(_07772_),
    .A2(net6177),
    .Y(_02570_),
    .B1(_07718_));
 sg13g2_o21ai_1 _23453_ (.B1(net6552),
    .Y(_07719_),
    .A1(net6176),
    .A2(net2175));
 sg13g2_a21oi_1 _23454_ (.A1(_07771_),
    .A2(net6177),
    .Y(_02571_),
    .B1(_07719_));
 sg13g2_o21ai_1 _23455_ (.B1(net6551),
    .Y(_07720_),
    .A1(net6177),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ));
 sg13g2_a21oi_1 _23456_ (.A1(_07770_),
    .A2(net6177),
    .Y(_02572_),
    .B1(_07720_));
 sg13g2_o21ai_1 _23457_ (.B1(net6552),
    .Y(_07721_),
    .A1(net2521),
    .A2(net6177));
 sg13g2_a21oi_1 _23458_ (.A1(_07769_),
    .A2(net6177),
    .Y(_02573_),
    .B1(_07721_));
 sg13g2_nor2b_2 _23459_ (.A(_08486_),
    .B_N(net2009),
    .Y(_07722_));
 sg13g2_nand2b_2 _23460_ (.Y(_07723_),
    .B(net2009),
    .A_N(_08486_));
 sg13g2_nor2_1 _23461_ (.A(_07884_),
    .B(net2106),
    .Y(_07724_));
 sg13g2_o21ai_1 _23462_ (.B1(net6069),
    .Y(_07725_),
    .A1(net665),
    .A2(_07723_));
 sg13g2_a21oi_1 _23463_ (.A1(_07776_),
    .A2(_07723_),
    .Y(_02574_),
    .B1(net666));
 sg13g2_o21ai_1 _23464_ (.B1(net6069),
    .Y(_07726_),
    .A1(net921),
    .A2(_07723_));
 sg13g2_a21oi_1 _23465_ (.A1(_07775_),
    .A2(_07723_),
    .Y(_02575_),
    .B1(_07726_));
 sg13g2_o21ai_1 _23466_ (.B1(net6069),
    .Y(_07727_),
    .A1(net921),
    .A2(net5024));
 sg13g2_a21oi_1 _23467_ (.A1(_07773_),
    .A2(net5024),
    .Y(_02576_),
    .B1(_07727_));
 sg13g2_o21ai_1 _23468_ (.B1(net6069),
    .Y(_07728_),
    .A1(net1018),
    .A2(net5024));
 sg13g2_a21oi_1 _23469_ (.A1(_07772_),
    .A2(net5024),
    .Y(_02577_),
    .B1(net1019));
 sg13g2_o21ai_1 _23470_ (.B1(net6069),
    .Y(_07729_),
    .A1(net746),
    .A2(_07723_));
 sg13g2_a21oi_1 _23471_ (.A1(_07772_),
    .A2(_07723_),
    .Y(_02578_),
    .B1(net747));
 sg13g2_o21ai_1 _23472_ (.B1(net6069),
    .Y(_07730_),
    .A1(net1417),
    .A2(_07723_));
 sg13g2_a21oi_1 _23473_ (.A1(_07771_),
    .A2(_07723_),
    .Y(_02579_),
    .B1(_07730_));
 sg13g2_o21ai_1 _23474_ (.B1(net6069),
    .Y(_07731_),
    .A1(net1417),
    .A2(net5024));
 sg13g2_a21oi_1 _23475_ (.A1(_07769_),
    .A2(net5024),
    .Y(_02580_),
    .B1(_07731_));
 sg13g2_o21ai_1 _23476_ (.B1(_07724_),
    .Y(_07732_),
    .A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ),
    .A2(_07722_));
 sg13g2_a21oi_1 _23477_ (.A1(_07767_),
    .A2(_07722_),
    .Y(_02581_),
    .B1(_07732_));
 sg13g2_nand3_1 _23478_ (.B(_07900_),
    .C(net6069),
    .A(_07777_),
    .Y(_07733_));
 sg13g2_nor2_1 _23479_ (.A(net2089),
    .B(net5024),
    .Y(_07734_));
 sg13g2_and2_1 _23480_ (.A(net2089),
    .B(net5024),
    .X(_07735_));
 sg13g2_nor3_1 _23481_ (.A(_07733_),
    .B(_07734_),
    .C(_07735_),
    .Y(_02582_));
 sg13g2_nor2_1 _23482_ (.A(net2420),
    .B(_07735_),
    .Y(_07736_));
 sg13g2_and2_1 _23483_ (.A(net2420),
    .B(_07735_),
    .X(_07737_));
 sg13g2_nor3_1 _23484_ (.A(_07733_),
    .B(_07736_),
    .C(_07737_),
    .Y(_02583_));
 sg13g2_a21oi_1 _23485_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .A2(_07735_),
    .Y(_07738_),
    .B1(net824));
 sg13g2_and3_1 _23486_ (.X(_07739_),
    .A(net824),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .C(_07735_));
 sg13g2_nor3_1 _23487_ (.A(_07733_),
    .B(net825),
    .C(_07739_),
    .Y(_02584_));
 sg13g2_xnor2_1 _23488_ (.Y(_07740_),
    .A(net1888),
    .B(_07739_));
 sg13g2_nor2_1 _23489_ (.A(_07733_),
    .B(net1889),
    .Y(_02585_));
 sg13g2_o21ai_1 _23490_ (.B1(net6553),
    .Y(_07741_),
    .A1(net303),
    .A2(_08477_));
 sg13g2_a21oi_1 _23491_ (.A1(_07763_),
    .A2(_08446_),
    .Y(_02586_),
    .B1(_07741_));
 sg13g2_nor3_1 _23492_ (.A(net6178),
    .B(net1842),
    .C(net2009),
    .Y(_07742_));
 sg13g2_nor2b_1 _23493_ (.A(net2890),
    .B_N(_07742_),
    .Y(_07743_));
 sg13g2_nor2b_1 _23494_ (.A(_07742_),
    .B_N(net2890),
    .Y(_07744_));
 sg13g2_nor3_1 _23495_ (.A(net5049),
    .B(_07743_),
    .C(_07744_),
    .Y(_02587_));
 sg13g2_and2_1 _23496_ (.A(net2986),
    .B(_07744_),
    .X(_07745_));
 sg13g2_nor2_1 _23497_ (.A(net2986),
    .B(_07744_),
    .Y(_07746_));
 sg13g2_nor3_1 _23498_ (.A(net5049),
    .B(_07745_),
    .C(_07746_),
    .Y(_02588_));
 sg13g2_and2_1 _23499_ (.A(net3049),
    .B(_07745_),
    .X(_07747_));
 sg13g2_nor2_1 _23500_ (.A(net3049),
    .B(_07745_),
    .Y(_07748_));
 sg13g2_nor3_1 _23501_ (.A(net5049),
    .B(_07747_),
    .C(_07748_),
    .Y(_02589_));
 sg13g2_and2_1 _23502_ (.A(net3041),
    .B(_07747_),
    .X(_07749_));
 sg13g2_nor2_1 _23503_ (.A(net3041),
    .B(_07747_),
    .Y(_07750_));
 sg13g2_nor3_1 _23504_ (.A(net5049),
    .B(_07749_),
    .C(net3042),
    .Y(_02590_));
 sg13g2_and2_1 _23505_ (.A(net2982),
    .B(_07749_),
    .X(_07751_));
 sg13g2_nor2_1 _23506_ (.A(net2982),
    .B(_07749_),
    .Y(_07752_));
 sg13g2_nor3_1 _23507_ (.A(net5049),
    .B(_07751_),
    .C(net2983),
    .Y(_02591_));
 sg13g2_o21ai_1 _23508_ (.B1(_08488_),
    .Y(_07753_),
    .A1(net1645),
    .A2(_07751_));
 sg13g2_a21oi_1 _23509_ (.A1(net1645),
    .A2(_07751_),
    .Y(_02592_),
    .B1(_07753_));
 sg13g2_a21oi_1 _23510_ (.A1(net1645),
    .A2(_07751_),
    .Y(_07754_),
    .B1(net2886));
 sg13g2_and3_2 _23511_ (.X(_07755_),
    .A(net2886),
    .B(net1645),
    .C(_07751_));
 sg13g2_nor3_1 _23512_ (.A(net5049),
    .B(net2887),
    .C(_07755_),
    .Y(_02593_));
 sg13g2_xnor2_1 _23513_ (.Y(_07756_),
    .A(net2976),
    .B(_07755_));
 sg13g2_nor2_1 _23514_ (.A(_08487_),
    .B(_07756_),
    .Y(_02594_));
 sg13g2_a21oi_1 _23515_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .A2(_07755_),
    .Y(_07757_),
    .B1(net1742));
 sg13g2_and3_1 _23516_ (.X(_07758_),
    .A(net1742),
    .B(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .C(_07755_));
 sg13g2_nor3_1 _23517_ (.A(_08487_),
    .B(net1743),
    .C(_07758_),
    .Y(_02595_));
 sg13g2_a21oi_1 _23518_ (.A1(net2932),
    .A2(_07758_),
    .Y(_07759_),
    .B1(_08487_));
 sg13g2_o21ai_1 _23519_ (.B1(_07759_),
    .Y(_07760_),
    .A1(net2932),
    .A2(_07758_));
 sg13g2_inv_1 _23520_ (.Y(_02596_),
    .A(net2933));
 sg13g2_a21oi_1 _23521_ (.A1(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .A2(net8),
    .Y(_07761_),
    .B1(_07884_));
 sg13g2_o21ai_1 _23522_ (.B1(_07761_),
    .Y(_02597_),
    .A1(_07764_),
    .A2(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ));
 sg13g2_a21oi_1 _23523_ (.A1(net738),
    .A2(net799),
    .Y(_07762_),
    .B1(_07884_));
 sg13g2_o21ai_1 _23524_ (.B1(_07762_),
    .Y(_02598_),
    .A1(_07763_),
    .A2(net799));
 sg13g2_xor2_1 _23525_ (.B(\soc_inst.spi_inst.state[0] ),
    .A(net850),
    .X(\soc_inst.spi_inst.next_state[1] ));
 sg13g2_dfrbpq_1 _23526_ (.RESET_B(net6572),
    .D(net2248),
    .Q(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23527_ (.RESET_B(net6573),
    .D(net2174),
    .Q(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23528_ (.RESET_B(net6584),
    .D(_00323_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23529_ (.RESET_B(net6572),
    .D(_00324_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _23530_ (.RESET_B(net6562),
    .D(_00325_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _23531_ (.RESET_B(net6561),
    .D(_00326_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _23532_ (.RESET_B(net6551),
    .D(_00327_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _23533_ (.RESET_B(net6562),
    .D(_00328_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _23534_ (.RESET_B(net6561),
    .D(_00329_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _23535_ (.RESET_B(net6559),
    .D(_00330_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _23536_ (.RESET_B(net6561),
    .D(_00331_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _23537_ (.RESET_B(net6561),
    .D(net2552),
    .Q(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _23538_ (.RESET_B(net6559),
    .D(_00333_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _23539_ (.RESET_B(net6554),
    .D(_00334_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _23540_ (.RESET_B(net6554),
    .D(_00335_),
    .Q(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _23541_ (.RESET_B(net6564),
    .D(net2581),
    .Q(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _23542_ (.RESET_B(net6589),
    .D(net2654),
    .Q(\soc_inst.spi_inst.spi_sclk ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _23543_ (.RESET_B(net6589),
    .D(net1444),
    .Q(\soc_inst.spi_inst.spi_mosi ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _23544_ (.RESET_B(net6586),
    .D(net722),
    .Q(\soc_inst.spi_inst.start_pending ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _23545_ (.RESET_B(net6613),
    .D(_00138_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[0] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23546_ (.RESET_B(net6614),
    .D(net188),
    .Q(\soc_inst.spi_inst.tx_shift_reg[1] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _23547_ (.RESET_B(net6617),
    .D(net190),
    .Q(\soc_inst.spi_inst.tx_shift_reg[2] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _23548_ (.RESET_B(net6613),
    .D(_00163_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[3] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _23549_ (.RESET_B(net6613),
    .D(net287),
    .Q(\soc_inst.spi_inst.tx_shift_reg[4] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23550_ (.RESET_B(net6613),
    .D(net156),
    .Q(\soc_inst.spi_inst.tx_shift_reg[5] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _23551_ (.RESET_B(net6613),
    .D(_00166_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[6] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _23552_ (.RESET_B(net6613),
    .D(net331),
    .Q(\soc_inst.spi_inst.tx_shift_reg[7] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23553_ (.RESET_B(net6613),
    .D(net175),
    .Q(\soc_inst.spi_inst.tx_shift_reg[8] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23554_ (.RESET_B(net6605),
    .D(net164),
    .Q(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _23555_ (.RESET_B(net6604),
    .D(net597),
    .Q(\soc_inst.spi_inst.tx_shift_reg[10] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23556_ (.RESET_B(net6604),
    .D(net414),
    .Q(\soc_inst.spi_inst.tx_shift_reg[11] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23557_ (.RESET_B(net6604),
    .D(_00141_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[12] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23558_ (.RESET_B(net6604),
    .D(net159),
    .Q(\soc_inst.spi_inst.tx_shift_reg[13] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _23559_ (.RESET_B(net6600),
    .D(_00143_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[14] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _23560_ (.RESET_B(net6557),
    .D(net205),
    .Q(\soc_inst.spi_inst.tx_shift_reg[15] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _23561_ (.RESET_B(net6556),
    .D(_00145_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[16] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _23562_ (.RESET_B(net6556),
    .D(_00146_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[17] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_1 _23563_ (.RESET_B(net6556),
    .D(net308),
    .Q(\soc_inst.spi_inst.tx_shift_reg[18] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _23564_ (.RESET_B(net6557),
    .D(net201),
    .Q(\soc_inst.spi_inst.tx_shift_reg[19] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_1 _23565_ (.RESET_B(net6557),
    .D(net1494),
    .Q(\soc_inst.spi_inst.tx_shift_reg[20] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _23566_ (.RESET_B(net6558),
    .D(_00151_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[21] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_1 _23567_ (.RESET_B(net6558),
    .D(net1336),
    .Q(\soc_inst.spi_inst.tx_shift_reg[22] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_1 _23568_ (.RESET_B(net6558),
    .D(net1104),
    .Q(\soc_inst.spi_inst.tx_shift_reg[23] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_1 _23569_ (.RESET_B(net6557),
    .D(net250),
    .Q(\soc_inst.spi_inst.tx_shift_reg[24] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _23570_ (.RESET_B(net6554),
    .D(net211),
    .Q(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _23571_ (.RESET_B(net6562),
    .D(_00156_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[26] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23572_ (.RESET_B(net6584),
    .D(_00157_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[27] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23573_ (.RESET_B(net6587),
    .D(net230),
    .Q(\soc_inst.spi_inst.tx_shift_reg[28] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _23574_ (.RESET_B(net6635),
    .D(_00159_),
    .Q(\soc_inst.spi_inst.tx_shift_reg[29] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23575_ (.RESET_B(net6584),
    .D(net263),
    .Q(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _23576_ (.RESET_B(net6585),
    .D(net366),
    .Q(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _23577_ (.RESET_B(net6586),
    .D(_00338_),
    .Q(\soc_inst.spi_inst.bit_counter[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _23578_ (.RESET_B(net6586),
    .D(net2085),
    .Q(\soc_inst.spi_inst.bit_counter[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _23579_ (.RESET_B(net6586),
    .D(net2608),
    .Q(\soc_inst.spi_inst.bit_counter[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _23580_ (.RESET_B(net6587),
    .D(net2430),
    .Q(\soc_inst.spi_inst.bit_counter[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _23581_ (.RESET_B(net6587),
    .D(_00342_),
    .Q(\soc_inst.spi_inst.bit_counter[4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _23582_ (.RESET_B(net6586),
    .D(_00343_),
    .Q(\soc_inst.spi_inst.bit_counter[5] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23583_ (.RESET_B(net6586),
    .D(net185),
    .Q(\soc_inst.spi_inst.state[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _23584_ (.RESET_B(net6593),
    .D(net851),
    .Q(\soc_inst.spi_inst.state[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _23585_ (.RESET_B(net6631),
    .D(_00344_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23586_ (.RESET_B(net6611),
    .D(_00345_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23587_ (.RESET_B(net6633),
    .D(_00346_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23588_ (.RESET_B(net6633),
    .D(_00347_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23589_ (.RESET_B(net6633),
    .D(_00348_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23590_ (.RESET_B(net6641),
    .D(_00349_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23591_ (.RESET_B(net6633),
    .D(_00350_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _23592_ (.RESET_B(net6633),
    .D(_00351_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _23593_ (.RESET_B(net6641),
    .D(_00352_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23594_ (.RESET_B(net6611),
    .D(_00353_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23595_ (.RESET_B(net6610),
    .D(_00354_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _23596_ (.RESET_B(net6610),
    .D(_00355_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _23597_ (.RESET_B(net6611),
    .D(_00356_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _23598_ (.RESET_B(net6641),
    .D(_00357_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23599_ (.RESET_B(net6641),
    .D(_00358_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23600_ (.RESET_B(net6641),
    .D(_00359_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _23601_ (.RESET_B(net6630),
    .D(_00360_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[16] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _23602_ (.RESET_B(net6630),
    .D(_00361_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _23603_ (.RESET_B(net6631),
    .D(_00362_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _23604_ (.RESET_B(net6630),
    .D(_00363_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _23605_ (.RESET_B(net6630),
    .D(_00364_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _23606_ (.RESET_B(net6630),
    .D(_00365_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23607_ (.RESET_B(net6630),
    .D(_00366_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _23608_ (.RESET_B(net6630),
    .D(_00367_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23609_ (.RESET_B(net6630),
    .D(_00368_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[24] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23610_ (.RESET_B(net6632),
    .D(_00369_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[25] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23611_ (.RESET_B(net6632),
    .D(_00370_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[26] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23612_ (.RESET_B(net6631),
    .D(_00371_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[27] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23613_ (.RESET_B(net6631),
    .D(_00372_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[28] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23614_ (.RESET_B(net6631),
    .D(_00373_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[29] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23615_ (.RESET_B(net6631),
    .D(_00374_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[30] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23616_ (.RESET_B(net6631),
    .D(_00375_),
    .Q(\soc_inst.spi_inst.rx_shift_reg[31] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23617_ (.RESET_B(net6584),
    .D(_00376_),
    .Q(\soc_inst.spi_inst.cpha ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _23618_ (.RESET_B(net6579),
    .D(_00377_),
    .Q(\soc_inst.spi_ena ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _23619_ (.RESET_B(net6588),
    .D(net2096),
    .Q(_00221_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _23620_ (.RESET_B(net6585),
    .D(_00379_),
    .Q(_00222_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _23621_ (.RESET_B(net6586),
    .D(net1206),
    .Q(_00223_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _23622_ (.RESET_B(net6588),
    .D(_00381_),
    .Q(_00224_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _23623_ (.RESET_B(net6586),
    .D(_00382_),
    .Q(_00225_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _23624_ (.RESET_B(net6584),
    .D(_00383_),
    .Q(\soc_inst.spi_inst.clock_divider[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _23625_ (.RESET_B(net6588),
    .D(_00384_),
    .Q(\soc_inst.spi_inst.clock_divider[6] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _23626_ (.RESET_B(net6584),
    .D(_00385_),
    .Q(\soc_inst.spi_inst.clock_divider[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23627_ (.RESET_B(net6593),
    .D(_00386_),
    .Q(\soc_inst.spi_inst.done ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23628_ (.RESET_B(net6562),
    .D(_00387_),
    .Q(\soc_inst.spi_inst.cpol ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _23629_ (.RESET_B(net6589),
    .D(_11837_[0]),
    .Q(\soc_inst.spi_inst.spi_clk_en ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _23630_ (.RESET_B(net6584),
    .D(_00127_),
    .Q(\soc_inst.spi_inst.busy ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23631_ (.RESET_B(net6576),
    .D(_00089_),
    .Q(\soc_inst.i2c_inst.clk_cnt[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23632_ (.RESET_B(net6576),
    .D(_00090_),
    .Q(\soc_inst.i2c_inst.clk_cnt[1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23633_ (.RESET_B(net6576),
    .D(net1232),
    .Q(\soc_inst.i2c_inst.clk_cnt[2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23634_ (.RESET_B(net6576),
    .D(_00092_),
    .Q(\soc_inst.i2c_inst.clk_cnt[3] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23635_ (.RESET_B(net6571),
    .D(_00093_),
    .Q(\soc_inst.i2c_inst.clk_cnt[4] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _23636_ (.RESET_B(net6571),
    .D(_00094_),
    .Q(\soc_inst.i2c_inst.clk_cnt[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23637_ (.RESET_B(net6571),
    .D(net2531),
    .Q(\soc_inst.i2c_inst.clk_cnt[6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _23638_ (.RESET_B(net6571),
    .D(_00096_),
    .Q(\soc_inst.i2c_inst.clk_cnt[7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _23639_ (.RESET_B(net6580),
    .D(net980),
    .Q(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23640_ (.RESET_B(net6570),
    .D(_00389_),
    .Q(\soc_inst.i2c_inst.ctrl_reg[2] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23641_ (.RESET_B(net6576),
    .D(_00390_),
    .Q(\soc_inst.i2c_inst.ack_enable ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23642_ (.RESET_B(net6569),
    .D(_00391_),
    .Q(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _23643_ (.RESET_B(net6576),
    .D(net113),
    .Q(\soc_inst.i2c_inst.arb_lost ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23644_ (.RESET_B(net6583),
    .D(_11836_[0]),
    .Q(\soc_inst.i2c_inst.start_pending ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _23645_ (.RESET_B(net6570),
    .D(net2251),
    .Q(\soc_inst.i2c_inst.data_reg[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _23646_ (.RESET_B(net6569),
    .D(net1719),
    .Q(\soc_inst.i2c_inst.data_reg[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23647_ (.RESET_B(net6567),
    .D(net1837),
    .Q(\soc_inst.i2c_inst.data_reg[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23648_ (.RESET_B(net6567),
    .D(net2018),
    .Q(\soc_inst.i2c_inst.data_reg[3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23649_ (.RESET_B(net6567),
    .D(net2087),
    .Q(\soc_inst.i2c_inst.data_reg[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23650_ (.RESET_B(net6568),
    .D(net2200),
    .Q(\soc_inst.i2c_inst.data_reg[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _23651_ (.RESET_B(net6568),
    .D(net1913),
    .Q(\soc_inst.i2c_inst.data_reg[6] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23652_ (.RESET_B(net6570),
    .D(net2050),
    .Q(\soc_inst.i2c_inst.data_reg[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23653_ (.RESET_B(net6570),
    .D(net1935),
    .Q(_00226_),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23654_ (.RESET_B(net6570),
    .D(net2307),
    .Q(_00227_),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23655_ (.RESET_B(net6570),
    .D(_00395_),
    .Q(_00228_),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _23656_ (.RESET_B(net6571),
    .D(_00396_),
    .Q(_00229_),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _23657_ (.RESET_B(net6567),
    .D(_00397_),
    .Q(_00230_),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23658_ (.RESET_B(net6567),
    .D(_00398_),
    .Q(\soc_inst.i2c_inst.prescale_reg[5] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23659_ (.RESET_B(net6571),
    .D(_00399_),
    .Q(\soc_inst.i2c_inst.prescale_reg[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23660_ (.RESET_B(net6570),
    .D(_00400_),
    .Q(_00231_),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23661_ (.RESET_B(net6576),
    .D(net595),
    .Q(\soc_inst.i2c_inst.restart_pending ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23662_ (.RESET_B(net6571),
    .D(_02599_),
    .Q(\soc_inst.i2c_inst.shift_reg[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _23663_ (.RESET_B(net6568),
    .D(_02600_),
    .Q(\soc_inst.i2c_inst.shift_reg[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _23664_ (.RESET_B(net6567),
    .D(_02601_),
    .Q(\soc_inst.i2c_inst.shift_reg[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23665_ (.RESET_B(net6567),
    .D(_02602_),
    .Q(\soc_inst.i2c_inst.shift_reg[3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23666_ (.RESET_B(net6567),
    .D(_02603_),
    .Q(\soc_inst.i2c_inst.shift_reg[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23667_ (.RESET_B(net6568),
    .D(_02604_),
    .Q(\soc_inst.i2c_inst.shift_reg[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23668_ (.RESET_B(net6568),
    .D(_02605_),
    .Q(\soc_inst.i2c_inst.shift_reg[6] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _23669_ (.RESET_B(net6575),
    .D(_02606_),
    .Q(\soc_inst.i2c_inst.shift_reg[7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _23670_ (.RESET_B(net6577),
    .D(net3122),
    .Q(\soc_inst.i2c_inst.bit_cnt[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _23671_ (.RESET_B(net6577),
    .D(_00402_),
    .Q(\soc_inst.i2c_inst.bit_cnt[1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _23672_ (.RESET_B(net6577),
    .D(net1015),
    .Q(\soc_inst.i2c_inst.bit_cnt[2] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _23673_ (.RESET_B(net6578),
    .D(_00404_),
    .Q(\soc_inst.i2c_inst.bit_cnt[3] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _23674_ (.RESET_B(net6577),
    .D(_00405_),
    .Q(_00232_),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _23675_ (.RESET_B(net6576),
    .D(net1567),
    .Q(\soc_inst.i2c_inst.stop_pending ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23676_ (.RESET_B(net6578),
    .D(_00406_),
    .Q(_00233_),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23677_ (.RESET_B(net6569),
    .D(_00106_),
    .Q(\soc_inst.i2c_inst.transfer_done ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _23678_ (.RESET_B(net6572),
    .D(_00111_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23679_ (.RESET_B(net6572),
    .D(_00118_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23680_ (.RESET_B(net6572),
    .D(net2640),
    .Q(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _23681_ (.RESET_B(net6572),
    .D(_00120_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _23682_ (.RESET_B(net6550),
    .D(net2527),
    .Q(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _23683_ (.RESET_B(net6551),
    .D(_00122_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _23684_ (.RESET_B(net6552),
    .D(_00123_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _23685_ (.RESET_B(net6561),
    .D(net2931),
    .Q(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _23686_ (.RESET_B(net6561),
    .D(_00125_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _23687_ (.RESET_B(net6561),
    .D(_00126_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _23688_ (.RESET_B(net6555),
    .D(net2473),
    .Q(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _23689_ (.RESET_B(net6555),
    .D(_00113_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23690_ (.RESET_B(net6554),
    .D(_00114_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23691_ (.RESET_B(net6554),
    .D(_00115_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23692_ (.RESET_B(net6554),
    .D(_00116_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _23693_ (.RESET_B(net6555),
    .D(_00117_),
    .Q(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _23694_ (.RESET_B(net6590),
    .D(net2539),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[0] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _23695_ (.RESET_B(net6590),
    .D(net2323),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _23696_ (.RESET_B(net6572),
    .D(net2144),
    .Q(_00234_),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23697_ (.RESET_B(net6573),
    .D(net2182),
    .Q(_00235_),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _23698_ (.RESET_B(net6572),
    .D(_00411_),
    .Q(_00236_),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _23699_ (.RESET_B(net6573),
    .D(_00412_),
    .Q(_00237_),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _23700_ (.RESET_B(net6550),
    .D(_00413_),
    .Q(_00238_),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _23701_ (.RESET_B(net6551),
    .D(_00414_),
    .Q(_00239_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _23702_ (.RESET_B(net6562),
    .D(_00415_),
    .Q(_00240_),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _23703_ (.RESET_B(net6562),
    .D(_00416_),
    .Q(_00241_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _23704_ (.RESET_B(net6561),
    .D(_00417_),
    .Q(_00242_),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _23705_ (.RESET_B(net6562),
    .D(_00418_),
    .Q(_00243_),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _23706_ (.RESET_B(net6555),
    .D(_00419_),
    .Q(_00244_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23707_ (.RESET_B(net6554),
    .D(net1679),
    .Q(_00245_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _23708_ (.RESET_B(net6559),
    .D(_00421_),
    .Q(_00246_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _23709_ (.RESET_B(net6559),
    .D(_00422_),
    .Q(_00247_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _23710_ (.RESET_B(net6559),
    .D(_00423_),
    .Q(_00248_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23711_ (.RESET_B(net6559),
    .D(net2056),
    .Q(_00249_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _23712_ (.RESET_B(net6678),
    .D(_00023_),
    .Q(\soc_inst.cpu_core.csr_file.timer_interrupt ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _23713_ (.RESET_B(net6587),
    .D(net2025),
    .Q(\soc_inst.spi_inst.len_sel[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23714_ (.RESET_B(net6587),
    .D(_00426_),
    .Q(\soc_inst.spi_inst.len_sel[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23715_ (.RESET_B(net6580),
    .D(net93),
    .Q(\soc_inst.gpio_inst.gpio_sync2[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _23716_ (.RESET_B(net6589),
    .D(net81),
    .Q(\soc_inst.gpio_inst.gpio_sync2[1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23717_ (.RESET_B(net6595),
    .D(net83),
    .Q(\soc_inst.gpio_inst.gpio_sync2[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _23718_ (.RESET_B(net6595),
    .D(net88),
    .Q(\soc_inst.gpio_inst.gpio_sync2[3] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _23719_ (.RESET_B(net6595),
    .D(net87),
    .Q(\soc_inst.gpio_inst.gpio_sync2[4] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _23720_ (.RESET_B(net6590),
    .D(net84),
    .Q(\soc_inst.gpio_inst.gpio_sync2[5] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _23721_ (.RESET_B(net6579),
    .D(net86),
    .Q(\soc_inst.gpio_inst.gpio_sync2[6] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _23722_ (.RESET_B(net6843),
    .D(_00427_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _23723_ (.RESET_B(net6840),
    .D(_00428_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _23724_ (.RESET_B(net6835),
    .D(_00429_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][2] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _23725_ (.RESET_B(net6850),
    .D(_00430_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][3] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _23726_ (.RESET_B(net6879),
    .D(_00431_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][4] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _23727_ (.RESET_B(net6952),
    .D(_00432_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _23728_ (.RESET_B(net6906),
    .D(_00433_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][6] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _23729_ (.RESET_B(net6928),
    .D(_00434_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][7] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _23730_ (.RESET_B(net6897),
    .D(_00435_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][8] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _23731_ (.RESET_B(net6957),
    .D(_00436_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][9] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23732_ (.RESET_B(net6965),
    .D(_00437_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _23733_ (.RESET_B(net6894),
    .D(_00438_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][11] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _23734_ (.RESET_B(net6949),
    .D(_00439_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _23735_ (.RESET_B(net6936),
    .D(_00440_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][13] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _23736_ (.RESET_B(net6808),
    .D(_00441_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][14] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _23737_ (.RESET_B(net6942),
    .D(_00442_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _23738_ (.RESET_B(net6922),
    .D(_00443_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _23739_ (.RESET_B(net6865),
    .D(_00444_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _23740_ (.RESET_B(net6934),
    .D(_00445_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][18] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _23741_ (.RESET_B(net6872),
    .D(_00446_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][19] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _23742_ (.RESET_B(net6968),
    .D(_00447_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _23743_ (.RESET_B(net6911),
    .D(_00448_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][21] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _23744_ (.RESET_B(net6823),
    .D(_00449_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_2 _23745_ (.RESET_B(net6980),
    .D(_00450_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _23746_ (.RESET_B(net6859),
    .D(_00451_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][24] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _23747_ (.RESET_B(net6810),
    .D(_00452_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _23748_ (.RESET_B(net6918),
    .D(_00453_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][26] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _23749_ (.RESET_B(net6828),
    .D(_00454_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][27] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _23750_ (.RESET_B(net6875),
    .D(_00455_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _23751_ (.RESET_B(net6861),
    .D(_00456_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][29] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _23752_ (.RESET_B(net6976),
    .D(_00457_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23753_ (.RESET_B(net6953),
    .D(_00458_),
    .Q(\soc_inst.cpu_core.register_file.registers[31][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _23754_ (.RESET_B(net6581),
    .D(net815),
    .Q(\soc_inst.gpio_bidir_oe [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23755_ (.RESET_B(net6581),
    .D(net446),
    .Q(\soc_inst.gpio_bidir_out [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23756_ (.RESET_B(net6579),
    .D(net2298),
    .Q(\soc_inst.gpio_inst.gpio_out[0] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23757_ (.RESET_B(net6590),
    .D(net1988),
    .Q(\soc_inst.gpio_inst.gpio_out[1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23758_ (.RESET_B(net6579),
    .D(_00463_),
    .Q(\soc_inst.gpio_inst.gpio_out[2] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _23759_ (.RESET_B(net6582),
    .D(_00464_),
    .Q(\soc_inst.gpio_inst.gpio_out[3] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _23760_ (.RESET_B(net6574),
    .D(net1387),
    .Q(\soc_inst.gpio_inst.gpio_out[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _23761_ (.RESET_B(net6581),
    .D(net783),
    .Q(\soc_inst.gpio_inst.gpio_out[5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23762_ (.RESET_B(net6581),
    .D(net13),
    .Q(\soc_inst.gpio_inst.gpio_sync1[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _23763_ (.RESET_B(net6589),
    .D(net2),
    .Q(\soc_inst.gpio_inst.gpio_sync1[1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23764_ (.RESET_B(net6595),
    .D(net3),
    .Q(\soc_inst.gpio_inst.gpio_sync1[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _23765_ (.RESET_B(net6591),
    .D(net4),
    .Q(\soc_inst.gpio_inst.gpio_sync1[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23766_ (.RESET_B(net6595),
    .D(net5),
    .Q(\soc_inst.gpio_inst.gpio_sync1[4] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _23767_ (.RESET_B(net6590),
    .D(net6),
    .Q(\soc_inst.gpio_inst.gpio_sync1[5] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _23768_ (.RESET_B(net6581),
    .D(net7),
    .Q(\soc_inst.gpio_inst.gpio_sync1[6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _23769_ (.RESET_B(net6640),
    .D(_00088_),
    .Q(\soc_inst.cpu_core.csr_file.external_interrupt ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _23770_ (.RESET_B(net6579),
    .D(_00467_),
    .Q(\soc_inst.gpio_inst.int_en_reg[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23771_ (.RESET_B(net6579),
    .D(net2467),
    .Q(\soc_inst.gpio_inst.int_en_reg[1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23772_ (.RESET_B(net6591),
    .D(net2899),
    .Q(\soc_inst.gpio_inst.int_en_reg[2] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23773_ (.RESET_B(net6592),
    .D(_00470_),
    .Q(\soc_inst.gpio_inst.int_en_reg[3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _23774_ (.RESET_B(net6592),
    .D(_00471_),
    .Q(\soc_inst.gpio_inst.int_en_reg[4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _23775_ (.RESET_B(net6589),
    .D(_00472_),
    .Q(\soc_inst.gpio_inst.int_en_reg[5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _23776_ (.RESET_B(net6580),
    .D(_00473_),
    .Q(\soc_inst.gpio_inst.int_en_reg[6] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _23777_ (.RESET_B(net6644),
    .D(_00474_),
    .Q(\soc_inst.mem_ctrl.spi_data_len[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _23778_ (.RESET_B(net6684),
    .D(_00475_),
    .Q(\soc_inst.mem_ctrl.spi_data_len[4] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _23779_ (.RESET_B(net6644),
    .D(_00476_),
    .Q(\soc_inst.mem_ctrl.spi_data_len[5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _23780_ (.RESET_B(net6643),
    .D(net1813),
    .Q(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _23781_ (.RESET_B(net6622),
    .D(_00478_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _23782_ (.RESET_B(net6624),
    .D(_00479_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23783_ (.RESET_B(net6624),
    .D(net319),
    .Q(\soc_inst.mem_ctrl.spi_data_in[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23784_ (.RESET_B(net6616),
    .D(_00481_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[3] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_2 _23785_ (.RESET_B(net6605),
    .D(_00482_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[4] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _23786_ (.RESET_B(net6605),
    .D(_00483_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _23787_ (.RESET_B(net6622),
    .D(net419),
    .Q(\soc_inst.mem_ctrl.spi_data_in[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23788_ (.RESET_B(net6621),
    .D(net267),
    .Q(\soc_inst.mem_ctrl.spi_data_in[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _23789_ (.RESET_B(net6614),
    .D(_00486_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[8] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _23790_ (.RESET_B(net6614),
    .D(_00487_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[9] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _23791_ (.RESET_B(net6615),
    .D(net1100),
    .Q(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_2 _23792_ (.RESET_B(net6613),
    .D(_00489_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[11] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_2 _23793_ (.RESET_B(net6614),
    .D(_00490_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[12] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _23794_ (.RESET_B(net6605),
    .D(_00491_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[13] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _23795_ (.RESET_B(net6605),
    .D(net965),
    .Q(\soc_inst.mem_ctrl.spi_data_in[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _23796_ (.RESET_B(net6615),
    .D(net867),
    .Q(\soc_inst.mem_ctrl.spi_data_in[15] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _23797_ (.RESET_B(net6609),
    .D(net353),
    .Q(\soc_inst.mem_ctrl.spi_data_in[16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _23798_ (.RESET_B(net6609),
    .D(_00495_),
    .Q(\soc_inst.mem_ctrl.spi_data_in[17] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _23799_ (.RESET_B(net6609),
    .D(net310),
    .Q(\soc_inst.mem_ctrl.spi_data_in[18] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _23800_ (.RESET_B(net6611),
    .D(net380),
    .Q(\soc_inst.mem_ctrl.spi_data_in[19] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _23801_ (.RESET_B(net6609),
    .D(net702),
    .Q(\soc_inst.mem_ctrl.spi_data_in[20] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _23802_ (.RESET_B(net6609),
    .D(net432),
    .Q(\soc_inst.mem_ctrl.spi_data_in[21] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _23803_ (.RESET_B(net6609),
    .D(net899),
    .Q(\soc_inst.mem_ctrl.spi_data_in[22] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _23804_ (.RESET_B(net6611),
    .D(net343),
    .Q(\soc_inst.mem_ctrl.spi_data_in[23] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _23805_ (.RESET_B(net6632),
    .D(net306),
    .Q(\soc_inst.mem_ctrl.spi_data_in[24] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23806_ (.RESET_B(net6632),
    .D(net384),
    .Q(\soc_inst.mem_ctrl.spi_data_in[25] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23807_ (.RESET_B(net6642),
    .D(net203),
    .Q(\soc_inst.mem_ctrl.spi_data_in[26] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23808_ (.RESET_B(net6632),
    .D(net333),
    .Q(\soc_inst.mem_ctrl.spi_data_in[27] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23809_ (.RESET_B(net6632),
    .D(net357),
    .Q(\soc_inst.mem_ctrl.spi_data_in[28] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23810_ (.RESET_B(net6635),
    .D(net351),
    .Q(\soc_inst.mem_ctrl.spi_data_in[29] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23811_ (.RESET_B(net6635),
    .D(net182),
    .Q(\soc_inst.mem_ctrl.spi_data_in[30] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23812_ (.RESET_B(net6634),
    .D(net166),
    .Q(\soc_inst.mem_ctrl.spi_data_in[31] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23813_ (.RESET_B(net6646),
    .D(_00108_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.stop ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _23814_ (.RESET_B(net6721),
    .D(net621),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _23815_ (.RESET_B(net6715),
    .D(net575),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23816_ (.RESET_B(net6721),
    .D(net442),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _23817_ (.RESET_B(net6738),
    .D(net787),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _23818_ (.RESET_B(net6718),
    .D(net478),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _23819_ (.RESET_B(net6702),
    .D(_00058_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[0] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _23820_ (.RESET_B(net6739),
    .D(_00059_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[1] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _23821_ (.RESET_B(net6742),
    .D(_00060_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[2] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _23822_ (.RESET_B(net6737),
    .D(_00061_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[3] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _23823_ (.RESET_B(net6701),
    .D(_00062_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[4] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _23824_ (.RESET_B(net6580),
    .D(net242),
    .Q(\soc_inst.i2c_inst.ack_received ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23825_ (.RESET_B(net6737),
    .D(_00027_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23826_ (.RESET_B(net6700),
    .D(_00038_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _23827_ (.RESET_B(net6737),
    .D(_00049_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23828_ (.RESET_B(net6737),
    .D(_00051_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23829_ (.RESET_B(net6699),
    .D(_00052_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _23830_ (.RESET_B(net6679),
    .D(_00053_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _23831_ (.RESET_B(net6702),
    .D(_00054_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23832_ (.RESET_B(net6718),
    .D(_00055_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _23833_ (.RESET_B(net6679),
    .D(_00056_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _23834_ (.RESET_B(net6738),
    .D(_00057_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[9] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _23835_ (.RESET_B(net6720),
    .D(_00028_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[10] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _23836_ (.RESET_B(net6718),
    .D(_00029_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _23837_ (.RESET_B(net6720),
    .D(_00030_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[12] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _23838_ (.RESET_B(net6664),
    .D(_00031_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[13] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _23839_ (.RESET_B(net6662),
    .D(_00032_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[14] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _23840_ (.RESET_B(net6662),
    .D(_00033_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _23841_ (.RESET_B(net6711),
    .D(_00034_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[16] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _23842_ (.RESET_B(net6674),
    .D(_00035_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[17] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _23843_ (.RESET_B(net6710),
    .D(_00036_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[18] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _23844_ (.RESET_B(net6661),
    .D(_00037_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[19] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _23845_ (.RESET_B(net6661),
    .D(_00039_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[20] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _23846_ (.RESET_B(net6709),
    .D(_00040_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[21] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _23847_ (.RESET_B(net6675),
    .D(_00041_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[22] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _23848_ (.RESET_B(net6674),
    .D(_00042_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _23849_ (.RESET_B(net6662),
    .D(_00043_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[24] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _23850_ (.RESET_B(net6668),
    .D(_00044_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[25] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _23851_ (.RESET_B(net6662),
    .D(_00045_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _23852_ (.RESET_B(net6663),
    .D(_00046_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[27] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _23853_ (.RESET_B(net6663),
    .D(_00047_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[28] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _23854_ (.RESET_B(net6664),
    .D(_00048_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[29] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _23855_ (.RESET_B(net6673),
    .D(_00050_),
    .Q(\soc_inst.cpu_core.csr_file.mcause[30] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _23856_ (.RESET_B(net6700),
    .D(_00083_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _23857_ (.RESET_B(net6739),
    .D(_00084_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _23858_ (.RESET_B(net6737),
    .D(_00085_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _23859_ (.RESET_B(net6737),
    .D(net3102),
    .Q(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _23860_ (.RESET_B(net6700),
    .D(_00087_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _23861_ (.RESET_B(net6699),
    .D(_00516_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _23862_ (.RESET_B(net6702),
    .D(net2151),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _23863_ (.RESET_B(net6742),
    .D(_00518_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _23864_ (.RESET_B(net6737),
    .D(_00519_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[3] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _23865_ (.RESET_B(net6703),
    .D(_00520_),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[4] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _23866_ (.RESET_B(net6701),
    .D(_00521_),
    .Q(\soc_inst.core_instr_addr[0] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _23867_ (.RESET_B(net6739),
    .D(_00522_),
    .Q(\soc_inst.core_instr_addr[1] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _23868_ (.RESET_B(net6739),
    .D(_00523_),
    .Q(\soc_inst.core_instr_addr[2] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _23869_ (.RESET_B(net6701),
    .D(_00524_),
    .Q(\soc_inst.core_instr_addr[3] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _23870_ (.RESET_B(net6701),
    .D(net2960),
    .Q(\soc_inst.core_instr_addr[4] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _23871_ (.RESET_B(net6741),
    .D(_00526_),
    .Q(\soc_inst.core_instr_addr[5] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _23872_ (.RESET_B(net6740),
    .D(_00527_),
    .Q(\soc_inst.core_instr_addr[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _23873_ (.RESET_B(net6740),
    .D(_00528_),
    .Q(\soc_inst.core_instr_addr[7] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _23874_ (.RESET_B(net6719),
    .D(_00529_),
    .Q(\soc_inst.core_instr_addr[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _23875_ (.RESET_B(net6741),
    .D(net3045),
    .Q(\soc_inst.core_instr_addr[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _23876_ (.RESET_B(net6729),
    .D(net3011),
    .Q(\soc_inst.core_instr_addr[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _23877_ (.RESET_B(net6729),
    .D(net3226),
    .Q(\soc_inst.core_instr_addr[11] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _23878_ (.RESET_B(net6719),
    .D(_00533_),
    .Q(\soc_inst.core_instr_addr[12] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _23879_ (.RESET_B(net6717),
    .D(_00534_),
    .Q(\soc_inst.core_instr_addr[13] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _23880_ (.RESET_B(net6717),
    .D(_00535_),
    .Q(\soc_inst.core_instr_addr[14] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_2 _23881_ (.RESET_B(net6720),
    .D(net2705),
    .Q(\soc_inst.core_instr_addr[15] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _23882_ (.RESET_B(net6723),
    .D(net3139),
    .Q(\soc_inst.core_instr_addr[16] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _23883_ (.RESET_B(net6714),
    .D(_00538_),
    .Q(\soc_inst.core_instr_addr[17] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _23884_ (.RESET_B(net6722),
    .D(_00539_),
    .Q(\soc_inst.core_instr_addr[18] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _23885_ (.RESET_B(net6724),
    .D(_00540_),
    .Q(\soc_inst.core_instr_addr[19] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _23886_ (.RESET_B(net6723),
    .D(_00541_),
    .Q(\soc_inst.core_instr_addr[20] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _23887_ (.RESET_B(net6716),
    .D(_00542_),
    .Q(\soc_inst.core_instr_addr[21] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _23888_ (.RESET_B(net6710),
    .D(_00543_),
    .Q(\soc_inst.core_instr_addr[22] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_2 _23889_ (.RESET_B(net6716),
    .D(_00544_),
    .Q(\soc_inst.core_instr_addr[23] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _23890_ (.RESET_B(net6577),
    .D(net3218),
    .Q(\soc_inst.i2c_inst.state[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _23891_ (.RESET_B(net6577),
    .D(_00546_),
    .Q(\soc_inst.i2c_inst.state[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _23892_ (.RESET_B(net6577),
    .D(_00547_),
    .Q(\soc_inst.i2c_inst.state[2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _23893_ (.RESET_B(net6577),
    .D(_00548_),
    .Q(\soc_inst.i2c_inst.state[3] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _23894_ (.RESET_B(net6685),
    .D(net2950),
    .Q(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23895_ (.RESET_B(net6685),
    .D(net2905),
    .Q(\soc_inst.mem_ctrl.spi_addr[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23896_ (.RESET_B(net6686),
    .D(net3032),
    .Q(\soc_inst.mem_ctrl.spi_addr[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23897_ (.RESET_B(net6685),
    .D(net2832),
    .Q(\soc_inst.mem_ctrl.spi_addr[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23898_ (.RESET_B(net6686),
    .D(_00553_),
    .Q(\soc_inst.mem_ctrl.spi_addr[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23899_ (.RESET_B(net6686),
    .D(_00554_),
    .Q(\soc_inst.mem_ctrl.spi_addr[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _23900_ (.RESET_B(net6686),
    .D(_00555_),
    .Q(\soc_inst.mem_ctrl.spi_addr[6] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23901_ (.RESET_B(net6686),
    .D(_00556_),
    .Q(\soc_inst.mem_ctrl.spi_addr[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23902_ (.RESET_B(net6669),
    .D(_00557_),
    .Q(\soc_inst.mem_ctrl.spi_addr[8] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _23903_ (.RESET_B(net6667),
    .D(_00558_),
    .Q(\soc_inst.mem_ctrl.spi_addr[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23904_ (.RESET_B(net6669),
    .D(net2955),
    .Q(\soc_inst.mem_ctrl.spi_addr[10] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _23905_ (.RESET_B(net6667),
    .D(net3141),
    .Q(\soc_inst.mem_ctrl.spi_addr[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23906_ (.RESET_B(net6626),
    .D(net2821),
    .Q(\soc_inst.mem_ctrl.spi_addr[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23907_ (.RESET_B(net6626),
    .D(net3083),
    .Q(\soc_inst.mem_ctrl.spi_addr[13] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _23908_ (.RESET_B(net6624),
    .D(net2866),
    .Q(\soc_inst.mem_ctrl.spi_addr[14] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_2 _23909_ (.RESET_B(net6668),
    .D(net2658),
    .Q(\soc_inst.mem_ctrl.spi_addr[15] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _23910_ (.RESET_B(net6625),
    .D(_00565_),
    .Q(\soc_inst.mem_ctrl.spi_addr[16] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23911_ (.RESET_B(net6625),
    .D(_00566_),
    .Q(\soc_inst.mem_ctrl.spi_addr[17] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23912_ (.RESET_B(net6625),
    .D(_00567_),
    .Q(\soc_inst.mem_ctrl.spi_addr[18] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23913_ (.RESET_B(net6624),
    .D(net3055),
    .Q(\soc_inst.mem_ctrl.spi_addr[19] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _23914_ (.RESET_B(net6666),
    .D(net3097),
    .Q(\soc_inst.mem_ctrl.spi_addr[20] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _23915_ (.RESET_B(net6624),
    .D(_00570_),
    .Q(\soc_inst.mem_ctrl.spi_addr[21] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _23916_ (.RESET_B(net6666),
    .D(net3079),
    .Q(\soc_inst.mem_ctrl.spi_addr[22] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23917_ (.RESET_B(net6667),
    .D(net2798),
    .Q(\soc_inst.mem_ctrl.spi_addr[23] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23918_ (.RESET_B(net6694),
    .D(_00573_),
    .Q(\soc_inst.core_instr_data[0] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _23919_ (.RESET_B(net6693),
    .D(_00574_),
    .Q(\soc_inst.core_instr_data[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _23920_ (.RESET_B(net6704),
    .D(_00575_),
    .Q(\soc_inst.core_instr_data[2] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23921_ (.RESET_B(net6696),
    .D(_00576_),
    .Q(\soc_inst.core_instr_data[3] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23922_ (.RESET_B(net6693),
    .D(_00577_),
    .Q(\soc_inst.core_instr_data[4] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _23923_ (.RESET_B(net6705),
    .D(_00578_),
    .Q(\soc_inst.core_instr_data[5] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _23924_ (.RESET_B(net6695),
    .D(_00579_),
    .Q(\soc_inst.core_instr_data[6] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _23925_ (.RESET_B(net6696),
    .D(_00580_),
    .Q(\soc_inst.core_instr_data[7] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _23926_ (.RESET_B(net6704),
    .D(_00581_),
    .Q(\soc_inst.core_instr_data[8] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _23927_ (.RESET_B(net6704),
    .D(_00582_),
    .Q(\soc_inst.core_instr_data[9] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23928_ (.RESET_B(net6704),
    .D(_00583_),
    .Q(\soc_inst.core_instr_data[10] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _23929_ (.RESET_B(net6705),
    .D(_00584_),
    .Q(\soc_inst.core_instr_data[11] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _23930_ (.RESET_B(net6707),
    .D(_00585_),
    .Q(\soc_inst.core_instr_data[12] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _23931_ (.RESET_B(net6705),
    .D(_00586_),
    .Q(\soc_inst.core_instr_data[13] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _23932_ (.RESET_B(net6704),
    .D(_00587_),
    .Q(\soc_inst.core_instr_data[14] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23933_ (.RESET_B(net6707),
    .D(_00588_),
    .Q(\soc_inst.core_instr_data[15] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23934_ (.RESET_B(net6706),
    .D(net2668),
    .Q(\soc_inst.core_instr_data[16] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _23935_ (.RESET_B(net6706),
    .D(net2697),
    .Q(\soc_inst.core_instr_data[17] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _23936_ (.RESET_B(net6706),
    .D(_00591_),
    .Q(\soc_inst.core_instr_data[18] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _23937_ (.RESET_B(net6706),
    .D(net2646),
    .Q(\soc_inst.core_instr_data[19] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _23938_ (.RESET_B(net6696),
    .D(net2868),
    .Q(\soc_inst.core_instr_data[20] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _23939_ (.RESET_B(net6694),
    .D(net2542),
    .Q(\soc_inst.core_instr_data[21] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _23940_ (.RESET_B(net6704),
    .D(net2403),
    .Q(\soc_inst.core_instr_data[22] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _23941_ (.RESET_B(net6707),
    .D(net2454),
    .Q(\soc_inst.core_instr_data[23] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _23942_ (.RESET_B(net6696),
    .D(net2475),
    .Q(\soc_inst.core_instr_data[24] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _23943_ (.RESET_B(net6705),
    .D(net2437),
    .Q(\soc_inst.core_instr_data[25] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _23944_ (.RESET_B(net6706),
    .D(net2550),
    .Q(\soc_inst.core_instr_data[26] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23945_ (.RESET_B(net6705),
    .D(net2579),
    .Q(\soc_inst.core_instr_data[27] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _23946_ (.RESET_B(net6705),
    .D(net2577),
    .Q(\soc_inst.core_instr_data[28] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23947_ (.RESET_B(net6705),
    .D(net2504),
    .Q(\soc_inst.core_instr_data[29] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23948_ (.RESET_B(net6694),
    .D(net1849),
    .Q(\soc_inst.core_instr_data[30] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23949_ (.RESET_B(net6694),
    .D(net1447),
    .Q(\soc_inst.core_instr_data[31] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23950_ (.RESET_B(net6698),
    .D(_00605_),
    .Q(\soc_inst.core_mem_rdata[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _23951_ (.RESET_B(net6643),
    .D(net1986),
    .Q(\soc_inst.core_mem_rdata[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _23952_ (.RESET_B(net6644),
    .D(net1968),
    .Q(\soc_inst.core_mem_rdata[2] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _23953_ (.RESET_B(net6643),
    .D(_00608_),
    .Q(\soc_inst.core_mem_rdata[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _23954_ (.RESET_B(net6684),
    .D(_00609_),
    .Q(\soc_inst.core_mem_rdata[4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _23955_ (.RESET_B(net6687),
    .D(_00610_),
    .Q(\soc_inst.core_mem_rdata[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _23956_ (.RESET_B(net6644),
    .D(_00611_),
    .Q(\soc_inst.core_mem_rdata[6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _23957_ (.RESET_B(net6667),
    .D(_00612_),
    .Q(\soc_inst.core_mem_rdata[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23958_ (.RESET_B(net6685),
    .D(net2138),
    .Q(\soc_inst.core_mem_rdata[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23959_ (.RESET_B(net6685),
    .D(_00614_),
    .Q(\soc_inst.core_mem_rdata[9] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23960_ (.RESET_B(net6625),
    .D(_00615_),
    .Q(\soc_inst.core_mem_rdata[10] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23961_ (.RESET_B(net6621),
    .D(_00616_),
    .Q(\soc_inst.core_mem_rdata[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _23962_ (.RESET_B(net6621),
    .D(_00617_),
    .Q(\soc_inst.core_mem_rdata[12] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _23963_ (.RESET_B(net6659),
    .D(_00618_),
    .Q(\soc_inst.core_mem_rdata[13] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23964_ (.RESET_B(net6659),
    .D(_00619_),
    .Q(\soc_inst.core_mem_rdata[14] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _23965_ (.RESET_B(net6659),
    .D(_00620_),
    .Q(\soc_inst.core_mem_rdata[15] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _23966_ (.RESET_B(net6620),
    .D(net1999),
    .Q(\soc_inst.core_mem_rdata[16] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _23967_ (.RESET_B(net6624),
    .D(net2205),
    .Q(\soc_inst.core_mem_rdata[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23968_ (.RESET_B(net6666),
    .D(net2213),
    .Q(\soc_inst.core_mem_rdata[18] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23969_ (.RESET_B(net6624),
    .D(net2191),
    .Q(\soc_inst.core_mem_rdata[19] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23970_ (.RESET_B(net6686),
    .D(net1381),
    .Q(\soc_inst.core_mem_rdata[20] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _23971_ (.RESET_B(net6686),
    .D(net1021),
    .Q(\soc_inst.core_mem_rdata[21] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _23972_ (.RESET_B(net6624),
    .D(net2061),
    .Q(\soc_inst.core_mem_rdata[22] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23973_ (.RESET_B(net6687),
    .D(net1189),
    .Q(\soc_inst.core_mem_rdata[23] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _23974_ (.RESET_B(net6643),
    .D(net1225),
    .Q(\soc_inst.core_mem_rdata[24] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23975_ (.RESET_B(net6626),
    .D(net1959),
    .Q(\soc_inst.core_mem_rdata[25] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _23976_ (.RESET_B(net6643),
    .D(net2334),
    .Q(\soc_inst.core_mem_rdata[26] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _23977_ (.RESET_B(net6643),
    .D(net2380),
    .Q(\soc_inst.core_mem_rdata[27] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _23978_ (.RESET_B(net6643),
    .D(net2316),
    .Q(\soc_inst.core_mem_rdata[28] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _23979_ (.RESET_B(net6698),
    .D(net1149),
    .Q(\soc_inst.core_mem_rdata[29] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _23980_ (.RESET_B(net6684),
    .D(net1509),
    .Q(\soc_inst.core_mem_rdata[30] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _23981_ (.RESET_B(net6698),
    .D(net1120),
    .Q(\soc_inst.core_mem_rdata[31] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _23982_ (.RESET_B(net6642),
    .D(net1439),
    .Q(\soc_inst.mem_ctrl.spi_read_enable ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23983_ (.RESET_B(net6644),
    .D(_00638_),
    .Q(\soc_inst.cpu_core.i_mem_ready ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _23984_ (.RESET_B(net6644),
    .D(net3151),
    .Q(\soc_inst.mem_ctrl.instr_ready_reg ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _23985_ (.RESET_B(net6694),
    .D(net690),
    .Q(\soc_inst.mem_ctrl.next_instr_data[0] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _23986_ (.RESET_B(net6693),
    .D(net763),
    .Q(\soc_inst.mem_ctrl.next_instr_data[1] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _23987_ (.RESET_B(net6695),
    .D(net1115),
    .Q(\soc_inst.mem_ctrl.next_instr_data[2] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _23988_ (.RESET_B(net6695),
    .D(net469),
    .Q(\soc_inst.mem_ctrl.next_instr_data[3] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _23989_ (.RESET_B(net6693),
    .D(net616),
    .Q(\soc_inst.mem_ctrl.next_instr_data[4] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _23990_ (.RESET_B(net6689),
    .D(net823),
    .Q(\soc_inst.mem_ctrl.next_instr_data[5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _23991_ (.RESET_B(net6691),
    .D(net775),
    .Q(\soc_inst.mem_ctrl.next_instr_data[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _23992_ (.RESET_B(net6695),
    .D(net946),
    .Q(\soc_inst.mem_ctrl.next_instr_data[7] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _23993_ (.RESET_B(net6692),
    .D(net559),
    .Q(\soc_inst.mem_ctrl.next_instr_data[8] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _23994_ (.RESET_B(net6695),
    .D(net1227),
    .Q(\soc_inst.mem_ctrl.next_instr_data[9] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _23995_ (.RESET_B(net6691),
    .D(net1010),
    .Q(\soc_inst.mem_ctrl.next_instr_data[10] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _23996_ (.RESET_B(net6691),
    .D(net656),
    .Q(\soc_inst.mem_ctrl.next_instr_data[11] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _23997_ (.RESET_B(net6696),
    .D(net1066),
    .Q(\soc_inst.mem_ctrl.next_instr_data[12] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _23998_ (.RESET_B(net6689),
    .D(net1133),
    .Q(\soc_inst.mem_ctrl.next_instr_data[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _23999_ (.RESET_B(net6690),
    .D(net643),
    .Q(\soc_inst.mem_ctrl.next_instr_data[14] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _24000_ (.RESET_B(net6690),
    .D(net796),
    .Q(\soc_inst.mem_ctrl.next_instr_data[15] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _24001_ (.RESET_B(net6693),
    .D(net884),
    .Q(\soc_inst.mem_ctrl.next_instr_data[16] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _24002_ (.RESET_B(net6695),
    .D(net552),
    .Q(\soc_inst.mem_ctrl.next_instr_data[17] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _24003_ (.RESET_B(net6684),
    .D(net902),
    .Q(\soc_inst.mem_ctrl.next_instr_data[18] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _24004_ (.RESET_B(net6689),
    .D(net737),
    .Q(\soc_inst.mem_ctrl.next_instr_data[19] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _24005_ (.RESET_B(net6695),
    .D(net765),
    .Q(\soc_inst.mem_ctrl.next_instr_data[20] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _24006_ (.RESET_B(net6691),
    .D(net662),
    .Q(\soc_inst.mem_ctrl.next_instr_data[21] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _24007_ (.RESET_B(net6695),
    .D(net498),
    .Q(\soc_inst.mem_ctrl.next_instr_data[22] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _24008_ (.RESET_B(net6696),
    .D(net681),
    .Q(\soc_inst.mem_ctrl.next_instr_data[23] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _24009_ (.RESET_B(net6691),
    .D(net907),
    .Q(\soc_inst.mem_ctrl.next_instr_data[24] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _24010_ (.RESET_B(net6693),
    .D(net1032),
    .Q(\soc_inst.mem_ctrl.next_instr_data[25] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24011_ (.RESET_B(net6693),
    .D(net557),
    .Q(\soc_inst.mem_ctrl.next_instr_data[26] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _24012_ (.RESET_B(net6689),
    .D(net977),
    .Q(\soc_inst.mem_ctrl.next_instr_data[27] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _24013_ (.RESET_B(net6693),
    .D(net487),
    .Q(\soc_inst.mem_ctrl.next_instr_data[28] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24014_ (.RESET_B(net6692),
    .D(net725),
    .Q(\soc_inst.mem_ctrl.next_instr_data[29] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24015_ (.RESET_B(net6684),
    .D(net904),
    .Q(\soc_inst.mem_ctrl.next_instr_data[30] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _24016_ (.RESET_B(net6692),
    .D(net664),
    .Q(\soc_inst.mem_ctrl.next_instr_data[31] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _24017_ (.RESET_B(net6642),
    .D(_00672_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _24018_ (.RESET_B(net6642),
    .D(net1223),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24019_ (.RESET_B(net6640),
    .D(_00673_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.is_write_op ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24020_ (.RESET_B(net6637),
    .D(net312),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24021_ (.RESET_B(net6637),
    .D(_00675_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _24022_ (.RESET_B(net6637),
    .D(net364),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24023_ (.RESET_B(net6596),
    .D(net359),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _24024_ (.RESET_B(net6591),
    .D(net254),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24025_ (.RESET_B(net6591),
    .D(_00679_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24026_ (.RESET_B(net6591),
    .D(net563),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _24027_ (.RESET_B(net6591),
    .D(net339),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _24028_ (.RESET_B(net6595),
    .D(net355),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _24029_ (.RESET_B(net6595),
    .D(_00683_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24030_ (.RESET_B(net6595),
    .D(net389),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _24031_ (.RESET_B(net6596),
    .D(net145),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _24032_ (.RESET_B(net6648),
    .D(net1238),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24033_ (.RESET_B(net6640),
    .D(net1358),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _24034_ (.RESET_B(net6653),
    .D(_00688_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24035_ (.RESET_B(net6649),
    .D(net1040),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24036_ (.RESET_B(net6647),
    .D(net1416),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24037_ (.RESET_B(net6640),
    .D(net1746),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24038_ (.RESET_B(net6651),
    .D(net998),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24039_ (.RESET_B(net6649),
    .D(_00693_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24040_ (.RESET_B(net6646),
    .D(net1088),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24041_ (.RESET_B(net6648),
    .D(net1229),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24042_ (.RESET_B(net6653),
    .D(_00696_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24043_ (.RESET_B(net6652),
    .D(_00697_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24044_ (.RESET_B(net6647),
    .D(net675),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24045_ (.RESET_B(net6648),
    .D(net1123),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _24046_ (.RESET_B(net6653),
    .D(_00700_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24047_ (.RESET_B(net6652),
    .D(net1208),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24048_ (.RESET_B(net6647),
    .D(_00702_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24049_ (.RESET_B(net6648),
    .D(net938),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24050_ (.RESET_B(net6653),
    .D(net1064),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24051_ (.RESET_B(net6652),
    .D(net1061),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24052_ (.RESET_B(net6648),
    .D(net944),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24053_ (.RESET_B(net6648),
    .D(net1264),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24054_ (.RESET_B(net6653),
    .D(_00708_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24055_ (.RESET_B(net6652),
    .D(net916),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24056_ (.RESET_B(net6647),
    .D(net889),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24057_ (.RESET_B(net6649),
    .D(_00711_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _24058_ (.RESET_B(net6690),
    .D(net1290),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24059_ (.RESET_B(net6653),
    .D(_00713_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24060_ (.RESET_B(net6650),
    .D(net154),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _24061_ (.RESET_B(net6652),
    .D(net248),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _24062_ (.RESET_B(net6691),
    .D(net1118),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24063_ (.RESET_B(net6653),
    .D(net302),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24064_ (.RESET_B(net6639),
    .D(_00718_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24065_ (.RESET_B(net6626),
    .D(net1952),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _24066_ (.RESET_B(net6626),
    .D(net1930),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _24067_ (.RESET_B(net6622),
    .D(net2296),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _24068_ (.RESET_B(net6626),
    .D(net2064),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _24069_ (.RESET_B(net6623),
    .D(net1392),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _24070_ (.RESET_B(net6622),
    .D(net2361),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _24071_ (.RESET_B(net6621),
    .D(net909),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _24072_ (.RESET_B(net6623),
    .D(net2424),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _24073_ (.RESET_B(net6623),
    .D(net2118),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _24074_ (.RESET_B(net6623),
    .D(net2053),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _24075_ (.RESET_B(net6622),
    .D(net569),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _24076_ (.RESET_B(net6626),
    .D(net1076),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _24077_ (.RESET_B(net6623),
    .D(net2180),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _24078_ (.RESET_B(net6621),
    .D(net417),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _24079_ (.RESET_B(net6621),
    .D(net397),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _24080_ (.RESET_B(net6621),
    .D(net602),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _24081_ (.RESET_B(net6610),
    .D(net957),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _24082_ (.RESET_B(net6609),
    .D(net1808),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _24083_ (.RESET_B(net6610),
    .D(net584),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _24084_ (.RESET_B(net6623),
    .D(net1671),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24085_ (.RESET_B(net6610),
    .D(net2336),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24086_ (.RESET_B(net6609),
    .D(net1042),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _24087_ (.RESET_B(net6610),
    .D(net995),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _24088_ (.RESET_B(net6633),
    .D(net1191),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _24089_ (.RESET_B(net6634),
    .D(net2520),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _24090_ (.RESET_B(net6642),
    .D(net881),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _24091_ (.RESET_B(net6633),
    .D(net936),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _24092_ (.RESET_B(net6634),
    .D(net789),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _24093_ (.RESET_B(net6634),
    .D(_00747_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _24094_ (.RESET_B(net6634),
    .D(net2737),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _24095_ (.RESET_B(net6634),
    .D(net2826),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24096_ (.RESET_B(net6634),
    .D(net2664),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _24097_ (.RESET_B(net6649),
    .D(_00751_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24098_ (.RESET_B(net6647),
    .D(_00752_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24099_ (.RESET_B(net6650),
    .D(_00753_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24100_ (.RESET_B(net6646),
    .D(_00754_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24101_ (.RESET_B(net6646),
    .D(_00755_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24102_ (.RESET_B(net6646),
    .D(_00756_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24103_ (.RESET_B(net6650),
    .D(_00757_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24104_ (.RESET_B(net6650),
    .D(_00758_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24105_ (.RESET_B(net6650),
    .D(_00759_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24106_ (.RESET_B(net6650),
    .D(_00760_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24107_ (.RESET_B(net6651),
    .D(_00761_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24108_ (.RESET_B(net6651),
    .D(_00762_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24109_ (.RESET_B(net6650),
    .D(_00763_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24110_ (.RESET_B(net6651),
    .D(_00764_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24111_ (.RESET_B(net6690),
    .D(_00765_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24112_ (.RESET_B(net6652),
    .D(_00766_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24113_ (.RESET_B(net6646),
    .D(_00767_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24114_ (.RESET_B(net6648),
    .D(_00768_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24115_ (.RESET_B(net6690),
    .D(net2710),
    .Q(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24116_ (.RESET_B(net6648),
    .D(_00770_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24117_ (.RESET_B(net6646),
    .D(_00771_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24118_ (.RESET_B(net6647),
    .D(_00772_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24119_ (.RESET_B(net6689),
    .D(_00773_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24120_ (.RESET_B(net6652),
    .D(_00774_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24121_ (.RESET_B(net6650),
    .D(net2760),
    .Q(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _24122_ (.RESET_B(net6689),
    .D(net2603),
    .Q(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24123_ (.RESET_B(net6689),
    .D(_00777_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24124_ (.RESET_B(net6690),
    .D(_00778_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24125_ (.RESET_B(net6689),
    .D(_00779_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24126_ (.RESET_B(net6651),
    .D(_00780_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24127_ (.RESET_B(net6690),
    .D(net2642),
    .Q(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _24128_ (.RESET_B(net6690),
    .D(_00782_),
    .Q(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _24129_ (.RESET_B(net6578),
    .D(net96),
    .Q(\soc_inst.bus_spi_sclk ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24130_ (.RESET_B(net6582),
    .D(net75),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_latched ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _24131_ (.RESET_B(net6639),
    .D(net2142),
    .Q(_00250_),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24132_ (.RESET_B(net6640),
    .D(_00784_),
    .Q(\soc_inst.mem_ctrl.spi_done ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24133_ (.RESET_B(net6640),
    .D(net2875),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24134_ (.RESET_B(net6581),
    .D(_00109_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24135_ (.RESET_B(net6721),
    .D(net272),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _24136_ (.RESET_B(net6715),
    .D(net142),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _24137_ (.RESET_B(net6680),
    .D(net196),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _24138_ (.RESET_B(net6716),
    .D(net224),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _24139_ (.RESET_B(net6738),
    .D(net133),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _24140_ (.RESET_B(net6718),
    .D(net136),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _24141_ (.RESET_B(net6680),
    .D(net282),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[11] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _24142_ (.RESET_B(net6681),
    .D(net139),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24143_ (.RESET_B(net6677),
    .D(net425),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_1 _24144_ (.RESET_B(net6709),
    .D(net237),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _24145_ (.RESET_B(net6677),
    .D(net128),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _24146_ (.RESET_B(net6712),
    .D(net285),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24147_ (.RESET_B(net6709),
    .D(net728),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24148_ (.RESET_B(net6711),
    .D(net150),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _24149_ (.RESET_B(net6712),
    .D(net193),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24150_ (.RESET_B(net6712),
    .D(net171),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[20] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24151_ (.RESET_B(net6675),
    .D(net199),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _24152_ (.RESET_B(net6675),
    .D(net178),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24153_ (.RESET_B(net6675),
    .D(net279),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _24154_ (.RESET_B(net6671),
    .D(net750),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24155_ (.RESET_B(net6678),
    .D(net581),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[25] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24156_ (.RESET_B(net6671),
    .D(net554),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[26] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24157_ (.RESET_B(net6672),
    .D(net386),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_1 _24158_ (.RESET_B(net6673),
    .D(net1153),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[28] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24159_ (.RESET_B(net6672),
    .D(net483),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[29] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _24160_ (.RESET_B(net6673),
    .D(net542),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _24161_ (.RESET_B(net6678),
    .D(_00812_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[31] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _24162_ (.RESET_B(net6596),
    .D(_00813_),
    .Q(uio_oe[5]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24163_ (.RESET_B(net6639),
    .D(_00814_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.initialized ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24164_ (.RESET_B(net6582),
    .D(net2989),
    .Q(uio_out[1]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24165_ (.RESET_B(net6582),
    .D(net2992),
    .Q(uio_out[2]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24166_ (.RESET_B(net6581),
    .D(_00817_),
    .Q(uio_out[4]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _24167_ (.RESET_B(net6581),
    .D(net2863),
    .Q(uio_out[5]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _24168_ (.RESET_B(net6590),
    .D(net89),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d1 ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _24169_ (.RESET_B(net6641),
    .D(_00819_),
    .Q(\soc_inst.mem_ctrl.spi_is_instr ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24170_ (.RESET_B(net6640),
    .D(net1570),
    .Q(_00251_),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24171_ (.RESET_B(net6636),
    .D(_00000_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _24172_ (.RESET_B(net6639),
    .D(net438),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24173_ (.RESET_B(net6638),
    .D(net406),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24174_ (.RESET_B(net6639),
    .D(net2883),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24175_ (.RESET_B(net6636),
    .D(net2274),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _24176_ (.RESET_B(net6646),
    .D(net3192),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24177_ (.RESET_B(net6636),
    .D(net2660),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24178_ (.RESET_B(net6594),
    .D(_00017_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _24179_ (.RESET_B(net6636),
    .D(net1136),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _24180_ (.RESET_B(net6636),
    .D(net3368),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _24181_ (.RESET_B(net6639),
    .D(net228),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _24182_ (.RESET_B(net6639),
    .D(net1377),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24183_ (.RESET_B(net6636),
    .D(net1078),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24184_ (.RESET_B(net6647),
    .D(net2854),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _24185_ (.RESET_B(net6636),
    .D(_00005_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24186_ (.RESET_B(net6700),
    .D(_00820_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[0] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24187_ (.RESET_B(net6700),
    .D(_00821_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[1] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24188_ (.RESET_B(net6700),
    .D(_00822_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24189_ (.RESET_B(net6699),
    .D(_00823_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[4] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24190_ (.RESET_B(net71),
    .D(net2921),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _24191_ (.RESET_B(net70),
    .D(_00825_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _24192_ (.RESET_B(net6700),
    .D(_00826_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _24193_ (.RESET_B(net6702),
    .D(_00827_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24194_ (.RESET_B(net6737),
    .D(_00828_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _24195_ (.RESET_B(net6700),
    .D(_00829_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24196_ (.RESET_B(net6699),
    .D(_00830_),
    .Q(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24197_ (.RESET_B(net6637),
    .D(_00831_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _24198_ (.RESET_B(net6637),
    .D(net3376),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _24199_ (.RESET_B(net6637),
    .D(_00833_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24200_ (.RESET_B(net6638),
    .D(_00834_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _24201_ (.RESET_B(net6639),
    .D(_00835_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _24202_ (.RESET_B(net6590),
    .D(net85),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d2 ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _24203_ (.RESET_B(net6591),
    .D(net91),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d3 ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _24204_ (.RESET_B(net6636),
    .D(_00836_),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.write_mosi ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24205_ (.RESET_B(net6652),
    .D(net94),
    .Q(\soc_inst.cpu_core.csr_file.mip_eip ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24206_ (.RESET_B(net6781),
    .D(_00837_),
    .Q(\soc_inst.cpu_core.id_int_is_interrupt ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _24207_ (.RESET_B(net6791),
    .D(net1178),
    .Q(\soc_inst.cpu_core.ex_reg_we ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24208_ (.RESET_B(net6729),
    .D(_00839_),
    .Q(\soc_inst.cpu_core.csr_file.mret_trigger ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _24209_ (.RESET_B(net6733),
    .D(_00840_),
    .Q(\soc_inst.cpu_core.ex_is_ebreak ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24210_ (.RESET_B(net6574),
    .D(net378),
    .Q(\soc_inst.core_mem_wdata[0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _24211_ (.RESET_B(net6594),
    .D(net300),
    .Q(\soc_inst.core_mem_wdata[1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24212_ (.RESET_B(net6704),
    .D(net792),
    .Q(\soc_inst.core_mem_wdata[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24213_ (.RESET_B(net6574),
    .D(_00844_),
    .Q(\soc_inst.core_mem_wdata[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _24214_ (.RESET_B(net6594),
    .D(_00845_),
    .Q(\soc_inst.core_mem_wdata[4] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _24215_ (.RESET_B(net6596),
    .D(_00846_),
    .Q(\soc_inst.core_mem_wdata[5] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _24216_ (.RESET_B(net6594),
    .D(_00847_),
    .Q(\soc_inst.core_mem_wdata[6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _24217_ (.RESET_B(net6632),
    .D(_00848_),
    .Q(\soc_inst.core_mem_wdata[7] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24218_ (.RESET_B(net6627),
    .D(_00849_),
    .Q(\soc_inst.core_mem_wdata[8] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _24219_ (.RESET_B(net6610),
    .D(_00850_),
    .Q(\soc_inst.core_mem_wdata[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _24220_ (.RESET_B(net6666),
    .D(_00851_),
    .Q(\soc_inst.core_mem_wdata[10] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _24221_ (.RESET_B(net6604),
    .D(net1397),
    .Q(\soc_inst.core_mem_wdata[11] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24222_ (.RESET_B(net6621),
    .D(_00853_),
    .Q(\soc_inst.core_mem_wdata[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _24223_ (.RESET_B(net6559),
    .D(_00854_),
    .Q(\soc_inst.core_mem_wdata[13] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _24224_ (.RESET_B(net6557),
    .D(_00855_),
    .Q(\soc_inst.core_mem_wdata[14] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24225_ (.RESET_B(net6615),
    .D(_00856_),
    .Q(\soc_inst.core_mem_wdata[15] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_2 _24226_ (.RESET_B(net6618),
    .D(_00857_),
    .Q(\soc_inst.core_mem_wdata[16] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24227_ (.RESET_B(net6618),
    .D(_00858_),
    .Q(\soc_inst.core_mem_wdata[17] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24228_ (.RESET_B(net6658),
    .D(_00859_),
    .Q(\soc_inst.core_mem_wdata[18] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _24229_ (.RESET_B(net6619),
    .D(_00860_),
    .Q(\soc_inst.core_mem_wdata[19] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24230_ (.RESET_B(net6619),
    .D(_00861_),
    .Q(\soc_inst.core_mem_wdata[20] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24231_ (.RESET_B(net6657),
    .D(_00862_),
    .Q(\soc_inst.core_mem_wdata[21] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _24232_ (.RESET_B(net6657),
    .D(_00863_),
    .Q(\soc_inst.core_mem_wdata[22] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24233_ (.RESET_B(net6661),
    .D(_00864_),
    .Q(\soc_inst.core_mem_wdata[23] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24234_ (.RESET_B(net6618),
    .D(_00865_),
    .Q(\soc_inst.core_mem_wdata[24] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24235_ (.RESET_B(net6615),
    .D(_00866_),
    .Q(\soc_inst.core_mem_wdata[25] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_2 _24236_ (.RESET_B(net6659),
    .D(_00867_),
    .Q(\soc_inst.core_mem_wdata[26] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24237_ (.RESET_B(net6657),
    .D(_00868_),
    .Q(\soc_inst.core_mem_wdata[27] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24238_ (.RESET_B(net6604),
    .D(_00869_),
    .Q(\soc_inst.core_mem_wdata[28] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _24239_ (.RESET_B(net6604),
    .D(_00870_),
    .Q(\soc_inst.core_mem_wdata[29] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24240_ (.RESET_B(net6657),
    .D(_00871_),
    .Q(\soc_inst.core_mem_wdata[30] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24241_ (.RESET_B(net6659),
    .D(_00872_),
    .Q(\soc_inst.core_mem_wdata[31] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _24242_ (.RESET_B(net6733),
    .D(net2456),
    .Q(\soc_inst.cpu_core.ex_is_ecall ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24243_ (.RESET_B(net6638),
    .D(net897),
    .Q(\soc_inst.cpu_core.error_flag_reg ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24244_ (.RESET_B(net6748),
    .D(net1887),
    .Q(_00252_),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24245_ (.RESET_B(net6748),
    .D(net2014),
    .Q(_00253_),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24246_ (.RESET_B(net6748),
    .D(_00877_),
    .Q(\soc_inst.cpu_core.if_instr[2] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24247_ (.RESET_B(net6787),
    .D(_00878_),
    .Q(\soc_inst.cpu_core.if_instr[3] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _24248_ (.RESET_B(net6793),
    .D(net2878),
    .Q(_00254_),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24249_ (.RESET_B(net6794),
    .D(_00880_),
    .Q(\soc_inst.cpu_core.if_instr[5] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _24250_ (.RESET_B(net6793),
    .D(_00881_),
    .Q(\soc_inst.cpu_core.if_instr[6] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24251_ (.RESET_B(net6788),
    .D(_00882_),
    .Q(\soc_inst.cpu_core.if_instr[7] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _24252_ (.RESET_B(net6750),
    .D(_00883_),
    .Q(\soc_inst.cpu_core.if_instr[8] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _24253_ (.RESET_B(net6748),
    .D(net1266),
    .Q(\soc_inst.cpu_core.if_instr[9] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _24254_ (.RESET_B(net6750),
    .D(net874),
    .Q(\soc_inst.cpu_core.if_instr[10] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _24255_ (.RESET_B(net6750),
    .D(net1249),
    .Q(\soc_inst.cpu_core.if_instr[11] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _24256_ (.RESET_B(net6789),
    .D(net3015),
    .Q(\soc_inst.cpu_core.if_funct3[0] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24257_ (.RESET_B(net6787),
    .D(_00888_),
    .Q(\soc_inst.cpu_core.if_funct3[1] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24258_ (.RESET_B(net6795),
    .D(net2946),
    .Q(\soc_inst.cpu_core.if_funct3[2] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _24259_ (.RESET_B(net6749),
    .D(_00890_),
    .Q(\soc_inst.cpu_core.if_instr[15] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _24260_ (.RESET_B(net6741),
    .D(_00891_),
    .Q(\soc_inst.cpu_core.if_instr[16] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _24261_ (.RESET_B(net6749),
    .D(_00892_),
    .Q(\soc_inst.cpu_core.if_instr[17] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24262_ (.RESET_B(net6739),
    .D(_00893_),
    .Q(\soc_inst.cpu_core.if_instr[18] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24263_ (.RESET_B(net6743),
    .D(_00894_),
    .Q(\soc_inst.cpu_core.if_instr[19] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24264_ (.RESET_B(net6794),
    .D(_00895_),
    .Q(\soc_inst.cpu_core.if_imm12[0] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24265_ (.RESET_B(net6749),
    .D(_00896_),
    .Q(\soc_inst.cpu_core.if_imm12[1] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _24266_ (.RESET_B(net6794),
    .D(_00897_),
    .Q(\soc_inst.cpu_core.if_imm12[2] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _24267_ (.RESET_B(net6793),
    .D(_00898_),
    .Q(\soc_inst.cpu_core.if_imm12[3] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _24268_ (.RESET_B(net6748),
    .D(_00899_),
    .Q(\soc_inst.cpu_core.if_imm12[4] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24269_ (.RESET_B(net6743),
    .D(_00900_),
    .Q(\soc_inst.cpu_core.if_funct7[0] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24270_ (.RESET_B(net6743),
    .D(_00901_),
    .Q(\soc_inst.cpu_core.if_funct7[1] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24271_ (.RESET_B(net6741),
    .D(_00902_),
    .Q(\soc_inst.cpu_core.if_funct7[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24272_ (.RESET_B(net6746),
    .D(_00903_),
    .Q(\soc_inst.cpu_core.if_funct7[3] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24273_ (.RESET_B(net6748),
    .D(_00904_),
    .Q(\soc_inst.cpu_core.if_funct7[4] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24274_ (.RESET_B(net6743),
    .D(_00905_),
    .Q(\soc_inst.cpu_core.if_funct7[5] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24275_ (.RESET_B(net6706),
    .D(_00906_),
    .Q(\soc_inst.cpu_core.if_funct7[6] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24276_ (.RESET_B(net6743),
    .D(_00907_),
    .Q(\soc_inst.cpu_core.if_pc[0] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24277_ (.RESET_B(net6787),
    .D(_00908_),
    .Q(\soc_inst.cpu_core.if_pc[1] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24278_ (.RESET_B(net6790),
    .D(_00909_),
    .Q(\soc_inst.cpu_core.if_pc[2] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24279_ (.RESET_B(net6781),
    .D(_00910_),
    .Q(\soc_inst.cpu_core.if_pc[3] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24280_ (.RESET_B(net6741),
    .D(_00911_),
    .Q(\soc_inst.cpu_core.if_pc[4] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24281_ (.RESET_B(net6784),
    .D(_00912_),
    .Q(\soc_inst.cpu_core.if_pc[5] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _24282_ (.RESET_B(net6784),
    .D(_00913_),
    .Q(\soc_inst.cpu_core.if_pc[6] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _24283_ (.RESET_B(net6782),
    .D(_00914_),
    .Q(\soc_inst.cpu_core.if_pc[7] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _24284_ (.RESET_B(net6783),
    .D(_00915_),
    .Q(\soc_inst.cpu_core.if_pc[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24285_ (.RESET_B(net6783),
    .D(net2835),
    .Q(\soc_inst.cpu_core.if_pc[9] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _24286_ (.RESET_B(net6766),
    .D(net2768),
    .Q(\soc_inst.cpu_core.if_pc[10] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24287_ (.RESET_B(net6766),
    .D(net2343),
    .Q(\soc_inst.cpu_core.if_pc[11] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _24288_ (.RESET_B(net6728),
    .D(net2764),
    .Q(\soc_inst.cpu_core.if_pc[12] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_1 _24289_ (.RESET_B(net6728),
    .D(net2591),
    .Q(\soc_inst.cpu_core.if_pc[13] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24290_ (.RESET_B(net6730),
    .D(net2484),
    .Q(\soc_inst.cpu_core.if_pc[14] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24291_ (.RESET_B(net6730),
    .D(net2412),
    .Q(\soc_inst.cpu_core.if_pc[15] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24292_ (.RESET_B(net6725),
    .D(net2401),
    .Q(\soc_inst.cpu_core.if_pc[16] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24293_ (.RESET_B(net6725),
    .D(net2350),
    .Q(\soc_inst.cpu_core.if_pc[17] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_1 _24294_ (.RESET_B(net6725),
    .D(net2680),
    .Q(\soc_inst.cpu_core.if_pc[18] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24295_ (.RESET_B(net6725),
    .D(net2766),
    .Q(\soc_inst.cpu_core.if_pc[19] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24296_ (.RESET_B(net6758),
    .D(net2559),
    .Q(\soc_inst.cpu_core.if_pc[20] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24297_ (.RESET_B(net6760),
    .D(_00928_),
    .Q(\soc_inst.cpu_core.if_pc[21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _24298_ (.RESET_B(net6758),
    .D(net2383),
    .Q(\soc_inst.cpu_core.if_pc[22] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24299_ (.RESET_B(net6728),
    .D(net2948),
    .Q(\soc_inst.cpu_core.if_pc[23] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24300_ (.RESET_B(net6687),
    .D(_00026_),
    .Q(\soc_inst.cpu_core.mem_stall ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _24301_ (.RESET_B(net6789),
    .D(_00931_),
    .Q(\soc_inst.cpu_core.if_is_compressed ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _24302_ (.RESET_B(net6744),
    .D(_00932_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24303_ (.RESET_B(net6746),
    .D(_00933_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24304_ (.RESET_B(net6742),
    .D(net1739),
    .Q(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24305_ (.RESET_B(net6751),
    .D(_00935_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _24306_ (.RESET_B(net6744),
    .D(_00936_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24307_ (.RESET_B(net6750),
    .D(_00937_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _24308_ (.RESET_B(net6706),
    .D(_00938_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24309_ (.RESET_B(net6715),
    .D(_00939_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24310_ (.RESET_B(net6715),
    .D(_00940_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _24311_ (.RESET_B(net6742),
    .D(_00941_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24312_ (.RESET_B(net6718),
    .D(_00942_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24313_ (.RESET_B(net6715),
    .D(_00943_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24314_ (.RESET_B(net6681),
    .D(_00944_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_2 _24315_ (.RESET_B(net6677),
    .D(_00945_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _24316_ (.RESET_B(net6709),
    .D(_00946_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24317_ (.RESET_B(net6710),
    .D(_00947_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24318_ (.RESET_B(net6727),
    .D(_00948_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24319_ (.RESET_B(net6724),
    .D(_00949_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24320_ (.RESET_B(net6725),
    .D(_00950_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_2 _24321_ (.RESET_B(net6725),
    .D(_00951_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24322_ (.RESET_B(net6756),
    .D(_00952_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24323_ (.RESET_B(net6727),
    .D(_00953_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24324_ (.RESET_B(net6724),
    .D(_00954_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24325_ (.RESET_B(net6712),
    .D(_00955_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24326_ (.RESET_B(net6725),
    .D(_00956_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24327_ (.RESET_B(net6710),
    .D(_00957_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24328_ (.RESET_B(net6772),
    .D(_00958_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _24329_ (.RESET_B(net6724),
    .D(_00959_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24330_ (.RESET_B(net6757),
    .D(_00960_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _24331_ (.RESET_B(net6659),
    .D(net2673),
    .Q(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _24332_ (.RESET_B(net6714),
    .D(_00962_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24333_ (.RESET_B(net6765),
    .D(_00963_),
    .Q(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_2 _24334_ (.RESET_B(net6781),
    .D(_00964_),
    .Q(_00255_),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24335_ (.RESET_B(net6781),
    .D(_00965_),
    .Q(_00256_),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24336_ (.RESET_B(net6749),
    .D(_00966_),
    .Q(\soc_inst.cpu_core.id_instr[2] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24337_ (.RESET_B(net6749),
    .D(_00967_),
    .Q(\soc_inst.cpu_core.id_instr[3] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24338_ (.RESET_B(net6787),
    .D(_00968_),
    .Q(_00257_),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24339_ (.RESET_B(net6792),
    .D(_00969_),
    .Q(\soc_inst.cpu_core.id_instr[5] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24340_ (.RESET_B(net6792),
    .D(_00970_),
    .Q(\soc_inst.cpu_core.id_instr[6] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24341_ (.RESET_B(net6788),
    .D(_00971_),
    .Q(\soc_inst.cpu_core.id_instr[7] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _24342_ (.RESET_B(net6789),
    .D(_00972_),
    .Q(\soc_inst.cpu_core.id_instr[8] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _24343_ (.RESET_B(net6788),
    .D(_00973_),
    .Q(\soc_inst.cpu_core.id_instr[9] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _24344_ (.RESET_B(net6788),
    .D(_00974_),
    .Q(\soc_inst.cpu_core.id_instr[10] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _24345_ (.RESET_B(net6789),
    .D(_00975_),
    .Q(\soc_inst.cpu_core.id_instr[11] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _24346_ (.RESET_B(net6797),
    .D(_00976_),
    .Q(\soc_inst.cpu_core.id_funct3[0] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _24347_ (.RESET_B(net6796),
    .D(_00977_),
    .Q(\soc_inst.cpu_core.id_funct3[1] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24348_ (.RESET_B(net6780),
    .D(_00978_),
    .Q(\soc_inst.cpu_core.id_funct3[2] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _24349_ (.RESET_B(net6778),
    .D(_00979_),
    .Q(\soc_inst.cpu_core.id_instr[15] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _24350_ (.RESET_B(net6745),
    .D(_00980_),
    .Q(\soc_inst.cpu_core.id_instr[16] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24351_ (.RESET_B(net6762),
    .D(_00981_),
    .Q(\soc_inst.cpu_core.id_instr[17] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _24352_ (.RESET_B(net6747),
    .D(_00982_),
    .Q(\soc_inst.cpu_core.id_instr[18] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24353_ (.RESET_B(net6781),
    .D(_00983_),
    .Q(\soc_inst.cpu_core.id_instr[19] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24354_ (.RESET_B(net6763),
    .D(_00984_),
    .Q(\soc_inst.cpu_core.id_imm12[0] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24355_ (.RESET_B(net6761),
    .D(_00985_),
    .Q(\soc_inst.cpu_core.id_imm12[1] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _24356_ (.RESET_B(net6733),
    .D(_00986_),
    .Q(\soc_inst.cpu_core.id_imm12[2] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_2 _24357_ (.RESET_B(net6767),
    .D(_00987_),
    .Q(\soc_inst.cpu_core.id_imm12[3] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24358_ (.RESET_B(net6733),
    .D(_00988_),
    .Q(\soc_inst.cpu_core.id_imm12[4] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _24359_ (.RESET_B(net6732),
    .D(_00989_),
    .Q(\soc_inst.cpu_core.id_imm12[5] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _24360_ (.RESET_B(net6761),
    .D(_00990_),
    .Q(\soc_inst.cpu_core.id_imm12[6] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _24361_ (.RESET_B(net6732),
    .D(_00991_),
    .Q(\soc_inst.cpu_core.id_imm12[7] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _24362_ (.RESET_B(net6766),
    .D(_00992_),
    .Q(\soc_inst.cpu_core.id_imm12[8] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _24363_ (.RESET_B(net6762),
    .D(_00993_),
    .Q(\soc_inst.cpu_core.id_imm12[9] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24364_ (.RESET_B(net6732),
    .D(_00994_),
    .Q(\soc_inst.cpu_core.id_imm12[10] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _24365_ (.RESET_B(net6780),
    .D(_00995_),
    .Q(\soc_inst.cpu_core.id_imm12[11] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _24366_ (.RESET_B(net6588),
    .D(_00173_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _24367_ (.RESET_B(net6606),
    .D(_00184_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24368_ (.RESET_B(net6606),
    .D(_00195_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24369_ (.RESET_B(net6606),
    .D(net1180),
    .Q(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24370_ (.RESET_B(net6606),
    .D(net3256),
    .Q(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24371_ (.RESET_B(net6606),
    .D(_00216_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24372_ (.RESET_B(net6606),
    .D(net1091),
    .Q(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24373_ (.RESET_B(net6608),
    .D(net401),
    .Q(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24374_ (.RESET_B(net6608),
    .D(net3165),
    .Q(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24375_ (.RESET_B(net6608),
    .D(_00220_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24376_ (.RESET_B(net6602),
    .D(net989),
    .Q(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _24377_ (.RESET_B(net6602),
    .D(net1082),
    .Q(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _24378_ (.RESET_B(net6602),
    .D(_00176_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _24379_ (.RESET_B(net6601),
    .D(_00177_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _24380_ (.RESET_B(net6600),
    .D(net1246),
    .Q(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_2 _24381_ (.RESET_B(net6600),
    .D(_00179_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_2 _24382_ (.RESET_B(net6661),
    .D(net2465),
    .Q(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24383_ (.RESET_B(net6662),
    .D(_00181_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24384_ (.RESET_B(net6658),
    .D(net2718),
    .Q(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24385_ (.RESET_B(net6658),
    .D(net2791),
    .Q(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _24386_ (.RESET_B(net6658),
    .D(net2389),
    .Q(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _24387_ (.RESET_B(net6661),
    .D(_00186_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _24388_ (.RESET_B(net6657),
    .D(net2770),
    .Q(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _24389_ (.RESET_B(net6658),
    .D(_00188_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _24390_ (.RESET_B(net6661),
    .D(net2571),
    .Q(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _24391_ (.RESET_B(net6660),
    .D(net2518),
    .Q(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24392_ (.RESET_B(net6663),
    .D(net2076),
    .Q(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _24393_ (.RESET_B(net6663),
    .D(net2319),
    .Q(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24394_ (.RESET_B(net6663),
    .D(net1981),
    .Q(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _24395_ (.RESET_B(net6663),
    .D(_00194_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _24396_ (.RESET_B(net6664),
    .D(_00196_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_2 _24397_ (.RESET_B(net6663),
    .D(net2892),
    .Q(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _24398_ (.RESET_B(net6608),
    .D(net2136),
    .Q(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _24399_ (.RESET_B(net6607),
    .D(_00199_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24400_ (.RESET_B(net6606),
    .D(net3230),
    .Q(\soc_inst.cpu_core.csr_file.mtime[34] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24401_ (.RESET_B(net6607),
    .D(net1200),
    .Q(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24402_ (.RESET_B(net6607),
    .D(net1483),
    .Q(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24403_ (.RESET_B(net6607),
    .D(_00203_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _24404_ (.RESET_B(net6608),
    .D(net1332),
    .Q(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _24405_ (.RESET_B(net6608),
    .D(_00205_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24406_ (.RESET_B(net6608),
    .D(_00207_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _24407_ (.RESET_B(net6608),
    .D(net1373),
    .Q(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24408_ (.RESET_B(net6603),
    .D(net1170),
    .Q(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _24409_ (.RESET_B(net6603),
    .D(net942),
    .Q(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _24410_ (.RESET_B(net6602),
    .D(net628),
    .Q(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _24411_ (.RESET_B(net6601),
    .D(_00212_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _24412_ (.RESET_B(net6601),
    .D(_00213_),
    .Q(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _24413_ (.RESET_B(net6601),
    .D(net1141),
    .Q(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _24414_ (.RESET_B(net6793),
    .D(_00996_),
    .Q(\soc_inst.cpu_core.id_rs1_data[0] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24415_ (.RESET_B(net6804),
    .D(_00997_),
    .Q(\soc_inst.cpu_core.id_rs1_data[1] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24416_ (.RESET_B(net6804),
    .D(_00998_),
    .Q(\soc_inst.cpu_core.id_rs1_data[2] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24417_ (.RESET_B(net6787),
    .D(_00999_),
    .Q(\soc_inst.cpu_core.id_rs1_data[3] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24418_ (.RESET_B(net6793),
    .D(_01000_),
    .Q(\soc_inst.cpu_core.id_rs1_data[4] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24419_ (.RESET_B(net6793),
    .D(_01001_),
    .Q(\soc_inst.cpu_core.id_rs1_data[5] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24420_ (.RESET_B(net6791),
    .D(_01002_),
    .Q(\soc_inst.cpu_core.id_rs1_data[6] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24421_ (.RESET_B(net6791),
    .D(_01003_),
    .Q(\soc_inst.cpu_core.id_rs1_data[7] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _24422_ (.RESET_B(net6785),
    .D(_01004_),
    .Q(\soc_inst.cpu_core.id_rs1_data[8] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _24423_ (.RESET_B(net6784),
    .D(_01005_),
    .Q(\soc_inst.cpu_core.id_rs1_data[9] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _24424_ (.RESET_B(net6785),
    .D(_01006_),
    .Q(\soc_inst.cpu_core.id_rs1_data[10] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24425_ (.RESET_B(net6780),
    .D(_01007_),
    .Q(\soc_inst.cpu_core.id_rs1_data[11] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _24426_ (.RESET_B(net6766),
    .D(_01008_),
    .Q(\soc_inst.cpu_core.id_rs1_data[12] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24427_ (.RESET_B(net6761),
    .D(_01009_),
    .Q(\soc_inst.cpu_core.id_rs1_data[13] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24428_ (.RESET_B(net6765),
    .D(_01010_),
    .Q(\soc_inst.cpu_core.id_rs1_data[14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24429_ (.RESET_B(net6761),
    .D(_01011_),
    .Q(\soc_inst.cpu_core.id_rs1_data[15] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24430_ (.RESET_B(net6756),
    .D(_01012_),
    .Q(\soc_inst.cpu_core.id_rs1_data[16] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _24431_ (.RESET_B(net6769),
    .D(_01013_),
    .Q(\soc_inst.cpu_core.id_rs1_data[17] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24432_ (.RESET_B(net6771),
    .D(_01014_),
    .Q(\soc_inst.cpu_core.id_rs1_data[18] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _24433_ (.RESET_B(net6772),
    .D(_01015_),
    .Q(\soc_inst.cpu_core.id_rs1_data[19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24434_ (.RESET_B(net6770),
    .D(_01016_),
    .Q(\soc_inst.cpu_core.id_rs1_data[20] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24435_ (.RESET_B(net6769),
    .D(_01017_),
    .Q(\soc_inst.cpu_core.id_rs1_data[21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24436_ (.RESET_B(net6759),
    .D(_01018_),
    .Q(\soc_inst.cpu_core.id_rs1_data[22] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _24437_ (.RESET_B(net6757),
    .D(_01019_),
    .Q(\soc_inst.cpu_core.id_rs1_data[23] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _24438_ (.RESET_B(net6759),
    .D(_01020_),
    .Q(\soc_inst.cpu_core.id_rs1_data[24] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _24439_ (.RESET_B(net6773),
    .D(_01021_),
    .Q(\soc_inst.cpu_core.id_rs1_data[25] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _24440_ (.RESET_B(net6771),
    .D(net3251),
    .Q(\soc_inst.cpu_core.id_rs1_data[26] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _24441_ (.RESET_B(net6770),
    .D(_01023_),
    .Q(\soc_inst.cpu_core.id_rs1_data[27] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _24442_ (.RESET_B(net6770),
    .D(_01024_),
    .Q(\soc_inst.cpu_core.id_rs1_data[28] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24443_ (.RESET_B(net6811),
    .D(_01025_),
    .Q(\soc_inst.cpu_core.id_rs1_data[29] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _24444_ (.RESET_B(net6763),
    .D(_01026_),
    .Q(\soc_inst.cpu_core.id_rs1_data[30] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24445_ (.RESET_B(net6765),
    .D(net2712),
    .Q(\soc_inst.cpu_core.id_rs1_data[31] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _24446_ (.RESET_B(net6701),
    .D(net2302),
    .Q(_00258_),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _24447_ (.RESET_B(net6701),
    .D(net2583),
    .Q(_00259_),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24448_ (.RESET_B(net6701),
    .D(net1983),
    .Q(\soc_inst.cpu_core.mem_instr[2] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24449_ (.RESET_B(net6701),
    .D(net2276),
    .Q(\soc_inst.cpu_core.mem_instr[3] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24450_ (.RESET_B(net6745),
    .D(net1832),
    .Q(_00260_),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _24451_ (.RESET_B(net6781),
    .D(net2775),
    .Q(\soc_inst.cpu_core.mem_instr[5] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _24452_ (.RESET_B(net6744),
    .D(net3024),
    .Q(\soc_inst.cpu_core.mem_instr[6] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _24453_ (.RESET_B(net6801),
    .D(_01035_),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[4] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _24454_ (.RESET_B(net6747),
    .D(_01036_),
    .Q(\soc_inst.core_mem_flag[0] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _24455_ (.RESET_B(net6741),
    .D(_01037_),
    .Q(\soc_inst.core_mem_flag[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _24456_ (.RESET_B(net6744),
    .D(_01038_),
    .Q(\soc_inst.core_mem_flag[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24457_ (.RESET_B(net6729),
    .D(net1084),
    .Q(\soc_inst.cpu_core.mem_instr[15] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_1 _24458_ (.RESET_B(net6740),
    .D(net2385),
    .Q(\soc_inst.cpu_core.mem_instr[16] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24459_ (.RESET_B(net6730),
    .D(net1159),
    .Q(\soc_inst.cpu_core.mem_instr[17] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24460_ (.RESET_B(net6745),
    .D(net2283),
    .Q(\soc_inst.cpu_core.mem_instr[18] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _24461_ (.RESET_B(net6744),
    .D(net1405),
    .Q(\soc_inst.cpu_core.mem_instr[19] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24462_ (.RESET_B(net6731),
    .D(net604),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[0] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24463_ (.RESET_B(net6760),
    .D(net2488),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[1] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24464_ (.RESET_B(net6717),
    .D(net1282),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[2] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _24465_ (.RESET_B(net6763),
    .D(net2716),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[3] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_2 _24466_ (.RESET_B(net6730),
    .D(net2662),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[4] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _24467_ (.RESET_B(net6728),
    .D(net918),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[5] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _24468_ (.RESET_B(net6731),
    .D(_01050_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_2 _24469_ (.RESET_B(net6728),
    .D(net2394),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[7] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _24470_ (.RESET_B(net6681),
    .D(net2565),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _24471_ (.RESET_B(net6761),
    .D(_01053_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_2 _24472_ (.RESET_B(net6728),
    .D(net2099),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[10] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _24473_ (.RESET_B(net6764),
    .D(_01055_),
    .Q(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _24474_ (.RESET_B(net6833),
    .D(_01056_),
    .Q(\soc_inst.cpu_core.id_rs2_data[0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _24475_ (.RESET_B(net6804),
    .D(_01057_),
    .Q(\soc_inst.cpu_core.id_rs2_data[1] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24476_ (.RESET_B(net6803),
    .D(_01058_),
    .Q(\soc_inst.cpu_core.id_rs2_data[2] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _24477_ (.RESET_B(net6749),
    .D(net2896),
    .Q(\soc_inst.cpu_core.id_rs2_data[3] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24478_ (.RESET_B(net6793),
    .D(_01060_),
    .Q(\soc_inst.cpu_core.id_rs2_data[4] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24479_ (.RESET_B(net6802),
    .D(_01061_),
    .Q(\soc_inst.cpu_core.id_rs2_data[5] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24480_ (.RESET_B(net6801),
    .D(_01062_),
    .Q(\soc_inst.cpu_core.id_rs2_data[6] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24481_ (.RESET_B(net6791),
    .D(_01063_),
    .Q(\soc_inst.cpu_core.id_rs2_data[7] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _24482_ (.RESET_B(net6762),
    .D(_01064_),
    .Q(\soc_inst.cpu_core.id_rs2_data[8] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24483_ (.RESET_B(net6766),
    .D(_01065_),
    .Q(\soc_inst.cpu_core.id_rs2_data[9] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24484_ (.RESET_B(net6766),
    .D(_01066_),
    .Q(\soc_inst.cpu_core.id_rs2_data[10] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _24485_ (.RESET_B(net6804),
    .D(_01067_),
    .Q(\soc_inst.cpu_core.id_rs2_data[11] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _24486_ (.RESET_B(net6732),
    .D(_01068_),
    .Q(\soc_inst.cpu_core.id_rs2_data[12] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24487_ (.RESET_B(net6731),
    .D(_01069_),
    .Q(\soc_inst.cpu_core.id_rs2_data[13] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24488_ (.RESET_B(net6731),
    .D(_01070_),
    .Q(\soc_inst.cpu_core.id_rs2_data[14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24489_ (.RESET_B(net6761),
    .D(_01071_),
    .Q(\soc_inst.cpu_core.id_rs2_data[15] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24490_ (.RESET_B(net6806),
    .D(_01072_),
    .Q(\soc_inst.cpu_core.id_rs2_data[16] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _24491_ (.RESET_B(net6759),
    .D(_01073_),
    .Q(\soc_inst.cpu_core.id_rs2_data[17] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _24492_ (.RESET_B(net6770),
    .D(_01074_),
    .Q(\soc_inst.cpu_core.id_rs2_data[18] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24493_ (.RESET_B(net6769),
    .D(_01075_),
    .Q(\soc_inst.cpu_core.id_rs2_data[19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24494_ (.RESET_B(net6771),
    .D(_01076_),
    .Q(\soc_inst.cpu_core.id_rs2_data[20] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24495_ (.RESET_B(net6806),
    .D(_01077_),
    .Q(\soc_inst.cpu_core.id_rs2_data[21] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _24496_ (.RESET_B(net6806),
    .D(_01078_),
    .Q(\soc_inst.cpu_core.id_rs2_data[22] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _24497_ (.RESET_B(net6806),
    .D(_01079_),
    .Q(\soc_inst.cpu_core.id_rs2_data[23] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _24498_ (.RESET_B(net6815),
    .D(_01080_),
    .Q(\soc_inst.cpu_core.id_rs2_data[24] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _24499_ (.RESET_B(net6807),
    .D(_01081_),
    .Q(\soc_inst.cpu_core.id_rs2_data[25] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24500_ (.RESET_B(net6813),
    .D(_01082_),
    .Q(\soc_inst.cpu_core.id_rs2_data[26] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24501_ (.RESET_B(net6813),
    .D(_01083_),
    .Q(\soc_inst.cpu_core.id_rs2_data[27] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _24502_ (.RESET_B(net6813),
    .D(_01084_),
    .Q(\soc_inst.cpu_core.id_rs2_data[28] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _24503_ (.RESET_B(net6813),
    .D(_01085_),
    .Q(\soc_inst.cpu_core.id_rs2_data[29] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _24504_ (.RESET_B(net6807),
    .D(_01086_),
    .Q(\soc_inst.cpu_core.id_rs2_data[30] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24505_ (.RESET_B(net6774),
    .D(_01087_),
    .Q(\soc_inst.cpu_core.id_rs2_data[31] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _24506_ (.RESET_B(net6788),
    .D(_01088_),
    .Q(\soc_inst.cpu_core.id_imm[0] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24507_ (.RESET_B(net6787),
    .D(_01089_),
    .Q(\soc_inst.cpu_core.id_imm[1] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24508_ (.RESET_B(net6787),
    .D(_01090_),
    .Q(\soc_inst.cpu_core.id_imm[2] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24509_ (.RESET_B(net6793),
    .D(net2817),
    .Q(\soc_inst.cpu_core.id_imm[3] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24510_ (.RESET_B(net6794),
    .D(_01092_),
    .Q(\soc_inst.cpu_core.id_imm[4] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24511_ (.RESET_B(net6794),
    .D(_01093_),
    .Q(\soc_inst.cpu_core.id_imm[5] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _24512_ (.RESET_B(net6791),
    .D(net2795),
    .Q(\soc_inst.cpu_core.id_imm[6] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24513_ (.RESET_B(net6802),
    .D(_01095_),
    .Q(\soc_inst.cpu_core.id_imm[7] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _24514_ (.RESET_B(net6784),
    .D(net2427),
    .Q(\soc_inst.cpu_core.id_imm[8] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24515_ (.RESET_B(net6785),
    .D(_01097_),
    .Q(\soc_inst.cpu_core.id_imm[9] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24516_ (.RESET_B(net6785),
    .D(net2479),
    .Q(\soc_inst.cpu_core.id_imm[10] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _24517_ (.RESET_B(net6787),
    .D(_01099_),
    .Q(\soc_inst.cpu_core.id_imm[11] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24518_ (.RESET_B(net6766),
    .D(_01100_),
    .Q(\soc_inst.cpu_core.id_imm[12] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24519_ (.RESET_B(net6764),
    .D(net2907),
    .Q(\soc_inst.cpu_core.id_imm[13] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24520_ (.RESET_B(net6763),
    .D(_01102_),
    .Q(\soc_inst.cpu_core.id_imm[14] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24521_ (.RESET_B(net6767),
    .D(_01103_),
    .Q(\soc_inst.cpu_core.id_imm[15] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24522_ (.RESET_B(net6772),
    .D(_01104_),
    .Q(\soc_inst.cpu_core.id_imm[16] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _24523_ (.RESET_B(net6772),
    .D(_01105_),
    .Q(\soc_inst.cpu_core.id_imm[17] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _24524_ (.RESET_B(net6771),
    .D(_01106_),
    .Q(\soc_inst.cpu_core.id_imm[18] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_2 _24525_ (.RESET_B(net6770),
    .D(_01107_),
    .Q(\soc_inst.cpu_core.id_imm[19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_2 _24526_ (.RESET_B(net6760),
    .D(_01108_),
    .Q(\soc_inst.cpu_core.id_imm[20] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _24527_ (.RESET_B(net6774),
    .D(_01109_),
    .Q(\soc_inst.cpu_core.id_imm[21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24528_ (.RESET_B(net6771),
    .D(_01110_),
    .Q(\soc_inst.cpu_core.id_imm[22] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24529_ (.RESET_B(net6773),
    .D(_01111_),
    .Q(\soc_inst.cpu_core.id_imm[23] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _24530_ (.RESET_B(net6769),
    .D(_01112_),
    .Q(\soc_inst.cpu_core.id_imm[24] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24531_ (.RESET_B(net6769),
    .D(_01113_),
    .Q(\soc_inst.cpu_core.id_imm[25] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24532_ (.RESET_B(net6774),
    .D(_01114_),
    .Q(\soc_inst.cpu_core.id_imm[26] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _24533_ (.RESET_B(net6769),
    .D(_01115_),
    .Q(\soc_inst.cpu_core.id_imm[27] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _24534_ (.RESET_B(net6774),
    .D(_01116_),
    .Q(\soc_inst.cpu_core.id_imm[28] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24535_ (.RESET_B(net6774),
    .D(_01117_),
    .Q(\soc_inst.cpu_core.id_imm[29] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24536_ (.RESET_B(net6777),
    .D(_01118_),
    .Q(\soc_inst.cpu_core.id_imm[30] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24537_ (.RESET_B(net6776),
    .D(net2666),
    .Q(\soc_inst.cpu_core.id_imm[31] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24538_ (.RESET_B(net6832),
    .D(_01120_),
    .Q(\soc_inst.cpu_core.mem_reg_we ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _24539_ (.RESET_B(net6801),
    .D(_01121_),
    .Q(\soc_inst.cpu_core.alu.op[0] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24540_ (.RESET_B(net6801),
    .D(_01122_),
    .Q(\soc_inst.cpu_core.alu.op[1] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24541_ (.RESET_B(net6801),
    .D(_01123_),
    .Q(\soc_inst.cpu_core.alu.op[2] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _24542_ (.RESET_B(net6801),
    .D(_01124_),
    .Q(\soc_inst.cpu_core.alu.op[3] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24543_ (.RESET_B(net6832),
    .D(_01125_),
    .Q(\soc_inst.cpu_core.alu.a[0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _24544_ (.RESET_B(net6801),
    .D(_01126_),
    .Q(\soc_inst.cpu_core.alu.a[1] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24545_ (.RESET_B(net6802),
    .D(_01127_),
    .Q(\soc_inst.cpu_core.alu.a[2] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24546_ (.RESET_B(net6803),
    .D(_01128_),
    .Q(\soc_inst.cpu_core.alu.a[3] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _24547_ (.RESET_B(net6832),
    .D(_01129_),
    .Q(\soc_inst.cpu_core.alu.a[4] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _24548_ (.RESET_B(net6804),
    .D(_01130_),
    .Q(\soc_inst.cpu_core.alu.a[5] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24549_ (.RESET_B(net6802),
    .D(_01131_),
    .Q(\soc_inst.cpu_core.alu.a[6] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _24550_ (.RESET_B(net6802),
    .D(_01132_),
    .Q(\soc_inst.cpu_core.alu.a[7] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _24551_ (.RESET_B(net6797),
    .D(_01133_),
    .Q(\soc_inst.cpu_core.alu.a[8] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _24552_ (.RESET_B(net6799),
    .D(_01134_),
    .Q(\soc_inst.cpu_core.alu.a[9] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _24553_ (.RESET_B(net6799),
    .D(_01135_),
    .Q(\soc_inst.cpu_core.alu.a[10] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24554_ (.RESET_B(net6799),
    .D(_01136_),
    .Q(\soc_inst.cpu_core.alu.a[11] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24555_ (.RESET_B(net6778),
    .D(_01137_),
    .Q(\soc_inst.cpu_core.alu.a[12] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24556_ (.RESET_B(net6778),
    .D(_01138_),
    .Q(\soc_inst.cpu_core.alu.a[13] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24557_ (.RESET_B(net6778),
    .D(_01139_),
    .Q(\soc_inst.cpu_core.alu.a[14] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24558_ (.RESET_B(net6776),
    .D(_01140_),
    .Q(\soc_inst.cpu_core.alu.a[15] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _24559_ (.RESET_B(net6772),
    .D(_01141_),
    .Q(\soc_inst.cpu_core.alu.a[16] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _24560_ (.RESET_B(net6806),
    .D(_01142_),
    .Q(\soc_inst.cpu_core.alu.a[17] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_2 _24561_ (.RESET_B(net6806),
    .D(_01143_),
    .Q(\soc_inst.cpu_core.alu.a[18] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _24562_ (.RESET_B(net6806),
    .D(_01144_),
    .Q(\soc_inst.cpu_core.alu.a[19] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _24563_ (.RESET_B(net6807),
    .D(_01145_),
    .Q(\soc_inst.cpu_core.alu.a[20] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _24564_ (.RESET_B(net6777),
    .D(_01146_),
    .Q(\soc_inst.cpu_core.alu.a[21] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24565_ (.RESET_B(net6807),
    .D(_01147_),
    .Q(\soc_inst.cpu_core.alu.a[22] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _24566_ (.RESET_B(net6778),
    .D(_01148_),
    .Q(\soc_inst.cpu_core.alu.a[23] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24567_ (.RESET_B(net6813),
    .D(_01149_),
    .Q(\soc_inst.cpu_core.alu.a[24] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _24568_ (.RESET_B(net6813),
    .D(_01150_),
    .Q(\soc_inst.cpu_core.alu.a[25] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _24569_ (.RESET_B(net6814),
    .D(_01151_),
    .Q(\soc_inst.cpu_core.alu.a[26] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _24570_ (.RESET_B(net6814),
    .D(_01152_),
    .Q(\soc_inst.cpu_core.alu.a[27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _24571_ (.RESET_B(net6814),
    .D(_01153_),
    .Q(\soc_inst.cpu_core.alu.a[28] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _24572_ (.RESET_B(net6834),
    .D(_01154_),
    .Q(\soc_inst.cpu_core.alu.a[29] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24573_ (.RESET_B(net6833),
    .D(_01155_),
    .Q(\soc_inst.cpu_core.alu.a[30] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _24574_ (.RESET_B(net6813),
    .D(_01156_),
    .Q(\soc_inst.cpu_core.alu.a[31] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _24575_ (.RESET_B(net6832),
    .D(_01157_),
    .Q(\soc_inst.cpu_core.alu.b[0] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _24576_ (.RESET_B(net6832),
    .D(_01158_),
    .Q(\soc_inst.cpu_core.alu.b[1] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _24577_ (.RESET_B(net6803),
    .D(net3391),
    .Q(\soc_inst.cpu_core.alu.b[2] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _24578_ (.RESET_B(net6834),
    .D(_01160_),
    .Q(\soc_inst.cpu_core.alu.b[3] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _24579_ (.RESET_B(net6832),
    .D(_01161_),
    .Q(\soc_inst.cpu_core.alu.b[4] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _24580_ (.RESET_B(net6803),
    .D(_01162_),
    .Q(\soc_inst.cpu_core.alu.b[5] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24581_ (.RESET_B(net6801),
    .D(net2974),
    .Q(\soc_inst.cpu_core.alu.b[6] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24582_ (.RESET_B(net6802),
    .D(_01164_),
    .Q(\soc_inst.cpu_core.alu.b[7] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _24583_ (.RESET_B(net6798),
    .D(_01165_),
    .Q(\soc_inst.cpu_core.alu.b[8] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _24584_ (.RESET_B(net6798),
    .D(_01166_),
    .Q(\soc_inst.cpu_core.alu.b[9] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24585_ (.RESET_B(net6796),
    .D(_01167_),
    .Q(\soc_inst.cpu_core.alu.b[10] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _24586_ (.RESET_B(net6799),
    .D(_01168_),
    .Q(\soc_inst.cpu_core.alu.b[11] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _24587_ (.RESET_B(net6777),
    .D(_01169_),
    .Q(\soc_inst.cpu_core.alu.b[12] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24588_ (.RESET_B(net6776),
    .D(_01170_),
    .Q(\soc_inst.cpu_core.alu.b[13] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24589_ (.RESET_B(net6777),
    .D(_01171_),
    .Q(\soc_inst.cpu_core.alu.b[14] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24590_ (.RESET_B(net6776),
    .D(_01172_),
    .Q(\soc_inst.cpu_core.alu.b[15] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24591_ (.RESET_B(net6773),
    .D(_01173_),
    .Q(\soc_inst.cpu_core.alu.b[16] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _24592_ (.RESET_B(net6773),
    .D(_01174_),
    .Q(\soc_inst.cpu_core.alu.b[17] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _24593_ (.RESET_B(net6773),
    .D(net3157),
    .Q(\soc_inst.cpu_core.alu.b[18] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _24594_ (.RESET_B(net6773),
    .D(_01176_),
    .Q(\soc_inst.cpu_core.alu.b[19] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _24595_ (.RESET_B(net6799),
    .D(net2952),
    .Q(\soc_inst.cpu_core.alu.b[20] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _24596_ (.RESET_B(net6815),
    .D(_01178_),
    .Q(\soc_inst.cpu_core.alu.b[21] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_2 _24597_ (.RESET_B(net6815),
    .D(_01179_),
    .Q(\soc_inst.cpu_core.alu.b[22] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _24598_ (.RESET_B(net6815),
    .D(_01180_),
    .Q(\soc_inst.cpu_core.alu.b[23] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _24599_ (.RESET_B(net6815),
    .D(_01181_),
    .Q(\soc_inst.cpu_core.alu.b[24] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _24600_ (.RESET_B(net6815),
    .D(_01182_),
    .Q(\soc_inst.cpu_core.alu.b[25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_2 _24601_ (.RESET_B(net6815),
    .D(_01183_),
    .Q(\soc_inst.cpu_core.alu.b[26] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_2 _24602_ (.RESET_B(net6814),
    .D(_01184_),
    .Q(\soc_inst.cpu_core.alu.b[27] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _24603_ (.RESET_B(net6814),
    .D(_01185_),
    .Q(\soc_inst.cpu_core.alu.b[28] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24604_ (.RESET_B(net6824),
    .D(_01186_),
    .Q(\soc_inst.cpu_core.alu.b[29] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _24605_ (.RESET_B(net6834),
    .D(_01187_),
    .Q(\soc_inst.cpu_core.alu.b[30] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _24606_ (.RESET_B(net6799),
    .D(_01188_),
    .Q(\soc_inst.cpu_core.alu.b[31] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24607_ (.RESET_B(net6803),
    .D(net3197),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[0] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _24608_ (.RESET_B(net6803),
    .D(_01190_),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _24609_ (.RESET_B(net6803),
    .D(net1594),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _24610_ (.RESET_B(net6832),
    .D(_01192_),
    .Q(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _24611_ (.RESET_B(net6794),
    .D(_01193_),
    .Q(\soc_inst.cpu_core.id_is_compressed ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _24612_ (.RESET_B(net6746),
    .D(_01194_),
    .Q(_00261_),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _24613_ (.RESET_B(net6746),
    .D(_01195_),
    .Q(_00262_),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24614_ (.RESET_B(net6746),
    .D(_01196_),
    .Q(\soc_inst.cpu_core.ex_instr[2] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24615_ (.RESET_B(net6781),
    .D(net3052),
    .Q(\soc_inst.cpu_core.ex_instr[3] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _24616_ (.RESET_B(net6744),
    .D(net2419),
    .Q(_00263_),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24617_ (.RESET_B(net6784),
    .D(_01199_),
    .Q(\soc_inst.cpu_core.ex_instr[5] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _24618_ (.RESET_B(net6798),
    .D(net2588),
    .Q(\soc_inst.cpu_core.ex_instr[6] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _24619_ (.RESET_B(net6794),
    .D(net2417),
    .Q(\soc_inst.cpu_core.ex_instr[7] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24620_ (.RESET_B(net6788),
    .D(_01202_),
    .Q(\soc_inst.cpu_core.ex_instr[8] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _24621_ (.RESET_B(net6788),
    .D(net2154),
    .Q(\soc_inst.cpu_core.ex_instr[9] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24622_ (.RESET_B(net6788),
    .D(_01204_),
    .Q(\soc_inst.cpu_core.ex_instr[10] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24623_ (.RESET_B(net6794),
    .D(_01205_),
    .Q(\soc_inst.cpu_core.ex_instr[11] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _24624_ (.RESET_B(net6780),
    .D(net2979),
    .Q(\soc_inst.cpu_core.ex_funct3[0] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _24625_ (.RESET_B(net6796),
    .D(net3029),
    .Q(\soc_inst.cpu_core.ex_funct3[1] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _24626_ (.RESET_B(net6745),
    .D(_01208_),
    .Q(\soc_inst.cpu_core.ex_funct3[2] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _24627_ (.RESET_B(net6776),
    .D(net361),
    .Q(\soc_inst.cpu_core.ex_instr[15] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _24628_ (.RESET_B(net6745),
    .D(net1351),
    .Q(\soc_inst.cpu_core.ex_instr[16] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24629_ (.RESET_B(net6734),
    .D(_01211_),
    .Q(\soc_inst.cpu_core.ex_instr[17] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _24630_ (.RESET_B(net6747),
    .D(net1364),
    .Q(\soc_inst.cpu_core.ex_instr[18] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _24631_ (.RESET_B(net6747),
    .D(net1865),
    .Q(\soc_inst.cpu_core.ex_instr[19] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24632_ (.RESET_B(net6758),
    .D(_01214_),
    .Q(\soc_inst.cpu_core.ex_instr[20] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24633_ (.RESET_B(net6765),
    .D(_01215_),
    .Q(\soc_inst.cpu_core.ex_instr[21] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_1 _24634_ (.RESET_B(net6728),
    .D(_01216_),
    .Q(\soc_inst.cpu_core.ex_instr[22] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24635_ (.RESET_B(net6763),
    .D(_01217_),
    .Q(\soc_inst.cpu_core.ex_instr[23] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_1 _24636_ (.RESET_B(net6730),
    .D(net2287),
    .Q(\soc_inst.cpu_core.ex_instr[24] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24637_ (.RESET_B(net6733),
    .D(_01219_),
    .Q(\soc_inst.cpu_core.ex_funct7[0] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_1 _24638_ (.RESET_B(net6732),
    .D(net2339),
    .Q(\soc_inst.cpu_core.ex_funct7[1] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24639_ (.RESET_B(net6731),
    .D(_01221_),
    .Q(\soc_inst.cpu_core.ex_funct7[2] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _24640_ (.RESET_B(net6762),
    .D(net2842),
    .Q(\soc_inst.cpu_core.ex_funct7[3] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_2 _24641_ (.RESET_B(net6734),
    .D(net2372),
    .Q(\soc_inst.cpu_core.ex_funct7[4] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _24642_ (.RESET_B(net6731),
    .D(_01224_),
    .Q(\soc_inst.cpu_core.ex_funct7[5] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _24643_ (.RESET_B(net6733),
    .D(_01225_),
    .Q(\soc_inst.cpu_core.ex_funct7[6] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _24644_ (.RESET_B(net6746),
    .D(net1673),
    .Q(\soc_inst.cpu_core.ex_exception_pc[0] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24645_ (.RESET_B(net6784),
    .D(net2369),
    .Q(\soc_inst.cpu_core.ex_exception_pc[1] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _24646_ (.RESET_B(net6782),
    .D(net2357),
    .Q(\soc_inst.cpu_core.ex_exception_pc[2] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _24647_ (.RESET_B(net6782),
    .D(net1924),
    .Q(\soc_inst.cpu_core.ex_exception_pc[3] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _24648_ (.RESET_B(net6782),
    .D(net2220),
    .Q(\soc_inst.cpu_core.ex_exception_pc[4] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _24649_ (.RESET_B(net6745),
    .D(net1269),
    .Q(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _24650_ (.RESET_B(net6744),
    .D(net1385),
    .Q(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _24651_ (.RESET_B(net6752),
    .D(net1698),
    .Q(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24652_ (.RESET_B(net6747),
    .D(net1882),
    .Q(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24653_ (.RESET_B(net6745),
    .D(net2103),
    .Q(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24654_ (.RESET_B(net6733),
    .D(net1402),
    .Q(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24655_ (.RESET_B(net6780),
    .D(net2293),
    .Q(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24656_ (.RESET_B(net6734),
    .D(net1454),
    .Q(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24657_ (.RESET_B(net6728),
    .D(net1868),
    .Q(\soc_inst.cpu_core.ex_exception_pc[13] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24658_ (.RESET_B(net6726),
    .D(net1383),
    .Q(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24659_ (.RESET_B(net6723),
    .D(net1823),
    .Q(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _24660_ (.RESET_B(net6726),
    .D(net2232),
    .Q(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _24661_ (.RESET_B(net6726),
    .D(net1779),
    .Q(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _24662_ (.RESET_B(net6726),
    .D(net2644),
    .Q(\soc_inst.cpu_core.ex_exception_pc[18] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24663_ (.RESET_B(net6726),
    .D(net1765),
    .Q(\soc_inst.cpu_core.ex_exception_pc[19] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24664_ (.RESET_B(net6723),
    .D(net1563),
    .Q(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24665_ (.RESET_B(net6723),
    .D(net1802),
    .Q(\soc_inst.cpu_core.ex_exception_pc[21] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24666_ (.RESET_B(net6726),
    .D(net1854),
    .Q(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24667_ (.RESET_B(net6723),
    .D(net1669),
    .Q(\soc_inst.cpu_core.ex_exception_pc[23] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24668_ (.RESET_B(net6684),
    .D(_00024_),
    .Q(\soc_inst.core_mem_re ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24669_ (.RESET_B(net6748),
    .D(net645),
    .Q(\soc_inst.cpu_core.ex_rs1_data[0] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _24670_ (.RESET_B(net6746),
    .D(net395),
    .Q(\soc_inst.cpu_core.ex_rs1_data[1] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24671_ (.RESET_B(net6741),
    .D(net2044),
    .Q(\soc_inst.cpu_core.ex_rs1_data[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _24672_ (.RESET_B(net6748),
    .D(net317),
    .Q(\soc_inst.cpu_core.ex_rs1_data[3] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _24673_ (.RESET_B(net6744),
    .D(net258),
    .Q(\soc_inst.cpu_core.ex_rs1_data[4] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24674_ (.RESET_B(net6750),
    .D(net520),
    .Q(\soc_inst.cpu_core.ex_rs1_data[5] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _24675_ (.RESET_B(net6706),
    .D(net456),
    .Q(\soc_inst.cpu_core.ex_rs1_data[6] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24676_ (.RESET_B(net6739),
    .D(net1198),
    .Q(\soc_inst.cpu_core.ex_rs1_data[7] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _24677_ (.RESET_B(net6729),
    .D(net261),
    .Q(\soc_inst.cpu_core.ex_rs1_data[8] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_1 _24678_ (.RESET_B(net6743),
    .D(net207),
    .Q(\soc_inst.cpu_core.ex_rs1_data[9] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24679_ (.RESET_B(net6729),
    .D(net244),
    .Q(\soc_inst.cpu_core.ex_rs1_data[10] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24680_ (.RESET_B(net6729),
    .D(net327),
    .Q(\soc_inst.cpu_core.ex_rs1_data[11] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24681_ (.RESET_B(net6668),
    .D(net232),
    .Q(\soc_inst.cpu_core.ex_rs1_data[12] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24682_ (.RESET_B(net6681),
    .D(net289),
    .Q(\soc_inst.cpu_core.ex_rs1_data[13] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24683_ (.RESET_B(net6709),
    .D(net368),
    .Q(\soc_inst.cpu_core.ex_rs1_data[14] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24684_ (.RESET_B(net6716),
    .D(net730),
    .Q(\soc_inst.cpu_core.ex_rs1_data[15] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _24685_ (.RESET_B(net6727),
    .D(net276),
    .Q(\soc_inst.cpu_core.ex_rs1_data[16] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_1 _24686_ (.RESET_B(net6724),
    .D(net218),
    .Q(\soc_inst.cpu_core.ex_rs1_data[17] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24687_ (.RESET_B(net6756),
    .D(net1034),
    .Q(\soc_inst.cpu_core.ex_rs1_data[18] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _24688_ (.RESET_B(net6725),
    .D(net525),
    .Q(\soc_inst.cpu_core.ex_rs1_data[19] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_1 _24689_ (.RESET_B(net6756),
    .D(net892),
    .Q(\soc_inst.cpu_core.ex_rs1_data[20] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _24690_ (.RESET_B(net6756),
    .D(net2224),
    .Q(\soc_inst.cpu_core.ex_rs1_data[21] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _24691_ (.RESET_B(net6757),
    .D(net886),
    .Q(\soc_inst.cpu_core.ex_rs1_data[22] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _24692_ (.RESET_B(net6756),
    .D(net1369),
    .Q(\soc_inst.cpu_core.ex_rs1_data[23] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_2 _24693_ (.RESET_B(net6759),
    .D(net1280),
    .Q(\soc_inst.cpu_core.ex_rs1_data[24] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _24694_ (.RESET_B(net6726),
    .D(net733),
    .Q(\soc_inst.cpu_core.ex_rs1_data[25] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24695_ (.RESET_B(net6771),
    .D(net215),
    .Q(\soc_inst.cpu_core.ex_rs1_data[26] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _24696_ (.RESET_B(net6723),
    .D(net321),
    .Q(\soc_inst.cpu_core.ex_rs1_data[27] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24697_ (.RESET_B(net6756),
    .D(net329),
    .Q(\soc_inst.cpu_core.ex_rs1_data[28] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _24698_ (.RESET_B(net6756),
    .D(net2823),
    .Q(\soc_inst.cpu_core.ex_rs1_data[29] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24699_ (.RESET_B(net6723),
    .D(net375),
    .Q(\soc_inst.cpu_core.ex_rs1_data[30] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24700_ (.RESET_B(net6761),
    .D(net382),
    .Q(\soc_inst.cpu_core.ex_rs1_data[31] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _24701_ (.RESET_B(net6703),
    .D(_01282_),
    .Q(\soc_inst.core_mem_addr[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24702_ (.RESET_B(net6698),
    .D(_01283_),
    .Q(\soc_inst.core_mem_addr[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _24703_ (.RESET_B(net6687),
    .D(net3267),
    .Q(\soc_inst.core_mem_addr[2] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _24704_ (.RESET_B(net6684),
    .D(_01285_),
    .Q(\soc_inst.core_mem_addr[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24705_ (.RESET_B(net6698),
    .D(net2909),
    .Q(\soc_inst.pwm_inst.channel_idx [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _24706_ (.RESET_B(net6698),
    .D(_01287_),
    .Q(\soc_inst.core_mem_addr[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _24707_ (.RESET_B(net6698),
    .D(_01288_),
    .Q(\soc_inst.core_mem_addr[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _24708_ (.RESET_B(net6698),
    .D(_01289_),
    .Q(\soc_inst.core_mem_addr[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _24709_ (.RESET_B(net6678),
    .D(net1052),
    .Q(\soc_inst.core_mem_addr[8] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24710_ (.RESET_B(net6699),
    .D(net1928),
    .Q(\soc_inst.core_mem_addr[9] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24711_ (.RESET_B(net6678),
    .D(net1111),
    .Q(\soc_inst.core_mem_addr[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _24712_ (.RESET_B(net6669),
    .D(net1539),
    .Q(\soc_inst.core_mem_addr[11] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24713_ (.RESET_B(net6767),
    .D(net2801),
    .Q(\soc_inst.core_mem_addr[12] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24714_ (.RESET_B(net6666),
    .D(net3288),
    .Q(\soc_inst.core_mem_addr[13] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _24715_ (.RESET_B(net6666),
    .D(net3264),
    .Q(\soc_inst.core_mem_addr[14] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _24716_ (.RESET_B(net6669),
    .D(net2366),
    .Q(\soc_inst.core_mem_addr[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24717_ (.RESET_B(net6731),
    .D(_01298_),
    .Q(\soc_inst.core_mem_addr[16] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24718_ (.RESET_B(net6668),
    .D(net2857),
    .Q(\soc_inst.core_mem_addr[17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _24719_ (.RESET_B(net6668),
    .D(net2837),
    .Q(\soc_inst.core_mem_addr[18] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _24720_ (.RESET_B(net6659),
    .D(net2688),
    .Q(\soc_inst.core_mem_addr[19] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_2 _24721_ (.RESET_B(net6668),
    .D(net2806),
    .Q(\soc_inst.core_mem_addr[20] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _24722_ (.RESET_B(net6668),
    .D(_01303_),
    .Q(\soc_inst.core_mem_addr[21] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _24723_ (.RESET_B(net6666),
    .D(net2695),
    .Q(\soc_inst.core_mem_addr[22] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_2 _24724_ (.RESET_B(net6668),
    .D(net2903),
    .Q(\soc_inst.core_mem_addr[23] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _24725_ (.RESET_B(net6685),
    .D(net2732),
    .Q(\soc_inst.core_mem_addr[24] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _24726_ (.RESET_B(net6684),
    .D(net2848),
    .Q(\soc_inst.core_mem_addr[25] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _24727_ (.RESET_B(net6685),
    .D(net2734),
    .Q(\soc_inst.core_mem_addr[26] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24728_ (.RESET_B(net6685),
    .D(net2758),
    .Q(\soc_inst.core_mem_addr[27] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _24729_ (.RESET_B(net6679),
    .D(net2631),
    .Q(\soc_inst.core_mem_addr[28] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _24730_ (.RESET_B(net6699),
    .D(net2546),
    .Q(\soc_inst.core_mem_addr[29] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24731_ (.RESET_B(net6686),
    .D(net2702),
    .Q(\soc_inst.core_mem_addr[30] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24732_ (.RESET_B(net6699),
    .D(net404),
    .Q(\soc_inst.core_mem_addr[31] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _24733_ (.RESET_B(net6579),
    .D(_01314_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _24734_ (.RESET_B(net6594),
    .D(_01315_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _24735_ (.RESET_B(net6704),
    .D(_01316_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[2] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24736_ (.RESET_B(net6579),
    .D(net399),
    .Q(\soc_inst.cpu_core.ex_rs2_data[3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24737_ (.RESET_B(net6594),
    .D(net252),
    .Q(\soc_inst.cpu_core.ex_rs2_data[4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _24738_ (.RESET_B(net6596),
    .D(net639),
    .Q(\soc_inst.cpu_core.ex_rs2_data[5] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24739_ (.RESET_B(net6594),
    .D(net298),
    .Q(\soc_inst.cpu_core.ex_rs2_data[6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _24740_ (.RESET_B(net6633),
    .D(net858),
    .Q(\soc_inst.cpu_core.ex_rs2_data[7] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _24741_ (.RESET_B(net6626),
    .D(net256),
    .Q(\soc_inst.cpu_core.ex_rs2_data[8] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _24742_ (.RESET_B(net6610),
    .D(net927),
    .Q(\soc_inst.cpu_core.ex_rs2_data[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _24743_ (.RESET_B(net6667),
    .D(net294),
    .Q(\soc_inst.cpu_core.ex_rs2_data[10] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _24744_ (.RESET_B(net6604),
    .D(_01325_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[11] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _24745_ (.RESET_B(net6666),
    .D(net1800),
    .Q(\soc_inst.cpu_core.ex_rs2_data[12] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _24746_ (.RESET_B(net6564),
    .D(net240),
    .Q(\soc_inst.cpu_core.ex_rs2_data[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _24747_ (.RESET_B(net6559),
    .D(net337),
    .Q(\soc_inst.cpu_core.ex_rs2_data[14] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _24748_ (.RESET_B(net6663),
    .D(net1549),
    .Q(\soc_inst.cpu_core.ex_rs2_data[15] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _24749_ (.RESET_B(net6619),
    .D(net325),
    .Q(\soc_inst.cpu_core.ex_rs2_data[16] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24750_ (.RESET_B(net6619),
    .D(net567),
    .Q(\soc_inst.cpu_core.ex_rs2_data[17] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24751_ (.RESET_B(net6671),
    .D(net511),
    .Q(\soc_inst.cpu_core.ex_rs2_data[18] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _24752_ (.RESET_B(net6657),
    .D(net688),
    .Q(\soc_inst.cpu_core.ex_rs2_data[19] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24753_ (.RESET_B(net6657),
    .D(net1977),
    .Q(\soc_inst.cpu_core.ex_rs2_data[20] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24754_ (.RESET_B(net6661),
    .D(net523),
    .Q(\soc_inst.cpu_core.ex_rs2_data[21] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24755_ (.RESET_B(net6658),
    .D(net587),
    .Q(\soc_inst.cpu_core.ex_rs2_data[22] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24756_ (.RESET_B(net6661),
    .D(net274),
    .Q(\soc_inst.cpu_core.ex_rs2_data[23] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _24757_ (.RESET_B(net6620),
    .D(net348),
    .Q(\soc_inst.cpu_core.ex_rs2_data[24] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24758_ (.RESET_B(net6620),
    .D(net2574),
    .Q(\soc_inst.cpu_core.ex_rs2_data[25] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _24759_ (.RESET_B(net6660),
    .D(net209),
    .Q(\soc_inst.cpu_core.ex_rs2_data[26] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _24760_ (.RESET_B(net6660),
    .D(net473),
    .Q(\soc_inst.cpu_core.ex_rs2_data[27] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24761_ (.RESET_B(net6615),
    .D(_01342_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[28] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _24762_ (.RESET_B(net6615),
    .D(_01343_),
    .Q(\soc_inst.cpu_core.ex_rs2_data[29] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _24763_ (.RESET_B(net6657),
    .D(net1796),
    .Q(\soc_inst.cpu_core.ex_rs2_data[30] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24764_ (.RESET_B(net6659),
    .D(net427),
    .Q(\soc_inst.cpu_core.ex_rs2_data[31] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24765_ (.RESET_B(net6797),
    .D(net2815),
    .Q(\soc_inst.cpu_core.ex_alu_result[0] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _24766_ (.RESET_B(net6833),
    .D(net3206),
    .Q(\soc_inst.cpu_core.ex_alu_result[1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _24767_ (.RESET_B(net6804),
    .D(_01348_),
    .Q(\soc_inst.cpu_core.ex_alu_result[2] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24768_ (.RESET_B(net6834),
    .D(net3280),
    .Q(\soc_inst.cpu_core.ex_alu_result[3] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _24769_ (.RESET_B(net6834),
    .D(net3111),
    .Q(\soc_inst.cpu_core.ex_alu_result[4] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _24770_ (.RESET_B(net6749),
    .D(_01351_),
    .Q(\soc_inst.cpu_core.ex_alu_result[5] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24771_ (.RESET_B(net6749),
    .D(_01352_),
    .Q(\soc_inst.cpu_core.ex_alu_result[6] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _24772_ (.RESET_B(net6798),
    .D(_01353_),
    .Q(\soc_inst.cpu_core.ex_alu_result[7] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _24773_ (.RESET_B(net6796),
    .D(net3216),
    .Q(\soc_inst.cpu_core.ex_alu_result[8] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _24774_ (.RESET_B(net6797),
    .D(net3161),
    .Q(\soc_inst.cpu_core.ex_alu_result[9] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _24775_ (.RESET_B(net6799),
    .D(_01356_),
    .Q(\soc_inst.cpu_core.ex_alu_result[10] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _24776_ (.RESET_B(net6799),
    .D(net3211),
    .Q(\soc_inst.cpu_core.ex_alu_result[11] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _24777_ (.RESET_B(net6777),
    .D(_01358_),
    .Q(\soc_inst.cpu_core.ex_alu_result[12] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24778_ (.RESET_B(net6767),
    .D(net3292),
    .Q(\soc_inst.cpu_core.ex_alu_result[13] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24779_ (.RESET_B(net6778),
    .D(_01360_),
    .Q(\soc_inst.cpu_core.ex_alu_result[14] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_2 _24780_ (.RESET_B(net6762),
    .D(_01361_),
    .Q(\soc_inst.cpu_core.ex_alu_result[15] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _24781_ (.RESET_B(net6777),
    .D(_01362_),
    .Q(\soc_inst.cpu_core.ex_alu_result[16] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24782_ (.RESET_B(net6776),
    .D(_01363_),
    .Q(\soc_inst.cpu_core.ex_alu_result[17] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24783_ (.RESET_B(net6763),
    .D(_01364_),
    .Q(\soc_inst.cpu_core.ex_alu_result[18] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_2 _24784_ (.RESET_B(net6774),
    .D(_01365_),
    .Q(\soc_inst.cpu_core.ex_alu_result[19] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _24785_ (.RESET_B(net6763),
    .D(_01366_),
    .Q(\soc_inst.cpu_core.ex_alu_result[20] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24786_ (.RESET_B(net6765),
    .D(_01367_),
    .Q(\soc_inst.cpu_core.ex_alu_result[21] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24787_ (.RESET_B(net6764),
    .D(_01368_),
    .Q(\soc_inst.cpu_core.ex_alu_result[22] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _24788_ (.RESET_B(net6776),
    .D(_01369_),
    .Q(\soc_inst.cpu_core.ex_alu_result[23] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _24789_ (.RESET_B(net6740),
    .D(_01370_),
    .Q(\soc_inst.cpu_core.ex_alu_result[24] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24790_ (.RESET_B(net6733),
    .D(_01371_),
    .Q(\soc_inst.cpu_core.ex_alu_result[25] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _24791_ (.RESET_B(net6814),
    .D(_01372_),
    .Q(\soc_inst.cpu_core.ex_alu_result[26] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24792_ (.RESET_B(net6777),
    .D(_01373_),
    .Q(\soc_inst.cpu_core.ex_alu_result[27] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_2 _24793_ (.RESET_B(net6761),
    .D(_01374_),
    .Q(\soc_inst.cpu_core.ex_alu_result[28] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _24794_ (.RESET_B(net6747),
    .D(_01375_),
    .Q(\soc_inst.cpu_core.ex_alu_result[29] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24795_ (.RESET_B(net6796),
    .D(_01376_),
    .Q(\soc_inst.cpu_core.ex_alu_result[30] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24796_ (.RESET_B(net6780),
    .D(_01377_),
    .Q(\soc_inst.cpu_core.ex_alu_result[31] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _24797_ (.RESET_B(net6688),
    .D(_00025_),
    .Q(\soc_inst.core_mem_we ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24798_ (.RESET_B(net6781),
    .D(_01378_),
    .Q(\soc_inst.cpu_core.ex_mem_we ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24799_ (.RESET_B(net6790),
    .D(net1252),
    .Q(\soc_inst.cpu_core.ex_mem_re ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24800_ (.RESET_B(net6840),
    .D(_01380_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][0] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _24801_ (.RESET_B(net6842),
    .D(_01381_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _24802_ (.RESET_B(net6835),
    .D(_01382_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][2] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _24803_ (.RESET_B(net6821),
    .D(_01383_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][3] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _24804_ (.RESET_B(net6876),
    .D(_01384_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][4] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24805_ (.RESET_B(net6952),
    .D(_01385_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _24806_ (.RESET_B(net6905),
    .D(_01386_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _24807_ (.RESET_B(net6926),
    .D(_01387_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][7] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _24808_ (.RESET_B(net6899),
    .D(_01388_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][8] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _24809_ (.RESET_B(net6959),
    .D(_01389_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][9] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _24810_ (.RESET_B(net6969),
    .D(_01390_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _24811_ (.RESET_B(net6890),
    .D(_01391_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _24812_ (.RESET_B(net6949),
    .D(_01392_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][12] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _24813_ (.RESET_B(net6931),
    .D(_01393_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _24814_ (.RESET_B(net6808),
    .D(_01394_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][14] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _24815_ (.RESET_B(net6946),
    .D(_01395_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][15] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _24816_ (.RESET_B(net6916),
    .D(_01396_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][16] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _24817_ (.RESET_B(net6854),
    .D(_01397_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][17] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _24818_ (.RESET_B(net6937),
    .D(_01398_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][18] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _24819_ (.RESET_B(net6870),
    .D(_01399_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _24820_ (.RESET_B(net6979),
    .D(_01400_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][20] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24821_ (.RESET_B(net6912),
    .D(_01401_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][21] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _24822_ (.RESET_B(net6827),
    .D(_01402_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _24823_ (.RESET_B(net6980),
    .D(_01403_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][23] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24824_ (.RESET_B(net6859),
    .D(_01404_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][24] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _24825_ (.RESET_B(net6810),
    .D(_01405_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][25] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _24826_ (.RESET_B(net6918),
    .D(_01406_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][26] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _24827_ (.RESET_B(net6828),
    .D(_01407_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _24828_ (.RESET_B(net6856),
    .D(_01408_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _24829_ (.RESET_B(net6888),
    .D(_01409_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][29] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _24830_ (.RESET_B(net6974),
    .D(_01410_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][30] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _24831_ (.RESET_B(net6955),
    .D(_01411_),
    .Q(\soc_inst.cpu_core.register_file.registers[22][31] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _24832_ (.RESET_B(net6845),
    .D(_01412_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][0] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _24833_ (.RESET_B(net6843),
    .D(_01413_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _24834_ (.RESET_B(net6885),
    .D(_01414_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][2] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _24835_ (.RESET_B(net6821),
    .D(_01415_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][3] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _24836_ (.RESET_B(net6878),
    .D(_01416_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][4] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _24837_ (.RESET_B(net6901),
    .D(_01417_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _24838_ (.RESET_B(net6908),
    .D(_01418_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _24839_ (.RESET_B(net6929),
    .D(_01419_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][7] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _24840_ (.RESET_B(net6889),
    .D(_01420_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][8] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _24841_ (.RESET_B(net6961),
    .D(_01421_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][9] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _24842_ (.RESET_B(net6966),
    .D(_01422_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _24843_ (.RESET_B(net6895),
    .D(_01423_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][11] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _24844_ (.RESET_B(net6950),
    .D(_01424_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _24845_ (.RESET_B(net6935),
    .D(_01425_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _24846_ (.RESET_B(net6817),
    .D(_01426_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][14] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _24847_ (.RESET_B(net6946),
    .D(_01427_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][15] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _24848_ (.RESET_B(net6916),
    .D(_01428_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _24849_ (.RESET_B(net6854),
    .D(_01429_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _24850_ (.RESET_B(net6937),
    .D(_01430_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _24851_ (.RESET_B(net6869),
    .D(_01431_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][19] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _24852_ (.RESET_B(net6979),
    .D(_01432_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][20] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24853_ (.RESET_B(net6909),
    .D(_01433_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][21] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _24854_ (.RESET_B(net6827),
    .D(_01434_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _24855_ (.RESET_B(net6981),
    .D(_01435_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24856_ (.RESET_B(net6860),
    .D(_01436_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][24] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24857_ (.RESET_B(net6818),
    .D(_01437_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][25] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _24858_ (.RESET_B(net6924),
    .D(_01438_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _24859_ (.RESET_B(net6828),
    .D(_01439_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][27] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _24860_ (.RESET_B(net6856),
    .D(_01440_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][28] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _24861_ (.RESET_B(net6883),
    .D(_01441_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][29] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _24862_ (.RESET_B(net6976),
    .D(_01442_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _24863_ (.RESET_B(net6954),
    .D(_01443_),
    .Q(\soc_inst.cpu_core.register_file.registers[21][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _24864_ (.RESET_B(net6846),
    .D(_01444_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][0] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24865_ (.RESET_B(net6846),
    .D(_01445_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _24866_ (.RESET_B(net6837),
    .D(_01446_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _24867_ (.RESET_B(net6851),
    .D(_01447_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][3] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24868_ (.RESET_B(net6878),
    .D(_01448_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][4] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24869_ (.RESET_B(net6901),
    .D(_01449_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24870_ (.RESET_B(net6905),
    .D(_01450_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][6] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _24871_ (.RESET_B(net6926),
    .D(_01451_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][7] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _24872_ (.RESET_B(net6899),
    .D(_01452_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24873_ (.RESET_B(net6957),
    .D(_01453_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][9] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _24874_ (.RESET_B(net6965),
    .D(_01454_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][10] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24875_ (.RESET_B(net6892),
    .D(_01455_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][11] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _24876_ (.RESET_B(net6943),
    .D(_01456_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _24877_ (.RESET_B(net6940),
    .D(_01457_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][13] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24878_ (.RESET_B(net6819),
    .D(_01458_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][14] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _24879_ (.RESET_B(net6941),
    .D(_01459_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][15] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _24880_ (.RESET_B(net6922),
    .D(_01460_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][16] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24881_ (.RESET_B(net6867),
    .D(_01461_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][17] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _24882_ (.RESET_B(net6923),
    .D(_01462_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][18] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _24883_ (.RESET_B(net6873),
    .D(_01463_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24884_ (.RESET_B(net6968),
    .D(_01464_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _24885_ (.RESET_B(net6909),
    .D(_01465_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][21] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _24886_ (.RESET_B(net6826),
    .D(_01466_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _24887_ (.RESET_B(net6982),
    .D(_01467_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24888_ (.RESET_B(net6862),
    .D(_01468_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][24] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24889_ (.RESET_B(net6819),
    .D(_01469_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][25] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _24890_ (.RESET_B(net6919),
    .D(_01470_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][26] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _24891_ (.RESET_B(net6838),
    .D(_01471_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][27] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _24892_ (.RESET_B(net6863),
    .D(_01472_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24893_ (.RESET_B(net6882),
    .D(_01473_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][29] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _24894_ (.RESET_B(net6974),
    .D(_01474_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][30] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24895_ (.RESET_B(net6953),
    .D(_01475_),
    .Q(\soc_inst.cpu_core.register_file.registers[20][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _24896_ (.RESET_B(net6892),
    .D(_01476_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _24897_ (.RESET_B(net6843),
    .D(_01477_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _24898_ (.RESET_B(net6892),
    .D(_01478_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24899_ (.RESET_B(net6852),
    .D(_01479_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][3] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _24900_ (.RESET_B(net6876),
    .D(_01480_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][4] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _24901_ (.RESET_B(net6903),
    .D(_01481_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24902_ (.RESET_B(net6907),
    .D(_01482_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][6] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _24903_ (.RESET_B(net6926),
    .D(_01483_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _24904_ (.RESET_B(net6898),
    .D(_01484_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][8] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _24905_ (.RESET_B(net6959),
    .D(_01485_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][9] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _24906_ (.RESET_B(net6969),
    .D(_01486_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _24907_ (.RESET_B(net6894),
    .D(_01487_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][11] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _24908_ (.RESET_B(net6948),
    .D(_01488_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24909_ (.RESET_B(net6936),
    .D(_01489_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][13] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24910_ (.RESET_B(net6808),
    .D(_01490_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][14] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _24911_ (.RESET_B(net6942),
    .D(_01491_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24912_ (.RESET_B(net6920),
    .D(_01492_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][16] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _24913_ (.RESET_B(net6856),
    .D(_01493_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][17] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _24914_ (.RESET_B(net6933),
    .D(_01494_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][18] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24915_ (.RESET_B(net6869),
    .D(_01495_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][19] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _24916_ (.RESET_B(net6971),
    .D(_01496_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _24917_ (.RESET_B(net6913),
    .D(_01497_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][21] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _24918_ (.RESET_B(net6823),
    .D(_01498_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][22] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_2 _24919_ (.RESET_B(net6978),
    .D(_01499_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _24920_ (.RESET_B(net6877),
    .D(_01500_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][24] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24921_ (.RESET_B(net6818),
    .D(_01501_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][25] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _24922_ (.RESET_B(net6925),
    .D(_01502_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _24923_ (.RESET_B(net6828),
    .D(_01503_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][27] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _24924_ (.RESET_B(net6874),
    .D(_01504_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _24925_ (.RESET_B(net6861),
    .D(_01505_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][29] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _24926_ (.RESET_B(net6976),
    .D(_01506_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _24927_ (.RESET_B(net6956),
    .D(_01507_),
    .Q(\soc_inst.cpu_core.register_file.registers[27][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _24928_ (.RESET_B(net6846),
    .D(_01508_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][0] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24929_ (.RESET_B(net6844),
    .D(_01509_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][1] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _24930_ (.RESET_B(net6884),
    .D(_01510_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][2] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _24931_ (.RESET_B(net6821),
    .D(_01511_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][3] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _24932_ (.RESET_B(net6879),
    .D(_01512_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][4] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _24933_ (.RESET_B(net6903),
    .D(_01513_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24934_ (.RESET_B(net6907),
    .D(_01514_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][6] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _24935_ (.RESET_B(net6928),
    .D(_01515_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][7] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _24936_ (.RESET_B(net6898),
    .D(_01516_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][8] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _24937_ (.RESET_B(net6963),
    .D(_01517_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][9] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24938_ (.RESET_B(net6970),
    .D(_01518_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _24939_ (.RESET_B(net6894),
    .D(_01519_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][11] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _24940_ (.RESET_B(net6943),
    .D(_01520_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _24941_ (.RESET_B(net6931),
    .D(_01521_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _24942_ (.RESET_B(net6808),
    .D(_01522_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][14] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _24943_ (.RESET_B(net6941),
    .D(_01523_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][15] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _24944_ (.RESET_B(net6920),
    .D(_01524_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][16] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _24945_ (.RESET_B(net6855),
    .D(_01525_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][17] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24946_ (.RESET_B(net6933),
    .D(_01526_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][18] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24947_ (.RESET_B(net6870),
    .D(_01527_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _24948_ (.RESET_B(net6972),
    .D(_01528_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _24949_ (.RESET_B(net6913),
    .D(_01529_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][21] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _24950_ (.RESET_B(net6827),
    .D(_01530_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][22] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _24951_ (.RESET_B(net6982),
    .D(_01531_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24952_ (.RESET_B(net6859),
    .D(_01532_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][24] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _24953_ (.RESET_B(net6810),
    .D(_01533_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][25] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24954_ (.RESET_B(net6924),
    .D(_01534_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _24955_ (.RESET_B(net6824),
    .D(_01535_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][27] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _24956_ (.RESET_B(net6856),
    .D(_01536_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][28] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _24957_ (.RESET_B(net6883),
    .D(_01537_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][29] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _24958_ (.RESET_B(net6977),
    .D(_01538_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][30] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24959_ (.RESET_B(net6953),
    .D(_01539_),
    .Q(\soc_inst.cpu_core.register_file.registers[19][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _24960_ (.RESET_B(net6890),
    .D(_01540_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][0] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _24961_ (.RESET_B(net6845),
    .D(_01541_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _24962_ (.RESET_B(net6836),
    .D(_01542_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][2] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _24963_ (.RESET_B(net6821),
    .D(_01543_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _24964_ (.RESET_B(net6879),
    .D(_01544_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _24965_ (.RESET_B(net6901),
    .D(_01545_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][5] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _24966_ (.RESET_B(net6907),
    .D(_01546_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][6] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _24967_ (.RESET_B(net6929),
    .D(_01547_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][7] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24968_ (.RESET_B(net6898),
    .D(_01548_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][8] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _24969_ (.RESET_B(net6957),
    .D(_01549_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][9] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _24970_ (.RESET_B(net6965),
    .D(_01550_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _24971_ (.RESET_B(net6895),
    .D(_01551_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][11] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _24972_ (.RESET_B(net6943),
    .D(_01552_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _24973_ (.RESET_B(net6931),
    .D(_01553_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][13] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24974_ (.RESET_B(net6817),
    .D(_01554_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][14] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _24975_ (.RESET_B(net6942),
    .D(_01555_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][15] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _24976_ (.RESET_B(net6916),
    .D(_01556_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _24977_ (.RESET_B(net6854),
    .D(_01557_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _24978_ (.RESET_B(net6932),
    .D(_01558_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][18] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _24979_ (.RESET_B(net6871),
    .D(_01559_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][19] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24980_ (.RESET_B(net6967),
    .D(_01560_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _24981_ (.RESET_B(net6912),
    .D(_01561_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][21] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _24982_ (.RESET_B(net6826),
    .D(_01562_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _24983_ (.RESET_B(net6982),
    .D(_01563_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24984_ (.RESET_B(net6859),
    .D(_01564_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][24] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _24985_ (.RESET_B(net6818),
    .D(_01565_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][25] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _24986_ (.RESET_B(net6918),
    .D(_01566_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][26] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24987_ (.RESET_B(net6824),
    .D(_01567_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _24988_ (.RESET_B(net6863),
    .D(_01568_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][28] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _24989_ (.RESET_B(net6882),
    .D(_01569_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _24990_ (.RESET_B(net6975),
    .D(_01570_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _24991_ (.RESET_B(net6954),
    .D(_01571_),
    .Q(\soc_inst.cpu_core.register_file.registers[18][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _24992_ (.RESET_B(net6840),
    .D(_01572_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][0] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _24993_ (.RESET_B(net6842),
    .D(_01573_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _24994_ (.RESET_B(net6835),
    .D(_01574_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][2] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24995_ (.RESET_B(net6849),
    .D(_01575_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _24996_ (.RESET_B(net6900),
    .D(_01576_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][4] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _24997_ (.RESET_B(net6952),
    .D(_01577_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _24998_ (.RESET_B(net6907),
    .D(_01578_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _24999_ (.RESET_B(net6926),
    .D(_01579_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][7] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25000_ (.RESET_B(net6900),
    .D(_01580_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _25001_ (.RESET_B(net6959),
    .D(_01581_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][9] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25002_ (.RESET_B(net6966),
    .D(_01582_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25003_ (.RESET_B(net6891),
    .D(_01583_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][11] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _25004_ (.RESET_B(net6944),
    .D(_01584_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25005_ (.RESET_B(net6932),
    .D(_01585_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][13] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _25006_ (.RESET_B(net6808),
    .D(_01586_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][14] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25007_ (.RESET_B(net6942),
    .D(_01587_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _25008_ (.RESET_B(net6921),
    .D(_01588_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _25009_ (.RESET_B(net6854),
    .D(_01589_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25010_ (.RESET_B(net6934),
    .D(_01590_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][18] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _25011_ (.RESET_B(net6870),
    .D(_01591_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25012_ (.RESET_B(net6967),
    .D(_01592_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25013_ (.RESET_B(net6911),
    .D(_01593_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][21] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25014_ (.RESET_B(net6823),
    .D(_01594_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_2 _25015_ (.RESET_B(net6982),
    .D(_01595_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25016_ (.RESET_B(net6861),
    .D(_01596_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25017_ (.RESET_B(net6810),
    .D(_01597_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25018_ (.RESET_B(net6918),
    .D(_01598_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][26] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25019_ (.RESET_B(net6829),
    .D(_01599_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][27] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25020_ (.RESET_B(net6866),
    .D(_01600_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _25021_ (.RESET_B(net6883),
    .D(_01601_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][29] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _25022_ (.RESET_B(net6976),
    .D(_01602_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25023_ (.RESET_B(net6953),
    .D(_01603_),
    .Q(\soc_inst.cpu_core.register_file.registers[17][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _25024_ (.RESET_B(net6846),
    .D(_01604_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _25025_ (.RESET_B(net6843),
    .D(_01605_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25026_ (.RESET_B(net6835),
    .D(_01606_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][2] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _25027_ (.RESET_B(net6821),
    .D(_01607_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][3] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25028_ (.RESET_B(net6879),
    .D(_01608_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][4] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25029_ (.RESET_B(net6902),
    .D(_01609_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][5] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25030_ (.RESET_B(net6908),
    .D(_01610_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25031_ (.RESET_B(net6928),
    .D(_01611_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25032_ (.RESET_B(net6899),
    .D(_01612_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _25033_ (.RESET_B(net6958),
    .D(_01613_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][9] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25034_ (.RESET_B(net6969),
    .D(_01614_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25035_ (.RESET_B(net6891),
    .D(_01615_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][11] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _25036_ (.RESET_B(net6944),
    .D(_01616_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _25037_ (.RESET_B(net6935),
    .D(_01617_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _25038_ (.RESET_B(net6808),
    .D(_01618_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][14] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _25039_ (.RESET_B(net6947),
    .D(_01619_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25040_ (.RESET_B(net6922),
    .D(_01620_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25041_ (.RESET_B(net6865),
    .D(_01621_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25042_ (.RESET_B(net6933),
    .D(_01622_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][18] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25043_ (.RESET_B(net6869),
    .D(_01623_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][19] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _25044_ (.RESET_B(net6971),
    .D(_01624_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _25045_ (.RESET_B(net6912),
    .D(_01625_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][21] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25046_ (.RESET_B(net6851),
    .D(_01626_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][22] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25047_ (.RESET_B(net6980),
    .D(_01627_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25048_ (.RESET_B(net6860),
    .D(_01628_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][24] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25049_ (.RESET_B(net6816),
    .D(_01629_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][25] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _25050_ (.RESET_B(net6880),
    .D(_01630_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25051_ (.RESET_B(net6838),
    .D(_01631_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25052_ (.RESET_B(net6860),
    .D(_01632_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _25053_ (.RESET_B(net6887),
    .D(_01633_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][29] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25054_ (.RESET_B(net6962),
    .D(_01634_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][30] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _25055_ (.RESET_B(net6955),
    .D(_01635_),
    .Q(\soc_inst.cpu_core.register_file.registers[28][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _25056_ (.RESET_B(net6833),
    .D(_01636_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _25057_ (.RESET_B(net6842),
    .D(_01637_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][1] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _25058_ (.RESET_B(net6839),
    .D(_01638_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25059_ (.RESET_B(net6850),
    .D(_01639_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25060_ (.RESET_B(net6878),
    .D(_01640_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _25061_ (.RESET_B(net6910),
    .D(_01641_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][5] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25062_ (.RESET_B(net6907),
    .D(_01642_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25063_ (.RESET_B(net6926),
    .D(_01643_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][7] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25064_ (.RESET_B(net6898),
    .D(_01644_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][8] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25065_ (.RESET_B(net6957),
    .D(_01645_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][9] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25066_ (.RESET_B(net6972),
    .D(_01646_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25067_ (.RESET_B(net6893),
    .D(_01647_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _25068_ (.RESET_B(net6949),
    .D(_01648_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _25069_ (.RESET_B(net6936),
    .D(_01649_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _25070_ (.RESET_B(net6808),
    .D(_01650_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][14] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25071_ (.RESET_B(net6947),
    .D(_01651_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][15] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _25072_ (.RESET_B(net6917),
    .D(_01652_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _25073_ (.RESET_B(net6865),
    .D(_01653_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25074_ (.RESET_B(net6937),
    .D(_01654_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25075_ (.RESET_B(net6917),
    .D(_01655_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25076_ (.RESET_B(net6967),
    .D(_01656_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _25077_ (.RESET_B(net6910),
    .D(_01657_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][21] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25078_ (.RESET_B(net6823),
    .D(_01658_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][22] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_2 _25079_ (.RESET_B(net6982),
    .D(_01659_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25080_ (.RESET_B(net6861),
    .D(_01660_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _25081_ (.RESET_B(net6818),
    .D(_01661_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][25] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _25082_ (.RESET_B(net6918),
    .D(_01662_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][26] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25083_ (.RESET_B(net6824),
    .D(_01663_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25084_ (.RESET_B(net6867),
    .D(_01664_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][28] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25085_ (.RESET_B(net6882),
    .D(_01665_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][29] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25086_ (.RESET_B(net6961),
    .D(_01666_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][30] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25087_ (.RESET_B(net6956),
    .D(_01667_),
    .Q(\soc_inst.cpu_core.register_file.registers[16][31] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25088_ (.RESET_B(net6890),
    .D(_01668_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25089_ (.RESET_B(net6890),
    .D(_01669_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25090_ (.RESET_B(net6836),
    .D(_01670_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25091_ (.RESET_B(net6850),
    .D(_01671_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _25092_ (.RESET_B(net6904),
    .D(_01672_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _25093_ (.RESET_B(net6902),
    .D(_01673_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25094_ (.RESET_B(net6905),
    .D(_01674_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25095_ (.RESET_B(net6928),
    .D(_01675_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25096_ (.RESET_B(net6899),
    .D(_01676_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _25097_ (.RESET_B(net6957),
    .D(_01677_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _25098_ (.RESET_B(net6970),
    .D(_01678_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25099_ (.RESET_B(net6893),
    .D(_01679_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _25100_ (.RESET_B(net6948),
    .D(_01680_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _25101_ (.RESET_B(net6935),
    .D(_01681_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _25102_ (.RESET_B(net6817),
    .D(_01682_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _25103_ (.RESET_B(net6946),
    .D(_01683_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25104_ (.RESET_B(net6916),
    .D(_01684_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25105_ (.RESET_B(net6865),
    .D(_01685_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25106_ (.RESET_B(net6937),
    .D(_01686_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _25107_ (.RESET_B(net6869),
    .D(_01687_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _25108_ (.RESET_B(net6971),
    .D(_01688_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25109_ (.RESET_B(net6911),
    .D(_01689_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _25110_ (.RESET_B(net6826),
    .D(_01690_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _25111_ (.RESET_B(net6980),
    .D(_01691_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25112_ (.RESET_B(net6861),
    .D(_01692_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _25113_ (.RESET_B(net6821),
    .D(_01693_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_2 _25114_ (.RESET_B(net6918),
    .D(_01694_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25115_ (.RESET_B(net6829),
    .D(_01695_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25116_ (.RESET_B(net6866),
    .D(_01696_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25117_ (.RESET_B(net6887),
    .D(_01697_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25118_ (.RESET_B(net6961),
    .D(_01698_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25119_ (.RESET_B(net6953),
    .D(_01699_),
    .Q(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25120_ (.RESET_B(net6846),
    .D(_01700_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][0] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25121_ (.RESET_B(net6844),
    .D(_01701_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25122_ (.RESET_B(net6884),
    .D(_01702_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25123_ (.RESET_B(net6821),
    .D(_01703_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _25124_ (.RESET_B(net6876),
    .D(_01704_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][4] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _25125_ (.RESET_B(net6902),
    .D(_01705_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][5] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25126_ (.RESET_B(net6907),
    .D(_01706_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][6] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _25127_ (.RESET_B(net6927),
    .D(_01707_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][7] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25128_ (.RESET_B(net6899),
    .D(_01708_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][8] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _25129_ (.RESET_B(net6959),
    .D(_01709_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][9] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25130_ (.RESET_B(net6965),
    .D(_01710_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25131_ (.RESET_B(net6893),
    .D(_01711_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][11] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25132_ (.RESET_B(net6944),
    .D(_01712_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][12] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _25133_ (.RESET_B(net6931),
    .D(_01713_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25134_ (.RESET_B(net6816),
    .D(_01714_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][14] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _25135_ (.RESET_B(net6941),
    .D(_01715_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][15] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _25136_ (.RESET_B(net6920),
    .D(_01716_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _25137_ (.RESET_B(net6854),
    .D(_01717_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25138_ (.RESET_B(net6934),
    .D(_01718_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][18] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25139_ (.RESET_B(net6870),
    .D(_01719_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _25140_ (.RESET_B(net6967),
    .D(_01720_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][20] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _25141_ (.RESET_B(net6913),
    .D(_01721_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][21] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25142_ (.RESET_B(net6826),
    .D(_01722_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][22] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _25143_ (.RESET_B(net6982),
    .D(_01723_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25144_ (.RESET_B(net6858),
    .D(_01724_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][24] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _25145_ (.RESET_B(net6817),
    .D(_01725_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][25] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25146_ (.RESET_B(net6925),
    .D(_01726_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][26] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25147_ (.RESET_B(net6829),
    .D(_01727_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][27] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25148_ (.RESET_B(net6856),
    .D(_01728_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _25149_ (.RESET_B(net6883),
    .D(_01729_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _25150_ (.RESET_B(net6975),
    .D(_01730_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][30] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25151_ (.RESET_B(net6954),
    .D(_01731_),
    .Q(\soc_inst.cpu_core.register_file.registers[24][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25152_ (.RESET_B(net6890),
    .D(_01732_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25153_ (.RESET_B(net6845),
    .D(_01733_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25154_ (.RESET_B(net6884),
    .D(_01734_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25155_ (.RESET_B(net6849),
    .D(_01735_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25156_ (.RESET_B(net6901),
    .D(_01736_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25157_ (.RESET_B(net6903),
    .D(_01737_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25158_ (.RESET_B(net6906),
    .D(_01738_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25159_ (.RESET_B(net6928),
    .D(_01739_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25160_ (.RESET_B(net6900),
    .D(_01740_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _25161_ (.RESET_B(net6961),
    .D(_01741_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _25162_ (.RESET_B(net6969),
    .D(_01742_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25163_ (.RESET_B(net6893),
    .D(_01743_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][11] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _25164_ (.RESET_B(net6948),
    .D(_01744_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _25165_ (.RESET_B(net6935),
    .D(_01745_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25166_ (.RESET_B(net6817),
    .D(_01746_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][14] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25167_ (.RESET_B(net6946),
    .D(_01747_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25168_ (.RESET_B(net6920),
    .D(_01748_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _25169_ (.RESET_B(net6854),
    .D(_01749_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25170_ (.RESET_B(net6937),
    .D(_01750_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25171_ (.RESET_B(net6869),
    .D(_01751_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _25172_ (.RESET_B(net6972),
    .D(_01752_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25173_ (.RESET_B(net6960),
    .D(_01753_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25174_ (.RESET_B(net6852),
    .D(_01754_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _25175_ (.RESET_B(net6980),
    .D(_01755_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25176_ (.RESET_B(net6858),
    .D(_01756_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25177_ (.RESET_B(net6818),
    .D(_01757_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][25] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _25178_ (.RESET_B(net6872),
    .D(_01758_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][26] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25179_ (.RESET_B(net6827),
    .D(_01759_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _25180_ (.RESET_B(net6874),
    .D(_01760_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25181_ (.RESET_B(net6887),
    .D(_01761_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _25182_ (.RESET_B(net6963),
    .D(_01762_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25183_ (.RESET_B(net6956),
    .D(_01763_),
    .Q(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _25184_ (.RESET_B(net6846),
    .D(_01764_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][0] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25185_ (.RESET_B(net6841),
    .D(_01765_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25186_ (.RESET_B(net6838),
    .D(_01766_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][2] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _25187_ (.RESET_B(net6852),
    .D(_01767_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25188_ (.RESET_B(net6880),
    .D(_01768_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _25189_ (.RESET_B(net6902),
    .D(_01769_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][5] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _25190_ (.RESET_B(net6906),
    .D(_01770_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][6] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25191_ (.RESET_B(net6928),
    .D(_01771_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][7] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25192_ (.RESET_B(net6889),
    .D(_01772_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][8] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _25193_ (.RESET_B(net6961),
    .D(_01773_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][9] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _25194_ (.RESET_B(net6969),
    .D(_01774_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25195_ (.RESET_B(net6896),
    .D(_01775_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _25196_ (.RESET_B(net6948),
    .D(_01776_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][12] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25197_ (.RESET_B(net6938),
    .D(_01777_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25198_ (.RESET_B(net6811),
    .D(_01778_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][14] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25199_ (.RESET_B(net6942),
    .D(_01779_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _25200_ (.RESET_B(net6922),
    .D(_01780_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25201_ (.RESET_B(net6866),
    .D(_01781_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][17] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25202_ (.RESET_B(net6923),
    .D(_01782_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][18] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _25203_ (.RESET_B(net6872),
    .D(_01783_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _25204_ (.RESET_B(net6972),
    .D(_01784_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25205_ (.RESET_B(net6911),
    .D(_01785_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][21] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _25206_ (.RESET_B(net6823),
    .D(_01786_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][22] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25207_ (.RESET_B(net6978),
    .D(_01787_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25208_ (.RESET_B(net6859),
    .D(_01788_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25209_ (.RESET_B(net6810),
    .D(_01789_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25210_ (.RESET_B(net6919),
    .D(_01790_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][26] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25211_ (.RESET_B(net6828),
    .D(_01791_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25212_ (.RESET_B(net6856),
    .D(_01792_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][28] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25213_ (.RESET_B(net6887),
    .D(_01793_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][29] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25214_ (.RESET_B(net6974),
    .D(_01794_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][30] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25215_ (.RESET_B(net6955),
    .D(_01795_),
    .Q(\soc_inst.cpu_core.register_file.registers[29][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25216_ (.RESET_B(net6841),
    .D(_01796_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _25217_ (.RESET_B(net6840),
    .D(_01797_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25218_ (.RESET_B(net6836),
    .D(_01798_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25219_ (.RESET_B(net6850),
    .D(_01799_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _25220_ (.RESET_B(net6876),
    .D(_01800_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25221_ (.RESET_B(net6952),
    .D(_01801_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _25222_ (.RESET_B(net6906),
    .D(_01802_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25223_ (.RESET_B(net6926),
    .D(_01803_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25224_ (.RESET_B(net6889),
    .D(_01804_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25225_ (.RESET_B(net6963),
    .D(_01805_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _25226_ (.RESET_B(net6966),
    .D(_01806_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25227_ (.RESET_B(net6892),
    .D(_01807_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25228_ (.RESET_B(net6943),
    .D(_01808_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25229_ (.RESET_B(net6932),
    .D(_01809_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25230_ (.RESET_B(net6816),
    .D(_01810_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25231_ (.RESET_B(net6945),
    .D(_01811_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _25232_ (.RESET_B(net6922),
    .D(_01812_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25233_ (.RESET_B(net6866),
    .D(_01813_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25234_ (.RESET_B(net6922),
    .D(_01814_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][18] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25235_ (.RESET_B(net6872),
    .D(_01815_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25236_ (.RESET_B(net6967),
    .D(_01816_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25237_ (.RESET_B(net6909),
    .D(_01817_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25238_ (.RESET_B(net6823),
    .D(_01818_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _25239_ (.RESET_B(net6978),
    .D(_01819_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25240_ (.RESET_B(net6860),
    .D(_01820_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25241_ (.RESET_B(net6818),
    .D(_01821_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25242_ (.RESET_B(net6925),
    .D(_01822_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25243_ (.RESET_B(net6827),
    .D(_01823_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25244_ (.RESET_B(net6874),
    .D(_01824_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25245_ (.RESET_B(net6883),
    .D(_01825_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25246_ (.RESET_B(net6975),
    .D(_01826_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25247_ (.RESET_B(net6952),
    .D(_01827_),
    .Q(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _25248_ (.RESET_B(net6843),
    .D(_01828_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _25249_ (.RESET_B(net6842),
    .D(_01829_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _25250_ (.RESET_B(net6835),
    .D(_01830_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25251_ (.RESET_B(net6851),
    .D(_01831_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25252_ (.RESET_B(net6878),
    .D(_01832_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _25253_ (.RESET_B(net6902),
    .D(_01833_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][5] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _25254_ (.RESET_B(net6908),
    .D(_01834_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25255_ (.RESET_B(net6927),
    .D(_01835_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _25256_ (.RESET_B(net6900),
    .D(_01836_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25257_ (.RESET_B(net6958),
    .D(_01837_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25258_ (.RESET_B(net6965),
    .D(_01838_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25259_ (.RESET_B(net6891),
    .D(_01839_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25260_ (.RESET_B(net6943),
    .D(_01840_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _25261_ (.RESET_B(net6931),
    .D(_01841_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _25262_ (.RESET_B(net6809),
    .D(_01842_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][14] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _25263_ (.RESET_B(net6941),
    .D(_01843_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _25264_ (.RESET_B(net6916),
    .D(_01844_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25265_ (.RESET_B(net6865),
    .D(_01845_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _25266_ (.RESET_B(net6933),
    .D(_01846_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25267_ (.RESET_B(net6870),
    .D(_01847_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _25268_ (.RESET_B(net6967),
    .D(_01848_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _25269_ (.RESET_B(net6911),
    .D(_01849_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][21] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25270_ (.RESET_B(net6825),
    .D(_01850_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _25271_ (.RESET_B(net6976),
    .D(_01851_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25272_ (.RESET_B(net6861),
    .D(_01852_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _25273_ (.RESET_B(net6811),
    .D(_01853_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25274_ (.RESET_B(net6924),
    .D(_01854_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25275_ (.RESET_B(net6826),
    .D(_01855_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25276_ (.RESET_B(net6857),
    .D(_01856_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25277_ (.RESET_B(net6888),
    .D(_01857_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _25278_ (.RESET_B(net6975),
    .D(_01858_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25279_ (.RESET_B(net6955),
    .D(_01859_),
    .Q(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25280_ (.RESET_B(net6846),
    .D(_01860_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][0] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25281_ (.RESET_B(net6890),
    .D(_01861_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25282_ (.RESET_B(net6884),
    .D(_01862_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][2] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25283_ (.RESET_B(net6850),
    .D(_01863_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][3] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25284_ (.RESET_B(net6876),
    .D(_01864_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][4] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25285_ (.RESET_B(net6902),
    .D(_01865_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][5] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25286_ (.RESET_B(net6905),
    .D(_01866_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][6] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25287_ (.RESET_B(net6928),
    .D(_01867_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _25288_ (.RESET_B(net6898),
    .D(_01868_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][8] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25289_ (.RESET_B(net6957),
    .D(_01869_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25290_ (.RESET_B(net6970),
    .D(_01870_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25291_ (.RESET_B(net6894),
    .D(_01871_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][11] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _25292_ (.RESET_B(net6949),
    .D(_01872_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _25293_ (.RESET_B(net6935),
    .D(_01873_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25294_ (.RESET_B(net6816),
    .D(_01874_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][14] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25295_ (.RESET_B(net6946),
    .D(_01875_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _25296_ (.RESET_B(net6916),
    .D(_01876_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][16] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25297_ (.RESET_B(net6855),
    .D(_01877_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][17] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25298_ (.RESET_B(net6933),
    .D(_01878_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25299_ (.RESET_B(net6917),
    .D(_01879_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _25300_ (.RESET_B(net6978),
    .D(_01880_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][20] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25301_ (.RESET_B(net6911),
    .D(_01881_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][21] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25302_ (.RESET_B(net6826),
    .D(_01882_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25303_ (.RESET_B(net6979),
    .D(_01883_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25304_ (.RESET_B(net6861),
    .D(_01884_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][24] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25305_ (.RESET_B(net6819),
    .D(_01885_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][25] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25306_ (.RESET_B(net6872),
    .D(_01886_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][26] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25307_ (.RESET_B(net6828),
    .D(_01887_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][27] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25308_ (.RESET_B(net6875),
    .D(_01888_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][28] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25309_ (.RESET_B(net6882),
    .D(_01889_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][29] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25310_ (.RESET_B(net6974),
    .D(_01890_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25311_ (.RESET_B(net6954),
    .D(_01891_),
    .Q(\soc_inst.cpu_core.register_file.registers[25][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _25312_ (.RESET_B(net6842),
    .D(_01892_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _25313_ (.RESET_B(net6842),
    .D(_01893_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25314_ (.RESET_B(net6836),
    .D(_01894_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25315_ (.RESET_B(net6853),
    .D(_01895_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25316_ (.RESET_B(net6880),
    .D(_01896_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25317_ (.RESET_B(net6952),
    .D(_01897_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _25318_ (.RESET_B(net6914),
    .D(_01898_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25319_ (.RESET_B(net6927),
    .D(_01899_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25320_ (.RESET_B(net6898),
    .D(_01900_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _25321_ (.RESET_B(net6961),
    .D(_01901_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25322_ (.RESET_B(net6965),
    .D(_01902_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25323_ (.RESET_B(net6893),
    .D(_01903_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _25324_ (.RESET_B(net6943),
    .D(_01904_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _25325_ (.RESET_B(net6932),
    .D(_01905_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25326_ (.RESET_B(net6809),
    .D(_01906_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25327_ (.RESET_B(net6942),
    .D(_01907_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _25328_ (.RESET_B(net6917),
    .D(_01908_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25329_ (.RESET_B(net6868),
    .D(_01909_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _25330_ (.RESET_B(net6933),
    .D(_01910_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][18] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _25331_ (.RESET_B(net6917),
    .D(_01911_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _25332_ (.RESET_B(net6967),
    .D(_01912_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _25333_ (.RESET_B(net6909),
    .D(_01913_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][21] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25334_ (.RESET_B(net6823),
    .D(_01914_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25335_ (.RESET_B(net6977),
    .D(_01915_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25336_ (.RESET_B(net6861),
    .D(_01916_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25337_ (.RESET_B(net6818),
    .D(_01917_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25338_ (.RESET_B(net6924),
    .D(_01918_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25339_ (.RESET_B(net6824),
    .D(_01919_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25340_ (.RESET_B(net6866),
    .D(_01920_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25341_ (.RESET_B(net6888),
    .D(_01921_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25342_ (.RESET_B(net6975),
    .D(_01922_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25343_ (.RESET_B(net6956),
    .D(_01923_),
    .Q(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25344_ (.RESET_B(net6841),
    .D(_01924_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][0] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25345_ (.RESET_B(net6844),
    .D(_01925_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][1] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25346_ (.RESET_B(net6836),
    .D(_01926_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25347_ (.RESET_B(net6850),
    .D(_01927_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _25348_ (.RESET_B(net6878),
    .D(_01928_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][4] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25349_ (.RESET_B(net6904),
    .D(_01929_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][5] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25350_ (.RESET_B(net6905),
    .D(_01930_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][6] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25351_ (.RESET_B(net6926),
    .D(_01931_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][7] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25352_ (.RESET_B(net6898),
    .D(_01932_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][8] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _25353_ (.RESET_B(net6959),
    .D(_01933_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][9] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _25354_ (.RESET_B(net6969),
    .D(_01934_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25355_ (.RESET_B(net6893),
    .D(_01935_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][11] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _25356_ (.RESET_B(net6948),
    .D(_01936_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _25357_ (.RESET_B(net6939),
    .D(_01937_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][13] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25358_ (.RESET_B(net6817),
    .D(_01938_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][14] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _25359_ (.RESET_B(net6946),
    .D(_01939_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][15] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _25360_ (.RESET_B(net6922),
    .D(_01940_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25361_ (.RESET_B(net6866),
    .D(_01941_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][17] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25362_ (.RESET_B(net6938),
    .D(_01942_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25363_ (.RESET_B(net6872),
    .D(_01943_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][19] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25364_ (.RESET_B(net6971),
    .D(_01944_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _25365_ (.RESET_B(net6909),
    .D(_01945_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][21] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25366_ (.RESET_B(net6827),
    .D(_01946_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][22] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _25367_ (.RESET_B(net6978),
    .D(_01947_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _25368_ (.RESET_B(net6860),
    .D(_01948_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][24] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25369_ (.RESET_B(net6810),
    .D(_01949_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25370_ (.RESET_B(net6924),
    .D(_01950_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25371_ (.RESET_B(net6828),
    .D(_01951_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25372_ (.RESET_B(net6856),
    .D(_01952_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][28] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25373_ (.RESET_B(net6883),
    .D(_01953_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _25374_ (.RESET_B(net6976),
    .D(_01954_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25375_ (.RESET_B(net6954),
    .D(_01955_),
    .Q(\soc_inst.cpu_core.register_file.registers[30][31] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25376_ (.RESET_B(net6846),
    .D(_01956_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25377_ (.RESET_B(net6842),
    .D(_01957_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _25378_ (.RESET_B(net6836),
    .D(_01958_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _25379_ (.RESET_B(net6849),
    .D(_01959_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25380_ (.RESET_B(net6878),
    .D(_01960_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _25381_ (.RESET_B(net6902),
    .D(_01961_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25382_ (.RESET_B(net6908),
    .D(_01962_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25383_ (.RESET_B(net6926),
    .D(_01963_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25384_ (.RESET_B(net6898),
    .D(_01964_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _25385_ (.RESET_B(net6960),
    .D(_01965_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25386_ (.RESET_B(net6970),
    .D(_01966_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25387_ (.RESET_B(net6893),
    .D(_01967_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _25388_ (.RESET_B(net6950),
    .D(_01968_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _25389_ (.RESET_B(net6936),
    .D(_01969_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _25390_ (.RESET_B(net6809),
    .D(_01970_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25391_ (.RESET_B(net6946),
    .D(_01971_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25392_ (.RESET_B(net6920),
    .D(_01972_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25393_ (.RESET_B(net6855),
    .D(_01973_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25394_ (.RESET_B(net6938),
    .D(_01974_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _25395_ (.RESET_B(net6870),
    .D(_01975_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _25396_ (.RESET_B(net6971),
    .D(_01976_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _25397_ (.RESET_B(net6960),
    .D(_01977_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25398_ (.RESET_B(net6822),
    .D(_01978_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _25399_ (.RESET_B(net6979),
    .D(_01979_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25400_ (.RESET_B(net6858),
    .D(_01980_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25401_ (.RESET_B(net6811),
    .D(_01981_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_2 _25402_ (.RESET_B(net6918),
    .D(_01982_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25403_ (.RESET_B(net6825),
    .D(_01983_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25404_ (.RESET_B(net6874),
    .D(_01984_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25405_ (.RESET_B(net6887),
    .D(_01985_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25406_ (.RESET_B(net6962),
    .D(_01986_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _25407_ (.RESET_B(net6956),
    .D(_01987_),
    .Q(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _25408_ (.RESET_B(net6845),
    .D(_01988_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25409_ (.RESET_B(net6844),
    .D(_01989_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25410_ (.RESET_B(net6884),
    .D(_01990_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25411_ (.RESET_B(net6849),
    .D(_01991_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _25412_ (.RESET_B(net6879),
    .D(_01992_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25413_ (.RESET_B(net6901),
    .D(_01993_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _25414_ (.RESET_B(net6908),
    .D(_01994_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25415_ (.RESET_B(net6929),
    .D(_01995_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25416_ (.RESET_B(net6899),
    .D(_01996_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25417_ (.RESET_B(net6958),
    .D(_01997_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25418_ (.RESET_B(net6965),
    .D(_01998_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25419_ (.RESET_B(net6892),
    .D(_01999_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _25420_ (.RESET_B(net6949),
    .D(_02000_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25421_ (.RESET_B(net6936),
    .D(_02001_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25422_ (.RESET_B(net6816),
    .D(_02002_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _25423_ (.RESET_B(net6947),
    .D(_02003_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25424_ (.RESET_B(net6921),
    .D(_02004_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25425_ (.RESET_B(net6855),
    .D(_02005_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25426_ (.RESET_B(net6937),
    .D(_02006_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25427_ (.RESET_B(net6869),
    .D(_02007_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25428_ (.RESET_B(net6968),
    .D(_02008_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _25429_ (.RESET_B(net6912),
    .D(_02009_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25430_ (.RESET_B(net6858),
    .D(_02010_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][22] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _25431_ (.RESET_B(net6981),
    .D(_02011_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _25432_ (.RESET_B(net6858),
    .D(_02012_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][24] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25433_ (.RESET_B(net6822),
    .D(_02013_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_2 _25434_ (.RESET_B(net6880),
    .D(_02014_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25435_ (.RESET_B(net6828),
    .D(_02015_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25436_ (.RESET_B(net6874),
    .D(_02016_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][28] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25437_ (.RESET_B(net6885),
    .D(_02017_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _25438_ (.RESET_B(net6976),
    .D(_02018_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _25439_ (.RESET_B(net6955),
    .D(_02019_),
    .Q(\soc_inst.cpu_core.register_file.registers[9][31] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _25440_ (.RESET_B(net6833),
    .D(_02020_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _25441_ (.RESET_B(net6843),
    .D(_02021_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25442_ (.RESET_B(net6835),
    .D(_02022_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25443_ (.RESET_B(net6851),
    .D(_02023_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25444_ (.RESET_B(net6879),
    .D(_02024_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _25445_ (.RESET_B(net6902),
    .D(_02025_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25446_ (.RESET_B(net6908),
    .D(_02026_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _25447_ (.RESET_B(net6929),
    .D(_02027_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25448_ (.RESET_B(net6899),
    .D(_02028_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25449_ (.RESET_B(net6957),
    .D(_02029_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _25450_ (.RESET_B(net6970),
    .D(_02030_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25451_ (.RESET_B(net6891),
    .D(_02031_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _25452_ (.RESET_B(net6950),
    .D(_02032_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _25453_ (.RESET_B(net6935),
    .D(_02033_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _25454_ (.RESET_B(net6808),
    .D(_02034_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _25455_ (.RESET_B(net6946),
    .D(_02035_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25456_ (.RESET_B(net6917),
    .D(_02036_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25457_ (.RESET_B(net6855),
    .D(_02037_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25458_ (.RESET_B(net6934),
    .D(_02038_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25459_ (.RESET_B(net6872),
    .D(_02039_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25460_ (.RESET_B(net6972),
    .D(_02040_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _25461_ (.RESET_B(net6912),
    .D(_02041_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25462_ (.RESET_B(net6823),
    .D(_02042_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_2 _25463_ (.RESET_B(net6981),
    .D(_02043_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25464_ (.RESET_B(net6860),
    .D(_02044_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25465_ (.RESET_B(net6809),
    .D(_02045_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _25466_ (.RESET_B(net6924),
    .D(_02046_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25467_ (.RESET_B(net6824),
    .D(_02047_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _25468_ (.RESET_B(net6867),
    .D(_02048_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25469_ (.RESET_B(net6887),
    .D(_02049_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25470_ (.RESET_B(net6962),
    .D(_02050_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25471_ (.RESET_B(net6953),
    .D(_02051_),
    .Q(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _25472_ (.RESET_B(net6833),
    .D(_02052_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _25473_ (.RESET_B(net6842),
    .D(_02053_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25474_ (.RESET_B(net6837),
    .D(_02054_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _25475_ (.RESET_B(net6851),
    .D(_02055_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25476_ (.RESET_B(net6878),
    .D(_02056_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25477_ (.RESET_B(net6903),
    .D(_02057_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _25478_ (.RESET_B(net6908),
    .D(_02058_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25479_ (.RESET_B(net6929),
    .D(_02059_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _25480_ (.RESET_B(net6900),
    .D(_02060_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _25481_ (.RESET_B(net6959),
    .D(_02061_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25482_ (.RESET_B(net6970),
    .D(_02062_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25483_ (.RESET_B(net6895),
    .D(_02063_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _25484_ (.RESET_B(net6948),
    .D(_02064_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25485_ (.RESET_B(net6938),
    .D(_02065_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25486_ (.RESET_B(net6809),
    .D(_02066_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _25487_ (.RESET_B(net6941),
    .D(_02067_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25488_ (.RESET_B(net6920),
    .D(_02068_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25489_ (.RESET_B(net6857),
    .D(_02069_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25490_ (.RESET_B(net6933),
    .D(_02070_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25491_ (.RESET_B(net6873),
    .D(_02071_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _25492_ (.RESET_B(net6973),
    .D(_02072_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _25493_ (.RESET_B(net6912),
    .D(_02073_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25494_ (.RESET_B(net6826),
    .D(_02074_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _25495_ (.RESET_B(net6981),
    .D(_02075_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25496_ (.RESET_B(net6860),
    .D(_02076_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _25497_ (.RESET_B(net6810),
    .D(_02077_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25498_ (.RESET_B(net6925),
    .D(_02078_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25499_ (.RESET_B(net6824),
    .D(_02079_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25500_ (.RESET_B(net6866),
    .D(_02080_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _25501_ (.RESET_B(net6887),
    .D(_02081_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _25502_ (.RESET_B(net6975),
    .D(_02082_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _25503_ (.RESET_B(net6955),
    .D(_02083_),
    .Q(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25504_ (.RESET_B(net6845),
    .D(_02084_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25505_ (.RESET_B(net6844),
    .D(_02085_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25506_ (.RESET_B(net6884),
    .D(_02086_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25507_ (.RESET_B(net6851),
    .D(_02087_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25508_ (.RESET_B(net6876),
    .D(_02088_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25509_ (.RESET_B(net6903),
    .D(_02089_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _25510_ (.RESET_B(net6905),
    .D(_02090_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25511_ (.RESET_B(net6927),
    .D(_02091_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25512_ (.RESET_B(net6889),
    .D(_02092_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25513_ (.RESET_B(net6961),
    .D(_02093_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25514_ (.RESET_B(net6965),
    .D(_02094_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25515_ (.RESET_B(net6896),
    .D(_02095_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _25516_ (.RESET_B(net6948),
    .D(_02096_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25517_ (.RESET_B(net6935),
    .D(_02097_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25518_ (.RESET_B(net6820),
    .D(_02098_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25519_ (.RESET_B(net6942),
    .D(_02099_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25520_ (.RESET_B(net6922),
    .D(_02100_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _25521_ (.RESET_B(net6856),
    .D(_02101_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25522_ (.RESET_B(net6933),
    .D(_02102_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25523_ (.RESET_B(net6872),
    .D(_02103_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _25524_ (.RESET_B(net6971),
    .D(_02104_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25525_ (.RESET_B(net6911),
    .D(_02105_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25526_ (.RESET_B(net6826),
    .D(_02106_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _25527_ (.RESET_B(net6980),
    .D(_02107_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _25528_ (.RESET_B(net6862),
    .D(_02108_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25529_ (.RESET_B(net6819),
    .D(_02109_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25530_ (.RESET_B(net6924),
    .D(_02110_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25531_ (.RESET_B(net6838),
    .D(_02111_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25532_ (.RESET_B(net6863),
    .D(_02112_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _25533_ (.RESET_B(net6887),
    .D(_02113_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][29] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _25534_ (.RESET_B(net6974),
    .D(_02114_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _25535_ (.RESET_B(net6955),
    .D(_02115_),
    .Q(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _25536_ (.RESET_B(net6890),
    .D(_02116_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][0] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25537_ (.RESET_B(net6845),
    .D(_02117_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][1] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25538_ (.RESET_B(net6885),
    .D(_02118_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][2] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25539_ (.RESET_B(net6849),
    .D(_02119_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25540_ (.RESET_B(net6877),
    .D(_02120_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][4] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25541_ (.RESET_B(net6901),
    .D(_02121_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][5] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25542_ (.RESET_B(net6907),
    .D(_02122_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][6] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25543_ (.RESET_B(net6930),
    .D(_02123_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25544_ (.RESET_B(net6889),
    .D(_02124_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][8] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25545_ (.RESET_B(net6958),
    .D(_02125_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][9] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25546_ (.RESET_B(net6969),
    .D(_02126_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25547_ (.RESET_B(net6895),
    .D(_02127_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][11] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _25548_ (.RESET_B(net6948),
    .D(_02128_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _25549_ (.RESET_B(net6935),
    .D(_02129_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _25550_ (.RESET_B(net6817),
    .D(_02130_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][14] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _25551_ (.RESET_B(net6941),
    .D(_02131_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][15] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25552_ (.RESET_B(net6920),
    .D(_02132_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _25553_ (.RESET_B(net6865),
    .D(_02133_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][17] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25554_ (.RESET_B(net6934),
    .D(_02134_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][18] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25555_ (.RESET_B(net6870),
    .D(_02135_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _25556_ (.RESET_B(net6971),
    .D(_02136_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25557_ (.RESET_B(net6911),
    .D(_02137_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][21] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25558_ (.RESET_B(net6822),
    .D(_02138_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][22] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_2 _25559_ (.RESET_B(net6980),
    .D(_02139_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][23] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _25560_ (.RESET_B(net6859),
    .D(_02140_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][24] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25561_ (.RESET_B(net6818),
    .D(_02141_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][25] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _25562_ (.RESET_B(net6924),
    .D(_02142_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25563_ (.RESET_B(net6829),
    .D(_02143_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25564_ (.RESET_B(net6874),
    .D(_02144_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][28] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25565_ (.RESET_B(net6886),
    .D(_02145_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][29] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _25566_ (.RESET_B(net6975),
    .D(_02146_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][30] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25567_ (.RESET_B(net6954),
    .D(_02147_),
    .Q(\soc_inst.cpu_core.register_file.registers[23][31] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25568_ (.RESET_B(net6890),
    .D(_02148_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][0] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25569_ (.RESET_B(net6844),
    .D(_02149_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][1] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25570_ (.RESET_B(net6884),
    .D(_02150_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][2] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25571_ (.RESET_B(net6849),
    .D(_02151_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][3] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _25572_ (.RESET_B(net6879),
    .D(_02152_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25573_ (.RESET_B(net6909),
    .D(_02153_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25574_ (.RESET_B(net6906),
    .D(_02154_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25575_ (.RESET_B(net6929),
    .D(_02155_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25576_ (.RESET_B(net6889),
    .D(_02156_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][8] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25577_ (.RESET_B(net6959),
    .D(_02157_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25578_ (.RESET_B(net6970),
    .D(_02158_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25579_ (.RESET_B(net6894),
    .D(_02159_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _25580_ (.RESET_B(net6949),
    .D(_02160_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][12] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _25581_ (.RESET_B(net6936),
    .D(_02161_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25582_ (.RESET_B(net6816),
    .D(_02162_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _25583_ (.RESET_B(net6947),
    .D(_02163_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25584_ (.RESET_B(net6920),
    .D(_02164_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _25585_ (.RESET_B(net6854),
    .D(_02165_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25586_ (.RESET_B(net6937),
    .D(_02166_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _25587_ (.RESET_B(net6869),
    .D(_02167_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _25588_ (.RESET_B(net6971),
    .D(_02168_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _25589_ (.RESET_B(net6912),
    .D(_02169_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25590_ (.RESET_B(net6851),
    .D(_02170_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][22] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25591_ (.RESET_B(net6980),
    .D(_02171_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25592_ (.RESET_B(net6858),
    .D(_02172_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25593_ (.RESET_B(net6816),
    .D(_02173_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25594_ (.RESET_B(net6880),
    .D(_02174_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][26] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25595_ (.RESET_B(net6829),
    .D(_02175_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25596_ (.RESET_B(net6874),
    .D(_02176_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25597_ (.RESET_B(net6885),
    .D(_02177_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][29] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _25598_ (.RESET_B(net6962),
    .D(_02178_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][30] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25599_ (.RESET_B(net6956),
    .D(_02179_),
    .Q(\soc_inst.cpu_core.register_file.registers[5][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25600_ (.RESET_B(net6840),
    .D(_02180_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][0] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _25601_ (.RESET_B(net6840),
    .D(_02181_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25602_ (.RESET_B(net6836),
    .D(_02182_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][2] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _25603_ (.RESET_B(net6851),
    .D(_02183_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][3] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25604_ (.RESET_B(net6876),
    .D(_02184_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][4] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25605_ (.RESET_B(net6903),
    .D(_02185_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _25606_ (.RESET_B(net6906),
    .D(_02186_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25607_ (.RESET_B(net6929),
    .D(_02187_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25608_ (.RESET_B(net6888),
    .D(_02188_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _25609_ (.RESET_B(net6959),
    .D(_02189_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][9] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25610_ (.RESET_B(net6966),
    .D(_02190_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][10] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25611_ (.RESET_B(net6893),
    .D(_02191_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25612_ (.RESET_B(net6944),
    .D(_02192_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25613_ (.RESET_B(net6931),
    .D(_02193_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][13] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25614_ (.RESET_B(net6809),
    .D(_02194_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25615_ (.RESET_B(net6947),
    .D(_02195_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _25616_ (.RESET_B(net6921),
    .D(_02196_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25617_ (.RESET_B(net6865),
    .D(_02197_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _25618_ (.RESET_B(net6934),
    .D(_02198_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][18] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25619_ (.RESET_B(net6870),
    .D(_02199_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25620_ (.RESET_B(net6967),
    .D(_02200_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _25621_ (.RESET_B(net6910),
    .D(_02201_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25622_ (.RESET_B(net6852),
    .D(_02202_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25623_ (.RESET_B(net6978),
    .D(_02203_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][23] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25624_ (.RESET_B(net6862),
    .D(_02204_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _25625_ (.RESET_B(net6811),
    .D(_02205_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][25] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25626_ (.RESET_B(net6925),
    .D(_02206_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25627_ (.RESET_B(net6825),
    .D(_02207_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25628_ (.RESET_B(net6867),
    .D(_02208_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25629_ (.RESET_B(net6882),
    .D(_02209_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _25630_ (.RESET_B(net6974),
    .D(_02210_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25631_ (.RESET_B(net6952),
    .D(_02211_),
    .Q(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _25632_ (.RESET_B(net6840),
    .D(_02212_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _25633_ (.RESET_B(net6840),
    .D(_02213_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25634_ (.RESET_B(net6836),
    .D(_02214_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _25635_ (.RESET_B(net6850),
    .D(_02215_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][3] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _25636_ (.RESET_B(net6901),
    .D(_02216_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25637_ (.RESET_B(net6901),
    .D(_02217_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _25638_ (.RESET_B(net6905),
    .D(_02218_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25639_ (.RESET_B(net6925),
    .D(_02219_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25640_ (.RESET_B(net6888),
    .D(_02220_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][8] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _25641_ (.RESET_B(net6963),
    .D(_02221_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _25642_ (.RESET_B(net6969),
    .D(_02222_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25643_ (.RESET_B(net6894),
    .D(_02223_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _25644_ (.RESET_B(net6949),
    .D(_02224_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _25645_ (.RESET_B(net6936),
    .D(_02225_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25646_ (.RESET_B(net6816),
    .D(_02226_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _25647_ (.RESET_B(net6947),
    .D(_02227_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _25648_ (.RESET_B(net6916),
    .D(_02228_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _25649_ (.RESET_B(net6865),
    .D(_02229_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _25650_ (.RESET_B(net6937),
    .D(_02230_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][18] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25651_ (.RESET_B(net6871),
    .D(_02231_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][19] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _25652_ (.RESET_B(net6972),
    .D(_02232_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][20] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25653_ (.RESET_B(net6910),
    .D(_02233_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25654_ (.RESET_B(net6813),
    .D(_02234_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25655_ (.RESET_B(net6978),
    .D(_02235_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][23] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25656_ (.RESET_B(net6860),
    .D(_02236_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][24] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25657_ (.RESET_B(net6810),
    .D(_02237_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25658_ (.RESET_B(net6927),
    .D(_02238_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25659_ (.RESET_B(net6825),
    .D(_02239_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][27] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _25660_ (.RESET_B(net6875),
    .D(_02240_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25661_ (.RESET_B(net6882),
    .D(_02241_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _25662_ (.RESET_B(net6974),
    .D(_02242_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25663_ (.RESET_B(net6952),
    .D(_02243_),
    .Q(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25664_ (.RESET_B(net6892),
    .D(_02244_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _25665_ (.RESET_B(net6844),
    .D(_02245_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25666_ (.RESET_B(net6835),
    .D(_02246_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][2] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _25667_ (.RESET_B(net6849),
    .D(_02247_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _25668_ (.RESET_B(net6876),
    .D(_02248_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][4] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _25669_ (.RESET_B(net6903),
    .D(_02249_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][5] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25670_ (.RESET_B(net6907),
    .D(_02250_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][6] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _25671_ (.RESET_B(net6928),
    .D(_02251_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][7] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25672_ (.RESET_B(net6889),
    .D(_02252_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][8] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25673_ (.RESET_B(net6960),
    .D(_02253_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][9] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25674_ (.RESET_B(net6966),
    .D(_02254_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25675_ (.RESET_B(net6894),
    .D(_02255_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][11] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _25676_ (.RESET_B(net6943),
    .D(_02256_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][12] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25677_ (.RESET_B(net6931),
    .D(_02257_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][13] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25678_ (.RESET_B(net6820),
    .D(_02258_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][14] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_2 _25679_ (.RESET_B(net6941),
    .D(_02259_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][15] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25680_ (.RESET_B(net6916),
    .D(_02260_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25681_ (.RESET_B(net6866),
    .D(_02261_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][17] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25682_ (.RESET_B(net6923),
    .D(_02262_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][18] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25683_ (.RESET_B(net6873),
    .D(_02263_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25684_ (.RESET_B(net6968),
    .D(_02264_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][20] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25685_ (.RESET_B(net6960),
    .D(_02265_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][21] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25686_ (.RESET_B(net6858),
    .D(_02266_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][22] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _25687_ (.RESET_B(net6982),
    .D(_02267_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][23] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25688_ (.RESET_B(net6862),
    .D(_02268_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][24] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _25689_ (.RESET_B(net6819),
    .D(_02269_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _25690_ (.RESET_B(net6918),
    .D(_02270_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][26] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25691_ (.RESET_B(net6829),
    .D(_02271_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25692_ (.RESET_B(net6874),
    .D(_02272_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][28] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _25693_ (.RESET_B(net6883),
    .D(_02273_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][29] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25694_ (.RESET_B(net6975),
    .D(_02274_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][30] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25695_ (.RESET_B(net6954),
    .D(_02275_),
    .Q(\soc_inst.cpu_core.register_file.registers[26][31] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25696_ (.RESET_B(net6892),
    .D(_02276_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][0] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _25697_ (.RESET_B(net6844),
    .D(_02277_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25698_ (.RESET_B(net6884),
    .D(_02278_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _25699_ (.RESET_B(net6849),
    .D(_02279_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25700_ (.RESET_B(net6878),
    .D(_02280_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25701_ (.RESET_B(net6904),
    .D(_02281_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25702_ (.RESET_B(net6905),
    .D(_02282_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25703_ (.RESET_B(net6927),
    .D(_02283_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25704_ (.RESET_B(net6899),
    .D(_02284_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25705_ (.RESET_B(net6961),
    .D(_02285_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25706_ (.RESET_B(net6966),
    .D(_02286_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25707_ (.RESET_B(net6894),
    .D(_02287_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _25708_ (.RESET_B(net6943),
    .D(_02288_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _25709_ (.RESET_B(net6931),
    .D(_02289_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _25710_ (.RESET_B(net6817),
    .D(_02290_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_2 _25711_ (.RESET_B(net6941),
    .D(_02291_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25712_ (.RESET_B(net6921),
    .D(_02292_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25713_ (.RESET_B(net6854),
    .D(_02293_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _25714_ (.RESET_B(net6934),
    .D(_02294_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25715_ (.RESET_B(net6869),
    .D(_02295_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][19] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25716_ (.RESET_B(net6972),
    .D(_02296_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25717_ (.RESET_B(net6909),
    .D(_02297_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][21] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25718_ (.RESET_B(net6852),
    .D(_02298_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25719_ (.RESET_B(net6978),
    .D(_02299_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][23] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25720_ (.RESET_B(net6862),
    .D(_02300_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _25721_ (.RESET_B(net6821),
    .D(_02301_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25722_ (.RESET_B(net6927),
    .D(_02302_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25723_ (.RESET_B(net6829),
    .D(_02303_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25724_ (.RESET_B(net6875),
    .D(_02304_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25725_ (.RESET_B(net6882),
    .D(_02305_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25726_ (.RESET_B(net6974),
    .D(_02306_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25727_ (.RESET_B(net6954),
    .D(_02307_),
    .Q(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _25728_ (.RESET_B(net6832),
    .D(_02308_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _25729_ (.RESET_B(net6803),
    .D(_02309_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][1] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25730_ (.RESET_B(net6839),
    .D(_02310_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][2] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25731_ (.RESET_B(net6859),
    .D(_02311_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25732_ (.RESET_B(net6882),
    .D(_02312_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][4] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25733_ (.RESET_B(net6837),
    .D(_02313_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][5] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _25734_ (.RESET_B(net6833),
    .D(_02314_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][6] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _25735_ (.RESET_B(net6839),
    .D(_02315_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][7] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25736_ (.RESET_B(net6835),
    .D(_02316_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][8] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _25737_ (.RESET_B(net6839),
    .D(_02317_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][9] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25738_ (.RESET_B(net6839),
    .D(_02318_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][10] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _25739_ (.RESET_B(net6843),
    .D(_02319_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][11] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _25740_ (.RESET_B(net6814),
    .D(_02320_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][12] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _25741_ (.RESET_B(net6774),
    .D(_02321_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][13] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _25742_ (.RESET_B(net6771),
    .D(_02322_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][14] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _25743_ (.RESET_B(net6815),
    .D(_02323_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][15] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25744_ (.RESET_B(net6772),
    .D(_02324_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][16] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_2 _25745_ (.RESET_B(net6822),
    .D(_02325_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][17] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _25746_ (.RESET_B(net6772),
    .D(_02326_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][18] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _25747_ (.RESET_B(net6867),
    .D(_02327_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][19] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _25748_ (.RESET_B(net6953),
    .D(_02328_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25749_ (.RESET_B(net6909),
    .D(_02329_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][21] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25750_ (.RESET_B(net6807),
    .D(_02330_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][22] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25751_ (.RESET_B(net6957),
    .D(_02331_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][23] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _25752_ (.RESET_B(net6827),
    .D(_02332_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][24] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25753_ (.RESET_B(net6806),
    .D(_02333_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][25] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _25754_ (.RESET_B(net6880),
    .D(_02334_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][26] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25755_ (.RESET_B(net6824),
    .D(_02335_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][27] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25756_ (.RESET_B(net6858),
    .D(_02336_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][28] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25757_ (.RESET_B(net6838),
    .D(_02337_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][29] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _25758_ (.RESET_B(net6960),
    .D(_02338_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][30] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25759_ (.RESET_B(net6839),
    .D(_02339_),
    .Q(\soc_inst.cpu_core.register_file.registers[1][31] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25760_ (.RESET_B(net6679),
    .D(_02340_),
    .Q(\soc_inst.cpu_core.csr_file.mie[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _25761_ (.RESET_B(net6680),
    .D(_02341_),
    .Q(\soc_inst.cpu_core.csr_file.mie[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _25762_ (.RESET_B(net6747),
    .D(net2435),
    .Q(\soc_inst.cpu_core.ex_branch_target[0] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25763_ (.RESET_B(net6746),
    .D(_02343_),
    .Q(\soc_inst.cpu_core.ex_branch_target[1] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _25764_ (.RESET_B(net6782),
    .D(net1785),
    .Q(\soc_inst.cpu_core.ex_branch_target[2] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25765_ (.RESET_B(net6798),
    .D(net2915),
    .Q(\soc_inst.cpu_core.ex_branch_target[3] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25766_ (.RESET_B(net6798),
    .D(_02346_),
    .Q(\soc_inst.cpu_core.ex_branch_target[4] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25767_ (.RESET_B(net6800),
    .D(net3074),
    .Q(\soc_inst.cpu_core.ex_branch_target[5] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25768_ (.RESET_B(net6800),
    .D(net3037),
    .Q(\soc_inst.cpu_core.ex_branch_target[6] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25769_ (.RESET_B(net6784),
    .D(net2911),
    .Q(\soc_inst.cpu_core.ex_branch_target[7] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25770_ (.RESET_B(net6785),
    .D(net2840),
    .Q(\soc_inst.cpu_core.ex_branch_target[8] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25771_ (.RESET_B(net6780),
    .D(net2781),
    .Q(\soc_inst.cpu_core.ex_branch_target[9] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _25772_ (.RESET_B(net6780),
    .D(_02352_),
    .Q(\soc_inst.cpu_core.ex_branch_target[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _25773_ (.RESET_B(net6785),
    .D(net1514),
    .Q(\soc_inst.cpu_core.ex_branch_target[11] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _25774_ (.RESET_B(net6734),
    .D(net2742),
    .Q(\soc_inst.cpu_core.ex_branch_target[12] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25775_ (.RESET_B(net6732),
    .D(net2447),
    .Q(\soc_inst.cpu_core.ex_branch_target[13] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25776_ (.RESET_B(net6731),
    .D(net2819),
    .Q(\soc_inst.cpu_core.ex_branch_target[14] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _25777_ (.RESET_B(net6726),
    .D(net2860),
    .Q(\soc_inst.cpu_core.ex_branch_target[15] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _25778_ (.RESET_B(net6757),
    .D(_02358_),
    .Q(\soc_inst.cpu_core.ex_branch_target[16] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _25779_ (.RESET_B(net6727),
    .D(net3035),
    .Q(\soc_inst.cpu_core.ex_branch_target[17] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _25780_ (.RESET_B(net6759),
    .D(net2477),
    .Q(\soc_inst.cpu_core.ex_branch_target[18] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _25781_ (.RESET_B(net6760),
    .D(net2442),
    .Q(\soc_inst.cpu_core.ex_branch_target[19] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _25782_ (.RESET_B(net6759),
    .D(net2720),
    .Q(\soc_inst.cpu_core.ex_branch_target[20] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _25783_ (.RESET_B(net6760),
    .D(net2755),
    .Q(\soc_inst.cpu_core.ex_branch_target[21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _25784_ (.RESET_B(net6758),
    .D(_02364_),
    .Q(\soc_inst.cpu_core.ex_branch_target[22] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _25785_ (.RESET_B(net6758),
    .D(_02365_),
    .Q(\soc_inst.cpu_core.ex_branch_target[23] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _25786_ (.RESET_B(net6769),
    .D(net2524),
    .Q(\soc_inst.cpu_core.ex_branch_target[24] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_2 _25787_ (.RESET_B(net6769),
    .D(net2682),
    .Q(\soc_inst.cpu_core.ex_branch_target[25] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _25788_ (.RESET_B(net6770),
    .D(net2304),
    .Q(\soc_inst.cpu_core.ex_branch_target[26] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _25789_ (.RESET_B(net6775),
    .D(net3094),
    .Q(\soc_inst.cpu_core.ex_branch_target[27] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _25790_ (.RESET_B(net6774),
    .D(net2618),
    .Q(\soc_inst.cpu_core.ex_branch_target[28] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _25791_ (.RESET_B(net6770),
    .D(net2470),
    .Q(\soc_inst.cpu_core.ex_branch_target[29] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _25792_ (.RESET_B(net6776),
    .D(net2415),
    .Q(\soc_inst.cpu_core.ex_branch_target[30] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_2 _25793_ (.RESET_B(net6778),
    .D(net1905),
    .Q(\soc_inst.cpu_core.ex_branch_target[31] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25794_ (.RESET_B(net6637),
    .D(net3370),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _25795_ (.RESET_B(net6637),
    .D(net3346),
    .Q(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _25796_ (.RESET_B(net6718),
    .D(net2313),
    .Q(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25797_ (.RESET_B(net6738),
    .D(net1203),
    .Q(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _25798_ (.RESET_B(net6680),
    .D(net2265),
    .Q(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25799_ (.RESET_B(net6717),
    .D(_02379_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25800_ (.RESET_B(net6740),
    .D(_02380_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _25801_ (.RESET_B(net6717),
    .D(net2262),
    .Q(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25802_ (.RESET_B(net6715),
    .D(_02382_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _25803_ (.RESET_B(net6716),
    .D(net2459),
    .Q(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25804_ (.RESET_B(net6717),
    .D(_02384_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25805_ (.RESET_B(net6712),
    .D(_02385_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _25806_ (.RESET_B(net6710),
    .D(_02386_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25807_ (.RESET_B(net6714),
    .D(_02387_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _25808_ (.RESET_B(net6712),
    .D(_02388_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _25809_ (.RESET_B(net6716),
    .D(net772),
    .Q(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25810_ (.RESET_B(net6713),
    .D(_02390_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _25811_ (.RESET_B(net6713),
    .D(_02391_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_1 _25812_ (.RESET_B(net6709),
    .D(_02392_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25813_ (.RESET_B(net6675),
    .D(_02393_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25814_ (.RESET_B(net6712),
    .D(_02394_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_1 _25815_ (.RESET_B(net6673),
    .D(_02395_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _25816_ (.RESET_B(net6678),
    .D(_02396_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_2 _25817_ (.RESET_B(net6673),
    .D(_02397_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25818_ (.RESET_B(net6672),
    .D(_02398_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25819_ (.RESET_B(net6672),
    .D(_02399_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25820_ (.RESET_B(net6672),
    .D(_02400_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25821_ (.RESET_B(net6672),
    .D(_02401_),
    .Q(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25822_ (.RESET_B(net6679),
    .D(net3068),
    .Q(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _25823_ (.RESET_B(net6718),
    .D(net778),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _25824_ (.RESET_B(net6715),
    .D(net717),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _25825_ (.RESET_B(net6680),
    .D(net1195),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _25826_ (.RESET_B(net6717),
    .D(net502),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _25827_ (.RESET_B(net6740),
    .D(net1070),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _25828_ (.RESET_B(net6719),
    .D(net1058),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25829_ (.RESET_B(net6680),
    .D(net537),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[11] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25830_ (.RESET_B(net6681),
    .D(net695),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[12] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_2 _25831_ (.RESET_B(net6681),
    .D(net710),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[13] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25832_ (.RESET_B(net6709),
    .D(net518),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[14] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25833_ (.RESET_B(net6677),
    .D(net505),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[15] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25834_ (.RESET_B(net6713),
    .D(net1145),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[16] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_1 _25835_ (.RESET_B(net6709),
    .D(net1026),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[17] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _25836_ (.RESET_B(net6710),
    .D(net466),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[18] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25837_ (.RESET_B(net6713),
    .D(net613),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[19] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_1 _25838_ (.RESET_B(net6713),
    .D(net346),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[20] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _25839_ (.RESET_B(net6675),
    .D(net844),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_2 _25840_ (.RESET_B(net6674),
    .D(net1183),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[22] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _25841_ (.RESET_B(net6675),
    .D(net950),
    .Q(\soc_inst.cpu_core.csr_file.mtvec[23] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _25842_ (.RESET_B(net6740),
    .D(_02422_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _25843_ (.RESET_B(net6738),
    .D(_02423_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _25844_ (.RESET_B(net6715),
    .D(_02424_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25845_ (.RESET_B(net6718),
    .D(net1262),
    .Q(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25846_ (.RESET_B(net6740),
    .D(net1293),
    .Q(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25847_ (.RESET_B(net6719),
    .D(net1217),
    .Q(\soc_inst.cpu_core.csr_file.mepc[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25848_ (.RESET_B(net6729),
    .D(_02428_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[11] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25849_ (.RESET_B(net6716),
    .D(_02429_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[12] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25850_ (.RESET_B(net6717),
    .D(net2347),
    .Q(\soc_inst.cpu_core.csr_file.mepc[13] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_2 _25851_ (.RESET_B(net6714),
    .D(_02431_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[14] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _25852_ (.RESET_B(net6714),
    .D(_02432_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[15] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _25853_ (.RESET_B(net6724),
    .D(net2115),
    .Q(\soc_inst.cpu_core.csr_file.mepc[16] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _25854_ (.RESET_B(net6724),
    .D(_02434_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _25855_ (.RESET_B(net6710),
    .D(net2535),
    .Q(\soc_inst.cpu_core.csr_file.mepc[18] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _25856_ (.RESET_B(net6712),
    .D(_02436_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _25857_ (.RESET_B(net6713),
    .D(net1577),
    .Q(\soc_inst.cpu_core.csr_file.mepc[20] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _25858_ (.RESET_B(net6677),
    .D(_02438_),
    .Q(\soc_inst.cpu_core.csr_file.mepc[21] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25859_ (.RESET_B(net6677),
    .D(net2134),
    .Q(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _25860_ (.RESET_B(net6714),
    .D(net2461),
    .Q(\soc_inst.cpu_core.csr_file.mepc[23] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _25861_ (.RESET_B(net6678),
    .D(net3071),
    .Q(\soc_inst.cpu_core.csr_file.mcause[31] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _25862_ (.RESET_B(net6682),
    .D(net80),
    .Q(\soc_inst.cpu_core.csr_file.mip_tip ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _25863_ (.RESET_B(net6584),
    .D(net1106),
    .Q(\soc_inst.pwm_ena [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25864_ (.RESET_B(net6574),
    .D(\soc_inst.i2c_ena ),
    .Q(\soc_inst.i2c_inst.status_reg[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _25865_ (.RESET_B(net6574),
    .D(net92),
    .Q(\soc_inst.i2c_inst.status_reg[1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _25866_ (.RESET_B(net6570),
    .D(net90),
    .Q(\soc_inst.i2c_inst.status_reg[2] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25867_ (.RESET_B(net6573),
    .D(net82),
    .Q(\soc_inst.i2c_inst.status_reg[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _25868_ (.RESET_B(net6678),
    .D(_02443_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _25869_ (.RESET_B(net6680),
    .D(net2793),
    .Q(_00264_),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _25870_ (.RESET_B(net6681),
    .D(net2772),
    .Q(_00265_),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _25871_ (.RESET_B(net6580),
    .D(net705),
    .Q(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25872_ (.RESET_B(net6590),
    .D(net409),
    .Q(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25873_ (.RESET_B(net6593),
    .D(net246),
    .Q(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25874_ (.RESET_B(net6589),
    .D(net213),
    .Q(\soc_inst.gpio_inst.int_pend_reg[3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25875_ (.RESET_B(net6591),
    .D(net430),
    .Q(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25876_ (.RESET_B(net6589),
    .D(net292),
    .Q(\soc_inst.gpio_inst.int_pend_reg[1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _25877_ (.RESET_B(net6782),
    .D(net2810),
    .Q(\soc_inst.cpu_core.id_pc[0] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25878_ (.RESET_B(net6791),
    .D(net2094),
    .Q(\soc_inst.cpu_core.id_pc[1] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25879_ (.RESET_B(net6792),
    .D(net1317),
    .Q(\soc_inst.cpu_core.id_pc[2] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _25880_ (.RESET_B(net6784),
    .D(net2325),
    .Q(\soc_inst.cpu_core.id_pc[3] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _25881_ (.RESET_B(net6791),
    .D(net2047),
    .Q(\soc_inst.cpu_core.id_pc[4] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25882_ (.RESET_B(net6791),
    .D(net1749),
    .Q(\soc_inst.cpu_core.id_pc[5] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25883_ (.RESET_B(net6786),
    .D(net1947),
    .Q(\soc_inst.cpu_core.id_pc[6] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25884_ (.RESET_B(net6786),
    .D(net2272),
    .Q(\soc_inst.cpu_core.id_pc[7] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25885_ (.RESET_B(net6785),
    .D(net2259),
    .Q(\soc_inst.cpu_core.id_pc[8] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25886_ (.RESET_B(net6796),
    .D(_02461_),
    .Q(\soc_inst.cpu_core.id_pc[9] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25887_ (.RESET_B(net6796),
    .D(_02462_),
    .Q(\soc_inst.cpu_core.id_pc[10] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _25888_ (.RESET_B(net6796),
    .D(_02463_),
    .Q(\soc_inst.cpu_core.id_pc[11] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_2 _25889_ (.RESET_B(net6766),
    .D(_02464_),
    .Q(\soc_inst.cpu_core.id_pc[12] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_2 _25890_ (.RESET_B(net6765),
    .D(_02465_),
    .Q(\soc_inst.cpu_core.id_pc[13] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25891_ (.RESET_B(net6763),
    .D(_02466_),
    .Q(\soc_inst.cpu_core.id_pc[14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_2 _25892_ (.RESET_B(net6765),
    .D(_02467_),
    .Q(\soc_inst.cpu_core.id_pc[15] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_2 _25893_ (.RESET_B(net6771),
    .D(_02468_),
    .Q(\soc_inst.cpu_core.id_pc[16] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_2 _25894_ (.RESET_B(net6759),
    .D(_02469_),
    .Q(\soc_inst.cpu_core.id_pc[17] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _25895_ (.RESET_B(net6759),
    .D(_02470_),
    .Q(\soc_inst.cpu_core.id_pc[18] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _25896_ (.RESET_B(net6757),
    .D(_02471_),
    .Q(\soc_inst.cpu_core.id_pc[19] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_2 _25897_ (.RESET_B(net6773),
    .D(_02472_),
    .Q(\soc_inst.cpu_core.id_pc[20] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_2 _25898_ (.RESET_B(net6760),
    .D(net2079),
    .Q(\soc_inst.cpu_core.id_pc[21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _25899_ (.RESET_B(net6773),
    .D(_02474_),
    .Q(\soc_inst.cpu_core.id_pc[22] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_2 _25900_ (.RESET_B(net6760),
    .D(net2629),
    .Q(\soc_inst.cpu_core.id_pc[23] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_2 _25901_ (.RESET_B(net6680),
    .D(_00082_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _25902_ (.RESET_B(net6672),
    .D(_00063_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[13] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _25903_ (.RESET_B(net6683),
    .D(_00064_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[14] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _25904_ (.RESET_B(net6676),
    .D(_00065_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[15] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _25905_ (.RESET_B(net6676),
    .D(_00066_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[16] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _25906_ (.RESET_B(net6711),
    .D(_00067_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _25907_ (.RESET_B(net6710),
    .D(_00068_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[18] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _25908_ (.RESET_B(net6662),
    .D(_00069_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[19] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _25909_ (.RESET_B(net6671),
    .D(_00070_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _25910_ (.RESET_B(net6675),
    .D(_00071_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[21] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _25911_ (.RESET_B(net6676),
    .D(_00072_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[22] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _25912_ (.RESET_B(net6676),
    .D(_00073_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[23] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _25913_ (.RESET_B(net6671),
    .D(_00074_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[24] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _25914_ (.RESET_B(net6669),
    .D(_00075_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[25] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _25915_ (.RESET_B(net6671),
    .D(_00076_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[26] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _25916_ (.RESET_B(net6664),
    .D(_00077_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[27] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _25917_ (.RESET_B(net6672),
    .D(_00078_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[28] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _25918_ (.RESET_B(net6671),
    .D(_00079_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[29] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _25919_ (.RESET_B(net6671),
    .D(_00080_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[30] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _25920_ (.RESET_B(net6669),
    .D(_00081_),
    .Q(\soc_inst.cpu_core.csr_file.mstatus[31] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _25921_ (.RESET_B(net6642),
    .D(net2752),
    .Q(_00266_),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _25922_ (.RESET_B(net6641),
    .D(_00006_),
    .Q(\soc_inst.mem_ctrl.access_state[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _25923_ (.RESET_B(net6643),
    .D(net3282),
    .Q(\soc_inst.mem_ctrl.access_state[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _25924_ (.RESET_B(net6641),
    .D(_00008_),
    .Q(\soc_inst.mem_ctrl.access_state[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _25925_ (.RESET_B(net6644),
    .D(_00009_),
    .Q(\soc_inst.mem_ctrl.access_state[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _25926_ (.RESET_B(net6563),
    .D(net2038),
    .Q(_00267_),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _25927_ (.RESET_B(net6563),
    .D(net1704),
    .Q(_00268_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _25928_ (.RESET_B(net6564),
    .D(net2671),
    .Q(_00269_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25929_ (.RESET_B(net6563),
    .D(_02479_),
    .Q(_00270_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _25930_ (.RESET_B(net6563),
    .D(_02480_),
    .Q(_00271_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _25931_ (.RESET_B(net6563),
    .D(_02481_),
    .Q(_00272_),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _25932_ (.RESET_B(net6564),
    .D(_02482_),
    .Q(_00273_),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _25933_ (.RESET_B(net6564),
    .D(_02483_),
    .Q(_00274_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25934_ (.RESET_B(net6557),
    .D(_02484_),
    .Q(_00275_),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _25935_ (.RESET_B(net6558),
    .D(_02485_),
    .Q(_00276_),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _25936_ (.RESET_B(net6557),
    .D(_02486_),
    .Q(_00277_),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _25937_ (.RESET_B(net6602),
    .D(net2374),
    .Q(_00278_),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _25938_ (.RESET_B(net6602),
    .D(net1826),
    .Q(_00279_),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _25939_ (.RESET_B(net6557),
    .D(_02489_),
    .Q(_00280_),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _25940_ (.RESET_B(net6600),
    .D(_02490_),
    .Q(_00281_),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _25941_ (.RESET_B(net6600),
    .D(net2684),
    .Q(_00282_),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _25942_ (.RESET_B(net37),
    .D(net2387),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _25943_ (.RESET_B(net36),
    .D(net2513),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _25944_ (.RESET_B(net34),
    .D(net2195),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _25945_ (.RESET_B(net32),
    .D(net1995),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _25946_ (.RESET_B(net31),
    .D(net2016),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _25947_ (.RESET_B(net30),
    .D(net2970),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _25948_ (.RESET_B(net67),
    .D(_02498_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _25949_ (.RESET_B(net68),
    .D(_00019_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _25950_ (.RESET_B(net69),
    .D(net1843),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _25951_ (.RESET_B(net72),
    .D(_00021_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_1 _25952_ (.RESET_B(net29),
    .D(_00022_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _25953_ (.RESET_B(net6550),
    .D(_02499_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25954_ (.RESET_B(net6565),
    .D(net2161),
    .Q(_00283_),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _25955_ (.RESET_B(net6565),
    .D(net2111),
    .Q(_00284_),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _25956_ (.RESET_B(net6606),
    .D(net2003),
    .Q(_00285_),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _25957_ (.RESET_B(net6563),
    .D(_02503_),
    .Q(_00286_),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _25958_ (.RESET_B(net6563),
    .D(_02504_),
    .Q(_00287_),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _25959_ (.RESET_B(net6563),
    .D(_02505_),
    .Q(_00288_),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _25960_ (.RESET_B(net6564),
    .D(_02506_),
    .Q(_00289_),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25961_ (.RESET_B(net6564),
    .D(net1320),
    .Q(_00290_),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25962_ (.RESET_B(net6560),
    .D(_02508_),
    .Q(_00291_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _25963_ (.RESET_B(net6560),
    .D(net220),
    .Q(_00292_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _25964_ (.RESET_B(net6560),
    .D(_02510_),
    .Q(_00293_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _25965_ (.RESET_B(net6602),
    .D(net2228),
    .Q(_00294_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _25966_ (.RESET_B(net6602),
    .D(_02512_),
    .Q(_00295_),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _25967_ (.RESET_B(net6600),
    .D(_02513_),
    .Q(_00296_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _25968_ (.RESET_B(net6600),
    .D(net1458),
    .Q(_00297_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _25969_ (.RESET_B(net6600),
    .D(net1856),
    .Q(_00298_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _25970_ (.RESET_B(net6614),
    .D(net226),
    .Q(_00299_),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _25971_ (.RESET_B(net6614),
    .D(net161),
    .Q(_00300_),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _25972_ (.RESET_B(net6614),
    .D(net1273),
    .Q(_00301_),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _25973_ (.RESET_B(net6618),
    .D(net296),
    .Q(_00302_),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _25974_ (.RESET_B(net6618),
    .D(net549),
    .Q(_00303_),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _25975_ (.RESET_B(net6618),
    .D(net572),
    .Q(_00304_),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _25976_ (.RESET_B(net6618),
    .D(net1312),
    .Q(_00305_),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _25977_ (.RESET_B(net6618),
    .D(_02523_),
    .Q(_00306_),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_2 _25978_ (.RESET_B(net6616),
    .D(net269),
    .Q(_00307_),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _25979_ (.RESET_B(net6615),
    .D(net234),
    .Q(_00308_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _25980_ (.RESET_B(net6620),
    .D(net1017),
    .Q(_00309_),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _25981_ (.RESET_B(net6616),
    .D(net713),
    .Q(_00310_),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_2 _25982_ (.RESET_B(net6605),
    .D(net370),
    .Q(_00311_),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_2 _25983_ (.RESET_B(net6605),
    .D(net314),
    .Q(_00312_),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_2 _25984_ (.RESET_B(net6615),
    .D(net735),
    .Q(_00313_),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _25985_ (.RESET_B(net6616),
    .D(net855),
    .Q(_00314_),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _25986_ (.RESET_B(net6548),
    .D(_00172_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_en ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25987_ (.RESET_B(net6548),
    .D(net1649),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25988_ (.RESET_B(net6548),
    .D(net173),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _25989_ (.RESET_B(net6547),
    .D(_02534_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _25990_ (.RESET_B(net6548),
    .D(_02535_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _25991_ (.RESET_B(net6548),
    .D(_02536_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25992_ (.RESET_B(net6547),
    .D(_02537_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _25993_ (.RESET_B(net6547),
    .D(_02538_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _25994_ (.RESET_B(net6547),
    .D(_02539_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _25995_ (.RESET_B(net6550),
    .D(net2624),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25996_ (.RESET_B(net6551),
    .D(_00170_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_rx_break_reg ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25997_ (.RESET_B(net28),
    .D(net496),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _25998_ (.RESET_B(net26),
    .D(net2408),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _25999_ (.RESET_B(net24),
    .D(net1862),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _26000_ (.RESET_B(net22),
    .D(net2433),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _26001_ (.RESET_B(net20),
    .D(net2747),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _26002_ (.RESET_B(net18),
    .D(_02545_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _26003_ (.RESET_B(net16),
    .D(_02546_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _26004_ (.RESET_B(net14),
    .D(_02547_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _26005_ (.RESET_B(net73),
    .D(_02548_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _26006_ (.RESET_B(net65),
    .D(_02549_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _26007_ (.RESET_B(net64),
    .D(_02550_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _26008_ (.RESET_B(net62),
    .D(net1471),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _26009_ (.RESET_B(net60),
    .D(net2677),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _26010_ (.RESET_B(net58),
    .D(net2497),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_1 _26011_ (.RESET_B(net56),
    .D(_02554_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _26012_ (.RESET_B(net6553),
    .D(_02555_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _26013_ (.RESET_B(net6552),
    .D(_02556_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _26014_ (.RESET_B(net6548),
    .D(_02557_),
    .Q(_00315_),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _26015_ (.RESET_B(net6550),
    .D(_02558_),
    .Q(_00316_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _26016_ (.RESET_B(net6548),
    .D(_02559_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _26017_ (.RESET_B(net6552),
    .D(_02560_),
    .Q(_00317_),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _26018_ (.RESET_B(net6549),
    .D(_02561_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _26019_ (.RESET_B(net6549),
    .D(_02562_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _26020_ (.RESET_B(net6556),
    .D(_02563_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _26021_ (.RESET_B(net6554),
    .D(_02564_),
    .Q(_00318_),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _26022_ (.RESET_B(net46),
    .D(_02565_),
    .Q(\soc_inst.uart_tx [0]),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _26023_ (.RESET_B(net44),
    .D(net530),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _26024_ (.RESET_B(net42),
    .D(net1656),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _26025_ (.RESET_B(net41),
    .D(net922),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _26026_ (.RESET_B(net39),
    .D(net1993),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _26027_ (.RESET_B(net35),
    .D(net671),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _26028_ (.RESET_B(net27),
    .D(net2176),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _26029_ (.RESET_B(net23),
    .D(net1418),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _26030_ (.RESET_B(net19),
    .D(_02573_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _26031_ (.RESET_B(net15),
    .D(net667),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _26032_ (.RESET_B(net66),
    .D(net2010),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _26033_ (.RESET_B(net63),
    .D(_02576_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _26034_ (.RESET_B(net59),
    .D(_02577_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _26035_ (.RESET_B(net55),
    .D(net748),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _26036_ (.RESET_B(net53),
    .D(_02579_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _26037_ (.RESET_B(net51),
    .D(_02580_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _26038_ (.RESET_B(net49),
    .D(net304),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _26039_ (.RESET_B(net47),
    .D(net2090),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _26040_ (.RESET_B(net43),
    .D(_02583_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _26041_ (.RESET_B(net40),
    .D(net826),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _26042_ (.RESET_B(net33),
    .D(net1890),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _26043_ (.RESET_B(net21),
    .D(net1839),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _26044_ (.RESET_B(net74),
    .D(_02587_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26045_ (.RESET_B(net61),
    .D(_02588_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26046_ (.RESET_B(net54),
    .D(_02589_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _26047_ (.RESET_B(net50),
    .D(net3043),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _26048_ (.RESET_B(net45),
    .D(_02591_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26049_ (.RESET_B(net38),
    .D(net1646),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26050_ (.RESET_B(net17),
    .D(_02593_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26051_ (.RESET_B(net57),
    .D(_02594_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _26052_ (.RESET_B(net48),
    .D(net1744),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _26053_ (.RESET_B(net25),
    .D(_02596_),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_1 _26054_ (.RESET_B(net52),
    .D(net739),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _26055_ (.RESET_B(net76),
    .D(net800),
    .Q(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _26056_ (.RESET_B(net6593),
    .D(net168),
    .Q(\soc_inst.spi_inst.clk_counter[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _26057_ (.RESET_B(net6593),
    .D(net578),
    .Q(\soc_inst.spi_inst.clk_counter[1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _26058_ (.RESET_B(net6593),
    .D(net761),
    .Q(\soc_inst.spi_inst.clk_counter[2] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _26059_ (.RESET_B(net6593),
    .D(net1902),
    .Q(\soc_inst.spi_inst.clk_counter[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _26060_ (.RESET_B(net6593),
    .D(net2778),
    .Q(\soc_inst.spi_inst.clk_counter[4] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _26061_ (.RESET_B(net6592),
    .D(net2208),
    .Q(\soc_inst.spi_inst.clk_counter[5] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _26062_ (.RESET_B(net6585),
    .D(net2622),
    .Q(\soc_inst.spi_inst.clk_counter[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _26063_ (.RESET_B(net6585),
    .D(net463),
    .Q(\soc_inst.spi_inst.clk_counter[7] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_tiehi _26031__15 (.L_HI(net15));
 sg13g2_tiehi _26003__16 (.L_HI(net16));
 sg13g2_tiehi _26050__17 (.L_HI(net17));
 sg13g2_tiehi _26002__18 (.L_HI(net18));
 sg13g2_tiehi _26030__19 (.L_HI(net19));
 sg13g2_tiehi _26001__20 (.L_HI(net20));
 sg13g2_tiehi _26043__21 (.L_HI(net21));
 sg13g2_tiehi _26000__22 (.L_HI(net22));
 sg13g2_tiehi _26029__23 (.L_HI(net23));
 sg13g2_tiehi _25999__24 (.L_HI(net24));
 sg13g2_tiehi _26053__25 (.L_HI(net25));
 sg13g2_tiehi _25998__26 (.L_HI(net26));
 sg13g2_tiehi _26028__27 (.L_HI(net27));
 sg13g2_tiehi _25997__28 (.L_HI(net28));
 sg13g2_tiehi _25952__29 (.L_HI(net29));
 sg13g2_tiehi _25947__30 (.L_HI(net30));
 sg13g2_tiehi _25946__31 (.L_HI(net31));
 sg13g2_tiehi _25945__32 (.L_HI(net32));
 sg13g2_tiehi _26042__33 (.L_HI(net33));
 sg13g2_tiehi _25944__34 (.L_HI(net34));
 sg13g2_tiehi _26027__35 (.L_HI(net35));
 sg13g2_tiehi _25943__36 (.L_HI(net36));
 sg13g2_tiehi _25942__37 (.L_HI(net37));
 sg13g2_tiehi _26049__38 (.L_HI(net38));
 sg13g2_tiehi _26026__39 (.L_HI(net39));
 sg13g2_tiehi _26041__40 (.L_HI(net40));
 sg13g2_tiehi _26025__41 (.L_HI(net41));
 sg13g2_tiehi _26024__42 (.L_HI(net42));
 sg13g2_tiehi _26040__43 (.L_HI(net43));
 sg13g2_tiehi _26023__44 (.L_HI(net44));
 sg13g2_tiehi _26048__45 (.L_HI(net45));
 sg13g2_tiehi _26022__46 (.L_HI(net46));
 sg13g2_tiehi _26039__47 (.L_HI(net47));
 sg13g2_tiehi _26052__48 (.L_HI(net48));
 sg13g2_tiehi _26038__49 (.L_HI(net49));
 sg13g2_tiehi _26047__50 (.L_HI(net50));
 sg13g2_tiehi _26037__51 (.L_HI(net51));
 sg13g2_tiehi _26054__52 (.L_HI(net52));
 sg13g2_tiehi _26036__53 (.L_HI(net53));
 sg13g2_tiehi _26046__54 (.L_HI(net54));
 sg13g2_tiehi _26035__55 (.L_HI(net55));
 sg13g2_tiehi _26011__56 (.L_HI(net56));
 sg13g2_tiehi _26051__57 (.L_HI(net57));
 sg13g2_tiehi _26010__58 (.L_HI(net58));
 sg13g2_tiehi _26034__59 (.L_HI(net59));
 sg13g2_tiehi _26009__60 (.L_HI(net60));
 sg13g2_tiehi _26045__61 (.L_HI(net61));
 sg13g2_tiehi _26008__62 (.L_HI(net62));
 sg13g2_tiehi _26033__63 (.L_HI(net63));
 sg13g2_tiehi _26007__64 (.L_HI(net64));
 sg13g2_tiehi _26006__65 (.L_HI(net65));
 sg13g2_tiehi _26032__66 (.L_HI(net66));
 sg13g2_tiehi _25948__67 (.L_HI(net67));
 sg13g2_tiehi _25949__68 (.L_HI(net68));
 sg13g2_tiehi _25950__69 (.L_HI(net69));
 sg13g2_tiehi _24191__70 (.L_HI(net70));
 sg13g2_tiehi _24190__71 (.L_HI(net71));
 sg13g2_tiehi _25951__72 (.L_HI(net72));
 sg13g2_tiehi _26005__73 (.L_HI(net73));
 sg13g2_tiehi _26044__74 (.L_HI(net74));
 sg13g2_tiehi _24130__75 (.L_HI(net75));
 sg13g2_tiehi _26055__76 (.L_HI(net76));
 sg13g2_tiehi tt_um_SotaSoC_77 (.L_HI(net77));
 sg13g2_tiehi tt_um_SotaSoC_78 (.L_HI(net78));
 sg13g2_tiehi tt_um_SotaSoC_79 (.L_HI(net79));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _26130_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _26131_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_2 _26132_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_8 _26133_ (.A(\soc_inst.flash_cs_n ),
    .X(uio_out[0]));
 sg13g2_buf_1 _26134_ (.A(\soc_inst.bus_spi_sclk ),
    .X(uio_out[3]));
 sg13g2_buf_8 _26135_ (.A(\soc_inst.mem_ctrl.ram_cs_n ),
    .X(uio_out[6]));
 sg13g2_buf_8 _26136_ (.A(\soc_inst.uart_tx [0]),
    .X(uo_out[0]));
 sg13g2_buf_8 _26137_ (.A(\soc_inst.cpu_core.error_flag_reg ),
    .X(uo_out[1]));
 sg13g2_buf_1 _26138_ (.A(\soc_inst.gpio_inst.gpio_out[1] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _26139_ (.A(\soc_inst.gpio_inst.gpio_out[5] ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_8 fanout4690 (.A(net4693),
    .X(net4690));
 sg13g2_buf_8 fanout4691 (.A(net4692),
    .X(net4691));
 sg13g2_buf_8 fanout4692 (.A(net4693),
    .X(net4692));
 sg13g2_buf_8 fanout4693 (.A(_10720_),
    .X(net4693));
 sg13g2_buf_8 fanout4694 (.A(net4699),
    .X(net4694));
 sg13g2_buf_1 fanout4695 (.A(net4699),
    .X(net4695));
 sg13g2_buf_8 fanout4696 (.A(net4697),
    .X(net4696));
 sg13g2_buf_1 fanout4697 (.A(net4699),
    .X(net4697));
 sg13g2_buf_8 fanout4698 (.A(net4699),
    .X(net4698));
 sg13g2_buf_8 fanout4699 (.A(_10720_),
    .X(net4699));
 sg13g2_buf_8 fanout4700 (.A(net4704),
    .X(net4700));
 sg13g2_buf_8 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_8 fanout4702 (.A(net4704),
    .X(net4702));
 sg13g2_buf_8 fanout4703 (.A(net4704),
    .X(net4703));
 sg13g2_buf_8 fanout4704 (.A(_10195_),
    .X(net4704));
 sg13g2_buf_2 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(net4707),
    .X(net4706));
 sg13g2_buf_8 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_8 fanout4708 (.A(_10167_),
    .X(net4708));
 sg13g2_buf_8 fanout4709 (.A(net4710),
    .X(net4709));
 sg13g2_buf_1 fanout4710 (.A(net4711),
    .X(net4710));
 sg13g2_buf_1 fanout4711 (.A(net4712),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(_10167_),
    .X(net4712));
 sg13g2_buf_8 fanout4713 (.A(_06818_),
    .X(net4713));
 sg13g2_buf_1 fanout4714 (.A(_06818_),
    .X(net4714));
 sg13g2_buf_8 fanout4715 (.A(net4716),
    .X(net4715));
 sg13g2_buf_8 fanout4716 (.A(_06737_),
    .X(net4716));
 sg13g2_buf_8 fanout4717 (.A(net4718),
    .X(net4717));
 sg13g2_buf_8 fanout4718 (.A(_07434_),
    .X(net4718));
 sg13g2_buf_8 fanout4719 (.A(net4721),
    .X(net4719));
 sg13g2_buf_8 fanout4720 (.A(net4721),
    .X(net4720));
 sg13g2_buf_8 fanout4721 (.A(_11428_),
    .X(net4721));
 sg13g2_buf_8 fanout4722 (.A(_11428_),
    .X(net4722));
 sg13g2_buf_8 fanout4723 (.A(net4725),
    .X(net4723));
 sg13g2_buf_1 fanout4724 (.A(net4725),
    .X(net4724));
 sg13g2_buf_8 fanout4725 (.A(_11134_),
    .X(net4725));
 sg13g2_buf_8 fanout4726 (.A(net4727),
    .X(net4726));
 sg13g2_buf_8 fanout4727 (.A(_11133_),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(_11133_),
    .X(net4728));
 sg13g2_buf_8 fanout4729 (.A(net4730),
    .X(net4729));
 sg13g2_buf_8 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(net4732),
    .X(net4731));
 sg13g2_buf_8 fanout4732 (.A(_09946_),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(net4734),
    .X(net4733));
 sg13g2_buf_8 fanout4734 (.A(net4735),
    .X(net4734));
 sg13g2_buf_8 fanout4735 (.A(_09946_),
    .X(net4735));
 sg13g2_buf_1 fanout4736 (.A(net4738),
    .X(net4736));
 sg13g2_buf_8 fanout4737 (.A(net4738),
    .X(net4737));
 sg13g2_buf_8 fanout4738 (.A(_09046_),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(net4740),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(_08910_),
    .X(net4740));
 sg13g2_buf_8 fanout4741 (.A(net4742),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(_07433_),
    .X(net4742));
 sg13g2_buf_8 fanout4743 (.A(net4744),
    .X(net4743));
 sg13g2_buf_8 fanout4744 (.A(_07414_),
    .X(net4744));
 sg13g2_buf_1 fanout4745 (.A(_07414_),
    .X(net4745));
 sg13g2_buf_8 fanout4746 (.A(net4749),
    .X(net4746));
 sg13g2_buf_8 fanout4747 (.A(net4748),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(net4749),
    .X(net4748));
 sg13g2_buf_8 fanout4749 (.A(_07206_),
    .X(net4749));
 sg13g2_buf_8 fanout4750 (.A(net4752),
    .X(net4750));
 sg13g2_buf_8 fanout4751 (.A(net4752),
    .X(net4751));
 sg13g2_buf_2 fanout4752 (.A(_11427_),
    .X(net4752));
 sg13g2_buf_8 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_8 fanout4754 (.A(_11427_),
    .X(net4754));
 sg13g2_buf_8 fanout4755 (.A(_09924_),
    .X(net4755));
 sg13g2_buf_1 fanout4756 (.A(_09924_),
    .X(net4756));
 sg13g2_buf_8 fanout4757 (.A(net4758),
    .X(net4757));
 sg13g2_buf_8 fanout4758 (.A(net4759),
    .X(net4758));
 sg13g2_buf_8 fanout4759 (.A(_09924_),
    .X(net4759));
 sg13g2_buf_8 fanout4760 (.A(_09896_),
    .X(net4760));
 sg13g2_buf_8 fanout4761 (.A(_09059_),
    .X(net4761));
 sg13g2_buf_8 fanout4762 (.A(net4767),
    .X(net4762));
 sg13g2_buf_1 fanout4763 (.A(net4767),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(net4766),
    .X(net4764));
 sg13g2_buf_8 fanout4765 (.A(net4767),
    .X(net4765));
 sg13g2_buf_1 fanout4766 (.A(net4767),
    .X(net4766));
 sg13g2_buf_2 fanout4767 (.A(_09725_),
    .X(net4767));
 sg13g2_buf_8 fanout4768 (.A(net4769),
    .X(net4768));
 sg13g2_buf_8 fanout4769 (.A(net4771),
    .X(net4769));
 sg13g2_buf_8 fanout4770 (.A(net4771),
    .X(net4770));
 sg13g2_buf_2 fanout4771 (.A(net4772),
    .X(net4771));
 sg13g2_buf_8 fanout4772 (.A(_09698_),
    .X(net4772));
 sg13g2_buf_8 fanout4773 (.A(net4778),
    .X(net4773));
 sg13g2_buf_1 fanout4774 (.A(net4778),
    .X(net4774));
 sg13g2_buf_8 fanout4775 (.A(net4777),
    .X(net4775));
 sg13g2_buf_1 fanout4776 (.A(net4777),
    .X(net4776));
 sg13g2_buf_8 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_8 fanout4778 (.A(_09632_),
    .X(net4778));
 sg13g2_buf_8 fanout4779 (.A(net4783),
    .X(net4779));
 sg13g2_buf_2 fanout4780 (.A(net4783),
    .X(net4780));
 sg13g2_buf_8 fanout4781 (.A(net4783),
    .X(net4781));
 sg13g2_buf_8 fanout4782 (.A(net4783),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(_09603_),
    .X(net4783));
 sg13g2_buf_8 fanout4784 (.A(_09144_),
    .X(net4784));
 sg13g2_buf_8 fanout4785 (.A(_09144_),
    .X(net4785));
 sg13g2_buf_8 fanout4786 (.A(net4787),
    .X(net4786));
 sg13g2_buf_2 fanout4787 (.A(net4791),
    .X(net4787));
 sg13g2_buf_8 fanout4788 (.A(net4791),
    .X(net4788));
 sg13g2_buf_8 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_8 fanout4790 (.A(net4791),
    .X(net4790));
 sg13g2_buf_8 fanout4791 (.A(_09060_),
    .X(net4791));
 sg13g2_buf_8 fanout4792 (.A(_09038_),
    .X(net4792));
 sg13g2_buf_8 fanout4793 (.A(net4797),
    .X(net4793));
 sg13g2_buf_1 fanout4794 (.A(net4797),
    .X(net4794));
 sg13g2_buf_8 fanout4795 (.A(net4796),
    .X(net4795));
 sg13g2_buf_8 fanout4796 (.A(net4797),
    .X(net4796));
 sg13g2_buf_8 fanout4797 (.A(_11128_),
    .X(net4797));
 sg13g2_buf_2 fanout4798 (.A(net4799),
    .X(net4798));
 sg13g2_buf_1 fanout4799 (.A(net4801),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(net4801),
    .X(net4800));
 sg13g2_buf_1 fanout4801 (.A(net4802),
    .X(net4801));
 sg13g2_buf_8 fanout4802 (.A(net4809),
    .X(net4802));
 sg13g2_buf_8 fanout4803 (.A(net4805),
    .X(net4803));
 sg13g2_buf_8 fanout4804 (.A(net4805),
    .X(net4804));
 sg13g2_buf_8 fanout4805 (.A(net4809),
    .X(net4805));
 sg13g2_buf_2 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_1 fanout4807 (.A(net4808),
    .X(net4807));
 sg13g2_buf_1 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_2 fanout4809 (.A(_11023_),
    .X(net4809));
 sg13g2_buf_8 fanout4810 (.A(net4811),
    .X(net4810));
 sg13g2_buf_1 fanout4811 (.A(net4814),
    .X(net4811));
 sg13g2_buf_8 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_1 fanout4813 (.A(net4814),
    .X(net4813));
 sg13g2_buf_1 fanout4814 (.A(net4821),
    .X(net4814));
 sg13g2_buf_8 fanout4815 (.A(net4816),
    .X(net4815));
 sg13g2_buf_8 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_8 fanout4817 (.A(net4821),
    .X(net4817));
 sg13g2_buf_8 fanout4818 (.A(net4819),
    .X(net4818));
 sg13g2_buf_8 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_8 fanout4820 (.A(net4821),
    .X(net4820));
 sg13g2_buf_8 fanout4821 (.A(_09821_),
    .X(net4821));
 sg13g2_buf_8 fanout4822 (.A(net4825),
    .X(net4822));
 sg13g2_buf_8 fanout4823 (.A(net4825),
    .X(net4823));
 sg13g2_buf_1 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_8 fanout4825 (.A(net4826),
    .X(net4825));
 sg13g2_buf_8 fanout4826 (.A(_09807_),
    .X(net4826));
 sg13g2_buf_8 fanout4827 (.A(net4831),
    .X(net4827));
 sg13g2_buf_1 fanout4828 (.A(net4831),
    .X(net4828));
 sg13g2_buf_8 fanout4829 (.A(net4831),
    .X(net4829));
 sg13g2_buf_8 fanout4830 (.A(net4831),
    .X(net4830));
 sg13g2_buf_8 fanout4831 (.A(_09799_),
    .X(net4831));
 sg13g2_buf_8 fanout4832 (.A(net4835),
    .X(net4832));
 sg13g2_buf_8 fanout4833 (.A(net4834),
    .X(net4833));
 sg13g2_buf_8 fanout4834 (.A(net4835),
    .X(net4834));
 sg13g2_buf_8 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(_09791_),
    .X(net4836));
 sg13g2_buf_8 fanout4837 (.A(net4840),
    .X(net4837));
 sg13g2_buf_8 fanout4838 (.A(net4839),
    .X(net4838));
 sg13g2_buf_8 fanout4839 (.A(net4840),
    .X(net4839));
 sg13g2_buf_8 fanout4840 (.A(net4841),
    .X(net4840));
 sg13g2_buf_8 fanout4841 (.A(_09783_),
    .X(net4841));
 sg13g2_buf_8 fanout4842 (.A(_09775_),
    .X(net4842));
 sg13g2_buf_1 fanout4843 (.A(_09775_),
    .X(net4843));
 sg13g2_buf_8 fanout4844 (.A(net4845),
    .X(net4844));
 sg13g2_buf_2 fanout4845 (.A(net4846),
    .X(net4845));
 sg13g2_buf_8 fanout4846 (.A(_09775_),
    .X(net4846));
 sg13g2_buf_8 fanout4847 (.A(net4848),
    .X(net4847));
 sg13g2_buf_8 fanout4848 (.A(net4851),
    .X(net4848));
 sg13g2_buf_8 fanout4849 (.A(net4850),
    .X(net4849));
 sg13g2_buf_8 fanout4850 (.A(net4851),
    .X(net4850));
 sg13g2_buf_8 fanout4851 (.A(_09767_),
    .X(net4851));
 sg13g2_buf_8 fanout4852 (.A(net4856),
    .X(net4852));
 sg13g2_buf_1 fanout4853 (.A(_09759_),
    .X(net4853));
 sg13g2_buf_8 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_8 fanout4855 (.A(net4856),
    .X(net4855));
 sg13g2_buf_8 fanout4856 (.A(_09759_),
    .X(net4856));
 sg13g2_buf_8 fanout4857 (.A(net4861),
    .X(net4857));
 sg13g2_buf_1 fanout4858 (.A(net4861),
    .X(net4858));
 sg13g2_buf_8 fanout4859 (.A(net4860),
    .X(net4859));
 sg13g2_buf_8 fanout4860 (.A(net4861),
    .X(net4860));
 sg13g2_buf_8 fanout4861 (.A(_09751_),
    .X(net4861));
 sg13g2_buf_8 fanout4862 (.A(net4866),
    .X(net4862));
 sg13g2_buf_8 fanout4863 (.A(net4865),
    .X(net4863));
 sg13g2_buf_1 fanout4864 (.A(net4865),
    .X(net4864));
 sg13g2_buf_8 fanout4865 (.A(net4866),
    .X(net4865));
 sg13g2_buf_8 fanout4866 (.A(_09743_),
    .X(net4866));
 sg13g2_buf_8 fanout4867 (.A(_09734_),
    .X(net4867));
 sg13g2_buf_8 fanout4868 (.A(net4871),
    .X(net4868));
 sg13g2_buf_8 fanout4869 (.A(net4871),
    .X(net4869));
 sg13g2_buf_1 fanout4870 (.A(net4871),
    .X(net4870));
 sg13g2_buf_8 fanout4871 (.A(_09734_),
    .X(net4871));
 sg13g2_buf_8 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_1 fanout4873 (.A(net4877),
    .X(net4873));
 sg13g2_buf_8 fanout4874 (.A(net4876),
    .X(net4874));
 sg13g2_buf_1 fanout4875 (.A(net4876),
    .X(net4875));
 sg13g2_buf_8 fanout4876 (.A(net4877),
    .X(net4876));
 sg13g2_buf_8 fanout4877 (.A(_09716_),
    .X(net4877));
 sg13g2_buf_8 fanout4878 (.A(net4880),
    .X(net4878));
 sg13g2_buf_8 fanout4879 (.A(net4883),
    .X(net4879));
 sg13g2_buf_1 fanout4880 (.A(net4883),
    .X(net4880));
 sg13g2_buf_8 fanout4881 (.A(net4883),
    .X(net4881));
 sg13g2_buf_1 fanout4882 (.A(net4883),
    .X(net4882));
 sg13g2_buf_2 fanout4883 (.A(_09707_),
    .X(net4883));
 sg13g2_buf_8 fanout4884 (.A(net4888),
    .X(net4884));
 sg13g2_buf_8 fanout4885 (.A(net4887),
    .X(net4885));
 sg13g2_buf_1 fanout4886 (.A(net4887),
    .X(net4886));
 sg13g2_buf_8 fanout4887 (.A(net4888),
    .X(net4887));
 sg13g2_buf_8 fanout4888 (.A(_09689_),
    .X(net4888));
 sg13g2_buf_8 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_1 fanout4890 (.A(_09680_),
    .X(net4890));
 sg13g2_buf_8 fanout4891 (.A(net4893),
    .X(net4891));
 sg13g2_buf_8 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_8 fanout4893 (.A(_09680_),
    .X(net4893));
 sg13g2_buf_8 fanout4894 (.A(net4897),
    .X(net4894));
 sg13g2_buf_8 fanout4895 (.A(net4896),
    .X(net4895));
 sg13g2_buf_8 fanout4896 (.A(net4897),
    .X(net4896));
 sg13g2_buf_8 fanout4897 (.A(net4898),
    .X(net4897));
 sg13g2_buf_8 fanout4898 (.A(_09669_),
    .X(net4898));
 sg13g2_buf_8 fanout4899 (.A(net4903),
    .X(net4899));
 sg13g2_buf_1 fanout4900 (.A(net4903),
    .X(net4900));
 sg13g2_buf_8 fanout4901 (.A(net4903),
    .X(net4901));
 sg13g2_buf_1 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(net4904),
    .X(net4903));
 sg13g2_buf_8 fanout4904 (.A(_09641_),
    .X(net4904));
 sg13g2_buf_8 fanout4905 (.A(net4910),
    .X(net4905));
 sg13g2_buf_1 fanout4906 (.A(net4910),
    .X(net4906));
 sg13g2_buf_8 fanout4907 (.A(net4909),
    .X(net4907));
 sg13g2_buf_1 fanout4908 (.A(net4909),
    .X(net4908));
 sg13g2_buf_8 fanout4909 (.A(net4910),
    .X(net4909));
 sg13g2_buf_8 fanout4910 (.A(_09621_),
    .X(net4910));
 sg13g2_buf_8 fanout4911 (.A(net4915),
    .X(net4911));
 sg13g2_buf_2 fanout4912 (.A(net4915),
    .X(net4912));
 sg13g2_buf_8 fanout4913 (.A(net4914),
    .X(net4913));
 sg13g2_buf_8 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_8 fanout4915 (.A(_09612_),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4917),
    .X(net4916));
 sg13g2_buf_8 fanout4917 (.A(_09589_),
    .X(net4917));
 sg13g2_buf_8 fanout4918 (.A(net4919),
    .X(net4918));
 sg13g2_buf_8 fanout4919 (.A(_09589_),
    .X(net4919));
 sg13g2_buf_8 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_8 fanout4921 (.A(net4924),
    .X(net4921));
 sg13g2_buf_8 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_8 fanout4923 (.A(net4924),
    .X(net4923));
 sg13g2_buf_8 fanout4924 (.A(_09390_),
    .X(net4924));
 sg13g2_buf_8 fanout4925 (.A(net4928),
    .X(net4925));
 sg13g2_buf_8 fanout4926 (.A(net4927),
    .X(net4926));
 sg13g2_buf_2 fanout4927 (.A(net4928),
    .X(net4927));
 sg13g2_buf_8 fanout4928 (.A(net4930),
    .X(net4928));
 sg13g2_buf_8 fanout4929 (.A(net4930),
    .X(net4929));
 sg13g2_buf_8 fanout4930 (.A(_09142_),
    .X(net4930));
 sg13g2_buf_2 fanout4931 (.A(net4932),
    .X(net4931));
 sg13g2_buf_8 fanout4932 (.A(net4933),
    .X(net4932));
 sg13g2_buf_1 fanout4933 (.A(net4935),
    .X(net4933));
 sg13g2_buf_8 fanout4934 (.A(net4935),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(_09118_),
    .X(net4935));
 sg13g2_buf_8 fanout4936 (.A(_09043_),
    .X(net4936));
 sg13g2_buf_8 fanout4937 (.A(net4938),
    .X(net4937));
 sg13g2_buf_8 fanout4938 (.A(net4939),
    .X(net4938));
 sg13g2_buf_8 fanout4939 (.A(_08971_),
    .X(net4939));
 sg13g2_buf_8 fanout4940 (.A(net4941),
    .X(net4940));
 sg13g2_buf_2 fanout4941 (.A(net4942),
    .X(net4941));
 sg13g2_buf_8 fanout4942 (.A(_08971_),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_8 fanout4944 (.A(net4945),
    .X(net4944));
 sg13g2_buf_8 fanout4945 (.A(net4953),
    .X(net4945));
 sg13g2_buf_8 fanout4946 (.A(net4947),
    .X(net4946));
 sg13g2_buf_8 fanout4947 (.A(net4953),
    .X(net4947));
 sg13g2_buf_8 fanout4948 (.A(net4952),
    .X(net4948));
 sg13g2_buf_8 fanout4949 (.A(net4950),
    .X(net4949));
 sg13g2_buf_8 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_8 fanout4951 (.A(net4952),
    .X(net4951));
 sg13g2_buf_2 fanout4952 (.A(net4953),
    .X(net4952));
 sg13g2_buf_8 fanout4953 (.A(_08970_),
    .X(net4953));
 sg13g2_buf_8 fanout4954 (.A(net4955),
    .X(net4954));
 sg13g2_buf_8 fanout4955 (.A(net4958),
    .X(net4955));
 sg13g2_buf_8 fanout4956 (.A(net4957),
    .X(net4956));
 sg13g2_buf_8 fanout4957 (.A(net4958),
    .X(net4957));
 sg13g2_buf_8 fanout4958 (.A(_09659_),
    .X(net4958));
 sg13g2_buf_8 fanout4959 (.A(net4960),
    .X(net4959));
 sg13g2_buf_2 fanout4960 (.A(_09650_),
    .X(net4960));
 sg13g2_buf_8 fanout4961 (.A(net4963),
    .X(net4961));
 sg13g2_buf_1 fanout4962 (.A(net4963),
    .X(net4962));
 sg13g2_buf_8 fanout4963 (.A(_09650_),
    .X(net4963));
 sg13g2_buf_8 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_8 fanout4965 (.A(net4968),
    .X(net4965));
 sg13g2_buf_8 fanout4966 (.A(net4968),
    .X(net4966));
 sg13g2_buf_1 fanout4967 (.A(net4968),
    .X(net4967));
 sg13g2_buf_8 fanout4968 (.A(_09578_),
    .X(net4968));
 sg13g2_buf_8 fanout4969 (.A(net4970),
    .X(net4969));
 sg13g2_buf_8 fanout4970 (.A(net4973),
    .X(net4970));
 sg13g2_buf_8 fanout4971 (.A(net4972),
    .X(net4971));
 sg13g2_buf_8 fanout4972 (.A(net4973),
    .X(net4972));
 sg13g2_buf_2 fanout4973 (.A(_09569_),
    .X(net4973));
 sg13g2_buf_8 fanout4974 (.A(net4977),
    .X(net4974));
 sg13g2_buf_8 fanout4975 (.A(net4976),
    .X(net4975));
 sg13g2_buf_8 fanout4976 (.A(net4977),
    .X(net4976));
 sg13g2_buf_8 fanout4977 (.A(net4978),
    .X(net4977));
 sg13g2_buf_8 fanout4978 (.A(_09560_),
    .X(net4978));
 sg13g2_buf_8 fanout4979 (.A(net4980),
    .X(net4979));
 sg13g2_buf_8 fanout4980 (.A(net4982),
    .X(net4980));
 sg13g2_buf_8 fanout4981 (.A(net4982),
    .X(net4981));
 sg13g2_buf_2 fanout4982 (.A(net4983),
    .X(net4982));
 sg13g2_buf_8 fanout4983 (.A(_09551_),
    .X(net4983));
 sg13g2_buf_8 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_2 fanout4985 (.A(_09542_),
    .X(net4985));
 sg13g2_buf_8 fanout4986 (.A(net4988),
    .X(net4986));
 sg13g2_buf_8 fanout4987 (.A(net4988),
    .X(net4987));
 sg13g2_buf_8 fanout4988 (.A(_09542_),
    .X(net4988));
 sg13g2_buf_8 fanout4989 (.A(net4993),
    .X(net4989));
 sg13g2_buf_8 fanout4990 (.A(net4993),
    .X(net4990));
 sg13g2_buf_8 fanout4991 (.A(net4993),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(net4993),
    .X(net4992));
 sg13g2_buf_8 fanout4993 (.A(_09533_),
    .X(net4993));
 sg13g2_buf_8 fanout4994 (.A(net4997),
    .X(net4994));
 sg13g2_buf_8 fanout4995 (.A(net4997),
    .X(net4995));
 sg13g2_buf_8 fanout4996 (.A(net4997),
    .X(net4996));
 sg13g2_buf_8 fanout4997 (.A(net4998),
    .X(net4997));
 sg13g2_buf_8 fanout4998 (.A(_09524_),
    .X(net4998));
 sg13g2_buf_8 fanout4999 (.A(_08968_),
    .X(net4999));
 sg13g2_buf_1 fanout5000 (.A(_08968_),
    .X(net5000));
 sg13g2_buf_8 fanout5001 (.A(net5002),
    .X(net5001));
 sg13g2_buf_8 fanout5002 (.A(net5008),
    .X(net5002));
 sg13g2_buf_8 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_1 fanout5004 (.A(net5005),
    .X(net5004));
 sg13g2_buf_1 fanout5005 (.A(net5006),
    .X(net5005));
 sg13g2_buf_8 fanout5006 (.A(net5008),
    .X(net5006));
 sg13g2_buf_8 fanout5007 (.A(net5008),
    .X(net5007));
 sg13g2_buf_8 fanout5008 (.A(_08967_),
    .X(net5008));
 sg13g2_buf_8 fanout5009 (.A(net5010),
    .X(net5009));
 sg13g2_buf_8 fanout5010 (.A(net5011),
    .X(net5010));
 sg13g2_buf_2 fanout5011 (.A(_08703_),
    .X(net5011));
 sg13g2_buf_8 fanout5012 (.A(net5013),
    .X(net5012));
 sg13g2_buf_8 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_1 fanout5014 (.A(net5015),
    .X(net5014));
 sg13g2_buf_8 fanout5015 (.A(_08703_),
    .X(net5015));
 sg13g2_buf_8 fanout5016 (.A(net5017),
    .X(net5016));
 sg13g2_buf_8 fanout5017 (.A(net5023),
    .X(net5017));
 sg13g2_buf_8 fanout5018 (.A(net5022),
    .X(net5018));
 sg13g2_buf_8 fanout5019 (.A(net5020),
    .X(net5019));
 sg13g2_buf_1 fanout5020 (.A(net5021),
    .X(net5020));
 sg13g2_buf_8 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_8 fanout5022 (.A(net5023),
    .X(net5022));
 sg13g2_buf_8 fanout5023 (.A(_08703_),
    .X(net5023));
 sg13g2_buf_8 fanout5024 (.A(_07722_),
    .X(net5024));
 sg13g2_buf_8 fanout5025 (.A(net5026),
    .X(net5025));
 sg13g2_buf_8 fanout5026 (.A(net5029),
    .X(net5026));
 sg13g2_buf_8 fanout5027 (.A(net5028),
    .X(net5027));
 sg13g2_buf_8 fanout5028 (.A(net5029),
    .X(net5028));
 sg13g2_buf_2 fanout5029 (.A(_10782_),
    .X(net5029));
 sg13g2_buf_8 fanout5030 (.A(net5034),
    .X(net5030));
 sg13g2_buf_8 fanout5031 (.A(net5034),
    .X(net5031));
 sg13g2_buf_8 fanout5032 (.A(net5033),
    .X(net5032));
 sg13g2_buf_8 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_8 fanout5034 (.A(_10782_),
    .X(net5034));
 sg13g2_buf_8 fanout5035 (.A(net5036),
    .X(net5035));
 sg13g2_buf_8 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(_10266_),
    .X(net5037));
 sg13g2_buf_8 fanout5038 (.A(net5039),
    .X(net5038));
 sg13g2_buf_8 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_8 fanout5040 (.A(net5041),
    .X(net5040));
 sg13g2_buf_2 fanout5041 (.A(_10266_),
    .X(net5041));
 sg13g2_buf_8 fanout5042 (.A(net5044),
    .X(net5042));
 sg13g2_buf_8 fanout5043 (.A(net5044),
    .X(net5043));
 sg13g2_buf_8 fanout5044 (.A(_10266_),
    .X(net5044));
 sg13g2_buf_2 fanout5045 (.A(net5046),
    .X(net5045));
 sg13g2_buf_2 fanout5046 (.A(_08966_),
    .X(net5046));
 sg13g2_buf_8 fanout5047 (.A(net5048),
    .X(net5047));
 sg13g2_buf_8 fanout5048 (.A(_08966_),
    .X(net5048));
 sg13g2_buf_8 fanout5049 (.A(_08487_),
    .X(net5049));
 sg13g2_buf_8 fanout5050 (.A(net5051),
    .X(net5050));
 sg13g2_buf_1 fanout5051 (.A(net5052),
    .X(net5051));
 sg13g2_buf_8 fanout5052 (.A(_07706_),
    .X(net5052));
 sg13g2_buf_8 fanout5053 (.A(_07674_),
    .X(net5053));
 sg13g2_buf_8 fanout5054 (.A(_07619_),
    .X(net5054));
 sg13g2_buf_8 fanout5055 (.A(net5058),
    .X(net5055));
 sg13g2_buf_8 fanout5056 (.A(net5057),
    .X(net5056));
 sg13g2_buf_8 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_8 fanout5058 (.A(_10861_),
    .X(net5058));
 sg13g2_buf_2 fanout5059 (.A(net5060),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net5061),
    .X(net5060));
 sg13g2_buf_1 fanout5061 (.A(_10523_),
    .X(net5061));
 sg13g2_buf_8 fanout5062 (.A(net5064),
    .X(net5062));
 sg13g2_buf_8 fanout5063 (.A(net5064),
    .X(net5063));
 sg13g2_buf_8 fanout5064 (.A(_09994_),
    .X(net5064));
 sg13g2_buf_8 fanout5065 (.A(net5068),
    .X(net5065));
 sg13g2_buf_1 fanout5066 (.A(net5068),
    .X(net5066));
 sg13g2_buf_8 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_8 fanout5068 (.A(_09994_),
    .X(net5068));
 sg13g2_buf_8 fanout5069 (.A(_09811_),
    .X(net5069));
 sg13g2_buf_1 fanout5070 (.A(_09811_),
    .X(net5070));
 sg13g2_buf_8 fanout5071 (.A(net5073),
    .X(net5071));
 sg13g2_buf_1 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(_08963_),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(net5075),
    .X(net5074));
 sg13g2_buf_2 fanout5075 (.A(net5076),
    .X(net5075));
 sg13g2_buf_2 fanout5076 (.A(_08962_),
    .X(net5076));
 sg13g2_buf_8 fanout5077 (.A(net5078),
    .X(net5077));
 sg13g2_buf_8 fanout5078 (.A(net5088),
    .X(net5078));
 sg13g2_buf_2 fanout5079 (.A(net5080),
    .X(net5079));
 sg13g2_buf_2 fanout5080 (.A(net5081),
    .X(net5080));
 sg13g2_buf_1 fanout5081 (.A(net5088),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(net5084),
    .X(net5082));
 sg13g2_buf_1 fanout5083 (.A(net5084),
    .X(net5083));
 sg13g2_buf_2 fanout5084 (.A(net5086),
    .X(net5084));
 sg13g2_buf_2 fanout5085 (.A(net5086),
    .X(net5085));
 sg13g2_buf_1 fanout5086 (.A(net5087),
    .X(net5086));
 sg13g2_buf_1 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(_07641_),
    .X(net5088));
 sg13g2_buf_8 fanout5089 (.A(net5091),
    .X(net5089));
 sg13g2_buf_1 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(_07601_),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(net5093),
    .X(net5092));
 sg13g2_buf_8 fanout5093 (.A(_07601_),
    .X(net5093));
 sg13g2_buf_8 fanout5094 (.A(_05254_),
    .X(net5094));
 sg13g2_buf_8 fanout5095 (.A(net5096),
    .X(net5095));
 sg13g2_buf_8 fanout5096 (.A(_04397_),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(_04337_),
    .X(net5097));
 sg13g2_buf_8 fanout5098 (.A(net5099),
    .X(net5098));
 sg13g2_buf_8 fanout5099 (.A(_04287_),
    .X(net5099));
 sg13g2_buf_8 fanout5100 (.A(net5101),
    .X(net5100));
 sg13g2_buf_8 fanout5101 (.A(_04285_),
    .X(net5101));
 sg13g2_buf_8 fanout5102 (.A(net5104),
    .X(net5102));
 sg13g2_buf_8 fanout5103 (.A(net5104),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(_11761_),
    .X(net5104));
 sg13g2_buf_8 fanout5105 (.A(_11761_),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(_11761_),
    .X(net5106));
 sg13g2_buf_8 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_1 fanout5108 (.A(_11312_),
    .X(net5108));
 sg13g2_buf_8 fanout5109 (.A(net5111),
    .X(net5109));
 sg13g2_buf_1 fanout5110 (.A(net5111),
    .X(net5110));
 sg13g2_buf_1 fanout5111 (.A(net5112),
    .X(net5111));
 sg13g2_buf_8 fanout5112 (.A(net5113),
    .X(net5112));
 sg13g2_buf_8 fanout5113 (.A(_10879_),
    .X(net5113));
 sg13g2_buf_8 fanout5114 (.A(_10867_),
    .X(net5114));
 sg13g2_buf_1 fanout5115 (.A(_10867_),
    .X(net5115));
 sg13g2_buf_8 fanout5116 (.A(_10860_),
    .X(net5116));
 sg13g2_buf_8 fanout5117 (.A(net5118),
    .X(net5117));
 sg13g2_buf_8 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_8 fanout5119 (.A(_10854_),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(net5121),
    .X(net5120));
 sg13g2_buf_2 fanout5121 (.A(_10854_),
    .X(net5121));
 sg13g2_buf_8 fanout5122 (.A(_10853_),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(_10321_),
    .X(net5123));
 sg13g2_buf_2 fanout5124 (.A(net5125),
    .X(net5124));
 sg13g2_buf_2 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_8 fanout5126 (.A(_10309_),
    .X(net5126));
 sg13g2_buf_8 fanout5127 (.A(_10309_),
    .X(net5127));
 sg13g2_buf_8 fanout5128 (.A(net5129),
    .X(net5128));
 sg13g2_buf_8 fanout5129 (.A(_10307_),
    .X(net5129));
 sg13g2_buf_8 fanout5130 (.A(net5132),
    .X(net5130));
 sg13g2_buf_2 fanout5131 (.A(net5132),
    .X(net5131));
 sg13g2_buf_8 fanout5132 (.A(_09993_),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(net5134),
    .X(net5133));
 sg13g2_buf_8 fanout5134 (.A(_09443_),
    .X(net5134));
 sg13g2_buf_8 fanout5135 (.A(net5136),
    .X(net5135));
 sg13g2_buf_8 fanout5136 (.A(net5137),
    .X(net5136));
 sg13g2_buf_8 fanout5137 (.A(_09425_),
    .X(net5137));
 sg13g2_buf_8 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_1 fanout5139 (.A(net5141),
    .X(net5139));
 sg13g2_buf_8 fanout5140 (.A(net5141),
    .X(net5140));
 sg13g2_buf_8 fanout5141 (.A(_09368_),
    .X(net5141));
 sg13g2_buf_8 fanout5142 (.A(net5144),
    .X(net5142));
 sg13g2_buf_1 fanout5143 (.A(net5144),
    .X(net5143));
 sg13g2_buf_8 fanout5144 (.A(net5146),
    .X(net5144));
 sg13g2_buf_8 fanout5145 (.A(net5146),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(net5147),
    .X(net5146));
 sg13g2_buf_1 fanout5147 (.A(_09141_),
    .X(net5147));
 sg13g2_buf_8 fanout5148 (.A(net5150),
    .X(net5148));
 sg13g2_buf_8 fanout5149 (.A(_09141_),
    .X(net5149));
 sg13g2_buf_1 fanout5150 (.A(_09141_),
    .X(net5150));
 sg13g2_buf_8 fanout5151 (.A(net5153),
    .X(net5151));
 sg13g2_buf_1 fanout5152 (.A(net5153),
    .X(net5152));
 sg13g2_buf_8 fanout5153 (.A(net5154),
    .X(net5153));
 sg13g2_buf_8 fanout5154 (.A(_09022_),
    .X(net5154));
 sg13g2_buf_8 fanout5155 (.A(net5157),
    .X(net5155));
 sg13g2_buf_8 fanout5156 (.A(_09022_),
    .X(net5156));
 sg13g2_buf_2 fanout5157 (.A(_09022_),
    .X(net5157));
 sg13g2_buf_8 fanout5158 (.A(net5159),
    .X(net5158));
 sg13g2_buf_8 fanout5159 (.A(_08965_),
    .X(net5159));
 sg13g2_buf_8 fanout5160 (.A(net5161),
    .X(net5160));
 sg13g2_buf_2 fanout5161 (.A(net5162),
    .X(net5161));
 sg13g2_buf_1 fanout5162 (.A(net5163),
    .X(net5162));
 sg13g2_buf_8 fanout5163 (.A(_08964_),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(net5165),
    .X(net5164));
 sg13g2_buf_2 fanout5165 (.A(net5168),
    .X(net5165));
 sg13g2_buf_8 fanout5166 (.A(net5168),
    .X(net5166));
 sg13g2_buf_1 fanout5167 (.A(net5168),
    .X(net5167));
 sg13g2_buf_8 fanout5168 (.A(_08951_),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(_08950_),
    .X(net5169));
 sg13g2_buf_8 fanout5170 (.A(net5172),
    .X(net5170));
 sg13g2_buf_1 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(_08909_),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(_08909_),
    .X(net5173));
 sg13g2_buf_2 fanout5174 (.A(_08909_),
    .X(net5174));
 sg13g2_buf_8 fanout5175 (.A(_08822_),
    .X(net5175));
 sg13g2_buf_8 fanout5176 (.A(net5178),
    .X(net5176));
 sg13g2_buf_1 fanout5177 (.A(net5178),
    .X(net5177));
 sg13g2_buf_8 fanout5178 (.A(_08821_),
    .X(net5178));
 sg13g2_buf_8 fanout5179 (.A(net5180),
    .X(net5179));
 sg13g2_buf_8 fanout5180 (.A(net5185),
    .X(net5180));
 sg13g2_buf_8 fanout5181 (.A(net5183),
    .X(net5181));
 sg13g2_buf_8 fanout5182 (.A(net5183),
    .X(net5182));
 sg13g2_buf_8 fanout5183 (.A(net5184),
    .X(net5183));
 sg13g2_buf_8 fanout5184 (.A(net5185),
    .X(net5184));
 sg13g2_buf_8 fanout5185 (.A(net5187),
    .X(net5185));
 sg13g2_buf_8 fanout5186 (.A(net5187),
    .X(net5186));
 sg13g2_buf_8 fanout5187 (.A(_08678_),
    .X(net5187));
 sg13g2_buf_8 fanout5188 (.A(net5192),
    .X(net5188));
 sg13g2_buf_2 fanout5189 (.A(net5191),
    .X(net5189));
 sg13g2_buf_8 fanout5190 (.A(net5191),
    .X(net5190));
 sg13g2_buf_8 fanout5191 (.A(net5192),
    .X(net5191));
 sg13g2_buf_8 fanout5192 (.A(_08241_),
    .X(net5192));
 sg13g2_buf_8 fanout5193 (.A(_08241_),
    .X(net5193));
 sg13g2_buf_8 fanout5194 (.A(net5195),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(net5196),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(_08240_),
    .X(net5196));
 sg13g2_buf_8 fanout5197 (.A(_08240_),
    .X(net5197));
 sg13g2_buf_8 fanout5198 (.A(net5200),
    .X(net5198));
 sg13g2_buf_1 fanout5199 (.A(net5200),
    .X(net5199));
 sg13g2_buf_8 fanout5200 (.A(net5208),
    .X(net5200));
 sg13g2_buf_8 fanout5201 (.A(net5208),
    .X(net5201));
 sg13g2_buf_8 fanout5202 (.A(net5208),
    .X(net5202));
 sg13g2_buf_8 fanout5203 (.A(net5204),
    .X(net5203));
 sg13g2_buf_8 fanout5204 (.A(net5207),
    .X(net5204));
 sg13g2_buf_8 fanout5205 (.A(net5207),
    .X(net5205));
 sg13g2_buf_8 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_8 fanout5207 (.A(net5208),
    .X(net5207));
 sg13g2_buf_8 fanout5208 (.A(_06394_),
    .X(net5208));
 sg13g2_buf_8 fanout5209 (.A(net5210),
    .X(net5209));
 sg13g2_buf_8 fanout5210 (.A(net5213),
    .X(net5210));
 sg13g2_buf_8 fanout5211 (.A(net5213),
    .X(net5211));
 sg13g2_buf_8 fanout5212 (.A(net5213),
    .X(net5212));
 sg13g2_buf_8 fanout5213 (.A(_06328_),
    .X(net5213));
 sg13g2_buf_8 fanout5214 (.A(net5215),
    .X(net5214));
 sg13g2_buf_8 fanout5215 (.A(net5218),
    .X(net5215));
 sg13g2_buf_8 fanout5216 (.A(net5217),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(net5218),
    .X(net5217));
 sg13g2_buf_8 fanout5218 (.A(_06328_),
    .X(net5218));
 sg13g2_buf_8 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_8 fanout5220 (.A(net5223),
    .X(net5220));
 sg13g2_buf_8 fanout5221 (.A(net5223),
    .X(net5221));
 sg13g2_buf_8 fanout5222 (.A(net5223),
    .X(net5222));
 sg13g2_buf_8 fanout5223 (.A(net5229),
    .X(net5223));
 sg13g2_buf_8 fanout5224 (.A(net5226),
    .X(net5224));
 sg13g2_buf_1 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_8 fanout5226 (.A(net5229),
    .X(net5226));
 sg13g2_buf_8 fanout5227 (.A(net5228),
    .X(net5227));
 sg13g2_buf_8 fanout5228 (.A(net5229),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(_06229_),
    .X(net5229));
 sg13g2_buf_8 fanout5230 (.A(net5234),
    .X(net5230));
 sg13g2_buf_8 fanout5231 (.A(net5234),
    .X(net5231));
 sg13g2_buf_8 fanout5232 (.A(net5234),
    .X(net5232));
 sg13g2_buf_8 fanout5233 (.A(net5234),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(net5240),
    .X(net5234));
 sg13g2_buf_8 fanout5235 (.A(net5237),
    .X(net5235));
 sg13g2_buf_8 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(net5240),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(net5239),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(net5240),
    .X(net5239));
 sg13g2_buf_8 fanout5240 (.A(_06196_),
    .X(net5240));
 sg13g2_buf_8 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_8 fanout5242 (.A(_04556_),
    .X(net5242));
 sg13g2_buf_8 fanout5243 (.A(net5244),
    .X(net5243));
 sg13g2_buf_8 fanout5244 (.A(_04357_),
    .X(net5244));
 sg13g2_buf_8 fanout5245 (.A(net5246),
    .X(net5245));
 sg13g2_buf_8 fanout5246 (.A(net5247),
    .X(net5246));
 sg13g2_buf_8 fanout5247 (.A(_04331_),
    .X(net5247));
 sg13g2_buf_8 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(_04331_),
    .X(net5249));
 sg13g2_buf_8 fanout5250 (.A(_04266_),
    .X(net5250));
 sg13g2_buf_8 fanout5251 (.A(net5255),
    .X(net5251));
 sg13g2_buf_8 fanout5252 (.A(net5255),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5255),
    .X(net5254));
 sg13g2_buf_8 fanout5255 (.A(_03469_),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(net5260),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(net5260),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(net5259),
    .X(net5258));
 sg13g2_buf_8 fanout5259 (.A(net5260),
    .X(net5259));
 sg13g2_buf_8 fanout5260 (.A(_03468_),
    .X(net5260));
 sg13g2_buf_8 fanout5261 (.A(net5265),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(net5265),
    .X(net5262));
 sg13g2_buf_8 fanout5263 (.A(net5264),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5265),
    .X(net5264));
 sg13g2_buf_8 fanout5265 (.A(_03465_),
    .X(net5265));
 sg13g2_buf_8 fanout5266 (.A(net5270),
    .X(net5266));
 sg13g2_buf_8 fanout5267 (.A(net5270),
    .X(net5267));
 sg13g2_buf_8 fanout5268 (.A(net5269),
    .X(net5268));
 sg13g2_buf_8 fanout5269 (.A(net5270),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(_03461_),
    .X(net5270));
 sg13g2_buf_8 fanout5271 (.A(net5275),
    .X(net5271));
 sg13g2_buf_8 fanout5272 (.A(net5275),
    .X(net5272));
 sg13g2_buf_8 fanout5273 (.A(net5275),
    .X(net5273));
 sg13g2_buf_8 fanout5274 (.A(net5275),
    .X(net5274));
 sg13g2_buf_8 fanout5275 (.A(_03456_),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5280),
    .X(net5276));
 sg13g2_buf_8 fanout5277 (.A(net5280),
    .X(net5277));
 sg13g2_buf_8 fanout5278 (.A(net5279),
    .X(net5278));
 sg13g2_buf_8 fanout5279 (.A(net5280),
    .X(net5279));
 sg13g2_buf_8 fanout5280 (.A(_03450_),
    .X(net5280));
 sg13g2_buf_8 fanout5281 (.A(net5285),
    .X(net5281));
 sg13g2_buf_8 fanout5282 (.A(net5285),
    .X(net5282));
 sg13g2_buf_8 fanout5283 (.A(net5284),
    .X(net5283));
 sg13g2_buf_8 fanout5284 (.A(net5285),
    .X(net5284));
 sg13g2_buf_8 fanout5285 (.A(_03444_),
    .X(net5285));
 sg13g2_buf_8 fanout5286 (.A(net5290),
    .X(net5286));
 sg13g2_buf_8 fanout5287 (.A(net5290),
    .X(net5287));
 sg13g2_buf_8 fanout5288 (.A(net5289),
    .X(net5288));
 sg13g2_buf_8 fanout5289 (.A(net5290),
    .X(net5289));
 sg13g2_buf_8 fanout5290 (.A(_03437_),
    .X(net5290));
 sg13g2_buf_8 fanout5291 (.A(net5294),
    .X(net5291));
 sg13g2_buf_8 fanout5292 (.A(net5293),
    .X(net5292));
 sg13g2_buf_8 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_8 fanout5294 (.A(_03430_),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(_03430_),
    .X(net5295));
 sg13g2_buf_8 fanout5296 (.A(net5297),
    .X(net5296));
 sg13g2_buf_8 fanout5297 (.A(net5299),
    .X(net5297));
 sg13g2_buf_8 fanout5298 (.A(net5299),
    .X(net5298));
 sg13g2_buf_8 fanout5299 (.A(_02674_),
    .X(net5299));
 sg13g2_buf_8 fanout5300 (.A(net5304),
    .X(net5300));
 sg13g2_buf_8 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_8 fanout5302 (.A(net5303),
    .X(net5302));
 sg13g2_buf_8 fanout5303 (.A(net5304),
    .X(net5303));
 sg13g2_buf_8 fanout5304 (.A(net5311),
    .X(net5304));
 sg13g2_buf_8 fanout5305 (.A(net5307),
    .X(net5305));
 sg13g2_buf_1 fanout5306 (.A(net5307),
    .X(net5306));
 sg13g2_buf_8 fanout5307 (.A(net5311),
    .X(net5307));
 sg13g2_buf_8 fanout5308 (.A(net5310),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(net5310),
    .X(net5309));
 sg13g2_buf_8 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_8 fanout5311 (.A(_11391_),
    .X(net5311));
 sg13g2_buf_8 fanout5312 (.A(net5313),
    .X(net5312));
 sg13g2_buf_8 fanout5313 (.A(_11025_),
    .X(net5313));
 sg13g2_buf_8 fanout5314 (.A(net5318),
    .X(net5314));
 sg13g2_buf_8 fanout5315 (.A(net5317),
    .X(net5315));
 sg13g2_buf_1 fanout5316 (.A(net5317),
    .X(net5316));
 sg13g2_buf_1 fanout5317 (.A(net5318),
    .X(net5317));
 sg13g2_buf_8 fanout5318 (.A(_10863_),
    .X(net5318));
 sg13g2_buf_2 fanout5319 (.A(net5320),
    .X(net5319));
 sg13g2_buf_8 fanout5320 (.A(_10856_),
    .X(net5320));
 sg13g2_buf_8 fanout5321 (.A(net5322),
    .X(net5321));
 sg13g2_buf_2 fanout5322 (.A(net5323),
    .X(net5322));
 sg13g2_buf_1 fanout5323 (.A(net5325),
    .X(net5323));
 sg13g2_buf_8 fanout5324 (.A(net5325),
    .X(net5324));
 sg13g2_buf_1 fanout5325 (.A(_10169_),
    .X(net5325));
 sg13g2_buf_8 fanout5326 (.A(_09899_),
    .X(net5326));
 sg13g2_buf_8 fanout5327 (.A(_09836_),
    .X(net5327));
 sg13g2_buf_8 fanout5328 (.A(_09836_),
    .X(net5328));
 sg13g2_buf_8 fanout5329 (.A(net5330),
    .X(net5329));
 sg13g2_buf_8 fanout5330 (.A(_09672_),
    .X(net5330));
 sg13g2_buf_8 fanout5331 (.A(net5332),
    .X(net5331));
 sg13g2_buf_8 fanout5332 (.A(net5333),
    .X(net5332));
 sg13g2_buf_8 fanout5333 (.A(_09516_),
    .X(net5333));
 sg13g2_buf_8 fanout5334 (.A(_09516_),
    .X(net5334));
 sg13g2_buf_1 fanout5335 (.A(_09516_),
    .X(net5335));
 sg13g2_buf_8 fanout5336 (.A(_09367_),
    .X(net5336));
 sg13g2_buf_8 fanout5337 (.A(_09367_),
    .X(net5337));
 sg13g2_buf_8 fanout5338 (.A(net5339),
    .X(net5338));
 sg13g2_buf_2 fanout5339 (.A(net5340),
    .X(net5339));
 sg13g2_buf_8 fanout5340 (.A(net5341),
    .X(net5340));
 sg13g2_buf_8 fanout5341 (.A(_09116_),
    .X(net5341));
 sg13g2_buf_8 fanout5342 (.A(net5343),
    .X(net5342));
 sg13g2_buf_8 fanout5343 (.A(net5344),
    .X(net5343));
 sg13g2_buf_2 fanout5344 (.A(_09116_),
    .X(net5344));
 sg13g2_buf_8 fanout5345 (.A(net5349),
    .X(net5345));
 sg13g2_buf_1 fanout5346 (.A(net5349),
    .X(net5346));
 sg13g2_buf_8 fanout5347 (.A(net5349),
    .X(net5347));
 sg13g2_buf_8 fanout5348 (.A(net5349),
    .X(net5348));
 sg13g2_buf_8 fanout5349 (.A(_09057_),
    .X(net5349));
 sg13g2_buf_8 fanout5350 (.A(net5351),
    .X(net5350));
 sg13g2_buf_8 fanout5351 (.A(_09017_),
    .X(net5351));
 sg13g2_buf_8 fanout5352 (.A(_09017_),
    .X(net5352));
 sg13g2_buf_1 fanout5353 (.A(_09017_),
    .X(net5353));
 sg13g2_buf_8 fanout5354 (.A(_08955_),
    .X(net5354));
 sg13g2_buf_2 fanout5355 (.A(net5357),
    .X(net5355));
 sg13g2_buf_1 fanout5356 (.A(net5357),
    .X(net5356));
 sg13g2_buf_1 fanout5357 (.A(net5358),
    .X(net5357));
 sg13g2_buf_8 fanout5358 (.A(_08954_),
    .X(net5358));
 sg13g2_buf_8 fanout5359 (.A(net5361),
    .X(net5359));
 sg13g2_buf_2 fanout5360 (.A(net5361),
    .X(net5360));
 sg13g2_buf_8 fanout5361 (.A(_08954_),
    .X(net5361));
 sg13g2_buf_8 fanout5362 (.A(net5364),
    .X(net5362));
 sg13g2_buf_2 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_8 fanout5364 (.A(_08906_),
    .X(net5364));
 sg13g2_buf_8 fanout5365 (.A(_08857_),
    .X(net5365));
 sg13g2_buf_8 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_2 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_2 fanout5368 (.A(_08832_),
    .X(net5368));
 sg13g2_buf_8 fanout5369 (.A(net5370),
    .X(net5369));
 sg13g2_buf_8 fanout5370 (.A(_06710_),
    .X(net5370));
 sg13g2_buf_8 fanout5371 (.A(net5372),
    .X(net5371));
 sg13g2_buf_8 fanout5372 (.A(net5375),
    .X(net5372));
 sg13g2_buf_8 fanout5373 (.A(net5375),
    .X(net5373));
 sg13g2_buf_8 fanout5374 (.A(net5375),
    .X(net5374));
 sg13g2_buf_8 fanout5375 (.A(_06493_),
    .X(net5375));
 sg13g2_buf_8 fanout5376 (.A(net5377),
    .X(net5376));
 sg13g2_buf_8 fanout5377 (.A(net5380),
    .X(net5377));
 sg13g2_buf_8 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_8 fanout5379 (.A(net5380),
    .X(net5379));
 sg13g2_buf_8 fanout5380 (.A(_06493_),
    .X(net5380));
 sg13g2_buf_8 fanout5381 (.A(net5385),
    .X(net5381));
 sg13g2_buf_8 fanout5382 (.A(net5385),
    .X(net5382));
 sg13g2_buf_8 fanout5383 (.A(net5385),
    .X(net5383));
 sg13g2_buf_8 fanout5384 (.A(net5385),
    .X(net5384));
 sg13g2_buf_8 fanout5385 (.A(_06460_),
    .X(net5385));
 sg13g2_buf_8 fanout5386 (.A(net5390),
    .X(net5386));
 sg13g2_buf_8 fanout5387 (.A(net5390),
    .X(net5387));
 sg13g2_buf_8 fanout5388 (.A(net5390),
    .X(net5388));
 sg13g2_buf_8 fanout5389 (.A(net5390),
    .X(net5389));
 sg13g2_buf_8 fanout5390 (.A(_06460_),
    .X(net5390));
 sg13g2_buf_8 fanout5391 (.A(net5392),
    .X(net5391));
 sg13g2_buf_8 fanout5392 (.A(net5395),
    .X(net5392));
 sg13g2_buf_8 fanout5393 (.A(net5394),
    .X(net5393));
 sg13g2_buf_8 fanout5394 (.A(net5395),
    .X(net5394));
 sg13g2_buf_8 fanout5395 (.A(_06361_),
    .X(net5395));
 sg13g2_buf_8 fanout5396 (.A(net5397),
    .X(net5396));
 sg13g2_buf_8 fanout5397 (.A(net5400),
    .X(net5397));
 sg13g2_buf_8 fanout5398 (.A(net5400),
    .X(net5398));
 sg13g2_buf_8 fanout5399 (.A(net5400),
    .X(net5399));
 sg13g2_buf_8 fanout5400 (.A(_06361_),
    .X(net5400));
 sg13g2_buf_8 fanout5401 (.A(net5402),
    .X(net5401));
 sg13g2_buf_8 fanout5402 (.A(net5405),
    .X(net5402));
 sg13g2_buf_8 fanout5403 (.A(net5405),
    .X(net5403));
 sg13g2_buf_8 fanout5404 (.A(net5405),
    .X(net5404));
 sg13g2_buf_8 fanout5405 (.A(_06096_),
    .X(net5405));
 sg13g2_buf_8 fanout5406 (.A(net5407),
    .X(net5406));
 sg13g2_buf_8 fanout5407 (.A(net5410),
    .X(net5407));
 sg13g2_buf_8 fanout5408 (.A(net5409),
    .X(net5408));
 sg13g2_buf_8 fanout5409 (.A(net5410),
    .X(net5409));
 sg13g2_buf_8 fanout5410 (.A(_06096_),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(net5412),
    .X(net5411));
 sg13g2_buf_8 fanout5412 (.A(net5415),
    .X(net5412));
 sg13g2_buf_8 fanout5413 (.A(net5415),
    .X(net5413));
 sg13g2_buf_8 fanout5414 (.A(net5415),
    .X(net5414));
 sg13g2_buf_8 fanout5415 (.A(_05897_),
    .X(net5415));
 sg13g2_buf_8 fanout5416 (.A(net5417),
    .X(net5416));
 sg13g2_buf_8 fanout5417 (.A(net5420),
    .X(net5417));
 sg13g2_buf_8 fanout5418 (.A(net5420),
    .X(net5418));
 sg13g2_buf_8 fanout5419 (.A(net5420),
    .X(net5419));
 sg13g2_buf_8 fanout5420 (.A(_05897_),
    .X(net5420));
 sg13g2_buf_8 fanout5421 (.A(net5426),
    .X(net5421));
 sg13g2_buf_1 fanout5422 (.A(net5426),
    .X(net5422));
 sg13g2_buf_8 fanout5423 (.A(net5426),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(net5426),
    .X(net5424));
 sg13g2_buf_1 fanout5425 (.A(net5426),
    .X(net5425));
 sg13g2_buf_8 fanout5426 (.A(_05695_),
    .X(net5426));
 sg13g2_buf_8 fanout5427 (.A(net5431),
    .X(net5427));
 sg13g2_buf_8 fanout5428 (.A(net5431),
    .X(net5428));
 sg13g2_buf_8 fanout5429 (.A(net5431),
    .X(net5429));
 sg13g2_buf_8 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_8 fanout5431 (.A(_05695_),
    .X(net5431));
 sg13g2_buf_8 fanout5432 (.A(net5433),
    .X(net5432));
 sg13g2_buf_8 fanout5433 (.A(net5436),
    .X(net5433));
 sg13g2_buf_8 fanout5434 (.A(net5436),
    .X(net5434));
 sg13g2_buf_8 fanout5435 (.A(net5436),
    .X(net5435));
 sg13g2_buf_8 fanout5436 (.A(_05627_),
    .X(net5436));
 sg13g2_buf_8 fanout5437 (.A(net5441),
    .X(net5437));
 sg13g2_buf_8 fanout5438 (.A(net5441),
    .X(net5438));
 sg13g2_buf_8 fanout5439 (.A(net5440),
    .X(net5439));
 sg13g2_buf_8 fanout5440 (.A(net5441),
    .X(net5440));
 sg13g2_buf_8 fanout5441 (.A(_05627_),
    .X(net5441));
 sg13g2_buf_8 fanout5442 (.A(net5443),
    .X(net5442));
 sg13g2_buf_8 fanout5443 (.A(net5446),
    .X(net5443));
 sg13g2_buf_8 fanout5444 (.A(net5446),
    .X(net5444));
 sg13g2_buf_8 fanout5445 (.A(net5446),
    .X(net5445));
 sg13g2_buf_8 fanout5446 (.A(_05592_),
    .X(net5446));
 sg13g2_buf_8 fanout5447 (.A(net5451),
    .X(net5447));
 sg13g2_buf_8 fanout5448 (.A(net5451),
    .X(net5448));
 sg13g2_buf_8 fanout5449 (.A(net5451),
    .X(net5449));
 sg13g2_buf_8 fanout5450 (.A(net5451),
    .X(net5450));
 sg13g2_buf_8 fanout5451 (.A(_05592_),
    .X(net5451));
 sg13g2_buf_8 fanout5452 (.A(_05283_),
    .X(net5452));
 sg13g2_buf_8 fanout5453 (.A(_05096_),
    .X(net5453));
 sg13g2_buf_8 fanout5454 (.A(_04848_),
    .X(net5454));
 sg13g2_buf_8 fanout5455 (.A(_04814_),
    .X(net5455));
 sg13g2_buf_8 fanout5456 (.A(_04809_),
    .X(net5456));
 sg13g2_buf_2 fanout5457 (.A(_04809_),
    .X(net5457));
 sg13g2_buf_8 fanout5458 (.A(net5459),
    .X(net5458));
 sg13g2_buf_8 fanout5459 (.A(_04804_),
    .X(net5459));
 sg13g2_buf_8 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_8 fanout5461 (.A(_04796_),
    .X(net5461));
 sg13g2_buf_8 fanout5462 (.A(_04773_),
    .X(net5462));
 sg13g2_buf_8 fanout5463 (.A(_04335_),
    .X(net5463));
 sg13g2_buf_1 fanout5464 (.A(_04335_),
    .X(net5464));
 sg13g2_buf_8 fanout5465 (.A(net5466),
    .X(net5465));
 sg13g2_buf_8 fanout5466 (.A(_04257_),
    .X(net5466));
 sg13g2_buf_8 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(net5471),
    .X(net5468));
 sg13g2_buf_8 fanout5469 (.A(net5471),
    .X(net5469));
 sg13g2_buf_8 fanout5470 (.A(net5471),
    .X(net5470));
 sg13g2_buf_8 fanout5471 (.A(_03464_),
    .X(net5471));
 sg13g2_buf_8 fanout5472 (.A(net5476),
    .X(net5472));
 sg13g2_buf_8 fanout5473 (.A(net5476),
    .X(net5473));
 sg13g2_buf_8 fanout5474 (.A(net5475),
    .X(net5474));
 sg13g2_buf_8 fanout5475 (.A(net5476),
    .X(net5475));
 sg13g2_buf_8 fanout5476 (.A(_03459_),
    .X(net5476));
 sg13g2_buf_8 fanout5477 (.A(net5481),
    .X(net5477));
 sg13g2_buf_8 fanout5478 (.A(net5481),
    .X(net5478));
 sg13g2_buf_8 fanout5479 (.A(net5480),
    .X(net5479));
 sg13g2_buf_8 fanout5480 (.A(net5481),
    .X(net5480));
 sg13g2_buf_8 fanout5481 (.A(_03447_),
    .X(net5481));
 sg13g2_buf_8 fanout5482 (.A(net5486),
    .X(net5482));
 sg13g2_buf_8 fanout5483 (.A(net5486),
    .X(net5483));
 sg13g2_buf_8 fanout5484 (.A(net5485),
    .X(net5484));
 sg13g2_buf_8 fanout5485 (.A(net5486),
    .X(net5485));
 sg13g2_buf_8 fanout5486 (.A(_02651_),
    .X(net5486));
 sg13g2_buf_8 fanout5487 (.A(net5491),
    .X(net5487));
 sg13g2_buf_8 fanout5488 (.A(net5491),
    .X(net5488));
 sg13g2_buf_8 fanout5489 (.A(net5490),
    .X(net5489));
 sg13g2_buf_8 fanout5490 (.A(net5491),
    .X(net5490));
 sg13g2_buf_8 fanout5491 (.A(_02642_),
    .X(net5491));
 sg13g2_buf_8 fanout5492 (.A(net5496),
    .X(net5492));
 sg13g2_buf_8 fanout5493 (.A(net5496),
    .X(net5493));
 sg13g2_buf_8 fanout5494 (.A(net5495),
    .X(net5494));
 sg13g2_buf_8 fanout5495 (.A(net5496),
    .X(net5495));
 sg13g2_buf_8 fanout5496 (.A(_02639_),
    .X(net5496));
 sg13g2_buf_8 fanout5497 (.A(net5501),
    .X(net5497));
 sg13g2_buf_8 fanout5498 (.A(net5501),
    .X(net5498));
 sg13g2_buf_8 fanout5499 (.A(net5500),
    .X(net5499));
 sg13g2_buf_8 fanout5500 (.A(net5501),
    .X(net5500));
 sg13g2_buf_8 fanout5501 (.A(_02638_),
    .X(net5501));
 sg13g2_buf_8 fanout5502 (.A(net5506),
    .X(net5502));
 sg13g2_buf_8 fanout5503 (.A(net5506),
    .X(net5503));
 sg13g2_buf_8 fanout5504 (.A(net5505),
    .X(net5504));
 sg13g2_buf_8 fanout5505 (.A(net5506),
    .X(net5505));
 sg13g2_buf_8 fanout5506 (.A(_02636_),
    .X(net5506));
 sg13g2_buf_8 fanout5507 (.A(net5511),
    .X(net5507));
 sg13g2_buf_8 fanout5508 (.A(net5511),
    .X(net5508));
 sg13g2_buf_8 fanout5509 (.A(net5510),
    .X(net5509));
 sg13g2_buf_8 fanout5510 (.A(net5511),
    .X(net5510));
 sg13g2_buf_8 fanout5511 (.A(_02634_),
    .X(net5511));
 sg13g2_buf_8 fanout5512 (.A(net5516),
    .X(net5512));
 sg13g2_buf_8 fanout5513 (.A(net5516),
    .X(net5513));
 sg13g2_buf_8 fanout5514 (.A(net5515),
    .X(net5514));
 sg13g2_buf_8 fanout5515 (.A(net5516),
    .X(net5515));
 sg13g2_buf_8 fanout5516 (.A(_02628_),
    .X(net5516));
 sg13g2_buf_8 fanout5517 (.A(_11408_),
    .X(net5517));
 sg13g2_buf_8 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_8 fanout5519 (.A(_10775_),
    .X(net5519));
 sg13g2_buf_8 fanout5520 (.A(net5521),
    .X(net5520));
 sg13g2_buf_2 fanout5521 (.A(net5522),
    .X(net5521));
 sg13g2_buf_1 fanout5522 (.A(net5524),
    .X(net5522));
 sg13g2_buf_8 fanout5523 (.A(net5524),
    .X(net5523));
 sg13g2_buf_1 fanout5524 (.A(_10168_),
    .X(net5524));
 sg13g2_buf_8 fanout5525 (.A(net5527),
    .X(net5525));
 sg13g2_buf_1 fanout5526 (.A(net5527),
    .X(net5526));
 sg13g2_buf_8 fanout5527 (.A(_09671_),
    .X(net5527));
 sg13g2_buf_8 fanout5528 (.A(_09594_),
    .X(net5528));
 sg13g2_buf_8 fanout5529 (.A(_09591_),
    .X(net5529));
 sg13g2_buf_8 fanout5530 (.A(_09424_),
    .X(net5530));
 sg13g2_buf_8 fanout5531 (.A(_09068_),
    .X(net5531));
 sg13g2_buf_1 fanout5532 (.A(_09068_),
    .X(net5532));
 sg13g2_buf_8 fanout5533 (.A(net5535),
    .X(net5533));
 sg13g2_buf_8 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_8 fanout5535 (.A(_09068_),
    .X(net5535));
 sg13g2_buf_8 fanout5536 (.A(net5541),
    .X(net5536));
 sg13g2_buf_2 fanout5537 (.A(net5541),
    .X(net5537));
 sg13g2_buf_8 fanout5538 (.A(net5539),
    .X(net5538));
 sg13g2_buf_8 fanout5539 (.A(net5540),
    .X(net5539));
 sg13g2_buf_8 fanout5540 (.A(net5541),
    .X(net5540));
 sg13g2_buf_8 fanout5541 (.A(_09014_),
    .X(net5541));
 sg13g2_buf_8 fanout5542 (.A(net5544),
    .X(net5542));
 sg13g2_buf_2 fanout5543 (.A(net5544),
    .X(net5543));
 sg13g2_buf_8 fanout5544 (.A(_09013_),
    .X(net5544));
 sg13g2_buf_8 fanout5545 (.A(net5548),
    .X(net5545));
 sg13g2_buf_1 fanout5546 (.A(net5548),
    .X(net5546));
 sg13g2_buf_8 fanout5547 (.A(net5548),
    .X(net5547));
 sg13g2_buf_8 fanout5548 (.A(net5549),
    .X(net5548));
 sg13g2_buf_8 fanout5549 (.A(_08991_),
    .X(net5549));
 sg13g2_buf_8 fanout5550 (.A(net5552),
    .X(net5550));
 sg13g2_buf_8 fanout5551 (.A(net5552),
    .X(net5551));
 sg13g2_buf_8 fanout5552 (.A(_08990_),
    .X(net5552));
 sg13g2_buf_8 fanout5553 (.A(net5555),
    .X(net5553));
 sg13g2_buf_8 fanout5554 (.A(_08990_),
    .X(net5554));
 sg13g2_buf_1 fanout5555 (.A(_08990_),
    .X(net5555));
 sg13g2_buf_8 fanout5556 (.A(net5557),
    .X(net5556));
 sg13g2_buf_2 fanout5557 (.A(net5558),
    .X(net5557));
 sg13g2_buf_8 fanout5558 (.A(_08904_),
    .X(net5558));
 sg13g2_buf_8 fanout5559 (.A(net5560),
    .X(net5559));
 sg13g2_buf_2 fanout5560 (.A(_08904_),
    .X(net5560));
 sg13g2_buf_8 fanout5561 (.A(net5562),
    .X(net5561));
 sg13g2_buf_8 fanout5562 (.A(_08819_),
    .X(net5562));
 sg13g2_buf_8 fanout5563 (.A(net5564),
    .X(net5563));
 sg13g2_buf_8 fanout5564 (.A(_08819_),
    .X(net5564));
 sg13g2_buf_8 fanout5565 (.A(_08814_),
    .X(net5565));
 sg13g2_buf_8 fanout5566 (.A(_08673_),
    .X(net5566));
 sg13g2_buf_1 fanout5567 (.A(_08673_),
    .X(net5567));
 sg13g2_buf_8 fanout5568 (.A(_08418_),
    .X(net5568));
 sg13g2_buf_8 fanout5569 (.A(net5570),
    .X(net5569));
 sg13g2_buf_8 fanout5570 (.A(net5572),
    .X(net5570));
 sg13g2_buf_8 fanout5571 (.A(net5572),
    .X(net5571));
 sg13g2_buf_8 fanout5572 (.A(net5579),
    .X(net5572));
 sg13g2_buf_8 fanout5573 (.A(net5575),
    .X(net5573));
 sg13g2_buf_1 fanout5574 (.A(net5575),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_8 fanout5576 (.A(net5579),
    .X(net5576));
 sg13g2_buf_8 fanout5577 (.A(net5578),
    .X(net5577));
 sg13g2_buf_8 fanout5578 (.A(net5579),
    .X(net5578));
 sg13g2_buf_8 fanout5579 (.A(_06559_),
    .X(net5579));
 sg13g2_buf_8 fanout5580 (.A(net5590),
    .X(net5580));
 sg13g2_buf_8 fanout5581 (.A(net5590),
    .X(net5581));
 sg13g2_buf_8 fanout5582 (.A(net5583),
    .X(net5582));
 sg13g2_buf_8 fanout5583 (.A(net5590),
    .X(net5583));
 sg13g2_buf_8 fanout5584 (.A(net5586),
    .X(net5584));
 sg13g2_buf_8 fanout5585 (.A(net5586),
    .X(net5585));
 sg13g2_buf_8 fanout5586 (.A(net5590),
    .X(net5586));
 sg13g2_buf_8 fanout5587 (.A(net5589),
    .X(net5587));
 sg13g2_buf_1 fanout5588 (.A(net5589),
    .X(net5588));
 sg13g2_buf_8 fanout5589 (.A(net5590),
    .X(net5589));
 sg13g2_buf_8 fanout5590 (.A(_06526_),
    .X(net5590));
 sg13g2_buf_8 fanout5591 (.A(net5601),
    .X(net5591));
 sg13g2_buf_8 fanout5592 (.A(net5601),
    .X(net5592));
 sg13g2_buf_8 fanout5593 (.A(net5594),
    .X(net5593));
 sg13g2_buf_8 fanout5594 (.A(net5601),
    .X(net5594));
 sg13g2_buf_8 fanout5595 (.A(net5597),
    .X(net5595));
 sg13g2_buf_8 fanout5596 (.A(net5597),
    .X(net5596));
 sg13g2_buf_8 fanout5597 (.A(net5601),
    .X(net5597));
 sg13g2_buf_8 fanout5598 (.A(net5600),
    .X(net5598));
 sg13g2_buf_1 fanout5599 (.A(net5600),
    .X(net5599));
 sg13g2_buf_8 fanout5600 (.A(net5601),
    .X(net5600));
 sg13g2_buf_8 fanout5601 (.A(_06427_),
    .X(net5601));
 sg13g2_buf_8 fanout5602 (.A(net5604),
    .X(net5602));
 sg13g2_buf_8 fanout5603 (.A(net5604),
    .X(net5603));
 sg13g2_buf_8 fanout5604 (.A(net5612),
    .X(net5604));
 sg13g2_buf_8 fanout5605 (.A(net5612),
    .X(net5605));
 sg13g2_buf_8 fanout5606 (.A(net5607),
    .X(net5606));
 sg13g2_buf_8 fanout5607 (.A(net5611),
    .X(net5607));
 sg13g2_buf_8 fanout5608 (.A(net5610),
    .X(net5608));
 sg13g2_buf_8 fanout5609 (.A(net5610),
    .X(net5609));
 sg13g2_buf_8 fanout5610 (.A(net5611),
    .X(net5610));
 sg13g2_buf_8 fanout5611 (.A(net5612),
    .X(net5611));
 sg13g2_buf_8 fanout5612 (.A(_06295_),
    .X(net5612));
 sg13g2_buf_8 fanout5613 (.A(net5617),
    .X(net5613));
 sg13g2_buf_8 fanout5614 (.A(net5617),
    .X(net5614));
 sg13g2_buf_8 fanout5615 (.A(net5617),
    .X(net5615));
 sg13g2_buf_8 fanout5616 (.A(net5617),
    .X(net5616));
 sg13g2_buf_8 fanout5617 (.A(_06262_),
    .X(net5617));
 sg13g2_buf_8 fanout5618 (.A(net5620),
    .X(net5618));
 sg13g2_buf_8 fanout5619 (.A(net5620),
    .X(net5619));
 sg13g2_buf_8 fanout5620 (.A(net5623),
    .X(net5620));
 sg13g2_buf_8 fanout5621 (.A(net5622),
    .X(net5621));
 sg13g2_buf_8 fanout5622 (.A(net5623),
    .X(net5622));
 sg13g2_buf_8 fanout5623 (.A(_06262_),
    .X(net5623));
 sg13g2_buf_8 fanout5624 (.A(net5625),
    .X(net5624));
 sg13g2_buf_8 fanout5625 (.A(net5628),
    .X(net5625));
 sg13g2_buf_8 fanout5626 (.A(net5628),
    .X(net5626));
 sg13g2_buf_8 fanout5627 (.A(net5628),
    .X(net5627));
 sg13g2_buf_8 fanout5628 (.A(_06162_),
    .X(net5628));
 sg13g2_buf_8 fanout5629 (.A(net5633),
    .X(net5629));
 sg13g2_buf_8 fanout5630 (.A(net5633),
    .X(net5630));
 sg13g2_buf_8 fanout5631 (.A(net5632),
    .X(net5631));
 sg13g2_buf_8 fanout5632 (.A(net5633),
    .X(net5632));
 sg13g2_buf_8 fanout5633 (.A(_06162_),
    .X(net5633));
 sg13g2_buf_8 fanout5634 (.A(net5637),
    .X(net5634));
 sg13g2_buf_1 fanout5635 (.A(net5637),
    .X(net5635));
 sg13g2_buf_8 fanout5636 (.A(net5637),
    .X(net5636));
 sg13g2_buf_8 fanout5637 (.A(_06129_),
    .X(net5637));
 sg13g2_buf_8 fanout5638 (.A(net5641),
    .X(net5638));
 sg13g2_buf_1 fanout5639 (.A(net5641),
    .X(net5639));
 sg13g2_buf_8 fanout5640 (.A(net5641),
    .X(net5640));
 sg13g2_buf_8 fanout5641 (.A(net5645),
    .X(net5641));
 sg13g2_buf_8 fanout5642 (.A(net5645),
    .X(net5642));
 sg13g2_buf_1 fanout5643 (.A(net5645),
    .X(net5643));
 sg13g2_buf_8 fanout5644 (.A(net5645),
    .X(net5644));
 sg13g2_buf_8 fanout5645 (.A(_06129_),
    .X(net5645));
 sg13g2_buf_8 fanout5646 (.A(net5649),
    .X(net5646));
 sg13g2_buf_8 fanout5647 (.A(net5649),
    .X(net5647));
 sg13g2_buf_8 fanout5648 (.A(net5649),
    .X(net5648));
 sg13g2_buf_8 fanout5649 (.A(_06062_),
    .X(net5649));
 sg13g2_buf_8 fanout5650 (.A(net5651),
    .X(net5650));
 sg13g2_buf_8 fanout5651 (.A(net5655),
    .X(net5651));
 sg13g2_buf_8 fanout5652 (.A(net5655),
    .X(net5652));
 sg13g2_buf_1 fanout5653 (.A(net5655),
    .X(net5653));
 sg13g2_buf_8 fanout5654 (.A(net5655),
    .X(net5654));
 sg13g2_buf_8 fanout5655 (.A(_06062_),
    .X(net5655));
 sg13g2_buf_8 fanout5656 (.A(net5660),
    .X(net5656));
 sg13g2_buf_8 fanout5657 (.A(net5660),
    .X(net5657));
 sg13g2_buf_8 fanout5658 (.A(net5660),
    .X(net5658));
 sg13g2_buf_1 fanout5659 (.A(net5660),
    .X(net5659));
 sg13g2_buf_8 fanout5660 (.A(_06029_),
    .X(net5660));
 sg13g2_buf_8 fanout5661 (.A(net5665),
    .X(net5661));
 sg13g2_buf_8 fanout5662 (.A(net5665),
    .X(net5662));
 sg13g2_buf_8 fanout5663 (.A(net5664),
    .X(net5663));
 sg13g2_buf_8 fanout5664 (.A(net5665),
    .X(net5664));
 sg13g2_buf_8 fanout5665 (.A(_06029_),
    .X(net5665));
 sg13g2_buf_8 fanout5666 (.A(net5669),
    .X(net5666));
 sg13g2_buf_8 fanout5667 (.A(net5669),
    .X(net5667));
 sg13g2_buf_8 fanout5668 (.A(net5669),
    .X(net5668));
 sg13g2_buf_8 fanout5669 (.A(_05996_),
    .X(net5669));
 sg13g2_buf_8 fanout5670 (.A(net5674),
    .X(net5670));
 sg13g2_buf_8 fanout5671 (.A(net5674),
    .X(net5671));
 sg13g2_buf_8 fanout5672 (.A(net5674),
    .X(net5672));
 sg13g2_buf_8 fanout5673 (.A(net5674),
    .X(net5673));
 sg13g2_buf_8 fanout5674 (.A(_05996_),
    .X(net5674));
 sg13g2_buf_8 fanout5675 (.A(net5676),
    .X(net5675));
 sg13g2_buf_8 fanout5676 (.A(net5679),
    .X(net5676));
 sg13g2_buf_8 fanout5677 (.A(net5679),
    .X(net5677));
 sg13g2_buf_8 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_8 fanout5679 (.A(_05963_),
    .X(net5679));
 sg13g2_buf_8 fanout5680 (.A(net5681),
    .X(net5680));
 sg13g2_buf_8 fanout5681 (.A(net5684),
    .X(net5681));
 sg13g2_buf_8 fanout5682 (.A(net5683),
    .X(net5682));
 sg13g2_buf_8 fanout5683 (.A(net5684),
    .X(net5683));
 sg13g2_buf_8 fanout5684 (.A(_05963_),
    .X(net5684));
 sg13g2_buf_8 fanout5685 (.A(net5686),
    .X(net5685));
 sg13g2_buf_8 fanout5686 (.A(net5689),
    .X(net5686));
 sg13g2_buf_8 fanout5687 (.A(net5689),
    .X(net5687));
 sg13g2_buf_8 fanout5688 (.A(net5689),
    .X(net5688));
 sg13g2_buf_8 fanout5689 (.A(_05930_),
    .X(net5689));
 sg13g2_buf_8 fanout5690 (.A(net5691),
    .X(net5690));
 sg13g2_buf_8 fanout5691 (.A(net5694),
    .X(net5691));
 sg13g2_buf_8 fanout5692 (.A(net5693),
    .X(net5692));
 sg13g2_buf_8 fanout5693 (.A(net5694),
    .X(net5693));
 sg13g2_buf_8 fanout5694 (.A(_05930_),
    .X(net5694));
 sg13g2_buf_8 fanout5695 (.A(net5699),
    .X(net5695));
 sg13g2_buf_8 fanout5696 (.A(net5699),
    .X(net5696));
 sg13g2_buf_8 fanout5697 (.A(net5699),
    .X(net5697));
 sg13g2_buf_8 fanout5698 (.A(net5699),
    .X(net5698));
 sg13g2_buf_8 fanout5699 (.A(_05862_),
    .X(net5699));
 sg13g2_buf_8 fanout5700 (.A(net5701),
    .X(net5700));
 sg13g2_buf_8 fanout5701 (.A(net5705),
    .X(net5701));
 sg13g2_buf_1 fanout5702 (.A(net5705),
    .X(net5702));
 sg13g2_buf_8 fanout5703 (.A(net5704),
    .X(net5703));
 sg13g2_buf_8 fanout5704 (.A(net5705),
    .X(net5704));
 sg13g2_buf_8 fanout5705 (.A(_05862_),
    .X(net5705));
 sg13g2_buf_8 fanout5706 (.A(net5707),
    .X(net5706));
 sg13g2_buf_8 fanout5707 (.A(net5710),
    .X(net5707));
 sg13g2_buf_8 fanout5708 (.A(net5710),
    .X(net5708));
 sg13g2_buf_8 fanout5709 (.A(net5710),
    .X(net5709));
 sg13g2_buf_8 fanout5710 (.A(_05828_),
    .X(net5710));
 sg13g2_buf_8 fanout5711 (.A(net5715),
    .X(net5711));
 sg13g2_buf_8 fanout5712 (.A(net5715),
    .X(net5712));
 sg13g2_buf_8 fanout5713 (.A(net5714),
    .X(net5713));
 sg13g2_buf_8 fanout5714 (.A(net5715),
    .X(net5714));
 sg13g2_buf_8 fanout5715 (.A(_05828_),
    .X(net5715));
 sg13g2_buf_8 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_8 fanout5717 (.A(net5726),
    .X(net5717));
 sg13g2_buf_8 fanout5718 (.A(net5726),
    .X(net5718));
 sg13g2_buf_1 fanout5719 (.A(net5726),
    .X(net5719));
 sg13g2_buf_8 fanout5720 (.A(net5721),
    .X(net5720));
 sg13g2_buf_8 fanout5721 (.A(net5725),
    .X(net5721));
 sg13g2_buf_8 fanout5722 (.A(net5724),
    .X(net5722));
 sg13g2_buf_1 fanout5723 (.A(net5724),
    .X(net5723));
 sg13g2_buf_8 fanout5724 (.A(net5725),
    .X(net5724));
 sg13g2_buf_8 fanout5725 (.A(net5726),
    .X(net5725));
 sg13g2_buf_8 fanout5726 (.A(_05795_),
    .X(net5726));
 sg13g2_buf_8 fanout5727 (.A(net5728),
    .X(net5727));
 sg13g2_buf_8 fanout5728 (.A(net5731),
    .X(net5728));
 sg13g2_buf_8 fanout5729 (.A(net5731),
    .X(net5729));
 sg13g2_buf_8 fanout5730 (.A(net5731),
    .X(net5730));
 sg13g2_buf_8 fanout5731 (.A(_05762_),
    .X(net5731));
 sg13g2_buf_8 fanout5732 (.A(net5736),
    .X(net5732));
 sg13g2_buf_8 fanout5733 (.A(net5736),
    .X(net5733));
 sg13g2_buf_8 fanout5734 (.A(net5735),
    .X(net5734));
 sg13g2_buf_8 fanout5735 (.A(net5736),
    .X(net5735));
 sg13g2_buf_8 fanout5736 (.A(_05762_),
    .X(net5736));
 sg13g2_buf_8 fanout5737 (.A(net5738),
    .X(net5737));
 sg13g2_buf_8 fanout5738 (.A(net5746),
    .X(net5738));
 sg13g2_buf_8 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_8 fanout5740 (.A(net5746),
    .X(net5740));
 sg13g2_buf_8 fanout5741 (.A(net5743),
    .X(net5741));
 sg13g2_buf_1 fanout5742 (.A(net5743),
    .X(net5742));
 sg13g2_buf_8 fanout5743 (.A(net5746),
    .X(net5743));
 sg13g2_buf_8 fanout5744 (.A(net5745),
    .X(net5744));
 sg13g2_buf_8 fanout5745 (.A(net5746),
    .X(net5745));
 sg13g2_buf_8 fanout5746 (.A(_05729_),
    .X(net5746));
 sg13g2_buf_8 fanout5747 (.A(net5748),
    .X(net5747));
 sg13g2_buf_8 fanout5748 (.A(net5751),
    .X(net5748));
 sg13g2_buf_8 fanout5749 (.A(net5751),
    .X(net5749));
 sg13g2_buf_8 fanout5750 (.A(net5751),
    .X(net5750));
 sg13g2_buf_8 fanout5751 (.A(_05661_),
    .X(net5751));
 sg13g2_buf_8 fanout5752 (.A(net5756),
    .X(net5752));
 sg13g2_buf_8 fanout5753 (.A(net5756),
    .X(net5753));
 sg13g2_buf_8 fanout5754 (.A(net5756),
    .X(net5754));
 sg13g2_buf_8 fanout5755 (.A(net5756),
    .X(net5755));
 sg13g2_buf_8 fanout5756 (.A(_05661_),
    .X(net5756));
 sg13g2_buf_8 fanout5757 (.A(net5758),
    .X(net5757));
 sg13g2_buf_8 fanout5758 (.A(_04854_),
    .X(net5758));
 sg13g2_buf_8 fanout5759 (.A(net5760),
    .X(net5759));
 sg13g2_buf_8 fanout5760 (.A(_04853_),
    .X(net5760));
 sg13g2_buf_8 fanout5761 (.A(net5762),
    .X(net5761));
 sg13g2_buf_8 fanout5762 (.A(_04843_),
    .X(net5762));
 sg13g2_buf_8 fanout5763 (.A(net5764),
    .X(net5763));
 sg13g2_buf_8 fanout5764 (.A(net5765),
    .X(net5764));
 sg13g2_buf_8 fanout5765 (.A(_04842_),
    .X(net5765));
 sg13g2_buf_8 fanout5766 (.A(net5768),
    .X(net5766));
 sg13g2_buf_1 fanout5767 (.A(net5768),
    .X(net5767));
 sg13g2_buf_2 fanout5768 (.A(_04795_),
    .X(net5768));
 sg13g2_buf_8 fanout5769 (.A(_04786_),
    .X(net5769));
 sg13g2_buf_8 fanout5770 (.A(net5771),
    .X(net5770));
 sg13g2_buf_8 fanout5771 (.A(_04553_),
    .X(net5771));
 sg13g2_buf_8 fanout5772 (.A(net5773),
    .X(net5772));
 sg13g2_buf_8 fanout5773 (.A(net5774),
    .X(net5773));
 sg13g2_buf_8 fanout5774 (.A(_04552_),
    .X(net5774));
 sg13g2_buf_8 fanout5775 (.A(_04225_),
    .X(net5775));
 sg13g2_buf_8 fanout5776 (.A(net5778),
    .X(net5776));
 sg13g2_buf_1 fanout5777 (.A(net5778),
    .X(net5777));
 sg13g2_buf_8 fanout5778 (.A(_04224_),
    .X(net5778));
 sg13g2_buf_8 fanout5779 (.A(net5780),
    .X(net5779));
 sg13g2_buf_8 fanout5780 (.A(_04224_),
    .X(net5780));
 sg13g2_buf_8 fanout5781 (.A(net5785),
    .X(net5781));
 sg13g2_buf_8 fanout5782 (.A(net5785),
    .X(net5782));
 sg13g2_buf_8 fanout5783 (.A(net5784),
    .X(net5783));
 sg13g2_buf_8 fanout5784 (.A(net5785),
    .X(net5784));
 sg13g2_buf_8 fanout5785 (.A(_03472_),
    .X(net5785));
 sg13g2_buf_8 fanout5786 (.A(net5790),
    .X(net5786));
 sg13g2_buf_8 fanout5787 (.A(net5790),
    .X(net5787));
 sg13g2_buf_8 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_8 fanout5789 (.A(net5790),
    .X(net5789));
 sg13g2_buf_8 fanout5790 (.A(_03471_),
    .X(net5790));
 sg13g2_buf_8 fanout5791 (.A(net5792),
    .X(net5791));
 sg13g2_buf_8 fanout5792 (.A(net5795),
    .X(net5792));
 sg13g2_buf_8 fanout5793 (.A(net5795),
    .X(net5793));
 sg13g2_buf_8 fanout5794 (.A(net5795),
    .X(net5794));
 sg13g2_buf_8 fanout5795 (.A(_03467_),
    .X(net5795));
 sg13g2_buf_8 fanout5796 (.A(net5800),
    .X(net5796));
 sg13g2_buf_8 fanout5797 (.A(net5800),
    .X(net5797));
 sg13g2_buf_8 fanout5798 (.A(net5799),
    .X(net5798));
 sg13g2_buf_8 fanout5799 (.A(net5800),
    .X(net5799));
 sg13g2_buf_8 fanout5800 (.A(_03466_),
    .X(net5800));
 sg13g2_buf_8 fanout5801 (.A(net5805),
    .X(net5801));
 sg13g2_buf_8 fanout5802 (.A(net5805),
    .X(net5802));
 sg13g2_buf_8 fanout5803 (.A(net5804),
    .X(net5803));
 sg13g2_buf_8 fanout5804 (.A(net5805),
    .X(net5804));
 sg13g2_buf_8 fanout5805 (.A(_03463_),
    .X(net5805));
 sg13g2_buf_8 fanout5806 (.A(net5810),
    .X(net5806));
 sg13g2_buf_8 fanout5807 (.A(net5810),
    .X(net5807));
 sg13g2_buf_8 fanout5808 (.A(net5809),
    .X(net5808));
 sg13g2_buf_8 fanout5809 (.A(net5810),
    .X(net5809));
 sg13g2_buf_8 fanout5810 (.A(_03460_),
    .X(net5810));
 sg13g2_buf_8 fanout5811 (.A(net5815),
    .X(net5811));
 sg13g2_buf_8 fanout5812 (.A(net5815),
    .X(net5812));
 sg13g2_buf_8 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_8 fanout5814 (.A(net5815),
    .X(net5814));
 sg13g2_buf_8 fanout5815 (.A(_03458_),
    .X(net5815));
 sg13g2_buf_8 fanout5816 (.A(net5820),
    .X(net5816));
 sg13g2_buf_8 fanout5817 (.A(net5820),
    .X(net5817));
 sg13g2_buf_8 fanout5818 (.A(net5819),
    .X(net5818));
 sg13g2_buf_8 fanout5819 (.A(net5820),
    .X(net5819));
 sg13g2_buf_8 fanout5820 (.A(_03457_),
    .X(net5820));
 sg13g2_buf_8 fanout5821 (.A(net5825),
    .X(net5821));
 sg13g2_buf_8 fanout5822 (.A(net5825),
    .X(net5822));
 sg13g2_buf_8 fanout5823 (.A(net5824),
    .X(net5823));
 sg13g2_buf_8 fanout5824 (.A(net5825),
    .X(net5824));
 sg13g2_buf_8 fanout5825 (.A(_03455_),
    .X(net5825));
 sg13g2_buf_8 fanout5826 (.A(net5830),
    .X(net5826));
 sg13g2_buf_8 fanout5827 (.A(net5830),
    .X(net5827));
 sg13g2_buf_8 fanout5828 (.A(net5829),
    .X(net5828));
 sg13g2_buf_8 fanout5829 (.A(net5830),
    .X(net5829));
 sg13g2_buf_8 fanout5830 (.A(_03454_),
    .X(net5830));
 sg13g2_buf_8 fanout5831 (.A(net5835),
    .X(net5831));
 sg13g2_buf_8 fanout5832 (.A(net5835),
    .X(net5832));
 sg13g2_buf_8 fanout5833 (.A(net5835),
    .X(net5833));
 sg13g2_buf_8 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_8 fanout5835 (.A(_03453_),
    .X(net5835));
 sg13g2_buf_8 fanout5836 (.A(net5840),
    .X(net5836));
 sg13g2_buf_8 fanout5837 (.A(net5840),
    .X(net5837));
 sg13g2_buf_8 fanout5838 (.A(net5839),
    .X(net5838));
 sg13g2_buf_8 fanout5839 (.A(net5840),
    .X(net5839));
 sg13g2_buf_8 fanout5840 (.A(_03452_),
    .X(net5840));
 sg13g2_buf_8 fanout5841 (.A(net5845),
    .X(net5841));
 sg13g2_buf_8 fanout5842 (.A(net5845),
    .X(net5842));
 sg13g2_buf_8 fanout5843 (.A(net5844),
    .X(net5843));
 sg13g2_buf_8 fanout5844 (.A(net5845),
    .X(net5844));
 sg13g2_buf_8 fanout5845 (.A(_03451_),
    .X(net5845));
 sg13g2_buf_8 fanout5846 (.A(net5850),
    .X(net5846));
 sg13g2_buf_8 fanout5847 (.A(net5850),
    .X(net5847));
 sg13g2_buf_8 fanout5848 (.A(net5849),
    .X(net5848));
 sg13g2_buf_8 fanout5849 (.A(net5850),
    .X(net5849));
 sg13g2_buf_8 fanout5850 (.A(_03449_),
    .X(net5850));
 sg13g2_buf_8 fanout5851 (.A(net5855),
    .X(net5851));
 sg13g2_buf_8 fanout5852 (.A(net5855),
    .X(net5852));
 sg13g2_buf_8 fanout5853 (.A(net5854),
    .X(net5853));
 sg13g2_buf_8 fanout5854 (.A(net5855),
    .X(net5854));
 sg13g2_buf_8 fanout5855 (.A(_03445_),
    .X(net5855));
 sg13g2_buf_8 fanout5856 (.A(net5860),
    .X(net5856));
 sg13g2_buf_8 fanout5857 (.A(net5860),
    .X(net5857));
 sg13g2_buf_8 fanout5858 (.A(net5859),
    .X(net5858));
 sg13g2_buf_8 fanout5859 (.A(net5860),
    .X(net5859));
 sg13g2_buf_8 fanout5860 (.A(_03442_),
    .X(net5860));
 sg13g2_buf_8 fanout5861 (.A(net5865),
    .X(net5861));
 sg13g2_buf_8 fanout5862 (.A(net5865),
    .X(net5862));
 sg13g2_buf_8 fanout5863 (.A(net5864),
    .X(net5863));
 sg13g2_buf_8 fanout5864 (.A(net5865),
    .X(net5864));
 sg13g2_buf_8 fanout5865 (.A(_03441_),
    .X(net5865));
 sg13g2_buf_8 fanout5866 (.A(net5870),
    .X(net5866));
 sg13g2_buf_8 fanout5867 (.A(net5870),
    .X(net5867));
 sg13g2_buf_8 fanout5868 (.A(net5869),
    .X(net5868));
 sg13g2_buf_8 fanout5869 (.A(net5870),
    .X(net5869));
 sg13g2_buf_8 fanout5870 (.A(_03440_),
    .X(net5870));
 sg13g2_buf_8 fanout5871 (.A(net5875),
    .X(net5871));
 sg13g2_buf_8 fanout5872 (.A(net5875),
    .X(net5872));
 sg13g2_buf_8 fanout5873 (.A(net5874),
    .X(net5873));
 sg13g2_buf_8 fanout5874 (.A(net5875),
    .X(net5874));
 sg13g2_buf_8 fanout5875 (.A(_03433_),
    .X(net5875));
 sg13g2_buf_8 fanout5876 (.A(net5880),
    .X(net5876));
 sg13g2_buf_8 fanout5877 (.A(net5880),
    .X(net5877));
 sg13g2_buf_8 fanout5878 (.A(net5879),
    .X(net5878));
 sg13g2_buf_8 fanout5879 (.A(net5880),
    .X(net5879));
 sg13g2_buf_8 fanout5880 (.A(_02652_),
    .X(net5880));
 sg13g2_buf_8 fanout5881 (.A(net5885),
    .X(net5881));
 sg13g2_buf_8 fanout5882 (.A(net5885),
    .X(net5882));
 sg13g2_buf_8 fanout5883 (.A(net5884),
    .X(net5883));
 sg13g2_buf_8 fanout5884 (.A(net5885),
    .X(net5884));
 sg13g2_buf_8 fanout5885 (.A(_02650_),
    .X(net5885));
 sg13g2_buf_8 fanout5886 (.A(net5890),
    .X(net5886));
 sg13g2_buf_8 fanout5887 (.A(net5890),
    .X(net5887));
 sg13g2_buf_8 fanout5888 (.A(net5889),
    .X(net5888));
 sg13g2_buf_8 fanout5889 (.A(net5890),
    .X(net5889));
 sg13g2_buf_8 fanout5890 (.A(_02649_),
    .X(net5890));
 sg13g2_buf_8 fanout5891 (.A(net5895),
    .X(net5891));
 sg13g2_buf_8 fanout5892 (.A(net5895),
    .X(net5892));
 sg13g2_buf_8 fanout5893 (.A(net5894),
    .X(net5893));
 sg13g2_buf_8 fanout5894 (.A(net5895),
    .X(net5894));
 sg13g2_buf_8 fanout5895 (.A(_02648_),
    .X(net5895));
 sg13g2_buf_8 fanout5896 (.A(net5900),
    .X(net5896));
 sg13g2_buf_8 fanout5897 (.A(net5900),
    .X(net5897));
 sg13g2_buf_8 fanout5898 (.A(net5899),
    .X(net5898));
 sg13g2_buf_8 fanout5899 (.A(net5900),
    .X(net5899));
 sg13g2_buf_8 fanout5900 (.A(_02647_),
    .X(net5900));
 sg13g2_buf_8 fanout5901 (.A(net5905),
    .X(net5901));
 sg13g2_buf_8 fanout5902 (.A(net5905),
    .X(net5902));
 sg13g2_buf_8 fanout5903 (.A(net5904),
    .X(net5903));
 sg13g2_buf_8 fanout5904 (.A(net5905),
    .X(net5904));
 sg13g2_buf_8 fanout5905 (.A(_02646_),
    .X(net5905));
 sg13g2_buf_8 fanout5906 (.A(net5910),
    .X(net5906));
 sg13g2_buf_8 fanout5907 (.A(net5910),
    .X(net5907));
 sg13g2_buf_8 fanout5908 (.A(net5909),
    .X(net5908));
 sg13g2_buf_8 fanout5909 (.A(net5910),
    .X(net5909));
 sg13g2_buf_8 fanout5910 (.A(_02645_),
    .X(net5910));
 sg13g2_buf_8 fanout5911 (.A(net5915),
    .X(net5911));
 sg13g2_buf_8 fanout5912 (.A(net5915),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(net5914),
    .X(net5913));
 sg13g2_buf_8 fanout5914 (.A(net5915),
    .X(net5914));
 sg13g2_buf_8 fanout5915 (.A(_02644_),
    .X(net5915));
 sg13g2_buf_8 fanout5916 (.A(net5920),
    .X(net5916));
 sg13g2_buf_8 fanout5917 (.A(net5920),
    .X(net5917));
 sg13g2_buf_8 fanout5918 (.A(net5919),
    .X(net5918));
 sg13g2_buf_8 fanout5919 (.A(net5920),
    .X(net5919));
 sg13g2_buf_8 fanout5920 (.A(_02643_),
    .X(net5920));
 sg13g2_buf_8 fanout5921 (.A(net5922),
    .X(net5921));
 sg13g2_buf_2 fanout5922 (.A(net5926),
    .X(net5922));
 sg13g2_buf_8 fanout5923 (.A(net5924),
    .X(net5923));
 sg13g2_buf_8 fanout5924 (.A(net5926),
    .X(net5924));
 sg13g2_buf_8 fanout5925 (.A(net5926),
    .X(net5925));
 sg13g2_buf_8 fanout5926 (.A(_02641_),
    .X(net5926));
 sg13g2_buf_8 fanout5927 (.A(net5931),
    .X(net5927));
 sg13g2_buf_8 fanout5928 (.A(net5931),
    .X(net5928));
 sg13g2_buf_8 fanout5929 (.A(net5930),
    .X(net5929));
 sg13g2_buf_8 fanout5930 (.A(net5931),
    .X(net5930));
 sg13g2_buf_8 fanout5931 (.A(_02637_),
    .X(net5931));
 sg13g2_buf_8 fanout5932 (.A(net5936),
    .X(net5932));
 sg13g2_buf_8 fanout5933 (.A(net5936),
    .X(net5933));
 sg13g2_buf_8 fanout5934 (.A(net5935),
    .X(net5934));
 sg13g2_buf_8 fanout5935 (.A(net5936),
    .X(net5935));
 sg13g2_buf_8 fanout5936 (.A(_02633_),
    .X(net5936));
 sg13g2_buf_8 fanout5937 (.A(net5941),
    .X(net5937));
 sg13g2_buf_8 fanout5938 (.A(net5941),
    .X(net5938));
 sg13g2_buf_8 fanout5939 (.A(net5940),
    .X(net5939));
 sg13g2_buf_8 fanout5940 (.A(net5941),
    .X(net5940));
 sg13g2_buf_8 fanout5941 (.A(_02631_),
    .X(net5941));
 sg13g2_buf_8 fanout5942 (.A(net5946),
    .X(net5942));
 sg13g2_buf_8 fanout5943 (.A(net5946),
    .X(net5943));
 sg13g2_buf_8 fanout5944 (.A(net5945),
    .X(net5944));
 sg13g2_buf_8 fanout5945 (.A(net5946),
    .X(net5945));
 sg13g2_buf_8 fanout5946 (.A(_02630_),
    .X(net5946));
 sg13g2_buf_8 fanout5947 (.A(net5951),
    .X(net5947));
 sg13g2_buf_8 fanout5948 (.A(net5951),
    .X(net5948));
 sg13g2_buf_8 fanout5949 (.A(net5950),
    .X(net5949));
 sg13g2_buf_8 fanout5950 (.A(net5951),
    .X(net5950));
 sg13g2_buf_8 fanout5951 (.A(_02629_),
    .X(net5951));
 sg13g2_buf_8 fanout5952 (.A(net5956),
    .X(net5952));
 sg13g2_buf_8 fanout5953 (.A(net5956),
    .X(net5953));
 sg13g2_buf_8 fanout5954 (.A(net5955),
    .X(net5954));
 sg13g2_buf_8 fanout5955 (.A(net5956),
    .X(net5955));
 sg13g2_buf_8 fanout5956 (.A(_02626_),
    .X(net5956));
 sg13g2_buf_8 fanout5957 (.A(net5961),
    .X(net5957));
 sg13g2_buf_8 fanout5958 (.A(net5961),
    .X(net5958));
 sg13g2_buf_8 fanout5959 (.A(net5960),
    .X(net5959));
 sg13g2_buf_8 fanout5960 (.A(net5961),
    .X(net5960));
 sg13g2_buf_8 fanout5961 (.A(_02625_),
    .X(net5961));
 sg13g2_buf_8 fanout5962 (.A(net5966),
    .X(net5962));
 sg13g2_buf_8 fanout5963 (.A(net5966),
    .X(net5963));
 sg13g2_buf_8 fanout5964 (.A(net5966),
    .X(net5964));
 sg13g2_buf_8 fanout5965 (.A(net5966),
    .X(net5965));
 sg13g2_buf_8 fanout5966 (.A(_02624_),
    .X(net5966));
 sg13g2_buf_8 fanout5967 (.A(net5971),
    .X(net5967));
 sg13g2_buf_8 fanout5968 (.A(net5971),
    .X(net5968));
 sg13g2_buf_8 fanout5969 (.A(net5970),
    .X(net5969));
 sg13g2_buf_8 fanout5970 (.A(net5971),
    .X(net5970));
 sg13g2_buf_8 fanout5971 (.A(_02623_),
    .X(net5971));
 sg13g2_buf_8 fanout5972 (.A(net5976),
    .X(net5972));
 sg13g2_buf_8 fanout5973 (.A(net5976),
    .X(net5973));
 sg13g2_buf_8 fanout5974 (.A(net5975),
    .X(net5974));
 sg13g2_buf_8 fanout5975 (.A(net5976),
    .X(net5975));
 sg13g2_buf_8 fanout5976 (.A(_02622_),
    .X(net5976));
 sg13g2_buf_8 fanout5977 (.A(net5981),
    .X(net5977));
 sg13g2_buf_8 fanout5978 (.A(net5981),
    .X(net5978));
 sg13g2_buf_8 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_8 fanout5980 (.A(net5981),
    .X(net5980));
 sg13g2_buf_8 fanout5981 (.A(_02620_),
    .X(net5981));
 sg13g2_buf_8 fanout5982 (.A(net5986),
    .X(net5982));
 sg13g2_buf_8 fanout5983 (.A(net5986),
    .X(net5983));
 sg13g2_buf_8 fanout5984 (.A(net5985),
    .X(net5984));
 sg13g2_buf_8 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_8 fanout5986 (.A(_02617_),
    .X(net5986));
 sg13g2_buf_8 fanout5987 (.A(net5991),
    .X(net5987));
 sg13g2_buf_8 fanout5988 (.A(net5991),
    .X(net5988));
 sg13g2_buf_8 fanout5989 (.A(net5990),
    .X(net5989));
 sg13g2_buf_8 fanout5990 (.A(net5991),
    .X(net5990));
 sg13g2_buf_8 fanout5991 (.A(_02614_),
    .X(net5991));
 sg13g2_buf_8 fanout5992 (.A(net5996),
    .X(net5992));
 sg13g2_buf_8 fanout5993 (.A(net5996),
    .X(net5993));
 sg13g2_buf_8 fanout5994 (.A(net5995),
    .X(net5994));
 sg13g2_buf_8 fanout5995 (.A(net5996),
    .X(net5995));
 sg13g2_buf_8 fanout5996 (.A(_02612_),
    .X(net5996));
 sg13g2_buf_8 fanout5997 (.A(_11432_),
    .X(net5997));
 sg13g2_buf_8 fanout5998 (.A(_11411_),
    .X(net5998));
 sg13g2_buf_8 fanout5999 (.A(_11411_),
    .X(net5999));
 sg13g2_buf_8 fanout6000 (.A(net6001),
    .X(net6000));
 sg13g2_buf_8 fanout6001 (.A(net6002),
    .X(net6001));
 sg13g2_buf_8 fanout6002 (.A(_11410_),
    .X(net6002));
 sg13g2_buf_8 fanout6003 (.A(_11291_),
    .X(net6003));
 sg13g2_buf_8 fanout6004 (.A(net6006),
    .X(net6004));
 sg13g2_buf_1 fanout6005 (.A(net6006),
    .X(net6005));
 sg13g2_buf_2 fanout6006 (.A(_11024_),
    .X(net6006));
 sg13g2_buf_8 fanout6007 (.A(net6008),
    .X(net6007));
 sg13g2_buf_8 fanout6008 (.A(_11024_),
    .X(net6008));
 sg13g2_buf_8 fanout6009 (.A(net6010),
    .X(net6009));
 sg13g2_buf_8 fanout6010 (.A(_10850_),
    .X(net6010));
 sg13g2_buf_8 fanout6011 (.A(_10849_),
    .X(net6011));
 sg13g2_buf_8 fanout6012 (.A(_09962_),
    .X(net6012));
 sg13g2_buf_8 fanout6013 (.A(_09957_),
    .X(net6013));
 sg13g2_buf_2 fanout6014 (.A(_09957_),
    .X(net6014));
 sg13g2_buf_8 fanout6015 (.A(_09955_),
    .X(net6015));
 sg13g2_buf_8 fanout6016 (.A(_09921_),
    .X(net6016));
 sg13g2_buf_8 fanout6017 (.A(net6019),
    .X(net6017));
 sg13g2_buf_1 fanout6018 (.A(net6019),
    .X(net6018));
 sg13g2_buf_8 fanout6019 (.A(net6020),
    .X(net6019));
 sg13g2_buf_8 fanout6020 (.A(_09892_),
    .X(net6020));
 sg13g2_buf_8 fanout6021 (.A(net6023),
    .X(net6021));
 sg13g2_buf_1 fanout6022 (.A(net6023),
    .X(net6022));
 sg13g2_buf_8 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_8 fanout6024 (.A(_09593_),
    .X(net6024));
 sg13g2_buf_8 fanout6025 (.A(net6028),
    .X(net6025));
 sg13g2_buf_8 fanout6026 (.A(net6028),
    .X(net6026));
 sg13g2_buf_8 fanout6027 (.A(net6028),
    .X(net6027));
 sg13g2_buf_8 fanout6028 (.A(_09592_),
    .X(net6028));
 sg13g2_buf_8 fanout6029 (.A(net6031),
    .X(net6029));
 sg13g2_buf_8 fanout6030 (.A(net6031),
    .X(net6030));
 sg13g2_buf_8 fanout6031 (.A(_09512_),
    .X(net6031));
 sg13g2_buf_8 fanout6032 (.A(net6033),
    .X(net6032));
 sg13g2_buf_8 fanout6033 (.A(_09511_),
    .X(net6033));
 sg13g2_buf_8 fanout6034 (.A(net6038),
    .X(net6034));
 sg13g2_buf_8 fanout6035 (.A(net6038),
    .X(net6035));
 sg13g2_buf_8 fanout6036 (.A(net6038),
    .X(net6036));
 sg13g2_buf_1 fanout6037 (.A(net6038),
    .X(net6037));
 sg13g2_buf_8 fanout6038 (.A(_09509_),
    .X(net6038));
 sg13g2_buf_8 fanout6039 (.A(net6044),
    .X(net6039));
 sg13g2_buf_1 fanout6040 (.A(net6044),
    .X(net6040));
 sg13g2_buf_8 fanout6041 (.A(net6044),
    .X(net6041));
 sg13g2_buf_8 fanout6042 (.A(net6044),
    .X(net6042));
 sg13g2_buf_8 fanout6043 (.A(net6044),
    .X(net6043));
 sg13g2_buf_8 fanout6044 (.A(_09509_),
    .X(net6044));
 sg13g2_buf_8 fanout6045 (.A(_09066_),
    .X(net6045));
 sg13g2_buf_8 fanout6046 (.A(_08989_),
    .X(net6046));
 sg13g2_buf_8 fanout6047 (.A(net6049),
    .X(net6047));
 sg13g2_buf_8 fanout6048 (.A(net6049),
    .X(net6048));
 sg13g2_buf_8 fanout6049 (.A(_08905_),
    .X(net6049));
 sg13g2_buf_8 fanout6050 (.A(net6051),
    .X(net6050));
 sg13g2_buf_8 fanout6051 (.A(_08820_),
    .X(net6051));
 sg13g2_buf_8 fanout6052 (.A(net6054),
    .X(net6052));
 sg13g2_buf_1 fanout6053 (.A(net6054),
    .X(net6053));
 sg13g2_buf_8 fanout6054 (.A(net6055),
    .X(net6054));
 sg13g2_buf_8 fanout6055 (.A(_08820_),
    .X(net6055));
 sg13g2_buf_8 fanout6056 (.A(net6061),
    .X(net6056));
 sg13g2_buf_2 fanout6057 (.A(net6059),
    .X(net6057));
 sg13g2_buf_1 fanout6058 (.A(net6059),
    .X(net6058));
 sg13g2_buf_1 fanout6059 (.A(net6060),
    .X(net6059));
 sg13g2_buf_2 fanout6060 (.A(net6061),
    .X(net6060));
 sg13g2_buf_8 fanout6061 (.A(_08791_),
    .X(net6061));
 sg13g2_buf_2 fanout6062 (.A(net6064),
    .X(net6062));
 sg13g2_buf_1 fanout6063 (.A(net6064),
    .X(net6063));
 sg13g2_buf_8 fanout6064 (.A(_08670_),
    .X(net6064));
 sg13g2_buf_8 fanout6065 (.A(net6066),
    .X(net6065));
 sg13g2_buf_8 fanout6066 (.A(_08669_),
    .X(net6066));
 sg13g2_buf_8 fanout6067 (.A(_08669_),
    .X(net6067));
 sg13g2_buf_1 fanout6068 (.A(_08669_),
    .X(net6068));
 sg13g2_buf_8 fanout6069 (.A(_07724_),
    .X(net6069));
 sg13g2_buf_8 fanout6070 (.A(_05895_),
    .X(net6070));
 sg13g2_buf_1 fanout6071 (.A(_05895_),
    .X(net6071));
 sg13g2_buf_8 fanout6072 (.A(net6073),
    .X(net6072));
 sg13g2_buf_8 fanout6073 (.A(_04475_),
    .X(net6073));
 sg13g2_buf_8 fanout6074 (.A(_04475_),
    .X(net6074));
 sg13g2_buf_2 fanout6075 (.A(_04475_),
    .X(net6075));
 sg13g2_buf_8 fanout6076 (.A(net6077),
    .X(net6076));
 sg13g2_buf_8 fanout6077 (.A(_03429_),
    .X(net6077));
 sg13g2_buf_8 fanout6078 (.A(net6080),
    .X(net6078));
 sg13g2_buf_8 fanout6079 (.A(net6080),
    .X(net6079));
 sg13g2_buf_8 fanout6080 (.A(_03429_),
    .X(net6080));
 sg13g2_buf_8 fanout6081 (.A(net6085),
    .X(net6081));
 sg13g2_buf_8 fanout6082 (.A(net6085),
    .X(net6082));
 sg13g2_buf_8 fanout6083 (.A(net6084),
    .X(net6083));
 sg13g2_buf_8 fanout6084 (.A(net6085),
    .X(net6084));
 sg13g2_buf_8 fanout6085 (.A(_02640_),
    .X(net6085));
 sg13g2_buf_8 fanout6086 (.A(_11459_),
    .X(net6086));
 sg13g2_buf_8 fanout6087 (.A(net6088),
    .X(net6087));
 sg13g2_buf_8 fanout6088 (.A(_11455_),
    .X(net6088));
 sg13g2_buf_8 fanout6089 (.A(_10758_),
    .X(net6089));
 sg13g2_buf_8 fanout6090 (.A(_09988_),
    .X(net6090));
 sg13g2_buf_8 fanout6091 (.A(_09972_),
    .X(net6091));
 sg13g2_buf_8 fanout6092 (.A(_09951_),
    .X(net6092));
 sg13g2_buf_2 fanout6093 (.A(_09951_),
    .X(net6093));
 sg13g2_buf_8 fanout6094 (.A(_09950_),
    .X(net6094));
 sg13g2_buf_1 fanout6095 (.A(_09950_),
    .X(net6095));
 sg13g2_buf_2 fanout6096 (.A(_09504_),
    .X(net6096));
 sg13g2_buf_8 fanout6097 (.A(_09248_),
    .X(net6097));
 sg13g2_buf_8 fanout6098 (.A(_09244_),
    .X(net6098));
 sg13g2_buf_8 fanout6099 (.A(net6102),
    .X(net6099));
 sg13g2_buf_8 fanout6100 (.A(net6102),
    .X(net6100));
 sg13g2_buf_1 fanout6101 (.A(net6102),
    .X(net6101));
 sg13g2_buf_8 fanout6102 (.A(_09136_),
    .X(net6102));
 sg13g2_buf_8 fanout6103 (.A(_09065_),
    .X(net6103));
 sg13g2_buf_1 fanout6104 (.A(_09065_),
    .X(net6104));
 sg13g2_buf_8 fanout6105 (.A(_09049_),
    .X(net6105));
 sg13g2_buf_8 fanout6106 (.A(_08984_),
    .X(net6106));
 sg13g2_buf_8 fanout6107 (.A(_08983_),
    .X(net6107));
 sg13g2_buf_8 fanout6108 (.A(net6109),
    .X(net6108));
 sg13g2_buf_8 fanout6109 (.A(_08790_),
    .X(net6109));
 sg13g2_buf_8 fanout6110 (.A(_08423_),
    .X(net6110));
 sg13g2_buf_8 fanout6111 (.A(net6112),
    .X(net6111));
 sg13g2_buf_8 fanout6112 (.A(_08211_),
    .X(net6112));
 sg13g2_buf_8 fanout6113 (.A(net6115),
    .X(net6113));
 sg13g2_buf_1 fanout6114 (.A(net6115),
    .X(net6114));
 sg13g2_buf_8 fanout6115 (.A(_08210_),
    .X(net6115));
 sg13g2_buf_8 fanout6116 (.A(net6117),
    .X(net6116));
 sg13g2_buf_8 fanout6117 (.A(net6118),
    .X(net6117));
 sg13g2_buf_2 fanout6118 (.A(net6119),
    .X(net6118));
 sg13g2_buf_1 fanout6119 (.A(_08210_),
    .X(net6119));
 sg13g2_buf_8 fanout6120 (.A(net6126),
    .X(net6120));
 sg13g2_buf_8 fanout6121 (.A(net6122),
    .X(net6121));
 sg13g2_buf_8 fanout6122 (.A(net6126),
    .X(net6122));
 sg13g2_buf_8 fanout6123 (.A(net6125),
    .X(net6123));
 sg13g2_buf_8 fanout6124 (.A(net6125),
    .X(net6124));
 sg13g2_buf_8 fanout6125 (.A(net6126),
    .X(net6125));
 sg13g2_buf_8 fanout6126 (.A(_08208_),
    .X(net6126));
 sg13g2_buf_8 fanout6127 (.A(net6128),
    .X(net6127));
 sg13g2_buf_8 fanout6128 (.A(net6129),
    .X(net6128));
 sg13g2_buf_8 fanout6129 (.A(_08207_),
    .X(net6129));
 sg13g2_buf_8 fanout6130 (.A(net6134),
    .X(net6130));
 sg13g2_buf_8 fanout6131 (.A(net6132),
    .X(net6131));
 sg13g2_buf_1 fanout6132 (.A(net6133),
    .X(net6132));
 sg13g2_buf_1 fanout6133 (.A(net6134),
    .X(net6133));
 sg13g2_buf_2 fanout6134 (.A(_08207_),
    .X(net6134));
 sg13g2_buf_8 fanout6135 (.A(_08206_),
    .X(net6135));
 sg13g2_buf_8 fanout6136 (.A(_08206_),
    .X(net6136));
 sg13g2_buf_8 fanout6137 (.A(net6138),
    .X(net6137));
 sg13g2_buf_2 fanout6138 (.A(net6139),
    .X(net6138));
 sg13g2_buf_8 fanout6139 (.A(net6140),
    .X(net6139));
 sg13g2_buf_8 fanout6140 (.A(_08133_),
    .X(net6140));
 sg13g2_buf_8 fanout6141 (.A(_08131_),
    .X(net6141));
 sg13g2_buf_8 fanout6142 (.A(_07874_),
    .X(net6142));
 sg13g2_buf_8 fanout6143 (.A(net6145),
    .X(net6143));
 sg13g2_buf_1 fanout6144 (.A(net6145),
    .X(net6144));
 sg13g2_buf_8 fanout6145 (.A(net6158),
    .X(net6145));
 sg13g2_buf_8 fanout6146 (.A(net6148),
    .X(net6146));
 sg13g2_buf_1 fanout6147 (.A(net6148),
    .X(net6147));
 sg13g2_buf_8 fanout6148 (.A(net6151),
    .X(net6148));
 sg13g2_buf_8 fanout6149 (.A(net6150),
    .X(net6149));
 sg13g2_buf_8 fanout6150 (.A(net6151),
    .X(net6150));
 sg13g2_buf_8 fanout6151 (.A(net6158),
    .X(net6151));
 sg13g2_buf_8 fanout6152 (.A(net6154),
    .X(net6152));
 sg13g2_buf_1 fanout6153 (.A(net6154),
    .X(net6153));
 sg13g2_buf_2 fanout6154 (.A(net6155),
    .X(net6154));
 sg13g2_buf_8 fanout6155 (.A(net6157),
    .X(net6155));
 sg13g2_buf_8 fanout6156 (.A(net6157),
    .X(net6156));
 sg13g2_buf_8 fanout6157 (.A(net6158),
    .X(net6157));
 sg13g2_buf_8 fanout6158 (.A(_07872_),
    .X(net6158));
 sg13g2_buf_2 fanout6159 (.A(net6161),
    .X(net6159));
 sg13g2_buf_1 fanout6160 (.A(net6161),
    .X(net6160));
 sg13g2_buf_8 fanout6161 (.A(net6165),
    .X(net6161));
 sg13g2_buf_8 fanout6162 (.A(net6165),
    .X(net6162));
 sg13g2_buf_8 fanout6163 (.A(net6164),
    .X(net6163));
 sg13g2_buf_8 fanout6164 (.A(net6165),
    .X(net6164));
 sg13g2_buf_8 fanout6165 (.A(_07868_),
    .X(net6165));
 sg13g2_buf_8 fanout6166 (.A(_07810_),
    .X(net6166));
 sg13g2_buf_8 fanout6167 (.A(_07810_),
    .X(net6167));
 sg13g2_buf_8 fanout6168 (.A(_07809_),
    .X(net6168));
 sg13g2_buf_8 fanout6169 (.A(_07809_),
    .X(net6169));
 sg13g2_buf_8 fanout6170 (.A(net6174),
    .X(net6170));
 sg13g2_buf_1 fanout6171 (.A(net6174),
    .X(net6171));
 sg13g2_buf_8 fanout6172 (.A(net6174),
    .X(net6172));
 sg13g2_buf_2 fanout6173 (.A(net6174),
    .X(net6173));
 sg13g2_buf_8 fanout6174 (.A(_07808_),
    .X(net6174));
 sg13g2_buf_8 fanout6175 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .X(net6175));
 sg13g2_buf_8 fanout6176 (.A(net6177),
    .X(net6176));
 sg13g2_buf_8 fanout6177 (.A(net6178),
    .X(net6177));
 sg13g2_buf_8 fanout6178 (.A(net2332),
    .X(net6178));
 sg13g2_buf_8 fanout6179 (.A(net3372),
    .X(net6179));
 sg13g2_buf_8 fanout6180 (.A(net6192),
    .X(net6180));
 sg13g2_buf_8 fanout6181 (.A(net6192),
    .X(net6181));
 sg13g2_buf_2 fanout6182 (.A(net6192),
    .X(net6182));
 sg13g2_buf_1 fanout6183 (.A(net6192),
    .X(net6183));
 sg13g2_buf_8 fanout6184 (.A(net6191),
    .X(net6184));
 sg13g2_buf_1 fanout6185 (.A(net6191),
    .X(net6185));
 sg13g2_buf_2 fanout6186 (.A(net6187),
    .X(net6186));
 sg13g2_buf_1 fanout6187 (.A(net6191),
    .X(net6187));
 sg13g2_buf_8 fanout6188 (.A(net6190),
    .X(net6188));
 sg13g2_buf_8 fanout6189 (.A(net6190),
    .X(net6189));
 sg13g2_buf_2 fanout6190 (.A(net6191),
    .X(net6190));
 sg13g2_buf_1 fanout6191 (.A(net6192),
    .X(net6191));
 sg13g2_buf_8 fanout6192 (.A(\soc_inst.mem_ctrl.access_state[2] ),
    .X(net6192));
 sg13g2_buf_8 fanout6193 (.A(net6195),
    .X(net6193));
 sg13g2_buf_1 fanout6194 (.A(net6195),
    .X(net6194));
 sg13g2_buf_2 fanout6195 (.A(\soc_inst.mem_ctrl.access_state[1] ),
    .X(net6195));
 sg13g2_buf_8 fanout6196 (.A(net6200),
    .X(net6196));
 sg13g2_buf_8 fanout6197 (.A(net6198),
    .X(net6197));
 sg13g2_buf_1 fanout6198 (.A(net6200),
    .X(net6198));
 sg13g2_buf_8 fanout6199 (.A(net6200),
    .X(net6199));
 sg13g2_buf_8 fanout6200 (.A(\soc_inst.mem_ctrl.access_state[1] ),
    .X(net6200));
 sg13g2_buf_8 fanout6201 (.A(net3180),
    .X(net6201));
 sg13g2_buf_8 fanout6202 (.A(net3369),
    .X(net6202));
 sg13g2_buf_1 fanout6203 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .X(net6203));
 sg13g2_buf_8 fanout6204 (.A(net6205),
    .X(net6204));
 sg13g2_buf_8 fanout6205 (.A(net2615),
    .X(net6205));
 sg13g2_buf_8 fanout6206 (.A(net6209),
    .X(net6206));
 sg13g2_buf_8 fanout6207 (.A(net6208),
    .X(net6207));
 sg13g2_buf_8 fanout6208 (.A(net6209),
    .X(net6208));
 sg13g2_buf_8 fanout6209 (.A(net6210),
    .X(net6209));
 sg13g2_buf_8 fanout6210 (.A(\soc_inst.core_mem_addr[3] ),
    .X(net6210));
 sg13g2_buf_8 fanout6211 (.A(\soc_inst.core_mem_addr[2] ),
    .X(net6211));
 sg13g2_buf_8 fanout6212 (.A(\soc_inst.core_mem_re ),
    .X(net6212));
 sg13g2_buf_8 fanout6213 (.A(net2774),
    .X(net6213));
 sg13g2_buf_8 fanout6214 (.A(net6215),
    .X(net6214));
 sg13g2_buf_2 fanout6215 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .X(net6215));
 sg13g2_buf_8 fanout6216 (.A(net6217),
    .X(net6216));
 sg13g2_buf_2 fanout6217 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .X(net6217));
 sg13g2_buf_8 fanout6218 (.A(net6220),
    .X(net6218));
 sg13g2_buf_8 fanout6219 (.A(net6220),
    .X(net6219));
 sg13g2_buf_8 fanout6220 (.A(\soc_inst.cpu_core.alu.b[4] ),
    .X(net6220));
 sg13g2_buf_8 fanout6221 (.A(\soc_inst.cpu_core.alu.b[4] ),
    .X(net6221));
 sg13g2_buf_2 fanout6222 (.A(net3397),
    .X(net6222));
 sg13g2_buf_8 fanout6223 (.A(net6224),
    .X(net6223));
 sg13g2_buf_8 fanout6224 (.A(net6232),
    .X(net6224));
 sg13g2_buf_8 fanout6225 (.A(net6232),
    .X(net6225));
 sg13g2_buf_1 fanout6226 (.A(net6232),
    .X(net6226));
 sg13g2_buf_8 fanout6227 (.A(net6229),
    .X(net6227));
 sg13g2_buf_1 fanout6228 (.A(net6229),
    .X(net6228));
 sg13g2_buf_2 fanout6229 (.A(net6230),
    .X(net6229));
 sg13g2_buf_8 fanout6230 (.A(net6231),
    .X(net6230));
 sg13g2_buf_8 fanout6231 (.A(net6232),
    .X(net6231));
 sg13g2_buf_8 fanout6232 (.A(net3324),
    .X(net6232));
 sg13g2_buf_8 fanout6233 (.A(net6236),
    .X(net6233));
 sg13g2_buf_8 fanout6234 (.A(net6235),
    .X(net6234));
 sg13g2_buf_1 fanout6235 (.A(net6236),
    .X(net6235));
 sg13g2_buf_8 fanout6236 (.A(net6239),
    .X(net6236));
 sg13g2_buf_8 fanout6237 (.A(net6239),
    .X(net6237));
 sg13g2_buf_2 fanout6238 (.A(net6239),
    .X(net6238));
 sg13g2_buf_8 fanout6239 (.A(net3390),
    .X(net6239));
 sg13g2_buf_8 fanout6240 (.A(net6244),
    .X(net6240));
 sg13g2_buf_8 fanout6241 (.A(net6242),
    .X(net6241));
 sg13g2_buf_8 fanout6242 (.A(net6243),
    .X(net6242));
 sg13g2_buf_8 fanout6243 (.A(net6244),
    .X(net6243));
 sg13g2_buf_8 fanout6244 (.A(net6248),
    .X(net6244));
 sg13g2_buf_8 fanout6245 (.A(net6246),
    .X(net6245));
 sg13g2_buf_2 fanout6246 (.A(net6247),
    .X(net6246));
 sg13g2_buf_8 fanout6247 (.A(net6248),
    .X(net6247));
 sg13g2_buf_8 fanout6248 (.A(\soc_inst.cpu_core.alu.b[1] ),
    .X(net6248));
 sg13g2_buf_8 fanout6249 (.A(net6260),
    .X(net6249));
 sg13g2_buf_8 fanout6250 (.A(net6260),
    .X(net6250));
 sg13g2_buf_8 fanout6251 (.A(net6254),
    .X(net6251));
 sg13g2_buf_8 fanout6252 (.A(net6253),
    .X(net6252));
 sg13g2_buf_8 fanout6253 (.A(net6254),
    .X(net6253));
 sg13g2_buf_2 fanout6254 (.A(net6260),
    .X(net6254));
 sg13g2_buf_8 fanout6255 (.A(net6256),
    .X(net6255));
 sg13g2_buf_8 fanout6256 (.A(net6258),
    .X(net6256));
 sg13g2_buf_8 fanout6257 (.A(net6258),
    .X(net6257));
 sg13g2_buf_8 fanout6258 (.A(net6259),
    .X(net6258));
 sg13g2_buf_8 fanout6259 (.A(net6260),
    .X(net6259));
 sg13g2_buf_8 fanout6260 (.A(\soc_inst.cpu_core.alu.b[0] ),
    .X(net6260));
 sg13g2_buf_8 fanout6261 (.A(net6262),
    .X(net6261));
 sg13g2_buf_8 fanout6262 (.A(net3259),
    .X(net6262));
 sg13g2_buf_8 fanout6263 (.A(\soc_inst.cpu_core.alu.a[29] ),
    .X(net6263));
 sg13g2_buf_8 fanout6264 (.A(net3330),
    .X(net6264));
 sg13g2_buf_8 fanout6265 (.A(net3328),
    .X(net6265));
 sg13g2_buf_8 fanout6266 (.A(net3326),
    .X(net6266));
 sg13g2_buf_1 fanout6267 (.A(\soc_inst.cpu_core.alu.a[26] ),
    .X(net6267));
 sg13g2_buf_8 fanout6268 (.A(net3350),
    .X(net6268));
 sg13g2_buf_8 fanout6269 (.A(net3336),
    .X(net6269));
 sg13g2_buf_8 fanout6270 (.A(net3387),
    .X(net6270));
 sg13g2_buf_8 fanout6271 (.A(net3385),
    .X(net6271));
 sg13g2_buf_8 fanout6272 (.A(net3319),
    .X(net6272));
 sg13g2_buf_2 fanout6273 (.A(\soc_inst.cpu_core.alu.a[21] ),
    .X(net6273));
 sg13g2_buf_8 fanout6274 (.A(net3386),
    .X(net6274));
 sg13g2_buf_2 fanout6275 (.A(\soc_inst.cpu_core.alu.a[20] ),
    .X(net6275));
 sg13g2_buf_8 fanout6276 (.A(net3395),
    .X(net6276));
 sg13g2_buf_1 fanout6277 (.A(\soc_inst.cpu_core.alu.a[19] ),
    .X(net6277));
 sg13g2_buf_8 fanout6278 (.A(net3393),
    .X(net6278));
 sg13g2_buf_8 fanout6279 (.A(net6280),
    .X(net6279));
 sg13g2_buf_8 fanout6280 (.A(net3378),
    .X(net6280));
 sg13g2_buf_8 fanout6281 (.A(net6282),
    .X(net6281));
 sg13g2_buf_8 fanout6282 (.A(net3374),
    .X(net6282));
 sg13g2_buf_8 fanout6283 (.A(net3389),
    .X(net6283));
 sg13g2_buf_8 fanout6284 (.A(net3363),
    .X(net6284));
 sg13g2_buf_8 fanout6285 (.A(net3353),
    .X(net6285));
 sg13g2_buf_8 fanout6286 (.A(net6287),
    .X(net6286));
 sg13g2_buf_8 fanout6287 (.A(net6288),
    .X(net6287));
 sg13g2_buf_8 fanout6288 (.A(net3322),
    .X(net6288));
 sg13g2_buf_8 fanout6289 (.A(net6295),
    .X(net6289));
 sg13g2_buf_8 fanout6290 (.A(net6295),
    .X(net6290));
 sg13g2_buf_8 fanout6291 (.A(net6295),
    .X(net6291));
 sg13g2_buf_8 fanout6292 (.A(net6295),
    .X(net6292));
 sg13g2_buf_8 fanout6293 (.A(net6294),
    .X(net6293));
 sg13g2_buf_8 fanout6294 (.A(net6295),
    .X(net6294));
 sg13g2_buf_8 fanout6295 (.A(\soc_inst.core_mem_flag[2] ),
    .X(net6295));
 sg13g2_buf_8 fanout6296 (.A(net6299),
    .X(net6296));
 sg13g2_buf_8 fanout6297 (.A(net6299),
    .X(net6297));
 sg13g2_buf_8 fanout6298 (.A(net6300),
    .X(net6298));
 sg13g2_buf_2 fanout6299 (.A(net6300),
    .X(net6299));
 sg13g2_buf_1 fanout6300 (.A(\soc_inst.core_mem_flag[1] ),
    .X(net6300));
 sg13g2_buf_8 fanout6301 (.A(net6303),
    .X(net6301));
 sg13g2_buf_1 fanout6302 (.A(net6303),
    .X(net6302));
 sg13g2_buf_2 fanout6303 (.A(\soc_inst.core_mem_flag[1] ),
    .X(net6303));
 sg13g2_buf_8 fanout6304 (.A(net6305),
    .X(net6304));
 sg13g2_buf_8 fanout6305 (.A(net3030),
    .X(net6305));
 sg13g2_buf_8 fanout6306 (.A(net2587),
    .X(net6306));
 sg13g2_buf_8 fanout6307 (.A(net6309),
    .X(net6307));
 sg13g2_buf_1 fanout6308 (.A(net6309),
    .X(net6308));
 sg13g2_buf_8 fanout6309 (.A(net6428),
    .X(net6309));
 sg13g2_buf_8 fanout6310 (.A(net6311),
    .X(net6310));
 sg13g2_buf_2 fanout6311 (.A(net6312),
    .X(net6311));
 sg13g2_buf_8 fanout6312 (.A(net6313),
    .X(net6312));
 sg13g2_buf_8 fanout6313 (.A(net6428),
    .X(net6313));
 sg13g2_buf_8 fanout6314 (.A(net6319),
    .X(net6314));
 sg13g2_buf_8 fanout6315 (.A(net6316),
    .X(net6315));
 sg13g2_buf_2 fanout6316 (.A(net6318),
    .X(net6316));
 sg13g2_buf_8 fanout6317 (.A(net6318),
    .X(net6317));
 sg13g2_buf_2 fanout6318 (.A(net6319),
    .X(net6318));
 sg13g2_buf_2 fanout6319 (.A(net6332),
    .X(net6319));
 sg13g2_buf_8 fanout6320 (.A(net6321),
    .X(net6320));
 sg13g2_buf_8 fanout6321 (.A(net6332),
    .X(net6321));
 sg13g2_buf_8 fanout6322 (.A(net6325),
    .X(net6322));
 sg13g2_buf_8 fanout6323 (.A(net6324),
    .X(net6323));
 sg13g2_buf_8 fanout6324 (.A(net6325),
    .X(net6324));
 sg13g2_buf_8 fanout6325 (.A(net6332),
    .X(net6325));
 sg13g2_buf_8 fanout6326 (.A(net6330),
    .X(net6326));
 sg13g2_buf_8 fanout6327 (.A(net6329),
    .X(net6327));
 sg13g2_buf_8 fanout6328 (.A(net6329),
    .X(net6328));
 sg13g2_buf_8 fanout6329 (.A(net6330),
    .X(net6329));
 sg13g2_buf_8 fanout6330 (.A(net6331),
    .X(net6330));
 sg13g2_buf_8 fanout6331 (.A(net6332),
    .X(net6331));
 sg13g2_buf_8 fanout6332 (.A(net6428),
    .X(net6332));
 sg13g2_buf_8 fanout6333 (.A(net6335),
    .X(net6333));
 sg13g2_buf_1 fanout6334 (.A(net6335),
    .X(net6334));
 sg13g2_buf_8 fanout6335 (.A(net6358),
    .X(net6335));
 sg13g2_buf_8 fanout6336 (.A(net6358),
    .X(net6336));
 sg13g2_buf_8 fanout6337 (.A(net6338),
    .X(net6337));
 sg13g2_buf_8 fanout6338 (.A(net6347),
    .X(net6338));
 sg13g2_buf_8 fanout6339 (.A(net6347),
    .X(net6339));
 sg13g2_buf_8 fanout6340 (.A(net6347),
    .X(net6340));
 sg13g2_buf_8 fanout6341 (.A(net6342),
    .X(net6341));
 sg13g2_buf_8 fanout6342 (.A(net6346),
    .X(net6342));
 sg13g2_buf_8 fanout6343 (.A(net6346),
    .X(net6343));
 sg13g2_buf_8 fanout6344 (.A(net6346),
    .X(net6344));
 sg13g2_buf_8 fanout6345 (.A(net6346),
    .X(net6345));
 sg13g2_buf_8 fanout6346 (.A(net6347),
    .X(net6346));
 sg13g2_buf_8 fanout6347 (.A(net6358),
    .X(net6347));
 sg13g2_buf_8 fanout6348 (.A(net6350),
    .X(net6348));
 sg13g2_buf_8 fanout6349 (.A(net6350),
    .X(net6349));
 sg13g2_buf_8 fanout6350 (.A(net6357),
    .X(net6350));
 sg13g2_buf_8 fanout6351 (.A(net6357),
    .X(net6351));
 sg13g2_buf_8 fanout6352 (.A(net6357),
    .X(net6352));
 sg13g2_buf_1 fanout6353 (.A(net6357),
    .X(net6353));
 sg13g2_buf_8 fanout6354 (.A(net6356),
    .X(net6354));
 sg13g2_buf_8 fanout6355 (.A(net6356),
    .X(net6355));
 sg13g2_buf_8 fanout6356 (.A(net6357),
    .X(net6356));
 sg13g2_buf_8 fanout6357 (.A(net6358),
    .X(net6357));
 sg13g2_buf_8 fanout6358 (.A(net6427),
    .X(net6358));
 sg13g2_buf_8 fanout6359 (.A(net6360),
    .X(net6359));
 sg13g2_buf_8 fanout6360 (.A(net6361),
    .X(net6360));
 sg13g2_buf_1 fanout6361 (.A(net6380),
    .X(net6361));
 sg13g2_buf_8 fanout6362 (.A(net6380),
    .X(net6362));
 sg13g2_buf_1 fanout6363 (.A(net6380),
    .X(net6363));
 sg13g2_buf_8 fanout6364 (.A(net6365),
    .X(net6364));
 sg13g2_buf_8 fanout6365 (.A(net6366),
    .X(net6365));
 sg13g2_buf_8 fanout6366 (.A(net6380),
    .X(net6366));
 sg13g2_buf_8 fanout6367 (.A(net6372),
    .X(net6367));
 sg13g2_buf_1 fanout6368 (.A(net6372),
    .X(net6368));
 sg13g2_buf_8 fanout6369 (.A(net6372),
    .X(net6369));
 sg13g2_buf_8 fanout6370 (.A(net6372),
    .X(net6370));
 sg13g2_buf_8 fanout6371 (.A(net6372),
    .X(net6371));
 sg13g2_buf_8 fanout6372 (.A(net6380),
    .X(net6372));
 sg13g2_buf_8 fanout6373 (.A(net6374),
    .X(net6373));
 sg13g2_buf_8 fanout6374 (.A(net6379),
    .X(net6374));
 sg13g2_buf_8 fanout6375 (.A(net6376),
    .X(net6375));
 sg13g2_buf_8 fanout6376 (.A(net6379),
    .X(net6376));
 sg13g2_buf_8 fanout6377 (.A(net6378),
    .X(net6377));
 sg13g2_buf_8 fanout6378 (.A(net6379),
    .X(net6378));
 sg13g2_buf_8 fanout6379 (.A(net6380),
    .X(net6379));
 sg13g2_buf_8 fanout6380 (.A(net6427),
    .X(net6380));
 sg13g2_buf_8 fanout6381 (.A(net6384),
    .X(net6381));
 sg13g2_buf_8 fanout6382 (.A(net6384),
    .X(net6382));
 sg13g2_buf_8 fanout6383 (.A(net6384),
    .X(net6383));
 sg13g2_buf_8 fanout6384 (.A(net6387),
    .X(net6384));
 sg13g2_buf_8 fanout6385 (.A(net6386),
    .X(net6385));
 sg13g2_buf_8 fanout6386 (.A(net6387),
    .X(net6386));
 sg13g2_buf_2 fanout6387 (.A(net6403),
    .X(net6387));
 sg13g2_buf_8 fanout6388 (.A(net6390),
    .X(net6388));
 sg13g2_buf_2 fanout6389 (.A(net6390),
    .X(net6389));
 sg13g2_buf_8 fanout6390 (.A(net6392),
    .X(net6390));
 sg13g2_buf_8 fanout6391 (.A(net6392),
    .X(net6391));
 sg13g2_buf_8 fanout6392 (.A(net6403),
    .X(net6392));
 sg13g2_buf_8 fanout6393 (.A(net6394),
    .X(net6393));
 sg13g2_buf_8 fanout6394 (.A(net6396),
    .X(net6394));
 sg13g2_buf_8 fanout6395 (.A(net6396),
    .X(net6395));
 sg13g2_buf_8 fanout6396 (.A(net6403),
    .X(net6396));
 sg13g2_buf_8 fanout6397 (.A(net6398),
    .X(net6397));
 sg13g2_buf_8 fanout6398 (.A(net6399),
    .X(net6398));
 sg13g2_buf_8 fanout6399 (.A(net6403),
    .X(net6399));
 sg13g2_buf_8 fanout6400 (.A(net6401),
    .X(net6400));
 sg13g2_buf_8 fanout6401 (.A(net6402),
    .X(net6401));
 sg13g2_buf_2 fanout6402 (.A(net6403),
    .X(net6402));
 sg13g2_buf_8 fanout6403 (.A(net6427),
    .X(net6403));
 sg13g2_buf_8 fanout6404 (.A(net6408),
    .X(net6404));
 sg13g2_buf_1 fanout6405 (.A(net6408),
    .X(net6405));
 sg13g2_buf_8 fanout6406 (.A(net6407),
    .X(net6406));
 sg13g2_buf_8 fanout6407 (.A(net6408),
    .X(net6407));
 sg13g2_buf_8 fanout6408 (.A(net6421),
    .X(net6408));
 sg13g2_buf_8 fanout6409 (.A(net6410),
    .X(net6409));
 sg13g2_buf_8 fanout6410 (.A(net6421),
    .X(net6410));
 sg13g2_buf_8 fanout6411 (.A(net6412),
    .X(net6411));
 sg13g2_buf_2 fanout6412 (.A(net6421),
    .X(net6412));
 sg13g2_buf_8 fanout6413 (.A(net6420),
    .X(net6413));
 sg13g2_buf_8 fanout6414 (.A(net6420),
    .X(net6414));
 sg13g2_buf_8 fanout6415 (.A(net6416),
    .X(net6415));
 sg13g2_buf_1 fanout6416 (.A(net6420),
    .X(net6416));
 sg13g2_buf_8 fanout6417 (.A(net6419),
    .X(net6417));
 sg13g2_buf_8 fanout6418 (.A(net6419),
    .X(net6418));
 sg13g2_buf_8 fanout6419 (.A(net6420),
    .X(net6419));
 sg13g2_buf_8 fanout6420 (.A(net6421),
    .X(net6420));
 sg13g2_buf_8 fanout6421 (.A(net6427),
    .X(net6421));
 sg13g2_buf_8 fanout6422 (.A(net6423),
    .X(net6422));
 sg13g2_buf_1 fanout6423 (.A(net6424),
    .X(net6423));
 sg13g2_buf_1 fanout6424 (.A(net6425),
    .X(net6424));
 sg13g2_buf_8 fanout6425 (.A(net6426),
    .X(net6425));
 sg13g2_buf_8 fanout6426 (.A(net6427),
    .X(net6426));
 sg13g2_buf_8 fanout6427 (.A(net6428),
    .X(net6427));
 sg13g2_buf_8 fanout6428 (.A(net1255),
    .X(net6428));
 sg13g2_buf_8 fanout6429 (.A(net6430),
    .X(net6429));
 sg13g2_buf_2 fanout6430 (.A(net6431),
    .X(net6430));
 sg13g2_buf_8 fanout6431 (.A(net2647),
    .X(net6431));
 sg13g2_buf_8 fanout6432 (.A(net6433),
    .X(net6432));
 sg13g2_buf_8 fanout6433 (.A(net3018),
    .X(net6433));
 sg13g2_buf_8 fanout6434 (.A(net6435),
    .X(net6434));
 sg13g2_buf_8 fanout6435 (.A(net2845),
    .X(net6435));
 sg13g2_buf_8 fanout6436 (.A(net2829),
    .X(net6436));
 sg13g2_buf_1 fanout6437 (.A(\soc_inst.cpu_core.if_imm12[1] ),
    .X(net6437));
 sg13g2_buf_8 fanout6438 (.A(net3396),
    .X(net6438));
 sg13g2_buf_2 fanout6439 (.A(\soc_inst.cpu_core.if_imm12[0] ),
    .X(net6439));
 sg13g2_buf_8 fanout6440 (.A(net6441),
    .X(net6440));
 sg13g2_buf_8 fanout6441 (.A(net6442),
    .X(net6441));
 sg13g2_buf_2 fanout6442 (.A(net6443),
    .X(net6442));
 sg13g2_buf_8 fanout6443 (.A(net2281),
    .X(net6443));
 sg13g2_buf_8 fanout6444 (.A(net1492),
    .X(net6444));
 sg13g2_buf_8 fanout6445 (.A(net1841),
    .X(net6445));
 sg13g2_buf_8 fanout6446 (.A(net6447),
    .X(net6446));
 sg13g2_buf_1 fanout6447 (.A(net6448),
    .X(net6447));
 sg13g2_buf_8 fanout6448 (.A(net1512),
    .X(net6448));
 sg13g2_buf_8 fanout6449 (.A(net6450),
    .X(net6449));
 sg13g2_buf_8 fanout6450 (.A(net1858),
    .X(net6450));
 sg13g2_buf_8 fanout6451 (.A(net6452),
    .X(net6451));
 sg13g2_buf_8 fanout6452 (.A(net3236),
    .X(net6452));
 sg13g2_buf_8 fanout6453 (.A(net219),
    .X(net6453));
 sg13g2_buf_8 fanout6454 (.A(net1497),
    .X(net6454));
 sg13g2_buf_8 fanout6455 (.A(net1434),
    .X(net6455));
 sg13g2_buf_8 fanout6456 (.A(net1434),
    .X(net6456));
 sg13g2_buf_8 fanout6457 (.A(net1399),
    .X(net6457));
 sg13g2_buf_8 fanout6458 (.A(net1399),
    .X(net6458));
 sg13g2_buf_8 fanout6459 (.A(net1518),
    .X(net6459));
 sg13g2_buf_8 fanout6460 (.A(net1518),
    .X(net6460));
 sg13g2_buf_8 fanout6461 (.A(net6462),
    .X(net6461));
 sg13g2_buf_8 fanout6462 (.A(net245),
    .X(net6462));
 sg13g2_buf_8 fanout6463 (.A(net6464),
    .X(net6463));
 sg13g2_buf_8 fanout6464 (.A(net212),
    .X(net6464));
 sg13g2_buf_8 fanout6465 (.A(net6466),
    .X(net6465));
 sg13g2_buf_8 fanout6466 (.A(net6467),
    .X(net6466));
 sg13g2_buf_8 fanout6467 (.A(net3348),
    .X(net6467));
 sg13g2_buf_8 fanout6468 (.A(net6469),
    .X(net6468));
 sg13g2_buf_8 fanout6469 (.A(net3090),
    .X(net6469));
 sg13g2_buf_8 fanout6470 (.A(net6471),
    .X(net6470));
 sg13g2_buf_8 fanout6471 (.A(net2724),
    .X(net6471));
 sg13g2_buf_8 fanout6472 (.A(net6477),
    .X(net6472));
 sg13g2_buf_8 fanout6473 (.A(net6474),
    .X(net6473));
 sg13g2_buf_8 fanout6474 (.A(net6477),
    .X(net6474));
 sg13g2_buf_8 fanout6475 (.A(net6477),
    .X(net6475));
 sg13g2_buf_2 fanout6476 (.A(net6477),
    .X(net6476));
 sg13g2_buf_8 fanout6477 (.A(net3058),
    .X(net6477));
 sg13g2_buf_8 fanout6478 (.A(net6479),
    .X(net6478));
 sg13g2_buf_8 fanout6479 (.A(net6481),
    .X(net6479));
 sg13g2_buf_8 fanout6480 (.A(net6481),
    .X(net6480));
 sg13g2_buf_2 fanout6481 (.A(\soc_inst.cpu_core.id_int_is_interrupt ),
    .X(net6481));
 sg13g2_buf_8 fanout6482 (.A(net6483),
    .X(net6482));
 sg13g2_buf_8 fanout6483 (.A(\soc_inst.mem_ctrl.spi_mem_inst.write_mosi ),
    .X(net6483));
 sg13g2_buf_8 fanout6484 (.A(net3261),
    .X(net6484));
 sg13g2_buf_8 fanout6485 (.A(net3375),
    .X(net6485));
 sg13g2_buf_8 fanout6486 (.A(net3392),
    .X(net6486));
 sg13g2_buf_8 fanout6487 (.A(net3113),
    .X(net6487));
 sg13g2_buf_8 fanout6488 (.A(net1775),
    .X(net6488));
 sg13g2_buf_8 fanout6489 (.A(net6495),
    .X(net6489));
 sg13g2_buf_8 fanout6490 (.A(net6495),
    .X(net6490));
 sg13g2_buf_8 fanout6491 (.A(net6494),
    .X(net6491));
 sg13g2_buf_8 fanout6492 (.A(net6494),
    .X(net6492));
 sg13g2_buf_1 fanout6493 (.A(net6494),
    .X(net6493));
 sg13g2_buf_8 fanout6494 (.A(net6495),
    .X(net6494));
 sg13g2_buf_8 fanout6495 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[6] ),
    .X(net6495));
 sg13g2_buf_8 fanout6496 (.A(net6499),
    .X(net6496));
 sg13g2_buf_8 fanout6497 (.A(net6499),
    .X(net6497));
 sg13g2_buf_1 fanout6498 (.A(net6499),
    .X(net6498));
 sg13g2_buf_2 fanout6499 (.A(net6502),
    .X(net6499));
 sg13g2_buf_8 fanout6500 (.A(net6502),
    .X(net6500));
 sg13g2_buf_2 fanout6501 (.A(net6502),
    .X(net6501));
 sg13g2_buf_8 fanout6502 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[4] ),
    .X(net6502));
 sg13g2_buf_8 fanout6503 (.A(net3009),
    .X(net6503));
 sg13g2_buf_8 fanout6504 (.A(net6505),
    .X(net6504));
 sg13g2_buf_8 fanout6505 (.A(net3327),
    .X(net6505));
 sg13g2_buf_8 fanout6506 (.A(net97),
    .X(net6506));
 sg13g2_buf_8 fanout6507 (.A(net3190),
    .X(net6507));
 sg13g2_buf_8 fanout6508 (.A(net6509),
    .X(net6508));
 sg13g2_buf_8 fanout6509 (.A(net3347),
    .X(net6509));
 sg13g2_buf_8 fanout6510 (.A(net6511),
    .X(net6510));
 sg13g2_buf_8 fanout6511 (.A(net3381),
    .X(net6511));
 sg13g2_buf_8 fanout6512 (.A(net6514),
    .X(net6512));
 sg13g2_buf_8 fanout6513 (.A(net6514),
    .X(net6513));
 sg13g2_buf_8 fanout6514 (.A(net3394),
    .X(net6514));
 sg13g2_buf_8 fanout6515 (.A(net6516),
    .X(net6515));
 sg13g2_buf_2 fanout6516 (.A(net6517),
    .X(net6516));
 sg13g2_buf_8 fanout6517 (.A(\soc_inst.core_instr_data[12] ),
    .X(net6517));
 sg13g2_buf_8 fanout6518 (.A(net3323),
    .X(net6518));
 sg13g2_buf_8 fanout6519 (.A(\soc_inst.core_instr_data[11] ),
    .X(net6519));
 sg13g2_buf_8 fanout6520 (.A(net6521),
    .X(net6520));
 sg13g2_buf_8 fanout6521 (.A(net3365),
    .X(net6521));
 sg13g2_buf_8 fanout6522 (.A(net6523),
    .X(net6522));
 sg13g2_buf_8 fanout6523 (.A(net3307),
    .X(net6523));
 sg13g2_buf_8 fanout6524 (.A(net6525),
    .X(net6524));
 sg13g2_buf_8 fanout6525 (.A(net3364),
    .X(net6525));
 sg13g2_buf_8 fanout6526 (.A(net3373),
    .X(net6526));
 sg13g2_buf_8 fanout6527 (.A(\soc_inst.core_instr_data[6] ),
    .X(net6527));
 sg13g2_buf_8 fanout6528 (.A(net3341),
    .X(net6528));
 sg13g2_buf_8 fanout6529 (.A(net3343),
    .X(net6529));
 sg13g2_buf_8 fanout6530 (.A(net2799),
    .X(net6530));
 sg13g2_buf_8 fanout6531 (.A(net2761),
    .X(net6531));
 sg13g2_buf_8 fanout6532 (.A(net2739),
    .X(net6532));
 sg13g2_buf_8 fanout6533 (.A(net3349),
    .X(net6533));
 sg13g2_buf_8 fanout6534 (.A(net3240),
    .X(net6534));
 sg13g2_buf_8 fanout6535 (.A(net6536),
    .X(net6535));
 sg13g2_buf_2 fanout6536 (.A(net3352),
    .X(net6536));
 sg13g2_buf_8 fanout6537 (.A(net6538),
    .X(net6537));
 sg13g2_buf_1 fanout6538 (.A(net3384),
    .X(net6538));
 sg13g2_buf_8 fanout6539 (.A(net6540),
    .X(net6539));
 sg13g2_buf_8 fanout6540 (.A(net3217),
    .X(net6540));
 sg13g2_buf_8 fanout6541 (.A(net6542),
    .X(net6541));
 sg13g2_buf_8 fanout6542 (.A(net6543),
    .X(net6542));
 sg13g2_buf_8 fanout6543 (.A(net2853),
    .X(net6543));
 sg13g2_buf_8 fanout6544 (.A(net6545),
    .X(net6544));
 sg13g2_buf_8 fanout6545 (.A(net3355),
    .X(net6545));
 sg13g2_buf_8 fanout6546 (.A(net241),
    .X(net6546));
 sg13g2_buf_8 fanout6547 (.A(net6548),
    .X(net6547));
 sg13g2_buf_8 fanout6548 (.A(net6549),
    .X(net6548));
 sg13g2_buf_8 fanout6549 (.A(net6566),
    .X(net6549));
 sg13g2_buf_8 fanout6550 (.A(net6566),
    .X(net6550));
 sg13g2_buf_8 fanout6551 (.A(net6552),
    .X(net6551));
 sg13g2_buf_8 fanout6552 (.A(net6566),
    .X(net6552));
 sg13g2_buf_8 fanout6553 (.A(net6566),
    .X(net6553));
 sg13g2_buf_8 fanout6554 (.A(net6556),
    .X(net6554));
 sg13g2_buf_8 fanout6555 (.A(net6556),
    .X(net6555));
 sg13g2_buf_8 fanout6556 (.A(net6566),
    .X(net6556));
 sg13g2_buf_8 fanout6557 (.A(net6560),
    .X(net6557));
 sg13g2_buf_2 fanout6558 (.A(net6560),
    .X(net6558));
 sg13g2_buf_8 fanout6559 (.A(net6560),
    .X(net6559));
 sg13g2_buf_8 fanout6560 (.A(net6566),
    .X(net6560));
 sg13g2_buf_8 fanout6561 (.A(net6562),
    .X(net6561));
 sg13g2_buf_8 fanout6562 (.A(net6565),
    .X(net6562));
 sg13g2_buf_8 fanout6563 (.A(net6564),
    .X(net6563));
 sg13g2_buf_8 fanout6564 (.A(net6565),
    .X(net6564));
 sg13g2_buf_8 fanout6565 (.A(net6566),
    .X(net6565));
 sg13g2_buf_8 fanout6566 (.A(net6599),
    .X(net6566));
 sg13g2_buf_8 fanout6567 (.A(net6569),
    .X(net6567));
 sg13g2_buf_8 fanout6568 (.A(net6569),
    .X(net6568));
 sg13g2_buf_8 fanout6569 (.A(net6575),
    .X(net6569));
 sg13g2_buf_8 fanout6570 (.A(net6571),
    .X(net6570));
 sg13g2_buf_8 fanout6571 (.A(net6575),
    .X(net6571));
 sg13g2_buf_8 fanout6572 (.A(net6573),
    .X(net6572));
 sg13g2_buf_8 fanout6573 (.A(net6574),
    .X(net6573));
 sg13g2_buf_8 fanout6574 (.A(net6575),
    .X(net6574));
 sg13g2_buf_8 fanout6575 (.A(net6599),
    .X(net6575));
 sg13g2_buf_8 fanout6576 (.A(net6583),
    .X(net6576));
 sg13g2_buf_8 fanout6577 (.A(net6578),
    .X(net6577));
 sg13g2_buf_8 fanout6578 (.A(net6583),
    .X(net6578));
 sg13g2_buf_8 fanout6579 (.A(net6580),
    .X(net6579));
 sg13g2_buf_8 fanout6580 (.A(net6583),
    .X(net6580));
 sg13g2_buf_8 fanout6581 (.A(net6582),
    .X(net6581));
 sg13g2_buf_8 fanout6582 (.A(net6583),
    .X(net6582));
 sg13g2_buf_8 fanout6583 (.A(net6599),
    .X(net6583));
 sg13g2_buf_8 fanout6584 (.A(net6598),
    .X(net6584));
 sg13g2_buf_8 fanout6585 (.A(net6598),
    .X(net6585));
 sg13g2_buf_8 fanout6586 (.A(net6588),
    .X(net6586));
 sg13g2_buf_8 fanout6587 (.A(net6588),
    .X(net6587));
 sg13g2_buf_8 fanout6588 (.A(net6598),
    .X(net6588));
 sg13g2_buf_8 fanout6589 (.A(net6592),
    .X(net6589));
 sg13g2_buf_8 fanout6590 (.A(net6592),
    .X(net6590));
 sg13g2_buf_8 fanout6591 (.A(net6592),
    .X(net6591));
 sg13g2_buf_8 fanout6592 (.A(net6597),
    .X(net6592));
 sg13g2_buf_8 fanout6593 (.A(net6597),
    .X(net6593));
 sg13g2_buf_8 fanout6594 (.A(net6597),
    .X(net6594));
 sg13g2_buf_8 fanout6595 (.A(net6596),
    .X(net6595));
 sg13g2_buf_8 fanout6596 (.A(net6597),
    .X(net6596));
 sg13g2_buf_8 fanout6597 (.A(net6598),
    .X(net6597));
 sg13g2_buf_8 fanout6598 (.A(net6599),
    .X(net6598));
 sg13g2_buf_8 fanout6599 (.A(net6755),
    .X(net6599));
 sg13g2_buf_8 fanout6600 (.A(net6603),
    .X(net6600));
 sg13g2_buf_1 fanout6601 (.A(net6603),
    .X(net6601));
 sg13g2_buf_8 fanout6602 (.A(net6603),
    .X(net6602));
 sg13g2_buf_8 fanout6603 (.A(net6629),
    .X(net6603));
 sg13g2_buf_8 fanout6604 (.A(net6605),
    .X(net6604));
 sg13g2_buf_8 fanout6605 (.A(net6629),
    .X(net6605));
 sg13g2_buf_8 fanout6606 (.A(net6612),
    .X(net6606));
 sg13g2_buf_1 fanout6607 (.A(net6612),
    .X(net6607));
 sg13g2_buf_8 fanout6608 (.A(net6612),
    .X(net6608));
 sg13g2_buf_8 fanout6609 (.A(net6611),
    .X(net6609));
 sg13g2_buf_8 fanout6610 (.A(net6611),
    .X(net6610));
 sg13g2_buf_8 fanout6611 (.A(net6612),
    .X(net6611));
 sg13g2_buf_8 fanout6612 (.A(net6629),
    .X(net6612));
 sg13g2_buf_8 fanout6613 (.A(net6614),
    .X(net6613));
 sg13g2_buf_8 fanout6614 (.A(net6617),
    .X(net6614));
 sg13g2_buf_8 fanout6615 (.A(net6617),
    .X(net6615));
 sg13g2_buf_2 fanout6616 (.A(net6617),
    .X(net6616));
 sg13g2_buf_8 fanout6617 (.A(net6628),
    .X(net6617));
 sg13g2_buf_8 fanout6618 (.A(net6620),
    .X(net6618));
 sg13g2_buf_1 fanout6619 (.A(net6620),
    .X(net6619));
 sg13g2_buf_8 fanout6620 (.A(net6628),
    .X(net6620));
 sg13g2_buf_8 fanout6621 (.A(net6623),
    .X(net6621));
 sg13g2_buf_8 fanout6622 (.A(net6623),
    .X(net6622));
 sg13g2_buf_8 fanout6623 (.A(net6628),
    .X(net6623));
 sg13g2_buf_8 fanout6624 (.A(net6627),
    .X(net6624));
 sg13g2_buf_1 fanout6625 (.A(net6627),
    .X(net6625));
 sg13g2_buf_8 fanout6626 (.A(net6627),
    .X(net6626));
 sg13g2_buf_8 fanout6627 (.A(net6628),
    .X(net6627));
 sg13g2_buf_8 fanout6628 (.A(net6629),
    .X(net6628));
 sg13g2_buf_8 fanout6629 (.A(net6755),
    .X(net6629));
 sg13g2_buf_8 fanout6630 (.A(net6631),
    .X(net6630));
 sg13g2_buf_8 fanout6631 (.A(net6632),
    .X(net6631));
 sg13g2_buf_8 fanout6632 (.A(net6635),
    .X(net6632));
 sg13g2_buf_8 fanout6633 (.A(net6635),
    .X(net6633));
 sg13g2_buf_8 fanout6634 (.A(net6635),
    .X(net6634));
 sg13g2_buf_8 fanout6635 (.A(net6656),
    .X(net6635));
 sg13g2_buf_8 fanout6636 (.A(net6638),
    .X(net6636));
 sg13g2_buf_8 fanout6637 (.A(net6638),
    .X(net6637));
 sg13g2_buf_8 fanout6638 (.A(net6656),
    .X(net6638));
 sg13g2_buf_8 fanout6639 (.A(net6640),
    .X(net6639));
 sg13g2_buf_8 fanout6640 (.A(net6656),
    .X(net6640));
 sg13g2_buf_8 fanout6641 (.A(net6645),
    .X(net6641));
 sg13g2_buf_8 fanout6642 (.A(net6645),
    .X(net6642));
 sg13g2_buf_8 fanout6643 (.A(net6645),
    .X(net6643));
 sg13g2_buf_8 fanout6644 (.A(net6645),
    .X(net6644));
 sg13g2_buf_8 fanout6645 (.A(net6656),
    .X(net6645));
 sg13g2_buf_8 fanout6646 (.A(net6647),
    .X(net6646));
 sg13g2_buf_8 fanout6647 (.A(net6655),
    .X(net6647));
 sg13g2_buf_8 fanout6648 (.A(net6655),
    .X(net6648));
 sg13g2_buf_2 fanout6649 (.A(net6655),
    .X(net6649));
 sg13g2_buf_8 fanout6650 (.A(net6654),
    .X(net6650));
 sg13g2_buf_8 fanout6651 (.A(net6654),
    .X(net6651));
 sg13g2_buf_8 fanout6652 (.A(net6654),
    .X(net6652));
 sg13g2_buf_8 fanout6653 (.A(net6654),
    .X(net6653));
 sg13g2_buf_8 fanout6654 (.A(net6655),
    .X(net6654));
 sg13g2_buf_8 fanout6655 (.A(net6656),
    .X(net6655));
 sg13g2_buf_8 fanout6656 (.A(net6755),
    .X(net6656));
 sg13g2_buf_8 fanout6657 (.A(net6660),
    .X(net6657));
 sg13g2_buf_8 fanout6658 (.A(net6660),
    .X(net6658));
 sg13g2_buf_8 fanout6659 (.A(net6660),
    .X(net6659));
 sg13g2_buf_8 fanout6660 (.A(net6670),
    .X(net6660));
 sg13g2_buf_8 fanout6661 (.A(net6665),
    .X(net6661));
 sg13g2_buf_8 fanout6662 (.A(net6665),
    .X(net6662));
 sg13g2_buf_8 fanout6663 (.A(net6665),
    .X(net6663));
 sg13g2_buf_2 fanout6664 (.A(net6665),
    .X(net6664));
 sg13g2_buf_8 fanout6665 (.A(net6670),
    .X(net6665));
 sg13g2_buf_8 fanout6666 (.A(net6670),
    .X(net6666));
 sg13g2_buf_8 fanout6667 (.A(net6670),
    .X(net6667));
 sg13g2_buf_8 fanout6668 (.A(net6669),
    .X(net6668));
 sg13g2_buf_8 fanout6669 (.A(net6670),
    .X(net6669));
 sg13g2_buf_8 fanout6670 (.A(net6754),
    .X(net6670));
 sg13g2_buf_8 fanout6671 (.A(net6674),
    .X(net6671));
 sg13g2_buf_8 fanout6672 (.A(net6674),
    .X(net6672));
 sg13g2_buf_8 fanout6673 (.A(net6674),
    .X(net6673));
 sg13g2_buf_8 fanout6674 (.A(net6683),
    .X(net6674));
 sg13g2_buf_8 fanout6675 (.A(net6677),
    .X(net6675));
 sg13g2_buf_1 fanout6676 (.A(net6677),
    .X(net6676));
 sg13g2_buf_8 fanout6677 (.A(net6683),
    .X(net6677));
 sg13g2_buf_8 fanout6678 (.A(net6682),
    .X(net6678));
 sg13g2_buf_8 fanout6679 (.A(net6682),
    .X(net6679));
 sg13g2_buf_8 fanout6680 (.A(net6681),
    .X(net6680));
 sg13g2_buf_8 fanout6681 (.A(net6682),
    .X(net6681));
 sg13g2_buf_8 fanout6682 (.A(net6683),
    .X(net6682));
 sg13g2_buf_8 fanout6683 (.A(net6754),
    .X(net6683));
 sg13g2_buf_8 fanout6684 (.A(net6688),
    .X(net6684));
 sg13g2_buf_8 fanout6685 (.A(net6688),
    .X(net6685));
 sg13g2_buf_8 fanout6686 (.A(net6688),
    .X(net6686));
 sg13g2_buf_2 fanout6687 (.A(net6688),
    .X(net6687));
 sg13g2_buf_8 fanout6688 (.A(net6708),
    .X(net6688));
 sg13g2_buf_8 fanout6689 (.A(net6692),
    .X(net6689));
 sg13g2_buf_8 fanout6690 (.A(net6691),
    .X(net6690));
 sg13g2_buf_8 fanout6691 (.A(net6692),
    .X(net6691));
 sg13g2_buf_8 fanout6692 (.A(net6708),
    .X(net6692));
 sg13g2_buf_8 fanout6693 (.A(net6697),
    .X(net6693));
 sg13g2_buf_8 fanout6694 (.A(net6697),
    .X(net6694));
 sg13g2_buf_8 fanout6695 (.A(net6697),
    .X(net6695));
 sg13g2_buf_8 fanout6696 (.A(net6697),
    .X(net6696));
 sg13g2_buf_8 fanout6697 (.A(net6708),
    .X(net6697));
 sg13g2_buf_8 fanout6698 (.A(net6699),
    .X(net6698));
 sg13g2_buf_8 fanout6699 (.A(net6703),
    .X(net6699));
 sg13g2_buf_8 fanout6700 (.A(net6702),
    .X(net6700));
 sg13g2_buf_8 fanout6701 (.A(net6702),
    .X(net6701));
 sg13g2_buf_8 fanout6702 (.A(net6703),
    .X(net6702));
 sg13g2_buf_8 fanout6703 (.A(net6708),
    .X(net6703));
 sg13g2_buf_8 fanout6704 (.A(net6705),
    .X(net6704));
 sg13g2_buf_8 fanout6705 (.A(net6707),
    .X(net6705));
 sg13g2_buf_8 fanout6706 (.A(net6707),
    .X(net6706));
 sg13g2_buf_8 fanout6707 (.A(net6708),
    .X(net6707));
 sg13g2_buf_8 fanout6708 (.A(net6754),
    .X(net6708));
 sg13g2_buf_8 fanout6709 (.A(net6711),
    .X(net6709));
 sg13g2_buf_8 fanout6710 (.A(net6711),
    .X(net6710));
 sg13g2_buf_8 fanout6711 (.A(net6722),
    .X(net6711));
 sg13g2_buf_8 fanout6712 (.A(net6714),
    .X(net6712));
 sg13g2_buf_8 fanout6713 (.A(net6714),
    .X(net6713));
 sg13g2_buf_8 fanout6714 (.A(net6722),
    .X(net6714));
 sg13g2_buf_8 fanout6715 (.A(net6716),
    .X(net6715));
 sg13g2_buf_8 fanout6716 (.A(net6721),
    .X(net6716));
 sg13g2_buf_8 fanout6717 (.A(net6720),
    .X(net6717));
 sg13g2_buf_8 fanout6718 (.A(net6720),
    .X(net6718));
 sg13g2_buf_8 fanout6719 (.A(net6720),
    .X(net6719));
 sg13g2_buf_8 fanout6720 (.A(net6721),
    .X(net6720));
 sg13g2_buf_8 fanout6721 (.A(net6722),
    .X(net6721));
 sg13g2_buf_8 fanout6722 (.A(net6753),
    .X(net6722));
 sg13g2_buf_8 fanout6723 (.A(net6724),
    .X(net6723));
 sg13g2_buf_8 fanout6724 (.A(net6736),
    .X(net6724));
 sg13g2_buf_8 fanout6725 (.A(net6727),
    .X(net6725));
 sg13g2_buf_8 fanout6726 (.A(net6727),
    .X(net6726));
 sg13g2_buf_8 fanout6727 (.A(net6736),
    .X(net6727));
 sg13g2_buf_8 fanout6728 (.A(net6730),
    .X(net6728));
 sg13g2_buf_8 fanout6729 (.A(net6730),
    .X(net6729));
 sg13g2_buf_8 fanout6730 (.A(net6736),
    .X(net6730));
 sg13g2_buf_8 fanout6731 (.A(net6735),
    .X(net6731));
 sg13g2_buf_8 fanout6732 (.A(net6735),
    .X(net6732));
 sg13g2_buf_8 fanout6733 (.A(net6735),
    .X(net6733));
 sg13g2_buf_2 fanout6734 (.A(net6735),
    .X(net6734));
 sg13g2_buf_8 fanout6735 (.A(net6736),
    .X(net6735));
 sg13g2_buf_8 fanout6736 (.A(net6753),
    .X(net6736));
 sg13g2_buf_8 fanout6737 (.A(net6739),
    .X(net6737));
 sg13g2_buf_8 fanout6738 (.A(net6739),
    .X(net6738));
 sg13g2_buf_8 fanout6739 (.A(net6742),
    .X(net6739));
 sg13g2_buf_8 fanout6740 (.A(net6741),
    .X(net6740));
 sg13g2_buf_8 fanout6741 (.A(net6742),
    .X(net6741));
 sg13g2_buf_8 fanout6742 (.A(net6743),
    .X(net6742));
 sg13g2_buf_8 fanout6743 (.A(net6753),
    .X(net6743));
 sg13g2_buf_8 fanout6744 (.A(net6745),
    .X(net6744));
 sg13g2_buf_8 fanout6745 (.A(net6752),
    .X(net6745));
 sg13g2_buf_8 fanout6746 (.A(net6747),
    .X(net6746));
 sg13g2_buf_8 fanout6747 (.A(net6752),
    .X(net6747));
 sg13g2_buf_8 fanout6748 (.A(net6751),
    .X(net6748));
 sg13g2_buf_8 fanout6749 (.A(net6751),
    .X(net6749));
 sg13g2_buf_8 fanout6750 (.A(net6751),
    .X(net6750));
 sg13g2_buf_8 fanout6751 (.A(net6752),
    .X(net6751));
 sg13g2_buf_8 fanout6752 (.A(net6753),
    .X(net6752));
 sg13g2_buf_8 fanout6753 (.A(net6754),
    .X(net6753));
 sg13g2_buf_8 fanout6754 (.A(net6755),
    .X(net6754));
 sg13g2_buf_8 fanout6755 (.A(rst_n),
    .X(net6755));
 sg13g2_buf_8 fanout6756 (.A(net6758),
    .X(net6756));
 sg13g2_buf_8 fanout6757 (.A(net6758),
    .X(net6757));
 sg13g2_buf_8 fanout6758 (.A(net6779),
    .X(net6758));
 sg13g2_buf_8 fanout6759 (.A(net6760),
    .X(net6759));
 sg13g2_buf_8 fanout6760 (.A(net6779),
    .X(net6760));
 sg13g2_buf_8 fanout6761 (.A(net6768),
    .X(net6761));
 sg13g2_buf_8 fanout6762 (.A(net6768),
    .X(net6762));
 sg13g2_buf_8 fanout6763 (.A(net6764),
    .X(net6763));
 sg13g2_buf_8 fanout6764 (.A(net6765),
    .X(net6764));
 sg13g2_buf_8 fanout6765 (.A(net6768),
    .X(net6765));
 sg13g2_buf_8 fanout6766 (.A(net6768),
    .X(net6766));
 sg13g2_buf_2 fanout6767 (.A(net6768),
    .X(net6767));
 sg13g2_buf_8 fanout6768 (.A(net6779),
    .X(net6768));
 sg13g2_buf_8 fanout6769 (.A(net6770),
    .X(net6769));
 sg13g2_buf_8 fanout6770 (.A(net6779),
    .X(net6770));
 sg13g2_buf_8 fanout6771 (.A(net6772),
    .X(net6771));
 sg13g2_buf_8 fanout6772 (.A(net6775),
    .X(net6772));
 sg13g2_buf_8 fanout6773 (.A(net6775),
    .X(net6773));
 sg13g2_buf_8 fanout6774 (.A(net6775),
    .X(net6774));
 sg13g2_buf_8 fanout6775 (.A(net6779),
    .X(net6775));
 sg13g2_buf_8 fanout6776 (.A(net6777),
    .X(net6776));
 sg13g2_buf_8 fanout6777 (.A(net6778),
    .X(net6777));
 sg13g2_buf_8 fanout6778 (.A(net6779),
    .X(net6778));
 sg13g2_buf_8 fanout6779 (.A(net6986),
    .X(net6779));
 sg13g2_buf_8 fanout6780 (.A(net6783),
    .X(net6780));
 sg13g2_buf_8 fanout6781 (.A(net6783),
    .X(net6781));
 sg13g2_buf_8 fanout6782 (.A(net6783),
    .X(net6782));
 sg13g2_buf_8 fanout6783 (.A(net6786),
    .X(net6783));
 sg13g2_buf_8 fanout6784 (.A(net6785),
    .X(net6784));
 sg13g2_buf_8 fanout6785 (.A(net6786),
    .X(net6785));
 sg13g2_buf_8 fanout6786 (.A(net6805),
    .X(net6786));
 sg13g2_buf_8 fanout6787 (.A(net6790),
    .X(net6787));
 sg13g2_buf_8 fanout6788 (.A(net6790),
    .X(net6788));
 sg13g2_buf_2 fanout6789 (.A(net6790),
    .X(net6789));
 sg13g2_buf_8 fanout6790 (.A(net6805),
    .X(net6790));
 sg13g2_buf_8 fanout6791 (.A(net6792),
    .X(net6791));
 sg13g2_buf_2 fanout6792 (.A(net6795),
    .X(net6792));
 sg13g2_buf_8 fanout6793 (.A(net6795),
    .X(net6793));
 sg13g2_buf_8 fanout6794 (.A(net6795),
    .X(net6794));
 sg13g2_buf_8 fanout6795 (.A(net6805),
    .X(net6795));
 sg13g2_buf_8 fanout6796 (.A(net6798),
    .X(net6796));
 sg13g2_buf_2 fanout6797 (.A(net6798),
    .X(net6797));
 sg13g2_buf_8 fanout6798 (.A(net6800),
    .X(net6798));
 sg13g2_buf_8 fanout6799 (.A(net6800),
    .X(net6799));
 sg13g2_buf_8 fanout6800 (.A(net6805),
    .X(net6800));
 sg13g2_buf_8 fanout6801 (.A(net6802),
    .X(net6801));
 sg13g2_buf_8 fanout6802 (.A(net6805),
    .X(net6802));
 sg13g2_buf_8 fanout6803 (.A(net6804),
    .X(net6803));
 sg13g2_buf_8 fanout6804 (.A(net6805),
    .X(net6804));
 sg13g2_buf_8 fanout6805 (.A(net6986),
    .X(net6805));
 sg13g2_buf_8 fanout6806 (.A(net6812),
    .X(net6806));
 sg13g2_buf_8 fanout6807 (.A(net6812),
    .X(net6807));
 sg13g2_buf_8 fanout6808 (.A(net6809),
    .X(net6808));
 sg13g2_buf_8 fanout6809 (.A(net6812),
    .X(net6809));
 sg13g2_buf_8 fanout6810 (.A(net6811),
    .X(net6810));
 sg13g2_buf_8 fanout6811 (.A(net6812),
    .X(net6811));
 sg13g2_buf_8 fanout6812 (.A(net6831),
    .X(net6812));
 sg13g2_buf_8 fanout6813 (.A(net6814),
    .X(net6813));
 sg13g2_buf_8 fanout6814 (.A(net6831),
    .X(net6814));
 sg13g2_buf_8 fanout6815 (.A(net6831),
    .X(net6815));
 sg13g2_buf_8 fanout6816 (.A(net6820),
    .X(net6816));
 sg13g2_buf_8 fanout6817 (.A(net6820),
    .X(net6817));
 sg13g2_buf_8 fanout6818 (.A(net6820),
    .X(net6818));
 sg13g2_buf_8 fanout6819 (.A(net6820),
    .X(net6819));
 sg13g2_buf_8 fanout6820 (.A(net6830),
    .X(net6820));
 sg13g2_buf_8 fanout6821 (.A(net6830),
    .X(net6821));
 sg13g2_buf_2 fanout6822 (.A(net6830),
    .X(net6822));
 sg13g2_buf_8 fanout6823 (.A(net6825),
    .X(net6823));
 sg13g2_buf_8 fanout6824 (.A(net6825),
    .X(net6824));
 sg13g2_buf_8 fanout6825 (.A(net6830),
    .X(net6825));
 sg13g2_buf_8 fanout6826 (.A(net6827),
    .X(net6826));
 sg13g2_buf_8 fanout6827 (.A(net6830),
    .X(net6827));
 sg13g2_buf_8 fanout6828 (.A(net6829),
    .X(net6828));
 sg13g2_buf_8 fanout6829 (.A(net6830),
    .X(net6829));
 sg13g2_buf_8 fanout6830 (.A(net6831),
    .X(net6830));
 sg13g2_buf_8 fanout6831 (.A(net6848),
    .X(net6831));
 sg13g2_buf_8 fanout6832 (.A(net6833),
    .X(net6832));
 sg13g2_buf_8 fanout6833 (.A(net6834),
    .X(net6833));
 sg13g2_buf_8 fanout6834 (.A(net6848),
    .X(net6834));
 sg13g2_buf_8 fanout6835 (.A(net6837),
    .X(net6835));
 sg13g2_buf_8 fanout6836 (.A(net6837),
    .X(net6836));
 sg13g2_buf_8 fanout6837 (.A(net6838),
    .X(net6837));
 sg13g2_buf_8 fanout6838 (.A(net6839),
    .X(net6838));
 sg13g2_buf_8 fanout6839 (.A(net6848),
    .X(net6839));
 sg13g2_buf_8 fanout6840 (.A(net6841),
    .X(net6840));
 sg13g2_buf_8 fanout6841 (.A(net6847),
    .X(net6841));
 sg13g2_buf_8 fanout6842 (.A(net6843),
    .X(net6842));
 sg13g2_buf_8 fanout6843 (.A(net6847),
    .X(net6843));
 sg13g2_buf_8 fanout6844 (.A(net6847),
    .X(net6844));
 sg13g2_buf_8 fanout6845 (.A(net6847),
    .X(net6845));
 sg13g2_buf_8 fanout6846 (.A(net6847),
    .X(net6846));
 sg13g2_buf_8 fanout6847 (.A(net6848),
    .X(net6847));
 sg13g2_buf_8 fanout6848 (.A(net6986),
    .X(net6848));
 sg13g2_buf_8 fanout6849 (.A(net6850),
    .X(net6849));
 sg13g2_buf_8 fanout6850 (.A(net6853),
    .X(net6850));
 sg13g2_buf_8 fanout6851 (.A(net6853),
    .X(net6851));
 sg13g2_buf_8 fanout6852 (.A(net6853),
    .X(net6852));
 sg13g2_buf_8 fanout6853 (.A(net6864),
    .X(net6853));
 sg13g2_buf_8 fanout6854 (.A(net6855),
    .X(net6854));
 sg13g2_buf_8 fanout6855 (.A(net6857),
    .X(net6855));
 sg13g2_buf_8 fanout6856 (.A(net6857),
    .X(net6856));
 sg13g2_buf_8 fanout6857 (.A(net6864),
    .X(net6857));
 sg13g2_buf_8 fanout6858 (.A(net6859),
    .X(net6858));
 sg13g2_buf_8 fanout6859 (.A(net6864),
    .X(net6859));
 sg13g2_buf_8 fanout6860 (.A(net6863),
    .X(net6860));
 sg13g2_buf_8 fanout6861 (.A(net6863),
    .X(net6861));
 sg13g2_buf_8 fanout6862 (.A(net6863),
    .X(net6862));
 sg13g2_buf_8 fanout6863 (.A(net6864),
    .X(net6863));
 sg13g2_buf_8 fanout6864 (.A(net6985),
    .X(net6864));
 sg13g2_buf_8 fanout6865 (.A(net6868),
    .X(net6865));
 sg13g2_buf_8 fanout6866 (.A(net6868),
    .X(net6866));
 sg13g2_buf_8 fanout6867 (.A(net6868),
    .X(net6867));
 sg13g2_buf_8 fanout6868 (.A(net6881),
    .X(net6868));
 sg13g2_buf_8 fanout6869 (.A(net6871),
    .X(net6869));
 sg13g2_buf_8 fanout6870 (.A(net6871),
    .X(net6870));
 sg13g2_buf_8 fanout6871 (.A(net6873),
    .X(net6871));
 sg13g2_buf_8 fanout6872 (.A(net6873),
    .X(net6872));
 sg13g2_buf_8 fanout6873 (.A(net6881),
    .X(net6873));
 sg13g2_buf_8 fanout6874 (.A(net6877),
    .X(net6874));
 sg13g2_buf_2 fanout6875 (.A(net6877),
    .X(net6875));
 sg13g2_buf_8 fanout6876 (.A(net6877),
    .X(net6876));
 sg13g2_buf_8 fanout6877 (.A(net6881),
    .X(net6877));
 sg13g2_buf_8 fanout6878 (.A(net6880),
    .X(net6878));
 sg13g2_buf_8 fanout6879 (.A(net6880),
    .X(net6879));
 sg13g2_buf_8 fanout6880 (.A(net6881),
    .X(net6880));
 sg13g2_buf_8 fanout6881 (.A(net6985),
    .X(net6881));
 sg13g2_buf_8 fanout6882 (.A(net6883),
    .X(net6882));
 sg13g2_buf_8 fanout6883 (.A(net6886),
    .X(net6883));
 sg13g2_buf_8 fanout6884 (.A(net6886),
    .X(net6884));
 sg13g2_buf_8 fanout6885 (.A(net6886),
    .X(net6885));
 sg13g2_buf_8 fanout6886 (.A(net6897),
    .X(net6886));
 sg13g2_buf_8 fanout6887 (.A(net6888),
    .X(net6887));
 sg13g2_buf_8 fanout6888 (.A(net6889),
    .X(net6888));
 sg13g2_buf_8 fanout6889 (.A(net6897),
    .X(net6889));
 sg13g2_buf_8 fanout6890 (.A(net6897),
    .X(net6890));
 sg13g2_buf_8 fanout6891 (.A(net6892),
    .X(net6891));
 sg13g2_buf_8 fanout6892 (.A(net6897),
    .X(net6892));
 sg13g2_buf_8 fanout6893 (.A(net6896),
    .X(net6893));
 sg13g2_buf_8 fanout6894 (.A(net6896),
    .X(net6894));
 sg13g2_buf_1 fanout6895 (.A(net6896),
    .X(net6895));
 sg13g2_buf_8 fanout6896 (.A(net6897),
    .X(net6896));
 sg13g2_buf_8 fanout6897 (.A(net6915),
    .X(net6897));
 sg13g2_buf_8 fanout6898 (.A(net6900),
    .X(net6898));
 sg13g2_buf_8 fanout6899 (.A(net6900),
    .X(net6899));
 sg13g2_buf_8 fanout6900 (.A(net6915),
    .X(net6900));
 sg13g2_buf_8 fanout6901 (.A(net6904),
    .X(net6901));
 sg13g2_buf_8 fanout6902 (.A(net6903),
    .X(net6902));
 sg13g2_buf_8 fanout6903 (.A(net6904),
    .X(net6903));
 sg13g2_buf_8 fanout6904 (.A(net6915),
    .X(net6904));
 sg13g2_buf_8 fanout6905 (.A(net6906),
    .X(net6905));
 sg13g2_buf_8 fanout6906 (.A(net6914),
    .X(net6906));
 sg13g2_buf_8 fanout6907 (.A(net6908),
    .X(net6907));
 sg13g2_buf_8 fanout6908 (.A(net6914),
    .X(net6908));
 sg13g2_buf_8 fanout6909 (.A(net6913),
    .X(net6909));
 sg13g2_buf_2 fanout6910 (.A(net6913),
    .X(net6910));
 sg13g2_buf_8 fanout6911 (.A(net6912),
    .X(net6911));
 sg13g2_buf_8 fanout6912 (.A(net6913),
    .X(net6912));
 sg13g2_buf_8 fanout6913 (.A(net6914),
    .X(net6913));
 sg13g2_buf_8 fanout6914 (.A(net6915),
    .X(net6914));
 sg13g2_buf_8 fanout6915 (.A(net6985),
    .X(net6915));
 sg13g2_buf_8 fanout6916 (.A(net6917),
    .X(net6916));
 sg13g2_buf_8 fanout6917 (.A(net6919),
    .X(net6917));
 sg13g2_buf_8 fanout6918 (.A(net6919),
    .X(net6918));
 sg13g2_buf_8 fanout6919 (.A(net6951),
    .X(net6919));
 sg13g2_buf_8 fanout6920 (.A(net6923),
    .X(net6920));
 sg13g2_buf_1 fanout6921 (.A(net6923),
    .X(net6921));
 sg13g2_buf_8 fanout6922 (.A(net6923),
    .X(net6922));
 sg13g2_buf_8 fanout6923 (.A(net6951),
    .X(net6923));
 sg13g2_buf_8 fanout6924 (.A(net6930),
    .X(net6924));
 sg13g2_buf_8 fanout6925 (.A(net6930),
    .X(net6925));
 sg13g2_buf_8 fanout6926 (.A(net6927),
    .X(net6926));
 sg13g2_buf_8 fanout6927 (.A(net6930),
    .X(net6927));
 sg13g2_buf_8 fanout6928 (.A(net6929),
    .X(net6928));
 sg13g2_buf_8 fanout6929 (.A(net6930),
    .X(net6929));
 sg13g2_buf_8 fanout6930 (.A(net6951),
    .X(net6930));
 sg13g2_buf_8 fanout6931 (.A(net6932),
    .X(net6931));
 sg13g2_buf_8 fanout6932 (.A(net6940),
    .X(net6932));
 sg13g2_buf_8 fanout6933 (.A(net6934),
    .X(net6933));
 sg13g2_buf_8 fanout6934 (.A(net6940),
    .X(net6934));
 sg13g2_buf_8 fanout6935 (.A(net6936),
    .X(net6935));
 sg13g2_buf_8 fanout6936 (.A(net6939),
    .X(net6936));
 sg13g2_buf_8 fanout6937 (.A(net6939),
    .X(net6937));
 sg13g2_buf_2 fanout6938 (.A(net6939),
    .X(net6938));
 sg13g2_buf_8 fanout6939 (.A(net6940),
    .X(net6939));
 sg13g2_buf_8 fanout6940 (.A(net6951),
    .X(net6940));
 sg13g2_buf_8 fanout6941 (.A(net6942),
    .X(net6941));
 sg13g2_buf_8 fanout6942 (.A(net6945),
    .X(net6942));
 sg13g2_buf_8 fanout6943 (.A(net6945),
    .X(net6943));
 sg13g2_buf_8 fanout6944 (.A(net6945),
    .X(net6944));
 sg13g2_buf_8 fanout6945 (.A(net6951),
    .X(net6945));
 sg13g2_buf_8 fanout6946 (.A(net6947),
    .X(net6946));
 sg13g2_buf_8 fanout6947 (.A(net6950),
    .X(net6947));
 sg13g2_buf_8 fanout6948 (.A(net6949),
    .X(net6948));
 sg13g2_buf_8 fanout6949 (.A(net6950),
    .X(net6949));
 sg13g2_buf_8 fanout6950 (.A(net6951),
    .X(net6950));
 sg13g2_buf_8 fanout6951 (.A(net6985),
    .X(net6951));
 sg13g2_buf_8 fanout6952 (.A(net6953),
    .X(net6952));
 sg13g2_buf_8 fanout6953 (.A(net6956),
    .X(net6953));
 sg13g2_buf_8 fanout6954 (.A(net6955),
    .X(net6954));
 sg13g2_buf_8 fanout6955 (.A(net6956),
    .X(net6955));
 sg13g2_buf_8 fanout6956 (.A(net6964),
    .X(net6956));
 sg13g2_buf_8 fanout6957 (.A(net6958),
    .X(net6957));
 sg13g2_buf_8 fanout6958 (.A(net6964),
    .X(net6958));
 sg13g2_buf_8 fanout6959 (.A(net6960),
    .X(net6959));
 sg13g2_buf_8 fanout6960 (.A(net6964),
    .X(net6960));
 sg13g2_buf_8 fanout6961 (.A(net6963),
    .X(net6961));
 sg13g2_buf_1 fanout6962 (.A(net6963),
    .X(net6962));
 sg13g2_buf_8 fanout6963 (.A(net6964),
    .X(net6963));
 sg13g2_buf_8 fanout6964 (.A(net6984),
    .X(net6964));
 sg13g2_buf_8 fanout6965 (.A(net6973),
    .X(net6965));
 sg13g2_buf_8 fanout6966 (.A(net6973),
    .X(net6966));
 sg13g2_buf_8 fanout6967 (.A(net6968),
    .X(net6967));
 sg13g2_buf_8 fanout6968 (.A(net6973),
    .X(net6968));
 sg13g2_buf_8 fanout6969 (.A(net6970),
    .X(net6969));
 sg13g2_buf_8 fanout6970 (.A(net6973),
    .X(net6970));
 sg13g2_buf_8 fanout6971 (.A(net6972),
    .X(net6971));
 sg13g2_buf_8 fanout6972 (.A(net6973),
    .X(net6972));
 sg13g2_buf_8 fanout6973 (.A(net6984),
    .X(net6973));
 sg13g2_buf_8 fanout6974 (.A(net6977),
    .X(net6974));
 sg13g2_buf_8 fanout6975 (.A(net6976),
    .X(net6975));
 sg13g2_buf_8 fanout6976 (.A(net6977),
    .X(net6976));
 sg13g2_buf_8 fanout6977 (.A(net6984),
    .X(net6977));
 sg13g2_buf_8 fanout6978 (.A(net6983),
    .X(net6978));
 sg13g2_buf_2 fanout6979 (.A(net6983),
    .X(net6979));
 sg13g2_buf_8 fanout6980 (.A(net6983),
    .X(net6980));
 sg13g2_buf_1 fanout6981 (.A(net6982),
    .X(net6981));
 sg13g2_buf_8 fanout6982 (.A(net6983),
    .X(net6982));
 sg13g2_buf_8 fanout6983 (.A(net6984),
    .X(net6983));
 sg13g2_buf_8 fanout6984 (.A(net6985),
    .X(net6984));
 sg13g2_buf_8 fanout6985 (.A(net6986),
    .X(net6985));
 sg13g2_buf_8 fanout6986 (.A(rst_n),
    .X(net6986));
 sg13g2_buf_8 fanout6987 (.A(_08135_),
    .X(net6987));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tiehi _26004__14 (.L_HI(net14));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_8 clkbuf_leaf_314_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_8 clkbuf_leaf_315_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_8 clkbuf_leaf_316_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_8 clkbuf_leaf_317_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_8 clkbuf_6_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_8 clkbuf_6_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkbuf_6_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkbuf_6_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkbuf_6_4__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkbuf_6_5__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkbuf_6_6__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkbuf_6_7__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkbuf_6_8__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_8 clkbuf_6_9__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkbuf_6_10__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkbuf_6_11__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkbuf_6_12__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkbuf_6_13__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkbuf_6_14__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkbuf_6_15__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkbuf_6_16__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_8 clkbuf_6_17__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkbuf_6_18__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkbuf_6_19__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkbuf_6_20__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkbuf_6_21__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkbuf_6_22__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkbuf_6_23__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkbuf_6_24__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_8 clkbuf_6_25__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkbuf_6_26__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkbuf_6_27__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkbuf_6_28__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkbuf_6_29__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkbuf_6_30__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkbuf_6_31__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkbuf_6_32__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_8 clkbuf_6_33__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkbuf_6_34__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkbuf_6_35__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkbuf_6_36__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkbuf_6_37__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkbuf_6_38__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkbuf_6_39__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkbuf_6_40__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_8 clkbuf_6_41__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkbuf_6_42__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkbuf_6_43__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkbuf_6_44__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkbuf_6_45__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkbuf_6_46__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkbuf_6_47__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkbuf_6_48__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_8 clkbuf_6_49__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkbuf_6_50__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkbuf_6_51__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkbuf_6_52__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkbuf_6_53__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkbuf_6_54__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkbuf_6_55__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkbuf_6_56__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_8 clkbuf_6_57__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkbuf_6_58__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkbuf_6_59__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkbuf_6_60__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_8 clkbuf_6_61__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkbuf_6_62__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkbuf_6_63__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_317_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_121_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\soc_inst.cpu_core.csr_file.timer_interrupt ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold2 (.A(\soc_inst.gpio_inst.gpio_sync1[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold3 (.A(\soc_inst.i2c_inst.transfer_done ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold4 (.A(\soc_inst.gpio_inst.gpio_sync1[2] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold5 (.A(\soc_inst.gpio_inst.gpio_sync1[5] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold6 (.A(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d1 ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold7 (.A(\soc_inst.gpio_inst.gpio_sync1[6] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold8 (.A(\soc_inst.gpio_inst.gpio_sync1[4] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold9 (.A(\soc_inst.gpio_inst.gpio_sync1[3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold10 (.A(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold11 (.A(\soc_inst.i2c_inst.arb_lost ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold12 (.A(\soc_inst.mem_ctrl.spi_mem_inst.sample_trigger_d2 ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold13 (.A(\soc_inst.i2c_inst.ack_received ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold14 (.A(\soc_inst.gpio_inst.gpio_sync1[0] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold15 (.A(\soc_inst.cpu_core.csr_file.external_interrupt ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold16 (.A(\soc_inst.bus_spi_sclk ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold17 (.A(_00110_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold18 (.A(\soc_inst.mem_ctrl.spi_mem_inst.is_write_op ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold19 (.A(_08666_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold20 (.A(\soc_inst.cpu_core.csr_file.mcause[4] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold21 (.A(\soc_inst.cpu_core.csr_file.mcause[27] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold22 (.A(\soc_inst.cpu_core.csr_file.mcause[18] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold23 (.A(\soc_inst.cpu_core.csr_file.mcause[26] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold24 (.A(\soc_inst.cpu_core.csr_file.mcause[25] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold25 (.A(\soc_inst.cpu_core.csr_file.mcause[29] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold26 (.A(\soc_inst.cpu_core.csr_file.mcause[16] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold27 (.A(\soc_inst.cpu_core.csr_file.mcause[15] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold28 (.A(\soc_inst.cpu_core.csr_file.mcause[11] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold29 (.A(\soc_inst.cpu_core.csr_file.mcause[17] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold30 (.A(\soc_inst.cpu_core.csr_file.mcause[12] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold31 (.A(\soc_inst.cpu_core.csr_file.mcause[21] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold32 (.A(_00232_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold33 (.A(_09442_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold34 (.A(_00392_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold35 (.A(\soc_inst.cpu_core.csr_file.mcause[7] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold36 (.A(\soc_inst.cpu_core.csr_file.mcause[28] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold37 (.A(\soc_inst.cpu_core.csr_file.mcause[5] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold38 (.A(\soc_inst.cpu_core.csr_file.mcause[23] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold39 (.A(\soc_inst.cpu_core.csr_file.mstatus[19] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold40 (.A(\soc_inst.cpu_core.csr_file.mcause[24] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold41 (.A(\soc_inst.cpu_core.csr_file.mcause[8] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold42 (.A(\soc_inst.cpu_core.csr_file.mcause[14] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold43 (.A(\soc_inst.cpu_core.csr_file.mcause[9] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold44 (.A(\soc_inst.cpu_core.csr_file.mcause[22] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold45 (.A(\soc_inst.cpu_core.csr_file.mstatus[17] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold46 (.A(\soc_inst.cpu_core.csr_file.mstatus[18] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold47 (.A(\soc_inst.cpu_core.csr_file.mscratch[15] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold48 (.A(_11164_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold49 (.A(_00796_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold50 (.A(\soc_inst.cpu_core.csr_file.mcause[30] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold51 (.A(\soc_inst.cpu_core.csr_file.mcause[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold52 (.A(\soc_inst.cpu_core.csr_file.mscratch[9] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold53 (.A(_11143_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold54 (.A(_00790_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold55 (.A(\soc_inst.cpu_core.csr_file.mscratch[10] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold56 (.A(_11145_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold57 (.A(_00791_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold58 (.A(\soc_inst.cpu_core.csr_file.mscratch[12] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold59 (.A(_11152_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00793_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold61 (.A(\soc_inst.cpu_core.csr_file.mscratch[6] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold62 (.A(_11135_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold63 (.A(_00787_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold64 (.A(\soc_inst.cpu_core.csr_file.mstatus[27] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold65 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[11] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold66 (.A(_00685_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold67 (.A(\soc_inst.cpu_core.csr_file.mstatus[25] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold68 (.A(\soc_inst.cpu_core.csr_file.mcause[10] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold69 (.A(\soc_inst.cpu_core.csr_file.mscratch[18] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold70 (.A(_11176_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold71 (.A(_00799_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold72 (.A(\soc_inst.cpu_core.csr_file.mstatus[29] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold73 (.A(\soc_inst.cpu_core.csr_file.mcause[13] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold74 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[28] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00714_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold76 (.A(\soc_inst.spi_inst.tx_shift_reg[4] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00165_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold78 (.A(\soc_inst.cpu_core.csr_file.mcause[19] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold79 (.A(\soc_inst.spi_inst.tx_shift_reg[12] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold80 (.A(_00142_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold81 (.A(\soc_inst.core_mem_wdata[17] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold82 (.A(_02517_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold83 (.A(\soc_inst.cpu_core.csr_file.mscratch[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold84 (.A(\soc_inst.spi_inst.tx_shift_reg[8] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00169_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold86 (.A(\soc_inst.mem_ctrl.spi_data_in[31] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold87 (.A(_00509_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold88 (.A(\soc_inst.spi_inst.clk_counter[0] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00128_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold90 (.A(\soc_inst.cpu_core.csr_file.mscratch[20] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold91 (.A(_11184_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold92 (.A(_00801_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold93 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold94 (.A(_02533_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold95 (.A(\soc_inst.spi_inst.tx_shift_reg[7] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00168_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold97 (.A(\soc_inst.cpu_core.csr_file.mscratch[22] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold98 (.A(_11192_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold99 (.A(_00803_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold100 (.A(\soc_inst.cpu_core.csr_file.mstatus[28] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold101 (.A(\soc_inst.cpu_core.csr_file.mstatus[31] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold102 (.A(\soc_inst.mem_ctrl.spi_data_in[30] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold103 (.A(_00508_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold104 (.A(\soc_inst.spi_inst.start_pending ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold105 (.A(_09234_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold106 (.A(\soc_inst.spi_inst.next_state[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold107 (.A(\soc_inst.cpu_core.csr_file.mcause[20] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold108 (.A(\soc_inst.spi_inst.tx_shift_reg[0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold109 (.A(_00149_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold110 (.A(\soc_inst.spi_inst.tx_shift_reg[1] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold111 (.A(_00160_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold112 (.A(\soc_inst.cpu_core.csr_file.mscratch[19] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold113 (.A(_11180_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00800_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold115 (.A(\soc_inst.cpu_core.csr_file.mscratch[7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold116 (.A(_11138_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00788_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold118 (.A(\soc_inst.cpu_core.csr_file.mscratch[21] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold119 (.A(_11188_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold120 (.A(_00802_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold121 (.A(\soc_inst.spi_inst.tx_shift_reg[18] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00148_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold123 (.A(\soc_inst.mem_ctrl.spi_data_in[26] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold124 (.A(_00504_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold125 (.A(\soc_inst.spi_inst.tx_shift_reg[14] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold126 (.A(_00144_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold127 (.A(\soc_inst.cpu_core.ex_rs1_data[9] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold128 (.A(_01259_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold129 (.A(\soc_inst.cpu_core.ex_rs2_data[26] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold130 (.A(_01340_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold131 (.A(\soc_inst.spi_inst.tx_shift_reg[24] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold132 (.A(_00155_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold133 (.A(\soc_inst.core_mem_wdata[3] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold134 (.A(_02449_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold135 (.A(\soc_inst.cpu_core.ex_rs1_data[26] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold136 (.A(_01276_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold137 (.A(\soc_inst.i2c_inst.clk_cnt[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold138 (.A(\soc_inst.cpu_core.ex_rs1_data[17] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold139 (.A(_01267_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold140 (.A(\soc_inst.core_mem_wdata[9] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold141 (.A(_02509_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold142 (.A(\soc_inst.cpu_core.csr_file.mstatus[20] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold143 (.A(\soc_inst.cpu_core.csr_file.mscratch[8] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold144 (.A(_11141_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold145 (.A(_00789_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold146 (.A(\soc_inst.core_mem_wdata[16] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold147 (.A(_02516_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold148 (.A(\soc_inst.mem_ctrl.spi_mem_inst.ram_in_quad_mode ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold149 (.A(_00002_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold150 (.A(\soc_inst.spi_inst.tx_shift_reg[27] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold151 (.A(_00158_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold152 (.A(\soc_inst.cpu_core.ex_rs1_data[12] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold153 (.A(_01262_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold154 (.A(\soc_inst.core_mem_wdata[25] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold155 (.A(_02525_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold156 (.A(\soc_inst.cpu_core.csr_file.mscratch[14] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold157 (.A(_11160_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold158 (.A(_00795_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold159 (.A(\soc_inst.cpu_core.ex_rs2_data[13] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold160 (.A(_04532_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold161 (.A(_01327_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold162 (.A(\soc_inst.i2c_inst.ctrl_reg[2] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold163 (.A(_00515_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold164 (.A(\soc_inst.cpu_core.ex_rs1_data[10] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold165 (.A(_01260_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold166 (.A(\soc_inst.core_mem_wdata[4] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold167 (.A(_02448_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold168 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[29] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold169 (.A(_00715_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold170 (.A(\soc_inst.spi_inst.tx_shift_reg[23] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold171 (.A(_00154_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold172 (.A(\soc_inst.cpu_core.ex_rs2_data[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold173 (.A(_01318_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold174 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[4] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold175 (.A(_00678_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold176 (.A(\soc_inst.cpu_core.ex_rs2_data[8] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold177 (.A(_01322_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold178 (.A(\soc_inst.cpu_core.ex_rs1_data[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold179 (.A(_01254_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold180 (.A(\soc_inst.cpu_core.csr_file.mstatus[26] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold181 (.A(\soc_inst.cpu_core.ex_rs1_data[8] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold182 (.A(_01258_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold183 (.A(\soc_inst.spi_inst.tx_shift_reg[29] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold184 (.A(_00161_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold185 (.A(\soc_inst.pwm_inst.channel_counter[0][0] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold186 (.A(\soc_inst.cpu_core.csr_file.mstatus[23] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold187 (.A(\soc_inst.mem_ctrl.spi_data_in[7] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00485_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold189 (.A(\soc_inst.core_mem_wdata[24] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold190 (.A(_02524_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold191 (.A(\soc_inst.cpu_core.csr_file.mscratch[5] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold192 (.A(_11131_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold193 (.A(_00786_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold194 (.A(\soc_inst.cpu_core.ex_rs2_data[23] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold195 (.A(_01337_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold196 (.A(\soc_inst.cpu_core.ex_rs1_data[16] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold197 (.A(_01266_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold198 (.A(\soc_inst.cpu_core.csr_file.mscratch[23] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold199 (.A(_11196_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold200 (.A(_00804_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold201 (.A(\soc_inst.cpu_core.csr_file.mscratch[11] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold202 (.A(_11148_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold203 (.A(_00792_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold204 (.A(\soc_inst.cpu_core.csr_file.mscratch[16] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold205 (.A(_11168_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold206 (.A(_00797_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold207 (.A(\soc_inst.spi_inst.tx_shift_reg[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00164_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold209 (.A(\soc_inst.cpu_core.ex_rs1_data[13] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold210 (.A(_01263_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold211 (.A(\soc_inst.gpio_inst.int_pend_reg[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold212 (.A(_07588_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold213 (.A(_02451_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold214 (.A(\soc_inst.cpu_core.ex_rs2_data[10] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold215 (.A(_01324_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold216 (.A(\soc_inst.core_mem_wdata[19] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold217 (.A(_02519_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold218 (.A(\soc_inst.cpu_core.ex_rs2_data[6] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold219 (.A(_01320_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold220 (.A(\soc_inst.cpu_core.ex_rs2_data[1] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00842_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold222 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[31] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold223 (.A(_00717_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold224 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_sample ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold225 (.A(_02581_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold226 (.A(\soc_inst.mem_ctrl.spi_data_in[24] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold227 (.A(_00502_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold228 (.A(\soc_inst.spi_inst.tx_shift_reg[17] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold229 (.A(_00147_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold230 (.A(\soc_inst.mem_ctrl.spi_data_in[18] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold231 (.A(_00496_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold232 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[8] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold233 (.A(_00674_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold234 (.A(\soc_inst.core_mem_wdata[29] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold235 (.A(_02529_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold236 (.A(\soc_inst.core_mem_rdata[5] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold237 (.A(\soc_inst.cpu_core.ex_rs1_data[3] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold238 (.A(_01253_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold239 (.A(\soc_inst.mem_ctrl.spi_data_in[2] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold240 (.A(_00480_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold241 (.A(\soc_inst.cpu_core.ex_rs1_data[27] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold242 (.A(_01277_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold243 (.A(\soc_inst.cpu_core.csr_file.mstatus[24] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold244 (.A(\soc_inst.spi_inst.tx_shift_reg[16] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold245 (.A(\soc_inst.cpu_core.ex_rs2_data[16] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold246 (.A(_01330_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold247 (.A(\soc_inst.cpu_core.ex_rs1_data[11] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold248 (.A(_01261_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold249 (.A(\soc_inst.cpu_core.ex_rs1_data[28] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold250 (.A(_01278_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold251 (.A(\soc_inst.spi_inst.tx_shift_reg[6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold252 (.A(_00167_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold253 (.A(\soc_inst.mem_ctrl.spi_data_in[27] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold254 (.A(_00505_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold255 (.A(\soc_inst.cpu_core.csr_file.mstatus[16] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold256 (.A(\soc_inst.cpu_core.ex_rs2_data[14] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold257 (.A(_04533_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold258 (.A(_01328_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold259 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[7] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold260 (.A(_00681_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold261 (.A(\soc_inst.cpu_core.csr_file.mstatus[22] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold262 (.A(\soc_inst.mem_ctrl.spi_data_in[1] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold263 (.A(\soc_inst.mem_ctrl.spi_data_in[23] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold264 (.A(_00501_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold265 (.A(\soc_inst.cpu_core.csr_file.mtvec[20] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold266 (.A(_07429_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold267 (.A(_02418_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold268 (.A(\soc_inst.cpu_core.ex_rs2_data[24] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold269 (.A(_01338_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold270 (.A(\soc_inst.cpu_core.csr_file.mstatus[21] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold271 (.A(\soc_inst.mem_ctrl.spi_data_in[29] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold272 (.A(_00507_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold273 (.A(\soc_inst.mem_ctrl.spi_data_in[16] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold274 (.A(_00494_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold275 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[8] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold276 (.A(_00682_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold277 (.A(\soc_inst.mem_ctrl.spi_data_in[28] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold278 (.A(_00506_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold279 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold280 (.A(_00677_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold281 (.A(\soc_inst.cpu_core.id_instr[15] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold282 (.A(_01209_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold283 (.A(\soc_inst.cpu_core.register_file.registers[15][21] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold284 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00676_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold286 (.A(\soc_inst.spi_inst.tx_shift_reg[30] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00162_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold288 (.A(\soc_inst.cpu_core.ex_rs1_data[14] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold289 (.A(_01264_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold290 (.A(\soc_inst.core_mem_wdata[28] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold291 (.A(_02528_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold292 (.A(\soc_inst.cpu_core.csr_file.mstatus[30] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold293 (.A(\soc_inst.cpu_core.register_file.registers[18][24] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold294 (.A(\soc_inst.cpu_core.csr_file.mstatus[14] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold295 (.A(\soc_inst.cpu_core.ex_rs1_data[30] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold296 (.A(_01280_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold297 (.A(\soc_inst.mem_ctrl.spi_data_in[17] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold298 (.A(\soc_inst.cpu_core.ex_rs2_data[0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00841_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold300 (.A(\soc_inst.mem_ctrl.spi_data_in[19] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00497_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold302 (.A(\soc_inst.cpu_core.ex_rs1_data[31] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold303 (.A(_01281_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold304 (.A(\soc_inst.mem_ctrl.spi_data_in[25] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold305 (.A(_00503_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold306 (.A(\soc_inst.cpu_core.csr_file.mscratch[27] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold307 (.A(_00808_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold308 (.A(\soc_inst.cpu_core.register_file.registers[13][31] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold309 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[10] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00684_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold311 (.A(\soc_inst.cpu_core.register_file.registers[1][23] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold312 (.A(\soc_inst.cpu_core.csr_file.mstatus[15] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold313 (.A(\soc_inst.cpu_core.register_file.registers[1][19] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold314 (.A(\soc_inst.cpu_core.register_file.registers[2][12] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold315 (.A(\soc_inst.cpu_core.ex_rs1_data[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold316 (.A(_01251_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold317 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[14] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold318 (.A(_00733_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold319 (.A(\soc_inst.cpu_core.ex_rs2_data[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold320 (.A(_01317_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold321 (.A(\soc_inst.cpu_core.csr_file.mtime[7] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold322 (.A(_00218_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold323 (.A(\soc_inst.cpu_core.register_file.registers[8][17] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold324 (.A(\soc_inst.core_mem_addr[31] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold325 (.A(_01313_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold326 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[13] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00001_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold328 (.A(\soc_inst.gpio_inst.int_pend_reg[5] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold329 (.A(_07580_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold330 (.A(_02447_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold331 (.A(\soc_inst.cpu_core.register_file.registers[17][6] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold332 (.A(\soc_inst.cpu_core.register_file.registers[16][20] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold333 (.A(\soc_inst.cpu_core.register_file.registers[24][11] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold334 (.A(\soc_inst.spi_inst.tx_shift_reg[10] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold335 (.A(_00140_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold336 (.A(\soc_inst.mem_ctrl.spi_data_in[5] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold337 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[13] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold338 (.A(_00732_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold339 (.A(\soc_inst.mem_ctrl.spi_data_in[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold340 (.A(_00484_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold341 (.A(\soc_inst.cpu_core.register_file.registers[20][20] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold342 (.A(\soc_inst.cpu_core.i_mem_ready ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold343 (.A(\soc_inst.cpu_core.register_file.registers[14][0] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold344 (.A(\soc_inst.cpu_core.csr_file.mscratch[13] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold345 (.A(_11156_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold346 (.A(_00794_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold347 (.A(\soc_inst.cpu_core.ex_rs2_data[31] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold348 (.A(_01345_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold349 (.A(\soc_inst.gpio_inst.int_pend_reg[2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold350 (.A(_07586_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold351 (.A(_02450_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold352 (.A(\soc_inst.mem_ctrl.spi_data_in[21] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold353 (.A(_00499_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold354 (.A(\soc_inst.cpu_core.register_file.registers[2][22] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold355 (.A(\soc_inst.cpu_core.register_file.registers[11][22] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold356 (.A(\soc_inst.cpu_core.register_file.registers[2][27] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold357 (.A(\soc_inst.mem_ctrl.spi_mem_inst.flash_in_cont_mode ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold358 (.A(_08664_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00012_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold360 (.A(\soc_inst.cpu_core.register_file.registers[24][10] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold361 (.A(\soc_inst.cpu_core.csr_file.mstatus[8] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold362 (.A(_09906_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00512_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold364 (.A(\soc_inst.cpu_core.register_file.registers[20][7] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold365 (.A(\soc_inst.cpu_core.register_file.registers[1][4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold366 (.A(\soc_inst.gpio_bidir_out [0]),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold367 (.A(_00460_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold368 (.A(\soc_inst.cpu_core.register_file.registers[14][9] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold369 (.A(\soc_inst.cpu_core.register_file.registers[8][9] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold370 (.A(\soc_inst.cpu_core.register_file.registers[13][26] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold371 (.A(\soc_inst.cpu_core.register_file.registers[16][7] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold372 (.A(\soc_inst.cpu_core.register_file.registers[20][28] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold373 (.A(\soc_inst.cpu_core.register_file.registers[2][3] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold374 (.A(\soc_inst.cpu_core.register_file.registers[4][26] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold375 (.A(\soc_inst.cpu_core.register_file.registers[2][8] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold376 (.A(\soc_inst.cpu_core.ex_rs1_data[6] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold377 (.A(_01256_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold378 (.A(\soc_inst.spi_inst.rx_shift_reg[31] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold379 (.A(_09422_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold380 (.A(\soc_inst.cpu_core.register_file.registers[20][9] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold381 (.A(\soc_inst.cpu_core.register_file.registers[16][17] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold382 (.A(\soc_inst.cpu_core.register_file.registers[2][7] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold383 (.A(\soc_inst.spi_inst.clk_counter[7] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold384 (.A(_00135_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold385 (.A(\soc_inst.cpu_core.csr_file.mtvec[18] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold386 (.A(_07427_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold387 (.A(_02416_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold388 (.A(\soc_inst.cpu_core.register_file.registers[8][7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold389 (.A(\soc_inst.mem_ctrl.next_instr_data[3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00643_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold391 (.A(\soc_inst.cpu_core.register_file.registers[24][27] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold392 (.A(\soc_inst.cpu_core.register_file.registers[11][26] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold393 (.A(\soc_inst.cpu_core.ex_rs2_data[27] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold394 (.A(_01341_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold395 (.A(\soc_inst.cpu_core.register_file.registers[15][17] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold396 (.A(\soc_inst.cpu_core.register_file.registers[24][24] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold397 (.A(\soc_inst.cpu_core.csr_file.mstatus[10] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold398 (.A(_09914_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold399 (.A(_00514_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold400 (.A(\soc_inst.cpu_core.register_file.registers[1][12] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold401 (.A(\soc_inst.cpu_core.register_file.registers[15][3] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold402 (.A(\soc_inst.cpu_core.register_file.registers[8][30] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold403 (.A(\soc_inst.cpu_core.csr_file.mscratch[29] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold404 (.A(_00810_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold405 (.A(\soc_inst.cpu_core.register_file.registers[1][28] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold406 (.A(\soc_inst.cpu_core.register_file.registers[15][11] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold407 (.A(\soc_inst.mem_ctrl.next_instr_data[28] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00668_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold409 (.A(\soc_inst.cpu_core.register_file.registers[1][8] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold410 (.A(\soc_inst.cpu_core.register_file.registers[11][7] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold411 (.A(\soc_inst.cpu_core.register_file.registers[11][29] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold412 (.A(\soc_inst.cpu_core.register_file.registers[13][2] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold413 (.A(\soc_inst.cpu_core.register_file.registers[4][24] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold414 (.A(\soc_inst.cpu_core.register_file.registers[20][0] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold415 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[7] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold416 (.A(_07676_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold417 (.A(_02540_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold418 (.A(\soc_inst.mem_ctrl.next_instr_data[22] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold419 (.A(_00662_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold420 (.A(\soc_inst.cpu_core.register_file.registers[13][27] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold421 (.A(\soc_inst.cpu_core.csr_file.mtvec[8] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold422 (.A(_07417_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold423 (.A(_02406_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold424 (.A(\soc_inst.cpu_core.csr_file.mtvec[15] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold425 (.A(_07424_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold426 (.A(_02413_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold427 (.A(\soc_inst.cpu_core.register_file.registers[24][7] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold428 (.A(\soc_inst.cpu_core.register_file.registers[1][2] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold429 (.A(\soc_inst.cpu_core.register_file.registers[4][31] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold430 (.A(\soc_inst.cpu_core.register_file.registers[11][15] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold431 (.A(\soc_inst.cpu_core.ex_rs2_data[18] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold432 (.A(_01332_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold433 (.A(\soc_inst.cpu_core.register_file.registers[8][15] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold434 (.A(\soc_inst.cpu_core.register_file.registers[11][24] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold435 (.A(\soc_inst.cpu_core.register_file.registers[13][11] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold436 (.A(\soc_inst.cpu_core.csr_file.mstatus[13] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold437 (.A(\soc_inst.cpu_core.csr_file.mtvec[14] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold438 (.A(_07423_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold439 (.A(_02412_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold440 (.A(\soc_inst.cpu_core.ex_rs1_data[5] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold441 (.A(_01255_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold442 (.A(\soc_inst.cpu_core.register_file.registers[20][14] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold443 (.A(\soc_inst.cpu_core.ex_rs2_data[21] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold444 (.A(_01335_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold445 (.A(\soc_inst.cpu_core.ex_rs1_data[19] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold446 (.A(_01269_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold447 (.A(\soc_inst.cpu_core.register_file.registers[16][4] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold448 (.A(\soc_inst.cpu_core.register_file.registers[2][10] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold449 (.A(\soc_inst.cpu_core.register_file.registers[11][20] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold450 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[0] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold451 (.A(_02566_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold452 (.A(\soc_inst.cpu_core.register_file.registers[2][24] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold453 (.A(\soc_inst.cpu_core.register_file.registers[15][31] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold454 (.A(\soc_inst.cpu_core.register_file.registers[14][2] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold455 (.A(\soc_inst.cpu_core.register_file.registers[13][22] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold456 (.A(\soc_inst.cpu_core.csr_file.mtvec[11] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold457 (.A(_07420_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold458 (.A(_02409_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold459 (.A(\soc_inst.cpu_core.register_file.registers[15][29] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold460 (.A(\soc_inst.cpu_core.register_file.registers[18][22] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold461 (.A(\soc_inst.cpu_core.register_file.registers[20][31] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold462 (.A(\soc_inst.cpu_core.csr_file.mscratch[30] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold463 (.A(_00811_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold464 (.A(\soc_inst.cpu_core.register_file.registers[8][10] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold465 (.A(\soc_inst.cpu_core.register_file.registers[15][27] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold466 (.A(\soc_inst.cpu_core.register_file.registers[8][28] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold467 (.A(\soc_inst.cpu_core.register_file.registers[8][29] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold468 (.A(\soc_inst.cpu_core.register_file.registers[17][28] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold469 (.A(\soc_inst.core_mem_wdata[20] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold470 (.A(_02520_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold471 (.A(\soc_inst.cpu_core.register_file.registers[13][20] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold472 (.A(\soc_inst.mem_ctrl.next_instr_data[17] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold473 (.A(_00657_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold474 (.A(\soc_inst.cpu_core.csr_file.mscratch[26] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold475 (.A(_00807_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold476 (.A(\soc_inst.cpu_core.register_file.registers[1][31] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold477 (.A(\soc_inst.mem_ctrl.next_instr_data[26] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold478 (.A(_00666_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold479 (.A(\soc_inst.mem_ctrl.next_instr_data[8] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00648_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold481 (.A(\soc_inst.cpu_core.register_file.registers[2][15] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold482 (.A(\soc_inst.cpu_core.register_file.registers[24][26] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold483 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[6] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold484 (.A(_00680_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold485 (.A(\soc_inst.cpu_core.register_file.registers[4][12] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold486 (.A(\soc_inst.cpu_core.register_file.registers[18][0] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold487 (.A(\soc_inst.cpu_core.ex_rs2_data[17] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold488 (.A(_01331_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold489 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[10] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold490 (.A(_00729_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold491 (.A(\soc_inst.cpu_core.register_file.registers[15][5] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold492 (.A(\soc_inst.core_mem_wdata[21] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold493 (.A(_02521_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold494 (.A(\soc_inst.cpu_core.csr_file.mstatus[6] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold495 (.A(_09902_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold496 (.A(_00511_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold497 (.A(\soc_inst.cpu_core.register_file.registers[8][31] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold498 (.A(\soc_inst.spi_inst.clk_counter[1] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold499 (.A(_00129_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold500 (.A(\soc_inst.cpu_core.register_file.registers[15][14] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold501 (.A(\soc_inst.cpu_core.csr_file.mscratch[25] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold502 (.A(_00806_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold503 (.A(\soc_inst.cpu_core.register_file.registers[20][23] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold504 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[18] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00737_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold506 (.A(\soc_inst.cpu_core.register_file.registers[17][29] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold507 (.A(\soc_inst.cpu_core.ex_rs2_data[22] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold508 (.A(_01336_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold509 (.A(\soc_inst.cpu_core.register_file.registers[20][10] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold510 (.A(\soc_inst.cpu_core.register_file.registers[15][28] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold511 (.A(\soc_inst.mem_ctrl.spi_data_in[13] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold512 (.A(\soc_inst.cpu_core.register_file.registers[17][7] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold513 (.A(\soc_inst.cpu_core.register_file.registers[4][30] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold514 (.A(\soc_inst.cpu_core.register_file.registers[14][6] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold515 (.A(\soc_inst.i2c_inst.restart_pending ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold516 (.A(_11835_[0]),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold517 (.A(\soc_inst.spi_inst.tx_shift_reg[9] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold518 (.A(_00139_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold519 (.A(\soc_inst.cpu_core.register_file.registers[13][14] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold520 (.A(\soc_inst.cpu_core.register_file.registers[20][3] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold521 (.A(\soc_inst.cpu_core.register_file.registers[24][12] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold522 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[15] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold523 (.A(_00734_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold524 (.A(\soc_inst.cpu_core.ex_instr[20] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold525 (.A(_01044_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold526 (.A(\soc_inst.mem_ctrl.spi_data_in[0] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold527 (.A(\soc_inst.cpu_core.register_file.registers[18][15] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold528 (.A(\soc_inst.cpu_core.register_file.registers[4][15] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold529 (.A(\soc_inst.cpu_core.register_file.registers[24][14] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold530 (.A(\soc_inst.cpu_core.register_file.registers[8][24] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold531 (.A(\soc_inst.cpu_core.register_file.registers[15][15] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold532 (.A(\soc_inst.cpu_core.csr_file.mtvec[19] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold533 (.A(_07428_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold534 (.A(_02417_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold535 (.A(\soc_inst.cpu_core.register_file.registers[14][15] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold536 (.A(\soc_inst.mem_ctrl.next_instr_data[4] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold537 (.A(_00644_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold538 (.A(\soc_inst.cpu_core.register_file.registers[18][9] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold539 (.A(\soc_inst.cpu_core.register_file.registers[2][20] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold540 (.A(\soc_inst.cpu_core.csr_file.mstatus[5] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold541 (.A(_09897_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold542 (.A(_00510_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold543 (.A(\soc_inst.cpu_core.register_file.registers[2][9] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold544 (.A(\soc_inst.cpu_core.register_file.registers[20][24] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold545 (.A(\soc_inst.cpu_core.register_file.registers[18][10] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold546 (.A(\soc_inst.cpu_core.register_file.registers[24][2] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold547 (.A(\soc_inst.cpu_core.register_file.registers[14][21] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold548 (.A(\soc_inst.cpu_core.csr_file.mtime[44] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold549 (.A(_00211_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold550 (.A(\soc_inst.cpu_core.register_file.registers[17][17] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold551 (.A(\soc_inst.cpu_core.id_imm12[0] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold552 (.A(\soc_inst.cpu_core.register_file.registers[24][16] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold553 (.A(\soc_inst.cpu_core.register_file.registers[13][16] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold554 (.A(\soc_inst.cpu_core.register_file.registers[4][7] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold555 (.A(\soc_inst.cpu_core.register_file.registers[18][2] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold556 (.A(\soc_inst.cpu_core.register_file.registers[1][22] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold557 (.A(\soc_inst.cpu_core.register_file.registers[8][3] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold558 (.A(\soc_inst.cpu_core.register_file.registers[14][18] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold559 (.A(\soc_inst.cpu_core.ex_rs2_data[5] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold560 (.A(_01319_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold561 (.A(\soc_inst.cpu_core.register_file.registers[13][25] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold562 (.A(\soc_inst.cpu_core.register_file.registers[1][15] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold563 (.A(\soc_inst.mem_ctrl.next_instr_data[14] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold564 (.A(_00654_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold565 (.A(\soc_inst.cpu_core.ex_rs1_data[0] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold566 (.A(_01250_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold567 (.A(\soc_inst.cpu_core.register_file.registers[15][10] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold568 (.A(\soc_inst.cpu_core.register_file.registers[2][26] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold569 (.A(\soc_inst.cpu_core.register_file.registers[15][22] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold570 (.A(\soc_inst.cpu_core.register_file.registers[14][27] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold571 (.A(\soc_inst.cpu_core.register_file.registers[4][3] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold572 (.A(\soc_inst.cpu_core.register_file.registers[4][21] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold573 (.A(\soc_inst.cpu_core.register_file.registers[8][16] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold574 (.A(\soc_inst.cpu_core.register_file.registers[24][25] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold575 (.A(\soc_inst.cpu_core.register_file.registers[24][5] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold576 (.A(\soc_inst.mem_ctrl.next_instr_data[11] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold577 (.A(_00651_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold578 (.A(\soc_inst.cpu_core.register_file.registers[14][22] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold579 (.A(\soc_inst.cpu_core.register_file.registers[2][30] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold580 (.A(\soc_inst.cpu_core.register_file.registers[11][8] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold581 (.A(\soc_inst.cpu_core.register_file.registers[17][3] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold582 (.A(\soc_inst.mem_ctrl.next_instr_data[21] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold583 (.A(_00661_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold584 (.A(\soc_inst.mem_ctrl.next_instr_data[31] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold585 (.A(_00671_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold586 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[1] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold587 (.A(_07725_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold588 (.A(_02574_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold589 (.A(\soc_inst.cpu_core.register_file.registers[17][16] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold590 (.A(\soc_inst.cpu_core.register_file.registers[24][19] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold591 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[4] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold592 (.A(_02570_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold593 (.A(\soc_inst.cpu_core.register_file.registers[14][17] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold594 (.A(\soc_inst.cpu_core.register_file.registers[1][9] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold595 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[12] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold596 (.A(_00698_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold597 (.A(\soc_inst.cpu_core.register_file.registers[13][17] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold598 (.A(\soc_inst.cpu_core.register_file.registers[20][30] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold599 (.A(\soc_inst.cpu_core.register_file.registers[11][25] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold600 (.A(\soc_inst.cpu_core.register_file.registers[2][1] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold601 (.A(\soc_inst.mem_ctrl.next_instr_data[23] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold602 (.A(_00663_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold603 (.A(\soc_inst.cpu_core.register_file.registers[24][9] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold604 (.A(\soc_inst.core_mem_rdata[13] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold605 (.A(\soc_inst.cpu_core.register_file.registers[1][10] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold606 (.A(\soc_inst.cpu_core.register_file.registers[24][23] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold607 (.A(\soc_inst.cpu_core.register_file.registers[18][20] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold608 (.A(\soc_inst.cpu_core.ex_rs2_data[19] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold609 (.A(_01333_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold610 (.A(\soc_inst.mem_ctrl.next_instr_data[0] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold611 (.A(_00640_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold612 (.A(\soc_inst.cpu_core.register_file.registers[18][18] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold613 (.A(\soc_inst.cpu_core.register_file.registers[2][6] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold614 (.A(\soc_inst.cpu_core.csr_file.mtvec[12] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold615 (.A(_07421_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold616 (.A(_02410_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold617 (.A(\soc_inst.cpu_core.register_file.registers[17][20] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold618 (.A(\soc_inst.cpu_core.register_file.registers[13][9] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold619 (.A(\soc_inst.cpu_core.register_file.registers[16][3] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold620 (.A(\soc_inst.cpu_core.register_file.registers[18][21] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold621 (.A(\soc_inst.cpu_core.register_file.registers[14][5] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold622 (.A(\soc_inst.mem_ctrl.spi_data_in[20] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00498_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold624 (.A(\soc_inst.gpio_inst.int_pend_reg[6] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold625 (.A(_07578_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold626 (.A(_02446_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold627 (.A(\soc_inst.cpu_core.register_file.registers[20][21] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold628 (.A(\soc_inst.cpu_core.register_file.registers[8][11] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold629 (.A(\soc_inst.cpu_core.csr_file.mtvec[13] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold630 (.A(_07422_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold631 (.A(_02411_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold632 (.A(\soc_inst.cpu_core.register_file.registers[14][30] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold633 (.A(\soc_inst.core_mem_wdata[27] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold634 (.A(_02527_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold635 (.A(\soc_inst.cpu_core.register_file.registers[20][25] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold636 (.A(\soc_inst.cpu_core.csr_file.mtvec[6] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold637 (.A(_07415_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold638 (.A(_02404_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold639 (.A(\soc_inst.cpu_core.csr_file.mtvec[3] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold640 (.A(\soc_inst.cpu_core.register_file.registers[14][11] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold641 (.A(\soc_inst.cpu_core.register_file.registers[4][29] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold642 (.A(\soc_inst.spi_inst.busy ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold643 (.A(_00137_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold644 (.A(\soc_inst.cpu_core.register_file.registers[13][28] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold645 (.A(\soc_inst.mem_ctrl.next_instr_data[29] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold646 (.A(_00669_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold647 (.A(\soc_inst.cpu_core.csr_file.mscratch[17] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold648 (.A(_11172_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold649 (.A(_00798_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold650 (.A(\soc_inst.cpu_core.ex_rs1_data[15] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold651 (.A(_01265_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold652 (.A(\soc_inst.cpu_core.register_file.registers[2][4] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold653 (.A(\soc_inst.cpu_core.ex_rs1_data[25] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold654 (.A(_01275_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold655 (.A(\soc_inst.core_mem_wdata[30] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold656 (.A(_02530_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold657 (.A(\soc_inst.mem_ctrl.next_instr_data[19] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold658 (.A(_00659_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold659 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg_0 ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold660 (.A(_02597_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold661 (.A(\soc_inst.cpu_core.register_file.registers[18][23] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold662 (.A(\soc_inst.cpu_core.register_file.registers[1][29] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold663 (.A(\soc_inst.cpu_core.register_file.registers[14][16] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold664 (.A(\soc_inst.cpu_core.register_file.registers[24][29] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold665 (.A(\soc_inst.cpu_core.register_file.registers[2][0] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold666 (.A(\soc_inst.mem_ctrl.spi_data_in[3] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold667 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[5] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold668 (.A(_07729_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold669 (.A(_02578_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold670 (.A(\soc_inst.cpu_core.csr_file.mscratch[24] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold671 (.A(_00805_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold672 (.A(\soc_inst.cpu_core.register_file.registers[4][23] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold673 (.A(\soc_inst.cpu_core.register_file.registers[17][31] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold674 (.A(\soc_inst.cpu_core.register_file.registers[17][24] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold675 (.A(\soc_inst.cpu_core.register_file.registers[8][21] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold676 (.A(\soc_inst.cpu_core.register_file.registers[18][26] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold677 (.A(\soc_inst.cpu_core.register_file.registers[4][11] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold678 (.A(\soc_inst.cpu_core.register_file.registers[11][28] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold679 (.A(\soc_inst.cpu_core.register_file.registers[2][18] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold680 (.A(\soc_inst.cpu_core.register_file.registers[17][30] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold681 (.A(\soc_inst.spi_inst.clk_counter[2] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold682 (.A(_00130_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold683 (.A(\soc_inst.mem_ctrl.next_instr_data[1] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold684 (.A(_00641_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold685 (.A(\soc_inst.mem_ctrl.next_instr_data[20] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold686 (.A(_00660_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold687 (.A(\soc_inst.cpu_core.register_file.registers[13][23] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold688 (.A(\soc_inst.cpu_core.register_file.registers[4][8] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold689 (.A(\soc_inst.cpu_core.register_file.registers[13][21] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold690 (.A(\soc_inst.cpu_core.register_file.registers[14][4] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold691 (.A(\soc_inst.cpu_core.csr_file.mtime[0] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold692 (.A(\soc_inst.cpu_core.csr_file.mtval[18] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold693 (.A(_02389_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold694 (.A(\soc_inst.core_mem_rdata[12] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold695 (.A(\soc_inst.mem_ctrl.next_instr_data[6] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00646_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold697 (.A(\soc_inst.cpu_core.csr_file.mtvec[5] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold698 (.A(_07413_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold699 (.A(_02403_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold700 (.A(\soc_inst.cpu_core.register_file.registers[17][14] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold701 (.A(\soc_inst.cpu_core.register_file.registers[17][15] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold702 (.A(\soc_inst.cpu_core.register_file.registers[2][11] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold703 (.A(\soc_inst.gpio_inst.gpio_out[5] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold704 (.A(_00466_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold705 (.A(\soc_inst.cpu_core.register_file.registers[13][19] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold706 (.A(\soc_inst.cpu_core.csr_file.mstatus[9] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold707 (.A(_09910_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold708 (.A(_00513_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold709 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[27] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold710 (.A(_00746_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold711 (.A(\soc_inst.cpu_core.register_file.registers[2][13] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold712 (.A(\soc_inst.cpu_core.ex_rs2_data[2] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00843_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold714 (.A(\soc_inst.cpu_core.register_file.registers[16][19] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold715 (.A(\soc_inst.cpu_core.register_file.registers[8][18] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold716 (.A(\soc_inst.mem_ctrl.next_instr_data[15] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold717 (.A(_00655_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold718 (.A(\soc_inst.cpu_core.register_file.registers[8][1] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold719 (.A(\soc_inst.cpu_core.register_file.registers[1][7] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold720 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_en ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold721 (.A(_02598_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold722 (.A(\soc_inst.cpu_core.register_file.registers[16][24] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold723 (.A(\soc_inst.mem_ctrl.spi_data_in[4] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold724 (.A(\soc_inst.cpu_core.register_file.registers[13][7] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold725 (.A(\soc_inst.cpu_core.register_file.registers[15][9] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold726 (.A(\soc_inst.cpu_core.register_file.registers[18][5] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold727 (.A(\soc_inst.cpu_core.register_file.registers[14][28] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold728 (.A(\soc_inst.cpu_core.register_file.registers[14][24] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold729 (.A(\soc_inst.cpu_core.register_file.registers[1][13] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold730 (.A(\soc_inst.cpu_core.register_file.registers[13][5] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold731 (.A(\soc_inst.cpu_core.register_file.registers[13][8] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold732 (.A(\soc_inst.cpu_core.register_file.registers[18][6] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold733 (.A(\soc_inst.cpu_core.register_file.registers[11][17] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold734 (.A(\soc_inst.cpu_core.register_file.registers[8][4] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold735 (.A(\soc_inst.gpio_bidir_oe [0]),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold736 (.A(_00459_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold737 (.A(\soc_inst.cpu_core.register_file.registers[1][30] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold738 (.A(\soc_inst.cpu_core.register_file.registers[16][30] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold739 (.A(\soc_inst.cpu_core.register_file.registers[24][0] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold740 (.A(\soc_inst.cpu_core.register_file.registers[13][4] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold741 (.A(\soc_inst.i2c_inst.start_pending ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold742 (.A(_09264_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold743 (.A(\soc_inst.mem_ctrl.next_instr_data[5] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold744 (.A(_00645_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold745 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[2] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold746 (.A(_07738_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold747 (.A(_02584_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold748 (.A(\soc_inst.cpu_core.register_file.registers[14][7] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold749 (.A(\soc_inst.cpu_core.register_file.registers[17][23] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold750 (.A(\soc_inst.cpu_core.register_file.registers[1][27] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold751 (.A(\soc_inst.cpu_core.register_file.registers[11][3] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold752 (.A(\soc_inst.cpu_core.register_file.registers[17][9] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold753 (.A(\soc_inst.cpu_core.register_file.registers[18][13] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold754 (.A(\soc_inst.cpu_core.register_file.registers[14][29] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold755 (.A(\soc_inst.cpu_core.register_file.registers[2][23] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold756 (.A(\soc_inst.cpu_core.register_file.registers[11][18] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold757 (.A(\soc_inst.cpu_core.register_file.registers[16][11] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold758 (.A(\soc_inst.cpu_core.register_file.registers[18][29] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold759 (.A(\soc_inst.cpu_core.register_file.registers[18][8] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold760 (.A(\soc_inst.cpu_core.register_file.registers[1][14] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold761 (.A(\soc_inst.cpu_core.register_file.registers[16][9] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold762 (.A(\soc_inst.mem_ctrl.spi_data_in[11] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold763 (.A(\soc_inst.cpu_core.csr_file.mtvec[21] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold764 (.A(_07430_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold765 (.A(_02419_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold766 (.A(\soc_inst.cpu_core.register_file.registers[16][8] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold767 (.A(\soc_inst.cpu_core.register_file.registers[24][6] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold768 (.A(\soc_inst.cpu_core.register_file.registers[11][4] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold769 (.A(\soc_inst.cpu_core.register_file.registers[18][19] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold770 (.A(\soc_inst.cpu_core.register_file.registers[2][19] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold771 (.A(\soc_inst.spi_inst.state[1] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold772 (.A(\soc_inst.spi_inst.next_state[1] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold773 (.A(\soc_inst.cpu_core.ex_rs2_data[29] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold774 (.A(\soc_inst.mem_ctrl.spi_data_in[8] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold775 (.A(\soc_inst.core_mem_wdata[31] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold776 (.A(_02531_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold777 (.A(\soc_inst.cpu_core.ex_rs2_data[7] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold778 (.A(_04527_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold779 (.A(_01321_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold780 (.A(\soc_inst.cpu_core.register_file.registers[14][20] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold781 (.A(\soc_inst.cpu_core.register_file.registers[11][12] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold782 (.A(\soc_inst.cpu_core.register_file.registers[20][12] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold783 (.A(\soc_inst.cpu_core.register_file.registers[20][5] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold784 (.A(\soc_inst.cpu_core.register_file.registers[15][0] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold785 (.A(\soc_inst.cpu_core.register_file.registers[14][12] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold786 (.A(\soc_inst.cpu_core.register_file.registers[8][12] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold787 (.A(\soc_inst.mem_ctrl.spi_data_in[15] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold788 (.A(_00493_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold789 (.A(\soc_inst.cpu_core.register_file.registers[20][11] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold790 (.A(\soc_inst.cpu_core.register_file.registers[16][18] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold791 (.A(\soc_inst.cpu_core.register_file.registers[11][31] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold792 (.A(\soc_inst.cpu_core.register_file.registers[4][22] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold793 (.A(\soc_inst.cpu_core.register_file.registers[14][31] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold794 (.A(\soc_inst.cpu_core.if_instr[10] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold795 (.A(_00885_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold796 (.A(\soc_inst.cpu_core.register_file.registers[16][25] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold797 (.A(\soc_inst.cpu_core.register_file.registers[13][29] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold798 (.A(\soc_inst.cpu_core.register_file.registers[16][10] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold799 (.A(\soc_inst.cpu_core.register_file.registers[1][21] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold800 (.A(\soc_inst.cpu_core.register_file.registers[20][22] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold801 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[25] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold802 (.A(_00744_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold803 (.A(\soc_inst.cpu_core.register_file.registers[17][25] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold804 (.A(\soc_inst.mem_ctrl.next_instr_data[16] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold805 (.A(_00656_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold806 (.A(\soc_inst.cpu_core.ex_rs1_data[22] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold807 (.A(_01272_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold808 (.A(\soc_inst.cpu_core.register_file.registers[4][17] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold809 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[24] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold810 (.A(_00710_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold811 (.A(\soc_inst.cpu_core.register_file.registers[4][10] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold812 (.A(\soc_inst.cpu_core.ex_rs1_data[20] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold813 (.A(_01270_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold814 (.A(\soc_inst.cpu_core.register_file.registers[24][13] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold815 (.A(\soc_inst.cpu_core.register_file.registers[17][12] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold816 (.A(\soc_inst.cpu_core.register_file.registers[2][21] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold817 (.A(\soc_inst.cpu_core.error_flag_reg ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold818 (.A(_00874_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold819 (.A(\soc_inst.mem_ctrl.spi_data_in[22] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold820 (.A(_00500_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold821 (.A(\soc_inst.cpu_core.register_file.registers[24][3] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold822 (.A(\soc_inst.mem_ctrl.next_instr_data[18] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold823 (.A(_00658_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold824 (.A(\soc_inst.mem_ctrl.next_instr_data[30] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold825 (.A(_00670_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold826 (.A(\soc_inst.cpu_core.register_file.registers[11][27] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold827 (.A(\soc_inst.mem_ctrl.next_instr_data[24] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00664_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold829 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[6] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold830 (.A(_00725_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold831 (.A(\soc_inst.cpu_core.register_file.registers[17][4] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold832 (.A(\soc_inst.cpu_core.register_file.registers[4][6] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold833 (.A(\soc_inst.cpu_core.register_file.registers[1][26] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold834 (.A(\soc_inst.cpu_core.register_file.registers[18][25] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold835 (.A(\soc_inst.cpu_core.register_file.registers[4][20] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold836 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[23] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold837 (.A(_00709_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold838 (.A(\soc_inst.cpu_core.ex_funct7[0] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold839 (.A(_01049_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold840 (.A(\soc_inst.cpu_core.register_file.registers[8][5] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold841 (.A(\soc_inst.cpu_core.register_file.registers[18][31] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold842 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[2] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold843 (.A(_02568_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold844 (.A(\soc_inst.cpu_core.register_file.registers[18][27] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold845 (.A(\soc_inst.cpu_core.register_file.registers[11][1] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold846 (.A(\soc_inst.cpu_core.register_file.registers[4][1] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold847 (.A(\soc_inst.cpu_core.ex_rs2_data[9] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold848 (.A(_01323_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold849 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[16] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold850 (.A(\soc_inst.cpu_core.register_file.registers[11][19] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold851 (.A(\soc_inst.cpu_core.register_file.registers[2][14] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold852 (.A(\soc_inst.mem_ctrl.spi_data_in[12] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold853 (.A(\soc_inst.cpu_core.register_file.registers[16][15] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold854 (.A(\soc_inst.cpu_core.register_file.registers[24][21] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold855 (.A(\soc_inst.cpu_core.register_file.registers[18][3] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold856 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[26] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold857 (.A(_00745_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold858 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[17] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold859 (.A(_00703_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold860 (.A(\soc_inst.cpu_core.register_file.registers[18][12] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold861 (.A(\soc_inst.cpu_core.register_file.registers[13][24] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold862 (.A(\soc_inst.cpu_core.csr_file.mtime[43] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold863 (.A(_00210_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold864 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[20] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold865 (.A(_00706_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold866 (.A(\soc_inst.mem_ctrl.next_instr_data[7] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold867 (.A(_00647_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold868 (.A(\soc_inst.cpu_core.register_file.registers[15][6] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold869 (.A(\soc_inst.cpu_core.csr_file.mtvec[23] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold870 (.A(_07432_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold871 (.A(_02421_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold872 (.A(\soc_inst.cpu_core.register_file.registers[2][16] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold873 (.A(\soc_inst.cpu_core.register_file.registers[13][10] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold874 (.A(\soc_inst.cpu_core.register_file.registers[24][17] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold875 (.A(\soc_inst.cpu_core.register_file.registers[17][0] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold876 (.A(\soc_inst.cpu_core.register_file.registers[16][14] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold877 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[16] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold878 (.A(_00735_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold879 (.A(\soc_inst.cpu_core.register_file.registers[15][7] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold880 (.A(\soc_inst.cpu_core.register_file.registers[17][5] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold881 (.A(\soc_inst.cpu_core.register_file.registers[16][23] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold882 (.A(\soc_inst.cpu_core.register_file.registers[16][31] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold883 (.A(\soc_inst.cpu_core.register_file.registers[11][16] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold884 (.A(\soc_inst.cpu_core.register_file.registers[15][24] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold885 (.A(\soc_inst.mem_ctrl.spi_data_in[14] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold886 (.A(_00492_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold887 (.A(\soc_inst.cpu_core.register_file.registers[2][2] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold888 (.A(\soc_inst.cpu_core.register_file.registers[15][25] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold889 (.A(\soc_inst.cpu_core.register_file.registers[20][19] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold890 (.A(\soc_inst.cpu_core.register_file.registers[20][18] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold891 (.A(\soc_inst.cpu_core.register_file.registers[16][22] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold892 (.A(\soc_inst.cpu_core.register_file.registers[17][11] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold893 (.A(\soc_inst.cpu_core.register_file.registers[20][2] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold894 (.A(\soc_inst.cpu_core.register_file.registers[15][20] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold895 (.A(\soc_inst.cpu_core.register_file.registers[8][25] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold896 (.A(\soc_inst.cpu_core.register_file.registers[24][4] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold897 (.A(\soc_inst.mem_ctrl.next_instr_data[27] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold898 (.A(_00667_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold899 (.A(\soc_inst.gpio_inst.int_pend_reg[0] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold900 (.A(_09437_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00388_),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold902 (.A(\soc_inst.core_mem_rdata[14] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold903 (.A(\soc_inst.cpu_core.register_file.registers[15][1] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold904 (.A(\soc_inst.cpu_core.register_file.registers[4][16] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold905 (.A(\soc_inst.cpu_core.register_file.registers[16][12] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold906 (.A(\soc_inst.cpu_core.register_file.registers[11][13] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold907 (.A(\soc_inst.cpu_core.register_file.registers[14][26] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold908 (.A(\soc_inst.cpu_core.register_file.registers[24][31] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold909 (.A(\soc_inst.cpu_core.csr_file.mtime[10] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold910 (.A(_00174_),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold911 (.A(\soc_inst.cpu_core.register_file.registers[14][3] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold912 (.A(\soc_inst.cpu_core.register_file.registers[1][11] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold913 (.A(\soc_inst.cpu_core.register_file.registers[13][15] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold914 (.A(\soc_inst.cpu_core.register_file.registers[16][1] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold915 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[22] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold916 (.A(_00741_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold917 (.A(\soc_inst.cpu_core.register_file.registers[24][8] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold918 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[6] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold919 (.A(_00692_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold920 (.A(\soc_inst.cpu_core.register_file.registers[11][5] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold921 (.A(\soc_inst.cpu_core.register_file.registers[14][14] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold922 (.A(\soc_inst.cpu_core.register_file.registers[4][27] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold923 (.A(\soc_inst.cpu_core.register_file.registers[2][28] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold924 (.A(\soc_inst.cpu_core.register_file.registers[8][6] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold925 (.A(\soc_inst.cpu_core.register_file.registers[16][2] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold926 (.A(\soc_inst.cpu_core.register_file.registers[24][1] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold927 (.A(\soc_inst.cpu_core.register_file.registers[13][3] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold928 (.A(\soc_inst.cpu_core.register_file.registers[24][20] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold929 (.A(\soc_inst.cpu_core.register_file.registers[16][0] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold930 (.A(\soc_inst.mem_ctrl.next_instr_data[10] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold931 (.A(_00650_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold932 (.A(\soc_inst.cpu_core.register_file.registers[15][2] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold933 (.A(\soc_inst.cpu_core.register_file.registers[15][30] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold934 (.A(\soc_inst.i2c_inst.bit_cnt[2] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold935 (.A(_09461_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold936 (.A(_00403_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold937 (.A(\soc_inst.core_mem_wdata[26] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold938 (.A(_02526_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold939 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[3] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold940 (.A(_07728_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold941 (.A(\soc_inst.core_mem_rdata[21] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold942 (.A(_00626_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold943 (.A(\soc_inst.cpu_core.register_file.registers[13][30] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold944 (.A(\soc_inst.cpu_core.register_file.registers[20][1] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold945 (.A(\soc_inst.cpu_core.csr_file.mtvec[17] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold946 (.A(_07426_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold947 (.A(_02415_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold948 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[7] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold949 (.A(_09366_),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold950 (.A(\soc_inst.cpu_core.register_file.registers[11][0] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold951 (.A(\soc_inst.cpu_core.register_file.registers[8][26] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold952 (.A(\soc_inst.mem_ctrl.next_instr_data[25] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold953 (.A(_00665_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold954 (.A(\soc_inst.cpu_core.ex_rs1_data[18] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold955 (.A(_01268_),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold956 (.A(\soc_inst.cpu_core.register_file.registers[13][12] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold957 (.A(\soc_inst.cpu_core.register_file.registers[1][18] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold958 (.A(\soc_inst.cpu_core.register_file.registers[2][25] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold959 (.A(\soc_inst.cpu_core.register_file.registers[17][10] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold960 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[3] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold961 (.A(_00689_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold962 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[21] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold963 (.A(_00740_),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold964 (.A(\soc_inst.cpu_core.register_file.registers[11][6] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold965 (.A(\soc_inst.cpu_core.register_file.registers[1][5] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold966 (.A(\soc_inst.cpu_core.register_file.registers[13][0] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold967 (.A(\soc_inst.cpu_core.register_file.registers[15][12] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold968 (.A(\soc_inst.cpu_core.register_file.registers[20][26] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold969 (.A(\soc_inst.cpu_core.register_file.registers[14][1] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold970 (.A(\soc_inst.cpu_core.register_file.registers[18][4] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold971 (.A(\soc_inst.cpu_core.register_file.registers[20][4] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold972 (.A(\soc_inst.core_mem_addr[8] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold973 (.A(_01290_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold974 (.A(\soc_inst.cpu_core.register_file.registers[11][14] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold975 (.A(\soc_inst.spi_inst.rx_shift_reg[30] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold976 (.A(_09421_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold977 (.A(\soc_inst.cpu_core.csr_file.mtvec[10] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold978 (.A(_07419_),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold979 (.A(_02408_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold980 (.A(\soc_inst.cpu_core.register_file.registers[17][19] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold981 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[19] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold982 (.A(_00705_),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold983 (.A(\soc_inst.cpu_core.register_file.registers[4][2] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold984 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[18] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold985 (.A(_00704_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold986 (.A(\soc_inst.mem_ctrl.next_instr_data[12] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold987 (.A(_00652_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold988 (.A(\soc_inst.cpu_core.register_file.registers[4][9] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold989 (.A(\soc_inst.cpu_core.csr_file.mtvec[9] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold990 (.A(_07418_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold991 (.A(_02407_),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold992 (.A(\soc_inst.pwm_inst.channel_counter[0][15] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold993 (.A(_08936_),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold994 (.A(\soc_inst.cpu_core.register_file.registers[15][18] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold995 (.A(\soc_inst.cpu_core.register_file.registers[11][30] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold996 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[11] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold997 (.A(_00730_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold998 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[5] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold999 (.A(_00003_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\soc_inst.cpu_core.register_file.registers[11][9] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\soc_inst.cpu_core.register_file.registers[18][16] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\soc_inst.cpu_core.csr_file.mtime[11] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold1003 (.A(_00175_),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\soc_inst.cpu_core.mem_instr[15] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold1005 (.A(_01039_),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\soc_inst.cpu_core.register_file.registers[24][28] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\soc_inst.mem_ctrl.spi_data_in[9] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[8] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_00694_),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\soc_inst.cpu_core.ex_rs2_data[28] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\soc_inst.cpu_core.csr_file.mtime[6] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_00217_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\soc_inst.cpu_core.register_file.registers[15][19] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[10] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\soc_inst.cpu_core.register_file.registers[1][6] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\soc_inst.cpu_core.register_file.registers[16][6] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\soc_inst.cpu_core.register_file.registers[8][20] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\soc_inst.cpu_core.register_file.registers[1][25] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\soc_inst.cpu_core.register_file.registers[24][18] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\soc_inst.mem_ctrl.spi_data_in[10] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_00488_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\soc_inst.cpu_core.register_file.registers[8][13] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\soc_inst.cpu_core.register_file.registers[15][8] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\soc_inst.spi_inst.tx_shift_reg[22] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_00153_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\soc_inst.pwm_ena [0]),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_02442_),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\soc_inst.cpu_core.register_file.registers[20][29] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\soc_inst.cpu_core.register_file.registers[4][25] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\soc_inst.cpu_core.register_file.registers[13][18] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\soc_inst.core_mem_addr[10] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_01292_),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\soc_inst.cpu_core.register_file.registers[16][26] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\soc_inst.cpu_core.register_file.registers[17][18] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\soc_inst.mem_ctrl.next_instr_data[2] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_00642_),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\soc_inst.cpu_core.register_file.registers[8][14] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[30] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold1039 (.A(_00716_),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\soc_inst.core_mem_rdata[31] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold1041 (.A(_00636_),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\soc_inst.cpu_core.id_imm12[5] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[13] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold1044 (.A(_00699_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\soc_inst.cpu_core.register_file.registers[17][13] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\soc_inst.spi_inst.rx_shift_reg[24] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_09415_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\soc_inst.cpu_core.register_file.registers[13][6] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\soc_inst.cpu_core.register_file.registers[16][29] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\soc_inst.cpu_core.register_file.registers[20][17] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\soc_inst.cpu_core.register_file.registers[8][8] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\soc_inst.cpu_core.register_file.registers[2][17] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\soc_inst.mem_ctrl.next_instr_data[13] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold1054 (.A(_00653_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[1] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold1056 (.A(_08637_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_00018_),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[2] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\soc_inst.cpu_core.register_file.registers[17][8] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\soc_inst.cpu_core.register_file.registers[1][1] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\soc_inst.cpu_core.csr_file.mtime[47] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold1062 (.A(_00214_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\soc_inst.cpu_core.register_file.registers[1][3] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\soc_inst.cpu_core.csr_file.mtvec[16] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold1065 (.A(_07425_),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_02414_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\soc_inst.spi_inst.rx_shift_reg[29] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_09420_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\soc_inst.core_mem_rdata[29] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_00634_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\soc_inst.cpu_core.register_file.registers[18][28] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\soc_inst.cpu_core.register_file.registers[17][27] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\soc_inst.cpu_core.csr_file.mscratch[28] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_00809_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\soc_inst.cpu_core.register_file.registers[16][16] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\soc_inst.cpu_core.register_file.registers[24][15] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\soc_inst.cpu_core.register_file.registers[4][19] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\soc_inst.cpu_core.register_file.registers[22][7] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\soc_inst.cpu_core.ex_instr[17] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_01041_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\soc_inst.spi_inst.rx_shift_reg[28] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_09419_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\soc_inst.spi_inst.rx_shift_reg[21] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_09412_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\soc_inst.cpu_core.register_file.registers[24][30] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\soc_inst.core_mem_rdata[10] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\soc_inst.cpu_core.csr_file.mtime[12] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold1088 (.A(_09324_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\soc_inst.cpu_core.register_file.registers[4][0] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\soc_inst.cpu_core.csr_file.mtime[42] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_00209_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\soc_inst.cpu_core.register_file.registers[18][17] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\soc_inst.cpu_core.register_file.registers[7][24] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\soc_inst.cpu_core.register_file.registers[11][23] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[27] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\soc_inst.cpu_core.register_file.registers[14][23] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\soc_inst.cpu_core.register_file.registers[16][5] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\soc_inst.cpu_core.ex_reg_we ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_00838_),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\soc_inst.cpu_core.csr_file.mtime[3] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_00206_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\soc_inst.cpu_core.csr_file.mtvec[22] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_07431_),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_02420_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\soc_inst.cpu_core.register_file.registers[14][13] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\soc_inst.cpu_core.register_file.registers[5][28] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\soc_inst.cpu_core.register_file.registers[8][2] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\soc_inst.cpu_core.register_file.registers[28][0] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\soc_inst.core_mem_rdata[23] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold1110 (.A(_00628_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[23] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_00742_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\soc_inst.cpu_core.register_file.registers[11][2] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\soc_inst.cpu_core.csr_file.mtvec[7] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_07416_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_02405_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\soc_inst.cpu_core.register_file.registers[1][17] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\soc_inst.cpu_core.ex_rs1_data[7] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold1119 (.A(_01257_),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\soc_inst.cpu_core.csr_file.mtime[35] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold1121 (.A(_00201_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\soc_inst.cpu_core.register_file.registers[18][11] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\soc_inst.cpu_core.csr_file.mtval[6] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_02377_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\soc_inst.cpu_core.register_file.registers[15][13] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_00223_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold1127 (.A(_00380_),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[15] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_00701_),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\soc_inst.cpu_core.register_file.registers[1][0] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\soc_inst.cpu_core.register_file.registers[9][24] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\soc_inst.cpu_core.register_file.registers[16][13] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\soc_inst.cpu_core.register_file.registers[3][5] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\soc_inst.cpu_core.register_file.registers[24][22] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\soc_inst.cpu_core.register_file.registers[20][6] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\soc_inst.gpio_inst.gpio_out[3] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\soc_inst.cpu_core.csr_file.mepc[10] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_02427_),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\soc_inst.cpu_core.register_file.registers[12][28] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\soc_inst.cpu_core.register_file.registers[11][21] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\soc_inst.cpu_core.register_file.registers[4][18] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\soc_inst.cpu_core.register_file.registers[22][8] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold1143 (.A(_00266_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_00107_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\soc_inst.core_mem_rdata[24] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold1146 (.A(_00629_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\soc_inst.mem_ctrl.next_instr_data[9] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold1148 (.A(_00649_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[9] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold1150 (.A(_00695_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\soc_inst.i2c_inst.clk_cnt[2] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold1152 (.A(_08860_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_00091_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\soc_inst.cpu_core.register_file.registers[12][27] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\soc_inst.cpu_core.register_file.registers[11][10] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\soc_inst.cpu_core.register_file.registers[16][28] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\soc_inst.cpu_core.register_file.registers[3][26] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[0] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold1159 (.A(_00686_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\soc_inst.cpu_core.register_file.registers[17][2] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\soc_inst.cpu_core.register_file.registers[9][17] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\soc_inst.cpu_core.register_file.registers[17][22] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\soc_inst.cpu_core.register_file.registers[2][31] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\soc_inst.cpu_core.register_file.registers[5][16] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\soc_inst.cpu_core.register_file.registers[10][30] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\soc_inst.cpu_core.csr_file.mtime[14] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_00178_),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\soc_inst.cpu_core.register_file.registers[15][23] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\soc_inst.cpu_core.if_instr[11] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold1170 (.A(_00886_),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\soc_inst.cpu_core.register_file.registers[19][17] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\soc_inst.cpu_core.ex_mem_re ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold1173 (.A(_01379_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\soc_inst.cpu_core.register_file.registers[2][5] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\soc_inst.cpu_core.register_file.registers[28][29] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\soc_inst.cpu_core.mem_stall ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\soc_inst.cpu_core.register_file.registers[13][1] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\soc_inst.cpu_core.register_file.registers[17][1] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\soc_inst.cpu_core.register_file.registers[15][16] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\soc_inst.cpu_core.register_file.registers[28][24] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\soc_inst.cpu_core.register_file.registers[8][27] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\soc_inst.cpu_core.csr_file.mepc[8] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_02425_),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[21] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00707_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\soc_inst.cpu_core.if_instr[9] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_00884_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\soc_inst.cpu_core.register_file.registers[17][26] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\soc_inst.cpu_core.ex_exception_pc[5] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold1190 (.A(_01231_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\soc_inst.cpu_core.if_instr[8] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\soc_inst.cpu_core.register_file.registers[12][18] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\soc_inst.core_mem_wdata[18] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_02518_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\soc_inst.cpu_core.register_file.registers[10][22] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\soc_inst.cpu_core.register_file.registers[22][11] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\soc_inst.cpu_core.register_file.registers[28][13] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\soc_inst.cpu_core.register_file.registers[9][2] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\soc_inst.cpu_core.register_file.registers[14][10] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\soc_inst.cpu_core.ex_rs1_data[24] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_01274_),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\soc_inst.cpu_core.ex_instr[22] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold1203 (.A(_01046_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\soc_inst.cpu_core.register_file.registers[29][17] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\soc_inst.cpu_core.register_file.registers[26][20] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\soc_inst.cpu_core.register_file.registers[2][29] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\soc_inst.cpu_core.register_file.registers[4][5] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\soc_inst.cpu_core.register_file.registers[4][28] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\soc_inst.cpu_core.register_file.registers[16][27] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[26] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold1211 (.A(_00712_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\soc_inst.cpu_core.id_rs2_data[2] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\soc_inst.cpu_core.csr_file.mepc[9] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_02426_),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\soc_inst.cpu_core.register_file.registers[18][30] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\soc_inst.cpu_core.register_file.registers[3][23] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\soc_inst.cpu_core.register_file.registers[8][22] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\soc_inst.cpu_core.register_file.registers[31][21] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\soc_inst.cpu_core.register_file.registers[8][23] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\soc_inst.cpu_core.mem_rs1_data[12] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\soc_inst.cpu_core.register_file.registers[6][30] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\soc_inst.spi_inst.rx_shift_reg[27] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_09418_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\soc_inst.cpu_core.register_file.registers[29][28] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\soc_inst.cpu_core.register_file.registers[1][24] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\soc_inst.cpu_core.register_file.registers[27][8] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\soc_inst.cpu_core.register_file.registers[23][31] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\soc_inst.cpu_core.register_file.registers[8][19] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\soc_inst.cpu_core.register_file.registers[23][9] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\soc_inst.mem_ctrl.spi_mem_inst.initialized ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\soc_inst.core_mem_rdata[11] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\soc_inst.core_mem_wdata[22] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_02522_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\soc_inst.cpu_core.register_file.registers[10][0] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\soc_inst.core_mem_rdata[0] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\soc_inst.cpu_core.register_file.registers[26][24] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\soc_inst.cpu_core.if_pc[2] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold1238 (.A(_02454_),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\soc_inst.cpu_core.id_rs2_data[28] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold1240 (.A(_00290_),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_02507_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\soc_inst.core_mem_wdata[13] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\soc_inst.cpu_core.register_file.registers[26][7] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\soc_inst.cpu_core.csr_file.mtime[13] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\soc_inst.cpu_core.register_file.registers[3][9] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\soc_inst.cpu_core.register_file.registers[11][11] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\soc_inst.cpu_core.register_file.registers[20][16] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\soc_inst.cpu_core.register_file.registers[27][6] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\soc_inst.cpu_core.register_file.registers[18][7] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\soc_inst.core_mem_wdata[23] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\soc_inst.cpu_core.register_file.registers[30][10] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\soc_inst.cpu_core.csr_file.mtime[38] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_00204_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\soc_inst.cpu_core.register_file.registers[27][22] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\soc_inst.cpu_core.register_file.registers[28][27] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\soc_inst.spi_inst.tx_shift_reg[21] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_00152_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\soc_inst.cpu_core.register_file.registers[7][18] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[22] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\soc_inst.cpu_core.register_file.registers[21][10] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\soc_inst.cpu_core.register_file.registers[9][10] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\soc_inst.spi_inst.tx_shift_reg[26] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\soc_inst.cpu_core.register_file.registers[27][2] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\soc_inst.cpu_core.id_rs2_data[29] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\soc_inst.cpu_core.register_file.registers[5][6] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\soc_inst.cpu_core.register_file.registers[21][30] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\soc_inst.cpu_core.register_file.registers[31][15] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\soc_inst.cpu_core.register_file.registers[7][20] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\soc_inst.cpu_core.mem_rs1_data[30] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\soc_inst.cpu_core.register_file.registers[7][7] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\soc_inst.cpu_core.id_instr[16] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold1272 (.A(_01210_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\soc_inst.cpu_core.register_file.registers[5][22] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\soc_inst.cpu_core.csr_file.mtime[1] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\soc_inst.cpu_core.register_file.registers[4][13] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\soc_inst.cpu_core.register_file.registers[28][31] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\soc_inst.cpu_core.register_file.registers[23][13] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[1] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_00687_),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\soc_inst.cpu_core.register_file.registers[25][16] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\soc_inst.cpu_core.register_file.registers[15][4] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\soc_inst.spi_inst.rx_shift_reg[20] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_09411_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\soc_inst.cpu_core.id_instr[18] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold1285 (.A(_01212_),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\soc_inst.spi_inst.rx_shift_reg[18] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_09409_),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\soc_inst.cpu_core.register_file.registers[14][8] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\soc_inst.cpu_core.ex_rs1_data[23] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_01273_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\soc_inst.cpu_core.register_file.registers[18][14] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\soc_inst.cpu_core.register_file.registers[17][21] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\soc_inst.cpu_core.csr_file.mtime[41] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold1294 (.A(_00208_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\soc_inst.cpu_core.register_file.registers[9][20] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[15] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_08628_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_00011_),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\soc_inst.cpu_core.mem_rs1_data[14] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\soc_inst.cpu_core.register_file.registers[22][6] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\soc_inst.core_mem_rdata[20] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_00625_),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\soc_inst.cpu_core.ex_exception_pc[14] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_01240_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\soc_inst.cpu_core.ex_exception_pc[6] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01232_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\soc_inst.gpio_inst.gpio_out[4] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_00465_),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[2] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\soc_inst.cpu_core.register_file.registers[27][18] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\soc_inst.cpu_core.register_file.registers[28][16] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[4] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_00723_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\soc_inst.cpu_core.register_file.registers[25][22] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\soc_inst.cpu_core.ex_alu_result[31] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\soc_inst.cpu_core.register_file.registers[9][15] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\soc_inst.cpu_core.ex_rs2_data[11] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold1318 (.A(_00852_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\soc_inst.cpu_core.mem_rs1_data[31] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\soc_inst.core_mem_wdata[6] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\soc_inst.cpu_core.register_file.registers[19][2] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\soc_inst.cpu_core.ex_exception_pc[10] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold1323 (.A(_01236_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\soc_inst.cpu_core.register_file.registers[9][7] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\soc_inst.cpu_core.mem_instr[19] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_01043_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\soc_inst.cpu_core.register_file.registers[10][20] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\soc_inst.cpu_core.register_file.registers[27][15] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\soc_inst.cpu_core.register_file.registers[28][22] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\soc_inst.cpu_core.register_file.registers[6][8] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\soc_inst.cpu_core.register_file.registers[21][2] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[25] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\soc_inst.cpu_core.register_file.registers[9][18] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\soc_inst.cpu_core.mem_rs1_data[8] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[7] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[4] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold1337 (.A(_00690_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[6] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_02572_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\soc_inst.cpu_core.register_file.registers[7][22] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\soc_inst.cpu_core.csr_file.mepc[6] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\soc_inst.cpu_core.register_file.registers[3][25] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\soc_inst.cpu_core.register_file.registers[6][16] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\soc_inst.cpu_core.register_file.registers[8][0] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\soc_inst.cpu_core.register_file.registers[29][23] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\soc_inst.cpu_core.register_file.registers[21][31] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\soc_inst.cpu_core.register_file.registers[21][21] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\soc_inst.cpu_core.register_file.registers[25][10] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\soc_inst.spi_inst.tx_shift_reg[11] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\soc_inst.cpu_core.register_file.registers[9][5] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\soc_inst.cpu_core.register_file.registers[31][11] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\soc_inst.cpu_core.register_file.registers[5][29] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\soc_inst.cpu_core.register_file.registers[28][21] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\soc_inst.cpu_core.register_file.registers[19][18] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\soc_inst.core_mem_wdata[7] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\soc_inst.cpu_core.register_file.registers[5][7] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\soc_inst.cpu_core.register_file.registers[9][28] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\soc_inst.cpu_core.register_file.registers[21][8] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\soc_inst.mem_ctrl.spi_read_enable ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold1360 (.A(_00637_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\soc_inst.cpu_core.register_file.registers[23][24] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\soc_inst.cpu_core.register_file.registers[10][16] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\soc_inst.spi_inst.tx_shift_reg[31] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold1364 (.A(_09378_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_00337_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\soc_inst.spi_inst.tx_shift_reg[2] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\soc_inst.core_instr_data[31] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_00604_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\soc_inst.cpu_core.register_file.registers[19][20] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\soc_inst.cpu_core.register_file.registers[3][16] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\soc_inst.cpu_core.register_file.registers[23][26] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\soc_inst.cpu_core.register_file.registers[19][23] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\soc_inst.cpu_core.mem_rs1_data[13] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\soc_inst.cpu_core.ex_exception_pc[12] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_01238_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\soc_inst.cpu_core.register_file.registers[29][27] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\soc_inst.cpu_core.mem_rs1_data[9] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold1378 (.A(_00297_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_02514_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\soc_inst.cpu_core.register_file.registers[3][21] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\soc_inst.cpu_core.register_file.registers[23][22] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\soc_inst.cpu_core.register_file.registers[19][24] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\soc_inst.cpu_core.register_file.registers[29][10] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\soc_inst.cpu_core.register_file.registers[30][3] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\soc_inst.cpu_core.register_file.registers[3][8] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\soc_inst.cpu_core.register_file.registers[23][16] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\soc_inst.cpu_core.id_rs2_data[1] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\soc_inst.spi_inst.rx_shift_reg[26] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold1389 (.A(_09417_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[6] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_07698_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold1392 (.A(_02551_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\soc_inst.cpu_core.register_file.registers[10][7] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\soc_inst.cpu_core.register_file.registers[28][25] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\soc_inst.cpu_core.register_file.registers[5][27] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\soc_inst.cpu_core.register_file.registers[6][9] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\soc_inst.cpu_core.register_file.registers[5][20] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\soc_inst.cpu_core.register_file.registers[21][13] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\soc_inst.cpu_core.register_file.registers[31][22] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\soc_inst.cpu_core.mem_rs1_data[10] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\soc_inst.spi_inst.done ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_09435_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\soc_inst.cpu_core.csr_file.mtime[36] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold1404 (.A(_00202_),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\soc_inst.cpu_core.register_file.registers[31][31] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\soc_inst.cpu_core.register_file.registers[21][29] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\soc_inst.cpu_core.register_file.registers[29][13] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\soc_inst.cpu_core.register_file.registers[7][27] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\soc_inst.cpu_core.csr_file.mscratch[0] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[14] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\soc_inst.cpu_core.register_file.registers[10][19] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\soc_inst.cpu_core.id_rs2_data[0] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\soc_inst.cpu_core.if_instr[18] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\soc_inst.spi_inst.tx_shift_reg[19] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_00150_),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\soc_inst.cpu_core.register_file.registers[22][24] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_00225_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\soc_inst.core_mem_wdata[8] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\soc_inst.cpu_core.register_file.registers[30][4] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\soc_inst.cpu_core.register_file.registers[19][16] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\soc_inst.cpu_core.register_file.registers[25][9] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\soc_inst.cpu_core.register_file.registers[30][29] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\soc_inst.cpu_core.register_file.registers[5][25] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\soc_inst.core_mem_wdata[14] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\soc_inst.cpu_core.mem_rs1_data[26] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\soc_inst.cpu_core.register_file.registers[30][16] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\soc_inst.cpu_core.register_file.registers[6][1] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\soc_inst.cpu_core.register_file.registers[5][15] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\soc_inst.core_mem_rdata[30] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold1430 (.A(_00635_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\soc_inst.cpu_core.register_file.registers[26][26] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\soc_inst.cpu_core.register_file.registers[26][27] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\soc_inst.cpu_core.if_instr[16] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\soc_inst.cpu_core.ex_branch_target[11] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_02353_),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\soc_inst.cpu_core.register_file.registers[27][26] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\soc_inst.cpu_core.register_file.registers[23][6] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\soc_inst.cpu_core.register_file.registers[16][21] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\soc_inst.core_mem_wdata[5] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\soc_inst.cpu_core.register_file.registers[27][13] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\soc_inst.cpu_core.register_file.registers[14][25] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\soc_inst.cpu_core.register_file.registers[27][23] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\soc_inst.cpu_core.register_file.registers[4][14] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\soc_inst.cpu_core.register_file.registers[5][2] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\soc_inst.cpu_core.register_file.registers[6][3] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\soc_inst.cpu_core.register_file.registers[9][9] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\soc_inst.spi_inst.tx_shift_reg[5] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\soc_inst.cpu_core.register_file.registers[22][17] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\soc_inst.cpu_core.register_file.registers[21][6] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\soc_inst.cpu_core.register_file.registers[10][4] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\soc_inst.cpu_core.register_file.registers[14][19] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\soc_inst.cpu_core.register_file.registers[5][17] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\soc_inst.cpu_core.register_file.registers[27][17] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\soc_inst.core_mem_wdata[10] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\soc_inst.cpu_core.register_file.registers[4][4] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\soc_inst.cpu_core.register_file.registers[9][11] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\soc_inst.cpu_core.register_file.registers[27][31] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\soc_inst.cpu_core.register_file.registers[26][6] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\soc_inst.core_mem_addr[11] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01293_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\soc_inst.cpu_core.register_file.registers[7][3] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\soc_inst.cpu_core.register_file.registers[21][27] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\soc_inst.spi_inst.rx_shift_reg[25] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\soc_inst.cpu_core.register_file.registers[26][13] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\soc_inst.cpu_core.register_file.registers[12][6] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\soc_inst.cpu_core.id_instr[17] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\soc_inst.cpu_core.register_file.registers[25][14] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\soc_inst.cpu_core.register_file.registers[21][25] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\soc_inst.cpu_core.ex_rs2_data[15] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold1470 (.A(_01329_),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\soc_inst.cpu_core.register_file.registers[7][31] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\soc_inst.cpu_core.register_file.registers[5][8] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\soc_inst.cpu_core.register_file.registers[20][27] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\soc_inst.cpu_core.register_file.registers[10][21] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\soc_inst.cpu_core.register_file.registers[9][22] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\soc_inst.cpu_core.register_file.registers[22][13] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\soc_inst.core_mem_rdata[15] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\soc_inst.spi_inst.rx_shift_reg[16] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold1479 (.A(_09407_),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\soc_inst.cpu_core.register_file.registers[23][27] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\soc_inst.gpio_inst.gpio_out[2] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\soc_inst.cpu_core.register_file.registers[30][15] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\soc_inst.cpu_core.ex_exception_pc[20] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_01246_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\soc_inst.cpu_core.register_file.registers[12][4] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\soc_inst.i2c_inst.stop_pending ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold1487 (.A(_08796_),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_00105_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\soc_inst.mem_ctrl.spi_mem_inst.start ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_08294_),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold1491 (.A(_00319_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\soc_inst.cpu_core.register_file.registers[3][24] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\soc_inst.cpu_core.register_file.registers[28][9] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\soc_inst.cpu_core.register_file.registers[9][13] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\soc_inst.cpu_core.register_file.registers[28][17] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\soc_inst.cpu_core.register_file.registers[22][2] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\soc_inst.cpu_core.csr_file.mepc[20] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold1498 (.A(_02437_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\soc_inst.cpu_core.register_file.registers[6][24] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\soc_inst.cpu_core.register_file.registers[28][20] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\soc_inst.cpu_core.register_file.registers[12][11] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\soc_inst.cpu_core.register_file.registers[3][11] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\soc_inst.cpu_core.mem_rs1_data[11] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\soc_inst.cpu_core.register_file.registers[31][24] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\soc_inst.cpu_core.register_file.registers[6][10] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\soc_inst.cpu_core.register_file.registers[6][21] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\soc_inst.cpu_core.register_file.registers[7][5] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\soc_inst.cpu_core.register_file.registers[25][1] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\soc_inst.cpu_core.register_file.registers[19][15] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\soc_inst.cpu_core.register_file.registers[22][20] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\soc_inst.cpu_core.register_file.registers[10][23] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\soc_inst.cpu_core.mem_rs1_data[27] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\soc_inst.cpu_core.register_file.registers[19][27] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[2] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_01191_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\soc_inst.cpu_core.register_file.registers[29][24] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\soc_inst.cpu_core.register_file.registers[30][7] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\soc_inst.cpu_core.register_file.registers[3][29] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\soc_inst.cpu_core.mem_rs1_data[3] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\soc_inst.cpu_core.register_file.registers[29][15] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\soc_inst.cpu_core.register_file.registers[7][25] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\soc_inst.cpu_core.register_file.registers[22][18] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\soc_inst.cpu_core.register_file.registers[12][13] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\soc_inst.cpu_core.register_file.registers[19][28] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\soc_inst.cpu_core.register_file.registers[12][20] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\soc_inst.cpu_core.register_file.registers[12][0] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\soc_inst.cpu_core.register_file.registers[12][5] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\soc_inst.cpu_core.register_file.registers[29][4] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\soc_inst.cpu_core.register_file.registers[19][13] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\soc_inst.cpu_core.register_file.registers[22][9] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\soc_inst.cpu_core.register_file.registers[27][19] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\soc_inst.cpu_core.register_file.registers[20][13] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\soc_inst.cpu_core.register_file.registers[25][28] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\soc_inst.cpu_core.register_file.registers[27][0] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\soc_inst.cpu_core.register_file.registers[28][7] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold1536 (.A(_00233_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\soc_inst.cpu_core.register_file.registers[31][17] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\soc_inst.cpu_core.register_file.registers[10][2] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\soc_inst.cpu_core.register_file.registers[28][4] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\soc_inst.cpu_core.register_file.registers[25][20] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\soc_inst.cpu_core.register_file.registers[25][15] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\soc_inst.cpu_core.register_file.registers[29][30] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\soc_inst.spi_inst.rx_shift_reg[19] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\soc_inst.cpu_core.register_file.registers[25][11] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\soc_inst.cpu_core.register_file.registers[12][26] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\soc_inst.cpu_core.register_file.registers[30][11] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\soc_inst.cpu_core.register_file.registers[6][26] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\soc_inst.cpu_core.mem_rs1_data[28] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\soc_inst.cpu_core.register_file.registers[10][5] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\soc_inst.cpu_core.register_file.registers[6][7] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\soc_inst.cpu_core.register_file.registers[10][25] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\soc_inst.cpu_core.register_file.registers[3][0] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\soc_inst.cpu_core.register_file.registers[27][12] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\soc_inst.cpu_core.register_file.registers[5][13] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\soc_inst.cpu_core.register_file.registers[20][15] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\soc_inst.cpu_core.register_file.registers[6][31] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\soc_inst.cpu_core.register_file.registers[12][10] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\soc_inst.cpu_core.register_file.registers[18][1] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[5] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold1560 (.A(_08643_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\soc_inst.cpu_core.register_file.registers[31][0] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_00274_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\soc_inst.cpu_core.register_file.registers[3][3] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\soc_inst.cpu_core.register_file.registers[7][28] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\soc_inst.cpu_core.register_file.registers[25][23] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[5] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_02592_),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\soc_inst.cpu_core.register_file.registers[5][23] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[0] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_02532_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\soc_inst.cpu_core.register_file.registers[25][6] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\soc_inst.cpu_core.register_file.registers[15][26] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\soc_inst.cpu_core.id_instr[10] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\soc_inst.cpu_core.register_file.registers[30][2] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\soc_inst.cpu_core.register_file.registers[9][16] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[1] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold1577 (.A(_02567_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\soc_inst.cpu_core.register_file.registers[3][31] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\soc_inst.cpu_core.register_file.registers[28][30] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\soc_inst.cpu_core.register_file.registers[6][25] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\soc_inst.cpu_core.register_file.registers[29][8] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\soc_inst.cpu_core.register_file.registers[6][14] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\soc_inst.cpu_core.register_file.registers[31][2] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\soc_inst.cpu_core.register_file.registers[6][13] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\soc_inst.cpu_core.mem_rs1_data[5] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\soc_inst.cpu_core.register_file.registers[12][2] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\soc_inst.cpu_core.register_file.registers[7][1] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\soc_inst.cpu_core.register_file.registers[3][30] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\soc_inst.cpu_core.ex_exception_pc[23] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold1590 (.A(_01249_),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[19] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold1592 (.A(_00738_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\soc_inst.cpu_core.ex_exception_pc[0] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_01226_),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\soc_inst.cpu_core.register_file.registers[26][12] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\soc_inst.cpu_core.register_file.registers[5][26] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\soc_inst.cpu_core.register_file.registers[27][24] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\soc_inst.i2c_inst.ctrl_reg[4] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00245_),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold1600 (.A(_00420_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\soc_inst.cpu_core.register_file.registers[7][12] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\soc_inst.cpu_core.register_file.registers[6][17] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\soc_inst.cpu_core.register_file.registers[6][12] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\soc_inst.cpu_core.register_file.registers[3][10] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\soc_inst.cpu_core.register_file.registers[20][8] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\soc_inst.cpu_core.register_file.registers[9][19] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\soc_inst.cpu_core.register_file.registers[25][21] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\soc_inst.cpu_core.register_file.registers[21][0] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\soc_inst.cpu_core.register_file.registers[31][10] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\soc_inst.cpu_core.register_file.registers[10][29] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\soc_inst.cpu_core.register_file.registers[5][31] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\soc_inst.cpu_core.register_file.registers[5][14] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\soc_inst.cpu_core.register_file.registers[3][15] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\soc_inst.cpu_core.register_file.registers[28][15] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\soc_inst.cpu_core.register_file.registers[31][6] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\soc_inst.cpu_core.register_file.registers[9][29] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[6] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\soc_inst.cpu_core.ex_exception_pc[7] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold1619 (.A(_01233_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\soc_inst.cpu_core.register_file.registers[6][23] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\soc_inst.cpu_core.register_file.registers[30][6] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\soc_inst.cpu_core.register_file.registers[21][20] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\soc_inst.cpu_core.register_file.registers[29][20] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold1624 (.A(_00268_),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_02477_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\soc_inst.cpu_core.register_file.registers[25][18] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\soc_inst.cpu_core.register_file.registers[6][6] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\soc_inst.cpu_core.register_file.registers[30][25] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\soc_inst.cpu_core.register_file.registers[21][1] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\soc_inst.cpu_core.csr_file.mscratch[31] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\soc_inst.cpu_core.register_file.registers[12][24] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\soc_inst.cpu_core.register_file.registers[9][21] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[5] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\soc_inst.cpu_core.register_file.registers[6][27] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\soc_inst.cpu_core.register_file.registers[23][28] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\soc_inst.cpu_core.register_file.registers[27][27] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\soc_inst.cpu_core.mem_rs1_data[17] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\soc_inst.cpu_core.register_file.registers[26][0] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\soc_inst.i2c_inst.shift_reg[1] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold1640 (.A(_00098_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\soc_inst.cpu_core.register_file.registers[27][28] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\soc_inst.cpu_core.register_file.registers[5][24] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\soc_inst.cpu_core.register_file.registers[10][31] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\soc_inst.spi_inst.rx_shift_reg[17] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\soc_inst.cpu_core.register_file.registers[3][1] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\soc_inst.cpu_core.register_file.registers[26][19] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\soc_inst.cpu_core.id_rs2_data[11] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\soc_inst.cpu_core.register_file.registers[19][30] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\soc_inst.cpu_core.register_file.registers[5][18] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\soc_inst.cpu_core.register_file.registers[19][21] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\soc_inst.pwm_inst.channel_duty[0][4] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\soc_inst.cpu_core.csr_file.mscratch[4] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\soc_inst.cpu_core.register_file.registers[25][7] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\soc_inst.cpu_core.register_file.registers[10][12] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\soc_inst.cpu_core.register_file.registers[1][16] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\soc_inst.cpu_core.register_file.registers[6][11] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\soc_inst.cpu_core.register_file.registers[22][29] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\soc_inst.spi_inst.tx_shift_reg[28] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\soc_inst.cpu_core.mem_rs1_data[2] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold1660 (.A(_00934_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\soc_inst.cpu_core.register_file.registers[31][9] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\soc_inst.cpu_core.register_file.registers[3][14] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[8] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold1664 (.A(_07757_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold1665 (.A(_02595_),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[5] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_00691_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\soc_inst.cpu_core.register_file.registers[12][9] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\soc_inst.cpu_core.if_pc[5] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold1670 (.A(_02457_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\soc_inst.cpu_core.register_file.registers[25][31] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\soc_inst.cpu_core.register_file.registers[31][25] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\soc_inst.cpu_core.register_file.registers[9][4] ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\soc_inst.cpu_core.register_file.registers[10][27] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\soc_inst.cpu_core.register_file.registers[5][3] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\soc_inst.cpu_core.register_file.registers[6][15] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\soc_inst.cpu_core.ex_funct3[2] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\soc_inst.cpu_core.register_file.registers[23][20] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold1679 (.A(_00289_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\soc_inst.cpu_core.register_file.registers[28][10] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold1681 (.A(_00241_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\soc_inst.cpu_core.register_file.registers[19][12] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\soc_inst.cpu_core.register_file.registers[21][28] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\soc_inst.cpu_core.register_file.registers[6][19] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\soc_inst.cpu_core.ex_exception_pc[19] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_01245_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\soc_inst.cpu_core.register_file.registers[25][19] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\soc_inst.cpu_core.register_file.registers[7][13] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\soc_inst.cpu_core.register_file.registers[12][14] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\soc_inst.spi_inst.tx_shift_reg[15] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\soc_inst.cpu_core.register_file.registers[30][19] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\soc_inst.cpu_core.register_file.registers[9][27] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\soc_inst.cpu_core.mem_rs1_data[19] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\soc_inst.cpu_core.register_file.registers[19][9] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\soc_inst.cpu_core.register_file.registers[19][0] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[10] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_08655_),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold1698 (.A(_00244_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\soc_inst.cpu_core.ex_exception_pc[17] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold1700 (.A(_01243_),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\soc_inst.cpu_core.register_file.registers[22][30] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\soc_inst.cpu_core.register_file.registers[22][22] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\soc_inst.cpu_core.register_file.registers[22][15] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\soc_inst.cpu_core.csr_file.mscratch[2] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\soc_inst.cpu_core.ex_branch_target[2] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_02344_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\soc_inst.cpu_core.mem_rs1_data[4] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\soc_inst.cpu_core.mem_rs1_data[16] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\soc_inst.cpu_core.register_file.registers[5][12] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\soc_inst.cpu_core.register_file.registers[12][23] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\soc_inst.cpu_core.register_file.registers[27][20] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\soc_inst.cpu_core.register_file.registers[3][6] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\soc_inst.cpu_core.register_file.registers[23][30] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\soc_inst.cpu_core.register_file.registers[6][22] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\soc_inst.cpu_core.register_file.registers[21][11] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\soc_inst.cpu_core.ex_rs2_data[30] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold1717 (.A(_01344_),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\soc_inst.cpu_core.register_file.registers[10][14] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\soc_inst.cpu_core.register_file.registers[25][13] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\soc_inst.cpu_core.ex_rs2_data[12] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_01326_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\soc_inst.cpu_core.ex_exception_pc[21] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_01247_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\soc_inst.cpu_core.register_file.registers[19][5] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\soc_inst.cpu_core.register_file.registers[10][10] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\soc_inst.cpu_core.csr_file.mscratch[1] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\soc_inst.cpu_core.register_file.registers[30][17] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[17] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_00736_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\soc_inst.cpu_core.register_file.registers[23][19] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\soc_inst.cpu_core.register_file.registers[3][7] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\soc_inst.cpu_core.register_file.registers[31][8] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold1734 (.A(_00477_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\soc_inst.cpu_core.register_file.registers[6][2] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\soc_inst.cpu_core.register_file.registers[29][7] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\soc_inst.cpu_core.register_file.registers[31][18] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\soc_inst.cpu_core.register_file.registers[26][29] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\soc_inst.cpu_core.register_file.registers[7][26] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\soc_inst.cpu_core.register_file.registers[21][18] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\soc_inst.cpu_core.register_file.registers[10][8] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\soc_inst.cpu_core.register_file.registers[26][8] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\soc_inst.cpu_core.ex_exception_pc[15] ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold1744 (.A(_01241_),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\soc_inst.cpu_core.register_file.registers[19][25] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\soc_inst.core_mem_wdata[12] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold1747 (.A(_02488_),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\soc_inst.cpu_core.register_file.registers[19][11] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\soc_inst.cpu_core.register_file.registers[21][9] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_00240_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\soc_inst.cpu_core.register_file.registers[21][16] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_00260_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold1753 (.A(_01032_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\soc_inst.cpu_core.register_file.registers[3][2] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\soc_inst.cpu_core.register_file.registers[26][30] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\soc_inst.cpu_core.id_instr[11] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\soc_inst.i2c_inst.shift_reg[2] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold1758 (.A(_00099_),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.rxd_reg ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold1760 (.A(_02586_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\soc_inst.cpu_core.register_file.registers[28][6] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\soc_inst.cpu_core.if_instr[17] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[2] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold1764 (.A(_00020_),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\soc_inst.cpu_core.register_file.registers[25][26] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\soc_inst.spi_inst.rx_shift_reg[22] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\soc_inst.cpu_core.register_file.registers[30][5] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\soc_inst.cpu_core.register_file.registers[22][19] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\soc_inst.core_instr_data[30] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold1770 (.A(_00603_),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\soc_inst.cpu_core.register_file.registers[19][7] ),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\soc_inst.cpu_core.register_file.registers[29][16] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\soc_inst.cpu_core.register_file.registers[21][3] ),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\soc_inst.cpu_core.ex_exception_pc[22] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold1775 (.A(_01248_),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold1776 (.A(_00298_),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold1777 (.A(_02515_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\soc_inst.cpu_core.csr_file.mtime[45] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\soc_inst.cpu_core.if_instr[15] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\soc_inst.cpu_core.register_file.registers[29][22] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[1] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold1782 (.A(_07682_),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold1783 (.A(_02542_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\soc_inst.cpu_core.register_file.registers[29][19] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\soc_inst.cpu_core.id_instr[19] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold1786 (.A(_01213_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\soc_inst.cpu_core.register_file.registers[28][12] ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\soc_inst.cpu_core.ex_exception_pc[13] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold1789 (.A(_01239_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\soc_inst.cpu_core.register_file.registers[28][11] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\soc_inst.cpu_core.register_file.registers[29][11] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\soc_inst.cpu_core.register_file.registers[29][6] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\soc_inst.cpu_core.register_file.registers[27][25] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\soc_inst.cpu_core.register_file.registers[26][4] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\soc_inst.cpu_core.register_file.registers[21][12] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\soc_inst.cpu_core.register_file.registers[30][31] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\soc_inst.cpu_core.register_file.registers[30][1] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\soc_inst.cpu_core.register_file.registers[7][4] ),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\soc_inst.cpu_core.register_file.registers[28][14] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\soc_inst.cpu_core.register_file.registers[3][18] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\soc_inst.cpu_core.register_file.registers[21][26] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\soc_inst.cpu_core.ex_exception_pc[8] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold1803 (.A(_01234_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\soc_inst.cpu_core.register_file.registers[30][20] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\soc_inst.cpu_core.register_file.registers[22][10] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\soc_inst.cpu_core.register_file.registers[9][25] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold1807 (.A(_00252_),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold1808 (.A(_00875_),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[3] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold1810 (.A(_07740_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold1811 (.A(_02585_),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\soc_inst.cpu_core.register_file.registers[21][7] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\soc_inst.cpu_core.register_file.registers[12][3] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\soc_inst.cpu_core.mem_rs1_data[1] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\soc_inst.cpu_core.register_file.registers[7][15] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\soc_inst.cpu_core.register_file.registers[3][17] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\soc_inst.cpu_core.register_file.registers[26][16] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\soc_inst.cpu_core.register_file.registers[7][29] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\soc_inst.cpu_core.register_file.registers[22][21] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\soc_inst.cpu_core.register_file.registers[7][16] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\soc_inst.cpu_core.register_file.registers[26][14] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\soc_inst.spi_inst.clk_counter[3] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_00131_),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\soc_inst.cpu_core.register_file.registers[27][5] ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\soc_inst.cpu_core.ex_branch_target[31] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_02373_),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\soc_inst.cpu_core.if_instr[7] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\soc_inst.cpu_core.register_file.registers[7][6] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\soc_inst.cpu_core.register_file.registers[26][18] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\soc_inst.cpu_core.register_file.registers[13][13] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold1831 (.A(_00239_),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\soc_inst.cpu_core.register_file.registers[25][30] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\soc_inst.i2c_inst.shift_reg[6] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold1834 (.A(_00103_),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\soc_inst.cpu_core.register_file.registers[3][13] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\soc_inst.cpu_core.register_file.registers[31][3] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\soc_inst.cpu_core.register_file.registers[31][1] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\soc_inst.cpu_core.register_file.registers[21][22] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\soc_inst.cpu_core.register_file.registers[3][27] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\soc_inst.cpu_core.register_file.registers[25][0] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\soc_inst.cpu_core.register_file.registers[30][14] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\soc_inst.cpu_core.register_file.registers[9][26] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\soc_inst.cpu_core.register_file.registers[21][15] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\soc_inst.cpu_core.ex_exception_pc[3] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold1845 (.A(_01229_),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\soc_inst.cpu_core.register_file.registers[23][21] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\soc_inst.cpu_core.register_file.registers[7][9] ),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\soc_inst.core_mem_addr[9] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold1849 (.A(_01291_),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[1] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold1851 (.A(_00720_),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold1852 (.A(_00306_),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\soc_inst.cpu_core.register_file.registers[26][9] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\soc_inst.cpu_core.register_file.registers[19][6] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold1855 (.A(_00226_),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold1856 (.A(_00393_),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\soc_inst.cpu_core.mem_rs1_data[0] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\soc_inst.cpu_core.register_file.registers[7][17] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\soc_inst.cpu_core.register_file.registers[19][26] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\soc_inst.cpu_core.register_file.registers[31][27] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\soc_inst.cpu_core.register_file.registers[27][10] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\soc_inst.cpu_core.register_file.registers[26][25] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\soc_inst.cpu_core.register_file.registers[25][2] ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\soc_inst.cpu_core.register_file.registers[9][30] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\soc_inst.cpu_core.register_file.registers[25][27] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\soc_inst.cpu_core.register_file.registers[12][29] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\soc_inst.cpu_core.if_pc[6] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold1868 (.A(_02458_),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\soc_inst.cpu_core.register_file.registers[29][25] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\soc_inst.cpu_core.register_file.registers[22][0] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\soc_inst.spi_inst.tx_shift_reg[20] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[0] ),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold1873 (.A(_00719_),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\soc_inst.cpu_core.register_file.registers[19][4] ),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\soc_inst.cpu_core.register_file.registers[12][12] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\soc_inst.cpu_core.register_file.registers[5][4] ),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\soc_inst.cpu_core.register_file.registers[23][25] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\soc_inst.cpu_core.register_file.registers[29][18] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\soc_inst.core_mem_rdata[25] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold1880 (.A(_00630_),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\soc_inst.cpu_core.register_file.registers[12][7] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\soc_inst.cpu_core.register_file.registers[31][28] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\soc_inst.cpu_core.register_file.registers[7][19] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\soc_inst.cpu_core.register_file.registers[23][1] ),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\soc_inst.cpu_core.register_file.registers[30][24] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\soc_inst.cpu_core.register_file.registers[12][25] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\soc_inst.cpu_core.csr_file.mepc[17] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\soc_inst.core_mem_rdata[2] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold1889 (.A(_00607_),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\soc_inst.cpu_core.register_file.registers[29][1] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\soc_inst.cpu_core.register_file.registers[23][2] ),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\soc_inst.cpu_core.register_file.registers[19][19] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\soc_inst.cpu_core.register_file.registers[19][8] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\soc_inst.cpu_core.register_file.registers[29][3] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\soc_inst.cpu_core.register_file.registers[25][12] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\soc_inst.cpu_core.register_file.registers[10][15] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\soc_inst.cpu_core.ex_rs2_data[20] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_01334_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\soc_inst.cpu_core.register_file.registers[27][29] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\soc_inst.cpu_core.register_file.registers[30][18] ),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\soc_inst.cpu_core.csr_file.mtime[28] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold1902 (.A(_00193_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\soc_inst.cpu_core.mem_instr[2] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_01030_),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\soc_inst.cpu_core.register_file.registers[28][19] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\soc_inst.core_mem_rdata[1] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_00606_),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\soc_inst.gpio_inst.gpio_out[1] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold1909 (.A(_00462_),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\soc_inst.cpu_core.register_file.registers[9][23] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\soc_inst.cpu_core.register_file.registers[5][11] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\soc_inst.cpu_core.register_file.registers[25][5] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[3] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold1914 (.A(_02569_),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[3] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold1916 (.A(_02495_),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold1917 (.A(_00295_),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\soc_inst.cpu_core.register_file.registers[5][9] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\soc_inst.core_mem_rdata[16] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold1920 (.A(_00621_),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\soc_inst.cpu_core.register_file.registers[6][20] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\soc_inst.cpu_core.register_file.registers[21][24] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold1923 (.A(_00285_),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold1924 (.A(_02502_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\soc_inst.cpu_core.register_file.registers[5][0] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\soc_inst.cpu_core.ex_branch_target[16] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\soc_inst.cpu_core.register_file.registers[25][25] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\soc_inst.cpu_core.register_file.registers[26][28] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\soc_inst.spi_inst.tx_shift_reg[25] ),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[1] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold1931 (.A(_02575_),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\soc_inst.cpu_core.csr_file.mtime[46] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\soc_inst.cpu_core.register_file.registers[7][2] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold1934 (.A(_00253_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold1935 (.A(_00876_),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[4] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold1937 (.A(_02496_),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\soc_inst.i2c_inst.shift_reg[3] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold1939 (.A(_00100_),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\soc_inst.cpu_core.register_file.registers[5][1] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\soc_inst.cpu_core.register_file.registers[25][3] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold1942 (.A(_00272_),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\soc_inst.cpu_core.ex_instr[10] ),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_in[11] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\soc_inst.spi_inst.len_sel[0] ),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold1946 (.A(_00425_),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\soc_inst.cpu_core.register_file.registers[6][0] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\soc_inst.cpu_core.register_file.registers[21][4] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\soc_inst.cpu_core.register_file.registers[10][28] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\soc_inst.cpu_core.register_file.registers[12][30] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold1951 (.A(_00228_),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\soc_inst.cpu_core.register_file.registers[27][3] ),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\soc_inst.cpu_core.register_file.registers[26][23] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\soc_inst.cpu_core.register_file.registers[31][4] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\soc_inst.cpu_core.register_file.registers[29][26] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\soc_inst.cpu_core.alu.a[2] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold1957 (.A(_00247_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold1958 (.A(_00267_),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_02476_),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold1960 (.A(_00246_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\soc_inst.cpu_core.register_file.registers[9][31] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\soc_inst.cpu_core.register_file.registers[10][6] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\soc_inst.cpu_core.register_file.registers[30][0] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\soc_inst.cpu_core.ex_rs1_data[2] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold1965 (.A(_01252_),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\soc_inst.cpu_core.register_file.registers[29][9] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\soc_inst.cpu_core.if_pc[4] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_02456_),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\soc_inst.cpu_core.register_file.registers[23][8] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\soc_inst.i2c_inst.shift_reg[7] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold1971 (.A(_00104_),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\soc_inst.cpu_core.register_file.registers[23][29] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[9] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold1974 (.A(_00728_),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\soc_inst.cpu_core.register_file.registers[29][5] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold1976 (.A(_00249_),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold1977 (.A(_00424_),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\soc_inst.cpu_core.register_file.registers[27][9] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\soc_inst.cpu_core.csr_file.mtime[37] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\soc_inst.cpu_core.register_file.registers[23][0] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\soc_inst.core_mem_rdata[22] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold1982 (.A(_00627_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold1983 (.A(_00237_),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[3] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1985 (.A(_00722_),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1986 (.A(_00224_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\soc_inst.cpu_core.register_file.registers[30][22] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\soc_inst.cpu_core.register_file.registers[9][1] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\soc_inst.cpu_core.register_file.registers[12][8] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\soc_inst.cpu_core.register_file.registers[26][3] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\soc_inst.cpu_core.register_file.registers[3][12] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\soc_inst.cpu_core.register_file.registers[22][31] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\soc_inst.cpu_core.alu.b[24] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\soc_inst.i2c_inst.clk_cnt[3] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_08862_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\soc_inst.cpu_core.csr_file.mtime[26] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1997 (.A(_00191_),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\soc_inst.cpu_core.csr_file.mepc[12] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\soc_inst.cpu_core.if_pc[21] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold2000 (.A(_02473_),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold2001 (.A(_00273_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\soc_inst.cpu_core.register_file.registers[3][20] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\soc_inst.cpu_core.register_file.registers[22][23] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\soc_inst.spi_inst.bit_counter[1] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold2005 (.A(_09380_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold2006 (.A(_00339_),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\soc_inst.i2c_inst.shift_reg[4] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold2008 (.A(_00101_),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\soc_inst.cpu_core.register_file.registers[27][30] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[0] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold2011 (.A(_02582_),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\soc_inst.cpu_core.register_file.registers[5][21] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\soc_inst.cpu_core.register_file.registers[28][26] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\soc_inst.cpu_core.if_pc[1] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold2015 (.A(_02453_),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold2016 (.A(_00221_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold2017 (.A(_00378_),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\soc_inst.cpu_core.register_file.registers[12][31] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\soc_inst.cpu_core.ex_funct7[5] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold2020 (.A(_01054_),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\soc_inst.cpu_core.register_file.registers[12][15] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\soc_inst.cpu_core.register_file.registers[25][8] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\soc_inst.cpu_core.ex_exception_pc[9] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold2024 (.A(_01235_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\soc_inst.cpu_core.register_file.registers[7][21] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\soc_inst.mem_ctrl.spi_data_out[28] ),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[0] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\soc_inst.cpu_core.register_file.registers[22][16] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\soc_inst.cpu_core.register_file.registers[19][14] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\soc_inst.cpu_core.register_file.registers[31][30] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold2031 (.A(_00284_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold2032 (.A(_02501_),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[3] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\soc_inst.cpu_core.mem_rs1_data[6] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\soc_inst.cpu_core.csr_file.mepc[16] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold2036 (.A(_02433_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\soc_inst.cpu_core.register_file.registers[12][19] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[8] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold2039 (.A(_00727_),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\soc_inst.cpu_core.register_file.registers[22][25] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\soc_inst.cpu_core.register_file.registers[27][11] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\soc_inst.cpu_core.register_file.registers[21][5] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_00238_),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\soc_inst.cpu_core.register_file.registers[22][27] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\soc_inst.cpu_core.register_file.registers[30][21] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\soc_inst.cpu_core.register_file.registers[31][29] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\soc_inst.cpu_core.register_file.registers[21][23] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\soc_inst.cpu_core.register_file.registers[26][5] ),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\soc_inst.cpu_core.ex_mem_we ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold2050 (.A(_05588_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\soc_inst.cpu_core.ex_instr[11] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\soc_inst.cpu_core.register_file.registers[27][1] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\soc_inst.cpu_core.register_file.registers[5][10] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\soc_inst.cpu_core.csr_file.mepc[22] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_02439_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\soc_inst.cpu_core.csr_file.mtime[32] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold2057 (.A(_00198_),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\soc_inst.core_mem_rdata[8] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold2059 (.A(_00613_),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\soc_inst.cpu_core.register_file.registers[26][10] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\soc_inst.cpu_core.register_file.registers[10][24] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold2062 (.A(_00250_),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold2063 (.A(_00783_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold2064 (.A(_00234_),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_00409_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\soc_inst.cpu_core.mem_rs1_data[25] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\soc_inst.cpu_core.register_file.registers[31][14] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\soc_inst.cpu_core.register_file.registers[10][17] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\soc_inst.cpu_core.register_file.registers[19][29] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\soc_inst.cpu_core.register_file.registers[12][1] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\soc_inst.cpu_core.csr_file.mtvec[1] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_00517_),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\soc_inst.cpu_core.register_file.registers[3][28] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\soc_inst.cpu_core.id_instr[9] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold2075 (.A(_01203_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\soc_inst.cpu_core.register_file.registers[6][18] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\soc_inst.spi_inst.rx_shift_reg[12] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold2078 (.A(_09403_),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold2079 (.A(_00231_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\soc_inst.cpu_core.register_file.registers[23][15] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold2081 (.A(_00283_),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold2082 (.A(_02500_),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\soc_inst.cpu_core.register_file.registers[30][30] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\soc_inst.cpu_core.register_file.registers[7][30] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\soc_inst.cpu_core.register_file.registers[26][15] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\soc_inst.cpu_core.register_file.registers[22][26] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\soc_inst.cpu_core.register_file.registers[31][12] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\soc_inst.cpu_core.register_file.registers[29][0] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\soc_inst.cpu_core.register_file.registers[27][7] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\soc_inst.cpu_core.register_file.registers[28][5] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\soc_inst.cpu_core.register_file.registers[5][30] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\soc_inst.cpu_core.register_file.registers[12][21] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\soc_inst.cpu_core.register_file.registers[30][26] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\soc_inst.pwm_inst.channel_duty[0][1] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_00322_),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[5] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold2097 (.A(_02571_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\soc_inst.cpu_core.register_file.registers[23][18] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\soc_inst.cpu_core.register_file.registers[9][12] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[12] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_00731_),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold2102 (.A(_00235_),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold2103 (.A(_00410_),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\soc_inst.cpu_core.register_file.registers[23][14] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\soc_inst.cpu_core.register_file.registers[22][4] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\soc_inst.cpu_core.register_file.registers[31][7] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\soc_inst.cpu_core.register_file.registers[21][19] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\soc_inst.cpu_core.register_file.registers[28][18] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\soc_inst.cpu_core.register_file.registers[10][18] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\soc_inst.cpu_core.register_file.registers[30][28] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\soc_inst.core_mem_rdata[19] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold2112 (.A(_00624_),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\soc_inst.i2c_inst.ack_enable ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold2114 (.A(_00288_),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[2] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold2116 (.A(_02494_),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\soc_inst.cpu_core.register_file.registers[31][20] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\soc_inst.cpu_core.register_file.registers[5][5] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\soc_inst.cpu_core.register_file.registers[19][22] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\soc_inst.i2c_inst.shift_reg[5] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold2121 (.A(_00102_),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\soc_inst.cpu_core.register_file.registers[27][16] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\soc_inst.cpu_core.register_file.registers[27][21] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\soc_inst.cpu_core.register_file.registers[7][14] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\soc_inst.core_mem_rdata[17] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold2126 (.A(_00622_),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\soc_inst.spi_inst.clk_counter[5] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold2128 (.A(_08784_),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold2129 (.A(_00133_),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\soc_inst.cpu_core.register_file.registers[12][17] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\soc_inst.cpu_core.register_file.registers[28][23] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\soc_inst.cpu_core.register_file.registers[10][11] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\soc_inst.core_mem_rdata[18] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold2134 (.A(_00623_),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\soc_inst.cpu_core.register_file.registers[3][19] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\soc_inst.cpu_core.register_file.registers[9][14] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\soc_inst.cpu_core.register_file.registers[28][28] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\soc_inst.cpu_core.register_file.registers[26][1] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\soc_inst.cpu_core.register_file.registers[29][21] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\soc_inst.cpu_core.ex_exception_pc[4] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold2141 (.A(_01230_),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\soc_inst.cpu_core.mem_rs1_data[15] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\soc_inst.cpu_core.register_file.registers[5][19] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\soc_inst.cpu_core.ex_rs1_data[21] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold2145 (.A(_01271_),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\soc_inst.cpu_core.register_file.registers[10][1] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\soc_inst.cpu_core.register_file.registers[7][11] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_00294_),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold2149 (.A(_02511_),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\soc_inst.spi_inst.rx_shift_reg[10] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold2151 (.A(_09401_),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\soc_inst.cpu_core.ex_exception_pc[16] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold2153 (.A(_01242_),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\soc_inst.cpu_core.register_file.registers[31][26] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\soc_inst.cpu_core.id_funct3[2] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold2156 (.A(_00270_),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\soc_inst.cpu_core.register_file.registers[10][13] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold2158 (.A(_00222_),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\soc_inst.cpu_core.ex_branch_target[23] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\soc_inst.cpu_core.register_file.registers[23][23] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\soc_inst.cpu_core.register_file.registers[22][5] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\soc_inst.cpu_core.register_file.registers[21][14] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\soc_inst.cpu_core.register_file.registers[3][22] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\soc_inst.cpu_core.register_file.registers[10][3] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\soc_inst.i2c_inst.clk_cnt[4] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\soc_inst.cpu_core.register_file.registers[31][5] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\soc_inst.spi_inst.tx_shift_reg[13] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\soc_inst.pwm_inst.channel_duty[0][0] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold2169 (.A(_00321_),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\soc_inst.pwm_inst.channel_duty[0][3] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\soc_inst.i2c_inst.shift_reg[0] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold2172 (.A(_00097_),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\soc_inst.cpu_core.csr_file.mtval[11] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\soc_inst.cpu_core.register_file.registers[30][27] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[1] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold2176 (.A(_07690_),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\soc_inst.cpu_core.csr_file.mepc[5] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\soc_inst.cpu_core.register_file.registers[7][10] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\soc_inst.cpu_core.if_pc[8] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_02460_),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\soc_inst.cpu_core.mem_rs1_data[20] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\soc_inst.cpu_core.csr_file.mtval[10] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold2183 (.A(_02381_),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\soc_inst.cpu_core.register_file.registers[12][22] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\soc_inst.cpu_core.csr_file.mtval[7] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold2186 (.A(_02378_),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\soc_inst.cpu_core.register_file.registers[31][16] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\soc_inst.cpu_core.register_file.registers[23][12] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\soc_inst.cpu_core.register_file.registers[9][3] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\soc_inst.cpu_core.register_file.registers[9][0] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\soc_inst.cpu_core.register_file.registers[26][17] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\soc_inst.cpu_core.if_pc[7] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold2193 (.A(_02459_),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[9] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold2195 (.A(_00014_),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\soc_inst.cpu_core.mem_instr[3] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold2197 (.A(_01031_),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\soc_inst.cpu_core.register_file.registers[23][11] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\soc_inst.cpu_core.register_file.registers[30][23] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold2200 (.A(_00287_),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\soc_inst.cpu_core.register_file.registers[9][6] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\soc_inst.cpu_core.if_instr[19] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\soc_inst.cpu_core.mem_instr[18] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold2204 (.A(_01042_),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold2205 (.A(_00286_),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\soc_inst.cpu_core.register_file.registers[22][28] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\soc_inst.cpu_core.id_imm12[4] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold2208 (.A(_01218_),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\soc_inst.cpu_core.register_file.registers[29][2] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\soc_inst.cpu_core.register_file.registers[27][4] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\soc_inst.cpu_core.register_file.registers[22][14] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\soc_inst.cpu_core.register_file.registers[10][26] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold2214 (.A(_01237_),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\soc_inst.cpu_core.register_file.registers[26][21] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[2] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold2217 (.A(_00721_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\soc_inst.gpio_inst.gpio_out[0] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold2219 (.A(_00461_),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\soc_inst.cpu_core.ex_alu_result[16] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\soc_inst.cpu_core.register_file.registers[28][3] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold2222 (.A(_00258_),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold2223 (.A(_01028_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\soc_inst.cpu_core.ex_branch_target[26] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold2225 (.A(_02368_),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\soc_inst.cpu_core.register_file.registers[26][2] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold2227 (.A(_00227_),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold2228 (.A(_00394_),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\soc_inst.cpu_core.register_file.registers[22][3] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold2230 (.A(_00271_),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold2231 (.A(_00296_),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\soc_inst.cpu_core.register_file.registers[22][1] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\soc_inst.cpu_core.csr_file.mtval[5] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold2234 (.A(_02376_),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\soc_inst.cpu_core.register_file.registers[25][29] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\soc_inst.core_mem_rdata[28] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold2237 (.A(_00633_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_00248_),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\soc_inst.cpu_core.csr_file.mtime[27] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold2240 (.A(_00192_),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\soc_inst.cpu_core.register_file.registers[6][29] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\soc_inst.cpu_core.register_file.registers[26][31] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[1] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold2244 (.A(_00408_),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\soc_inst.cpu_core.if_pc[3] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold2246 (.A(_02455_),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\soc_inst.cpu_core.register_file.registers[19][10] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\soc_inst.spi_inst.rx_shift_reg[4] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold2249 (.A(_09395_),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.uart_tx_data[4] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\soc_inst.cpu_core.register_file.registers[3][4] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\soc_inst.cpu_core.register_file.registers[30][8] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.fsm_state[3] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\soc_inst.core_mem_rdata[26] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold2255 (.A(_00631_),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[20] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold2257 (.A(_00739_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\soc_inst.cpu_core.mem_rs1_data[22] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\soc_inst.cpu_core.ex_funct7[1] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold2260 (.A(_01220_),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[2] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold2262 (.A(_07692_),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\soc_inst.cpu_core.if_pc[11] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold2264 (.A(_00918_),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\soc_inst.core_mem_rdata[9] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\soc_inst.cpu_core.id_instr[8] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\soc_inst.cpu_core.csr_file.mepc[13] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold2268 (.A(_02430_),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\soc_inst.pwm_inst.channel_duty[0][2] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\soc_inst.cpu_core.if_pc[17] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold2271 (.A(_00924_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\soc_inst.cpu_core.register_file.registers[23][17] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\soc_inst.cpu_core.register_file.registers[31][19] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\soc_inst.core_mem_rdata[6] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold2275 (.A(_10493_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\soc_inst.i2c_inst.data_reg[2] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\soc_inst.cpu_core.ex_exception_pc[2] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold2278 (.A(_01228_),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\soc_inst.cpu_core.id_rs2_data[31] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\soc_inst.cpu_core.register_file.registers[25][17] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[5] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold2282 (.A(_00724_),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold2283 (.A(_00293_),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold2284 (.A(_00276_),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\soc_inst.cpu_core.register_file.registers[31][13] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\soc_inst.core_mem_addr[15] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold2287 (.A(_01297_),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\soc_inst.cpu_core.register_file.registers[30][13] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\soc_inst.cpu_core.ex_exception_pc[1] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold2290 (.A(_01227_),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\soc_inst.cpu_core.register_file.registers[7][8] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\soc_inst.cpu_core.ex_funct7[4] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold2293 (.A(_01223_),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold2294 (.A(_00278_),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold2295 (.A(_02487_),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\soc_inst.i2c_inst.data_reg[3] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\soc_inst.cpu_core.register_file.registers[22][12] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\soc_inst.cpu_core.register_file.registers[28][2] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\soc_inst.i2c_inst.data_reg[7] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\soc_inst.core_mem_rdata[27] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold2301 (.A(_00632_),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\soc_inst.cpu_core.csr_file.mtvec[4] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\soc_inst.cpu_core.if_pc[22] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold2304 (.A(_00929_),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\soc_inst.cpu_core.mem_instr[16] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold2306 (.A(_01040_),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[0] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold2308 (.A(_02492_),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\soc_inst.cpu_core.csr_file.mtime[20] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold2310 (.A(_00185_),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\soc_inst.cpu_core.mem_rs1_data[7] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\soc_inst.spi_inst.rx_shift_reg[23] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\soc_inst.cpu_core.register_file.registers[25][24] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\soc_inst.cpu_core.ex_funct7[2] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold2315 (.A(_01051_),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\soc_inst.cpu_core.register_file.registers[6][4] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\soc_inst.cpu_core.csr_file.mtval[9] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\soc_inst.spi_inst.rx_shift_reg[9] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold2319 (.A(_09400_),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\soc_inst.cpu_core.register_file.registers[7][0] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\soc_inst.cpu_core.if_pc[16] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold2322 (.A(_00923_),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\soc_inst.core_instr_data[22] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold2324 (.A(_00595_),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\soc_inst.cpu_core.register_file.registers[6][5] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\soc_inst.pwm_inst.channel_duty[0][14] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[0] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold2328 (.A(_07678_),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold2329 (.A(_02541_),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\soc_inst.mem_ctrl.spi_data_out[26] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\soc_inst.mem_ctrl.spi_data_out[29] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\soc_inst.cpu_core.if_pc[15] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold2333 (.A(_00922_),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold2334 (.A(_00281_),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\soc_inst.cpu_core.ex_branch_target[30] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold2336 (.A(_02372_),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\soc_inst.cpu_core.id_instr[7] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold2338 (.A(_01201_),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold2339 (.A(_00263_),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold2340 (.A(_01198_),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.bit_counter[1] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\soc_inst.cpu_core.register_file.registers[26][22] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\soc_inst.cpu_core.register_file.registers[19][31] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[7] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold2345 (.A(_00726_),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\soc_inst.pwm_inst.channel_duty[0][7] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\soc_inst.cpu_core.id_imm[8] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold2348 (.A(_01096_),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\soc_inst.spi_inst.bit_counter[3] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold2350 (.A(_09384_),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold2351 (.A(_00341_),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\soc_inst.pwm_inst.channel_duty[0][13] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[2] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold2354 (.A(_02543_),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\soc_inst.cpu_core.ex_branch_target[0] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold2356 (.A(_02342_),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\soc_inst.core_instr_data[25] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold2358 (.A(_00598_),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\soc_inst.spi_inst.rx_shift_reg[6] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold2360 (.A(_09397_),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\soc_inst.cpu_core.register_file.registers[28][1] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\soc_inst.cpu_core.ex_branch_target[19] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold2363 (.A(_02361_),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\soc_inst.cpu_core.register_file.registers[29][12] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold2365 (.A(\soc_inst.cpu_core.csr_file.csr_addr[6] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\soc_inst.cpu_core.mem_rs1_data[21] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\soc_inst.cpu_core.ex_branch_target[13] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold2368 (.A(_02355_),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\soc_inst.cpu_core.register_file.registers[31][23] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\soc_inst.cpu_core.csr_file.mepc[15] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\soc_inst.cpu_core.register_file.registers[6][28] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\soc_inst.cpu_core.if_is_compressed ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold2373 (.A(_04468_),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\soc_inst.core_instr_data[23] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold2375 (.A(_00596_),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\soc_inst.cpu_core.ex_is_ecall ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold2377 (.A(_00873_),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\soc_inst.cpu_core.register_file.registers[23][7] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\soc_inst.cpu_core.csr_file.mtval[12] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold2380 (.A(_02383_),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold2381 (.A(\soc_inst.cpu_core.csr_file.mepc[23] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold2382 (.A(_02440_),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\soc_inst.core_mem_rdata[3] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold2384 (.A(_10413_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\soc_inst.cpu_core.csr_file.mtime[16] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold2386 (.A(_00180_),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\soc_inst.gpio_inst.int_en_reg[1] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold2388 (.A(_00468_),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\soc_inst.cpu_core.register_file.registers[19][3] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\soc_inst.cpu_core.ex_branch_target[29] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold2391 (.A(_02371_),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\soc_inst.pwm_inst.channel_counter[0][10] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold2393 (.A(_08927_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold2394 (.A(_00112_),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\soc_inst.core_instr_data[24] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold2396 (.A(_00597_),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\soc_inst.cpu_core.ex_branch_target[18] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold2398 (.A(_02360_),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\soc_inst.cpu_core.id_imm[10] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold2400 (.A(_01098_),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold2401 (.A(_00255_),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\soc_inst.spi_inst.rx_shift_reg[15] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold2403 (.A(_09406_),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\soc_inst.cpu_core.if_pc[14] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold2405 (.A(_00921_),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\soc_inst.spi_inst.rx_shift_reg[14] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold2407 (.A(_09405_),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\soc_inst.cpu_core.ex_instr[21] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold2409 (.A(_01045_),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.recieved_data[7] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\soc_inst.i2c_inst.data_reg[5] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\soc_inst.cpu_core.register_file.registers[19][1] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold2413 (.A(\soc_inst.core_instr_addr[3] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\soc_inst.core_instr_addr[8] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\soc_inst.cpu_core.register_file.registers[27][14] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[8] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold2417 (.A(_07702_),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold2418 (.A(_02553_),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\soc_inst.cpu_core.register_file.registers[23][5] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\soc_inst.gpio_inst.int_en_reg[5] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\soc_inst.cpu_core.register_file.registers[7][23] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\soc_inst.cpu_core.id_imm12[1] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\soc_inst.cpu_core.csr_file.mie[11] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold2424 (.A(\soc_inst.core_instr_data[29] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold2425 (.A(_00602_),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold2426 (.A(\soc_inst.gpio_inst.int_en_reg[6] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold2427 (.A(_00275_),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\soc_inst.mem_ctrl.spi_data_out[27] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[4] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold2430 (.A(_07696_),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\soc_inst.cpu_core.csr_file.mepc[14] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\soc_inst.cpu_core.register_file.registers[28][8] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[1] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold2434 (.A(_02493_),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\soc_inst.cpu_core.register_file.registers[30][9] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold2436 (.A(\soc_inst.spi_inst.rx_shift_reg[11] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\soc_inst.cpu_core.csr_file.mtime[25] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold2438 (.A(_09342_),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold2439 (.A(_00190_),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[24] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold2441 (.A(_00743_),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.uart_rx_data[7] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\soc_inst.cpu_core.register_file.registers[23][4] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\soc_inst.cpu_core.ex_branch_target[24] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold2445 (.A(_02366_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\soc_inst.pwm_inst.channel_counter[0][4] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold2447 (.A(_08917_),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold2448 (.A(_00121_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold2449 (.A(\soc_inst.cpu_core.ex_instr[8] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\soc_inst.i2c_inst.clk_cnt[6] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold2451 (.A(_08867_),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold2452 (.A(_00095_),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\soc_inst.cpu_core.id_rs1_data[6] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold2454 (.A(\soc_inst.mem_ctrl.spi_data_out[22] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\soc_inst.cpu_core.csr_file.mepc[18] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold2456 (.A(_02435_),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\soc_inst.gpio_inst.int_en_reg[4] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\soc_inst.cpu_core.register_file.registers[29][14] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\soc_inst.mem_ctrl.spi_mem_inst.boot_mode_reg[0] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold2460 (.A(_00407_),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold2461 (.A(_00280_),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\soc_inst.core_instr_data[21] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold2463 (.A(_00594_),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold2464 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[3] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\soc_inst.cpu_core.csr_file.mtvec[0] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\soc_inst.core_mem_addr[29] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold2467 (.A(_01311_),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\soc_inst.spi_inst.rx_shift_reg[5] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\soc_inst.cpu_core.register_file.registers[23][10] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\soc_inst.core_instr_data[26] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold2471 (.A(_00599_),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\soc_inst.pwm_inst.channel_duty[0][11] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold2473 (.A(_00332_),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold2474 (.A(_00291_),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold2475 (.A(\soc_inst.spi_inst.rx_shift_reg[8] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold2476 (.A(_09399_),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold2477 (.A(\soc_inst.cpu_core.id_imm12[2] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\soc_inst.cpu_core.alu.b[22] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\soc_inst.cpu_core.if_pc[20] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold2480 (.A(_00927_),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\soc_inst.i2c_inst.clk_cnt[7] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold2482 (.A(_08869_),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\soc_inst.cpu_core.ex_is_ebreak ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\soc_inst.i2c_inst.prescale_reg[6] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold2485 (.A(\soc_inst.cpu_core.csr_file.csr_addr[8] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold2486 (.A(_01052_),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold2487 (.A(\soc_inst.cpu_core.id_imm12[10] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\soc_inst.cpu_core.id_rs2_data[8] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\soc_inst.pwm_inst.channel_duty[0][8] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\soc_inst.i2c_inst.clk_cnt[5] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\soc_inst.cpu_core.csr_file.mtime[24] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold2492 (.A(_00189_),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold2493 (.A(\soc_inst.cpu_core.csr_file.csr_addr[9] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\soc_inst.cpu_core.ex_rs2_data[25] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold2495 (.A(_01339_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\soc_inst.cpu_core.register_file.registers[21][17] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\soc_inst.core_instr_data[28] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold2498 (.A(_00601_),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\soc_inst.core_instr_data[27] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold2500 (.A(_00600_),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\soc_inst.pwm_inst.channel_duty[0][15] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold2502 (.A(_00336_),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold2503 (.A(_00259_),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold2504 (.A(_01029_),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\soc_inst.i2c_inst.data_reg[4] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold2506 (.A(\soc_inst.cpu_core.register_file.registers[29][29] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\soc_inst.cpu_core.csr_file.mepc[21] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\soc_inst.cpu_core.id_instr[6] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold2509 (.A(_01200_),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\soc_inst.core_mem_rdata[7] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold2511 (.A(\soc_inst.cpu_core.if_pc[13] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold2512 (.A(_00920_),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold2513 (.A(_00277_),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold2514 (.A(_00229_),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\soc_inst.i2c_inst.clk_cnt[1] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold2516 (.A(_00236_),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold2517 (.A(\soc_inst.cpu_core.register_file.registers[23][3] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold2518 (.A(\soc_inst.cpu_core.id_rs1_data[4] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold2519 (.A(_00230_),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\soc_inst.cpu_core.mem_rs1_data[23] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\soc_inst.spi_inst.rx_shift_reg[7] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\soc_inst.pwm_inst.channel_duty[0][12] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\soc_inst.mem_ctrl.spi_data_out[25] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold2524 (.A(_00776_),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\soc_inst.cpu_core.register_file.registers[30][12] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\soc_inst.cpu_core.alu.b[25] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\soc_inst.spi_inst.bit_counter[2] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold2528 (.A(_09383_),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold2529 (.A(_00340_),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\soc_inst.cpu_core.id_imm12[9] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold2531 (.A(_11419_),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold2532 (.A(_11420_),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold2533 (.A(_11421_),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\soc_inst.cpu_core.id_imm12[7] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold2535 (.A(\soc_inst.cpu_core.register_file.registers[26][11] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\soc_inst.core_mem_we ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\soc_inst.cpu_core.register_file.registers[12][16] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold2538 (.A(\soc_inst.cpu_core.ex_branch_target[28] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold2539 (.A(_02370_),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\soc_inst.mem_ctrl.spi_data_out[31] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\soc_inst.spi_inst.clk_counter[6] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold2542 (.A(_08786_),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold2543 (.A(_00134_),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\soc_inst.uart_instances[0].uart_inst.uart_rx_valid_reg ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold2545 (.A(_00171_),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold2546 (.A(_00243_),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold2547 (.A(\soc_inst.cpu_core.csr_file.mstatus[7] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold2548 (.A(_07568_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\soc_inst.cpu_core.id_pc[23] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold2550 (.A(_02475_),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\soc_inst.core_mem_addr[28] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold2552 (.A(_01310_),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\soc_inst.cpu_core.csr_file.mtime[29] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold2554 (.A(\soc_inst.mem_ctrl.spi_data_out[10] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\soc_inst.cpu_core.register_file.registers[9][8] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\soc_inst.i2c_inst.prescale_reg[5] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\soc_inst.core_mem_rdata[4] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold2558 (.A(_10441_),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\soc_inst.pwm_inst.channel_counter[0][2] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold2560 (.A(_08913_),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold2561 (.A(_00119_),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\soc_inst.mem_ctrl.spi_data_out[30] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold2563 (.A(_00781_),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\soc_inst.cpu_core.ex_exception_pc[18] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold2565 (.A(_01244_),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\soc_inst.core_instr_data[19] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold2567 (.A(_00592_),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\soc_inst.cpu_core.if_imm12[4] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\soc_inst.cpu_core.id_imm[4] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\soc_inst.cpu_core.if_funct7[2] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\soc_inst.cpu_core.id_rs2_data[12] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold2572 (.A(_00242_),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold2573 (.A(\soc_inst.cpu_core.register_file.registers[25][4] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold2574 (.A(\soc_inst.spi_inst.spi_sclk ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold2575 (.A(_00136_),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\soc_inst.cpu_core.register_file.registers[29][31] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\soc_inst.cpu_core.ex_alu_result[7] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold2578 (.A(\soc_inst.mem_ctrl.spi_addr[15] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold2579 (.A(_00564_),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[11] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold2581 (.A(_00016_),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\soc_inst.cpu_core.ex_instr[24] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold2583 (.A(_01048_),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[31] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold2585 (.A(_00750_),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\soc_inst.cpu_core.id_imm[31] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold2587 (.A(_01119_),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\soc_inst.core_instr_data[16] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold2589 (.A(_00589_),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\soc_inst.cpu_core.id_rs2_data[10] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold2591 (.A(_00269_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold2592 (.A(_02478_),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\soc_inst.cpu_core.mem_rs1_data[29] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold2594 (.A(_00961_),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\soc_inst.cpu_core.mem_rs1_data[24] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[7] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold2597 (.A(_07700_),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold2598 (.A(_02552_),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\soc_inst.cpu_core.alu.b[23] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\soc_inst.cpu_core.if_pc[18] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold2601 (.A(_00925_),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold2602 (.A(\soc_inst.cpu_core.ex_branch_target[25] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold2603 (.A(_02367_),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold2604 (.A(_00282_),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold2605 (.A(_02491_),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold2606 (.A(\soc_inst.core_instr_addr[1] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\soc_inst.cpu_core.register_file.registers[10][9] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\soc_inst.core_mem_addr[19] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold2609 (.A(_01301_),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\soc_inst.spi_inst.rx_shift_reg[2] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold2611 (.A(_09393_),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\soc_inst.pwm_inst.channel_counter[0][5] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold2613 (.A(_08918_),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\soc_inst.core_instr_addr[21] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\soc_inst.core_mem_addr[22] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold2616 (.A(_01304_),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\soc_inst.core_instr_data[17] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold2618 (.A(_00590_),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold2619 (.A(\soc_inst.cpu_core.id_imm12[6] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold2620 (.A(_11767_),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\soc_inst.cpu_core.mem_rs1_data[18] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold2622 (.A(\soc_inst.core_mem_addr[30] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold2623 (.A(_01312_),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\soc_inst.core_instr_addr[5] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\soc_inst.core_instr_addr[15] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold2626 (.A(_00536_),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\soc_inst.cpu_core.csr_file.mepc[7] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold2628 (.A(\soc_inst.cpu_core.id_imm[7] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[0] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold2630 (.A(\soc_inst.mem_ctrl.spi_data_out[18] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold2631 (.A(_00769_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold2632 (.A(\soc_inst.cpu_core.id_rs1_data[31] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold2633 (.A(_01027_),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold2634 (.A(\soc_inst.core_instr_addr[6] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[3] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\soc_inst.cpu_core.ex_instr[23] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold2637 (.A(_01047_),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\soc_inst.cpu_core.csr_file.mtime[18] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold2639 (.A(_00182_),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\soc_inst.cpu_core.ex_branch_target[20] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold2641 (.A(_02362_),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\soc_inst.cpu_core.ex_branch_target[10] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold2643 (.A(\soc_inst.mem_ctrl.spi_data_out[23] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\soc_inst.cpu_core.csr_file.mstatus[0] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\soc_inst.core_mem_wdata[0] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold2646 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[5] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\soc_inst.cpu_core.id_imm12[11] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold2648 (.A(_02609_),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\soc_inst.cpu_core.id_rs1_data[30] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\soc_inst.cpu_core.if_funct7[4] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold2651 (.A(\soc_inst.spi_inst.rx_shift_reg[0] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\soc_inst.core_mem_addr[24] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold2653 (.A(_01306_),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\soc_inst.core_mem_addr[26] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold2655 (.A(_01308_),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\soc_inst.cpu_core.register_file.registers[1][20] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[29] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold2658 (.A(_00748_),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\soc_inst.core_instr_addr[4] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold2660 (.A(\soc_inst.core_instr_data[1] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold2661 (.A(\soc_inst.core_instr_data[18] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\soc_inst.cpu_core.ex_branch_target[12] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold2663 (.A(_02354_),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\soc_inst.cpu_core.if_funct7[5] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\soc_inst.cpu_core.csr_file.mtvec[2] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold2666 (.A(\soc_inst.cpu_core.csr_file.mstatus[1] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.bit_counter[3] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold2668 (.A(_02544_),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\soc_inst.cpu_core.id_rs2_data[17] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\soc_inst.pwm_inst.channel_duty[0][9] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\soc_inst.cpu_core.id_rs2_data[16] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\soc_inst.mem_ctrl.access_state[4] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold2673 (.A(_00320_),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold2674 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[6] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\soc_inst.cpu_core.ex_branch_target[21] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold2676 (.A(_02363_),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold2677 (.A(\soc_inst.spi_inst.rx_shift_reg[1] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold2678 (.A(\soc_inst.core_mem_addr[27] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold2679 (.A(_01309_),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\soc_inst.mem_ctrl.spi_data_out[24] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold2681 (.A(_00775_),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold2682 (.A(\soc_inst.core_instr_data[2] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold2683 (.A(_00261_),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\soc_inst.cpu_core.if_pc[12] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold2685 (.A(_00919_),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\soc_inst.cpu_core.if_pc[19] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold2687 (.A(_00926_),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold2688 (.A(\soc_inst.cpu_core.if_pc[10] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold2689 (.A(_00917_),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\soc_inst.cpu_core.csr_file.mtime[22] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold2691 (.A(_00187_),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold2692 (.A(_00265_),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold2693 (.A(_02445_),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold2694 (.A(\soc_inst.cpu_core.csr_file.mstatus[2] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\soc_inst.cpu_core.ex_instr[5] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold2696 (.A(_01033_),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold2697 (.A(\soc_inst.mem_ctrl.spi_data_out[21] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\soc_inst.spi_inst.clk_counter[4] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold2699 (.A(_00132_),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\soc_inst.mem_ctrl.spi_data_len[3] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold2701 (.A(\soc_inst.cpu_core.ex_branch_target[9] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold2702 (.A(_02351_),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold2703 (.A(\soc_inst.gpio_inst.int_en_reg[3] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\soc_inst.gpio_inst.int_en_reg[0] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold2705 (.A(\soc_inst.cpu_core.csr_file.mstatus[4] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\soc_inst.cpu_core.ex_funct7[6] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\soc_inst.cpu_core.csr_file.mtval[8] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\soc_inst.pwm_inst.channel_counter[0][11] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold2709 (.A(_08930_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\soc_inst.cpu_core.csr_file.mtime[19] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold2711 (.A(_09330_),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold2712 (.A(_00183_),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold2713 (.A(_00264_),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold2714 (.A(_02444_),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold2715 (.A(\soc_inst.cpu_core.id_imm[6] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold2716 (.A(_01094_),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\soc_inst.cpu_core.csr_file.mepc[19] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold2718 (.A(\soc_inst.mem_ctrl.spi_addr[23] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold2719 (.A(_00572_),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\soc_inst.core_instr_data[3] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold2721 (.A(\soc_inst.cpu_core.ex_alu_result[12] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold2722 (.A(_01294_),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold2723 (.A(\soc_inst.cpu_core.id_rs2_data[19] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\soc_inst.spi_inst.clock_divider[7] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold2725 (.A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\soc_inst.core_mem_addr[20] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold2727 (.A(_01302_),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\soc_inst.core_instr_addr[7] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold2729 (.A(\soc_inst.cpu_core.csr_file.csr_addr[11] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold2730 (.A(\soc_inst.cpu_core.if_pc[0] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold2731 (.A(_02452_),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold2732 (.A(\soc_inst.spi_inst.state[0] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[28] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold2734 (.A(_11005_),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\soc_inst.cpu_core.ex_alu_result[0] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold2736 (.A(_01346_),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\soc_inst.cpu_core.id_imm[3] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold2738 (.A(_01091_),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\soc_inst.cpu_core.ex_branch_target[14] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold2740 (.A(_02356_),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold2741 (.A(\soc_inst.mem_ctrl.spi_addr[12] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold2742 (.A(_00561_),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\soc_inst.cpu_core.ex_rs1_data[29] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold2744 (.A(_01279_),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold2745 (.A(\soc_inst.pwm_inst.channel_duty[0][10] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold2746 (.A(\soc_inst.mem_ctrl.spi_mem_inst.shift_reg_out[30] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold2747 (.A(_00749_),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold2748 (.A(\soc_inst.cpu_core.csr_file.mie[7] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold2749 (.A(\soc_inst.cpu_core.alu.b[11] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\soc_inst.cpu_core.if_imm12[1] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\soc_inst.cpu_core.ex_branch_target[22] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold2752 (.A(\soc_inst.mem_ctrl.spi_addr[3] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold2753 (.A(_00552_),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold2754 (.A(_00256_),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\soc_inst.cpu_core.if_pc[9] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold2756 (.A(_00916_),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold2757 (.A(\soc_inst.core_mem_addr[18] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold2758 (.A(_01300_),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\soc_inst.cpu_core.if_funct7[0] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\soc_inst.cpu_core.ex_branch_target[8] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold2761 (.A(_02350_),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\soc_inst.cpu_core.ex_funct7[3] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold2763 (.A(_01222_),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold2764 (.A(\soc_inst.spi_inst.bit_counter[0] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold2765 (.A(\soc_inst.pwm_inst.channel_duty[0][6] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\soc_inst.cpu_core.if_imm12[2] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\soc_inst.cpu_core.id_rs1_data[7] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\soc_inst.core_mem_addr[25] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold2769 (.A(_01307_),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\soc_inst.pwm_inst.channel_duty[0][5] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\soc_inst.spi_inst.rx_shift_reg[3] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold2772 (.A(\soc_inst.mem_ctrl.spi_data_len[5] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\soc_inst.cpu_core.id_rs1_data[24] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold2774 (.A(\soc_inst.mem_ctrl.spi_mem_inst.stop ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold2775 (.A(_00004_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\soc_inst.cpu_core.id_rs2_data[4] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold2777 (.A(\soc_inst.core_mem_addr[17] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold2778 (.A(_01299_),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\soc_inst.cpu_core.id_rs1_data[3] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold2780 (.A(\soc_inst.cpu_core.ex_branch_target[15] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold2781 (.A(_02357_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\soc_inst.core_mem_wdata[15] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold2783 (.A(uio_out[5]),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold2784 (.A(_00818_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold2785 (.A(\soc_inst.i2c_inst.data_reg[1] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold2786 (.A(\soc_inst.mem_ctrl.spi_addr[14] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold2787 (.A(_00563_),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\soc_inst.core_instr_data[20] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold2789 (.A(_00593_),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\soc_inst.cpu_core.id_rs2_data[15] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold2791 (.A(\soc_inst.mem_ctrl.spi_data_out[13] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\soc_inst.cpu_core.id_rs2_data[14] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold2793 (.A(\soc_inst.pwm_inst.channel_counter[0][3] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold2794 (.A(_08914_),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold2795 (.A(\soc_inst.mem_ctrl.spi_mem_inst.spi_clk_en ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold2796 (.A(_00785_),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\soc_inst.cpu_core.ex_branch_target[4] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold2798 (.A(_00254_),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold2799 (.A(_00879_),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold2800 (.A(\soc_inst.cpu_core.ex_alu_result[21] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold2801 (.A(\soc_inst.cpu_core.id_rs2_data[9] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold2802 (.A(\soc_inst.cpu_core.id_rs2_data[13] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold2803 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[3] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold2804 (.A(_00013_),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold2805 (.A(\soc_inst.cpu_core.alu.a[3] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold2806 (.A(\soc_inst.cpu_core.id_imm12[3] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[6] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold2808 (.A(_07754_),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold2809 (.A(_00262_),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold2810 (.A(\soc_inst.core_mem_addr[21] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[0] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\soc_inst.cpu_core.csr_file.mtime[31] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold2813 (.A(_00197_),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\soc_inst.cpu_core.id_imm12[8] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold2815 (.A(_11769_),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold2816 (.A(\soc_inst.cpu_core.id_rs2_data[3] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold2817 (.A(_01059_),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold2818 (.A(\soc_inst.spi_inst.bit_counter[4] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold2819 (.A(\soc_inst.gpio_inst.int_en_reg[2] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold2820 (.A(_00469_),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold2821 (.A(\soc_inst.cpu_core.ex_alu_result[6] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold2822 (.A(\soc_inst.cpu_core.id_rs1_data[18] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold2823 (.A(\soc_inst.core_mem_addr[23] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold2824 (.A(_01305_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\soc_inst.mem_ctrl.spi_addr[1] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold2826 (.A(_00550_),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold2827 (.A(\soc_inst.cpu_core.id_imm[13] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold2828 (.A(_01101_),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold2829 (.A(\soc_inst.pwm_inst.channel_idx [0]),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold2830 (.A(_01286_),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\soc_inst.cpu_core.ex_branch_target[7] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold2832 (.A(_02349_),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\soc_inst.cpu_core.id_rs1_data[25] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold2834 (.A(\soc_inst.spi_inst.clock_divider[6] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold2835 (.A(\soc_inst.cpu_core.ex_branch_target[3] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold2836 (.A(_02345_),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\soc_inst.mem_ctrl.spi_data_out[19] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\soc_inst.mem_ctrl.spi_data_len[4] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\soc_inst.spi_inst.bit_counter[5] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold2840 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[0] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold2841 (.A(_11296_),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold2842 (.A(_00824_),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold2843 (.A(\soc_inst.spi_inst.rx_shift_reg[13] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold2844 (.A(\soc_inst.cpu_core.alu.a[6] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold2845 (.A(\soc_inst.cpu_core.if_funct3[1] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold2846 (.A(\soc_inst.core_instr_addr[18] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold2847 (.A(\soc_inst.cpu_core.alu.a[1] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold2848 (.A(\soc_inst.core_instr_addr[0] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold2849 (.A(\soc_inst.cpu_core.id_pc[13] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold2850 (.A(\soc_inst.pwm_inst.channel_counter[0][7] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold2851 (.A(_08923_),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold2852 (.A(_00124_),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[9] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold2854 (.A(_07760_),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold2855 (.A(\soc_inst.cpu_core.csr_file.mtime[21] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold2856 (.A(_09334_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold2857 (.A(\soc_inst.cpu_core.if_instr[2] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold2858 (.A(\soc_inst.cpu_core.id_rs2_data[5] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\soc_inst.cpu_core.ex_alu_result[5] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold2860 (.A(\soc_inst.cpu_core.id_rs1_data[20] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold2861 (.A(\soc_inst.pwm_inst.channel_counter[0][8] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold2862 (.A(_08924_),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\soc_inst.cpu_core.alu.b[27] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold2864 (.A(\soc_inst.cpu_core.alu.b[7] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold2865 (.A(_04417_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold2866 (.A(\soc_inst.cpu_core.if_funct3[2] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold2867 (.A(_00889_),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold2868 (.A(\soc_inst.cpu_core.if_pc[23] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold2869 (.A(_00930_),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\soc_inst.mem_ctrl.next_instr_addr[0] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold2871 (.A(_00549_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\soc_inst.cpu_core.alu.b[20] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold2873 (.A(_01177_),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold2874 (.A(\soc_inst.cpu_core.id_rs1_data[13] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold2875 (.A(\soc_inst.mem_ctrl.spi_addr[10] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold2876 (.A(_00559_),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold2877 (.A(\soc_inst.cpu_core.id_rs2_data[18] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold2878 (.A(\soc_inst.mem_ctrl.spi_data_out[16] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold2879 (.A(\soc_inst.core_mem_addr[6] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold2880 (.A(\soc_inst.cpu_core.csr_file.mepc[4] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold2881 (.A(_00525_),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold2882 (.A(\soc_inst.cpu_core.id_imm[30] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold2883 (.A(_04319_),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold2884 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[9] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold2885 (.A(\soc_inst.cpu_core.ex_alu_result[23] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold2886 (.A(\soc_inst.i2c_inst.bit_cnt[1] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold2887 (.A(_09457_),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\soc_inst.mem_ctrl.spi_addr[4] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold2889 (.A(\soc_inst.mem_ctrl.spi_addr[8] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold2890 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[6] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold2891 (.A(_02497_),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\soc_inst.cpu_core.id_rs1_data[27] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold2893 (.A(\soc_inst.cpu_core.alu.b[6] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold2894 (.A(_04415_),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold2895 (.A(_01163_),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\soc_inst.cpu_core.alu.b[30] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold2897 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[7] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\soc_inst.cpu_core.id_rs1_data[0] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold2899 (.A(\soc_inst.cpu_core.ex_funct3[0] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold2900 (.A(_01206_),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\soc_inst.cpu_core.csr_file.mtime[23] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold2902 (.A(\soc_inst.mem_ctrl.spi_data_out[20] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold2903 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[4] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold2904 (.A(_07752_),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold2905 (.A(\soc_inst.i2c_inst.data_reg[6] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\soc_inst.i2c_inst.data_reg[0] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold2907 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[1] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold2908 (.A(\soc_inst.cpu_core.id_rs1_data[9] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold2909 (.A(uio_out[1]),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold2910 (.A(_00815_),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold2911 (.A(\soc_inst.cpu_core.id_rs2_data[7] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold2912 (.A(uio_out[2]),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold2913 (.A(_00816_),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold2914 (.A(\soc_inst.cpu_core.ex_alu_result[28] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold2915 (.A(\soc_inst.pwm_inst.channel_counter[0][13] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold2916 (.A(_08934_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold2917 (.A(\soc_inst.spi_inst.clock_divider[5] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold2918 (.A(_00318_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold2919 (.A(\soc_inst.cpu_core.alu.b[10] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold2920 (.A(_04423_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold2921 (.A(\soc_inst.cpu_core.id_rs1_data[10] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold2922 (.A(\soc_inst.cpu_core.ex_alu_result[20] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold2923 (.A(\soc_inst.mem_ctrl.spi_data_out[2] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold2924 (.A(\soc_inst.cpu_core.alu.b[21] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold2925 (.A(\soc_inst.mem_ctrl.spi_addr[21] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold2926 (.A(\soc_inst.mem_ctrl.spi_data_out[6] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold2927 (.A(\soc_inst.mem_ctrl.spi_data_out[17] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold2928 (.A(\soc_inst.cpu_core.id_rs1_data[23] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold2929 (.A(\soc_inst.cpu_core.id_pc[18] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold2930 (.A(_00251_),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold2931 (.A(\soc_inst.core_instr_addr[10] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold2932 (.A(_00531_),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold2933 (.A(\soc_inst.cpu_core.ex_branch_target[1] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold2934 (.A(\soc_inst.pwm_inst.channel_counter[0][6] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold2935 (.A(\soc_inst.cpu_core.if_funct3[0] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold2936 (.A(_00887_),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold2937 (.A(\soc_inst.cpu_core.id_instr[2] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold2938 (.A(\soc_inst.cpu_core.ex_instr[2] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold2939 (.A(\soc_inst.cpu_core.if_imm12[3] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold2940 (.A(\soc_inst.cpu_core.alu.a[4] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold2941 (.A(\soc_inst.cpu_core.id_rs1_data[12] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold2942 (.A(\soc_inst.cpu_core.csr_file.mepc[0] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold2943 (.A(\soc_inst.pwm_inst.channel_counter[0][12] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold2944 (.A(\soc_inst.cpu_core.mem_instr[6] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold2945 (.A(_01034_),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold2946 (.A(\soc_inst.pwm_inst.channel_counter[0][1] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold2947 (.A(\soc_inst.cpu_core.csr_file.mtval[4] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold2948 (.A(_09182_),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold2949 (.A(\soc_inst.cpu_core.ex_funct3[1] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold2950 (.A(_01207_),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold2951 (.A(\soc_inst.core_mem_flag[0] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold2952 (.A(\soc_inst.mem_ctrl.spi_addr[2] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold2953 (.A(_00551_),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold2954 (.A(\soc_inst.cpu_core.ex_alu_result[18] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold2955 (.A(\soc_inst.cpu_core.ex_branch_target[17] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold2956 (.A(_02359_),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold2957 (.A(\soc_inst.cpu_core.ex_branch_target[6] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold2958 (.A(_02348_),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold2959 (.A(\soc_inst.core_mem_addr[5] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold2960 (.A(\soc_inst.cpu_core.id_rs2_data[6] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold2961 (.A(\soc_inst.cpu_core.alu.b[12] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold2962 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[3] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold2963 (.A(_07750_),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold2964 (.A(_02590_),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold2965 (.A(\soc_inst.core_instr_addr[9] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold2966 (.A(_00530_),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold2967 (.A(\soc_inst.mem_ctrl.spi_data_out[9] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold2968 (.A(\soc_inst.cpu_core.id_imm[0] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold2969 (.A(\soc_inst.cpu_core.id_imm[28] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold2970 (.A(\soc_inst.uart_instances[0].uart_inst.uart_receiver.cycle_counter[2] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold2971 (.A(_00257_),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold2972 (.A(\soc_inst.cpu_core.id_instr[3] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold2973 (.A(_01197_),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold2974 (.A(\soc_inst.cpu_core.id_pc[19] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold2975 (.A(\soc_inst.mem_ctrl.spi_addr[19] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold2976 (.A(_00568_),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold2977 (.A(\soc_inst.cpu_core.id_pc[9] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold2978 (.A(\soc_inst.mem_ctrl.spi_data_out[12] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold2979 (.A(\soc_inst.cpu_core.csr_file.mret_trigger ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold2980 (.A(\soc_inst.cpu_core.id_rs1_data[17] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold2981 (.A(\soc_inst.cpu_core.id_imm[22] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold2982 (.A(\soc_inst.cpu_core.alu.b[28] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold2983 (.A(\soc_inst.cpu_core.id_imm[25] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold2984 (.A(\soc_inst.cpu_core.alu.b[5] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold2985 (.A(\soc_inst.cpu_core.ex_alu_result[22] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold2986 (.A(\soc_inst.cpu_core.if_instr[3] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold2987 (.A(uio_out[4]),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold2988 (.A(\soc_inst.cpu_core.csr_file.mtval[31] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold2989 (.A(_02402_),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold2990 (.A(\soc_inst.mem_ctrl.spi_data_out[11] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold2991 (.A(\soc_inst.cpu_core.csr_file.mcause[31] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold2992 (.A(_02441_),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold2993 (.A(\soc_inst.cpu_core.id_rs1_data[14] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold2994 (.A(\soc_inst.cpu_core.ex_branch_target[5] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold2995 (.A(_02347_),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold2996 (.A(\soc_inst.cpu_core.id_pc[11] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold2997 (.A(\soc_inst.core_instr_addr[2] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold2998 (.A(\soc_inst.cpu_core.alu.a[29] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold2999 (.A(\soc_inst.mem_ctrl.spi_addr[22] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold3000 (.A(_00571_),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold3001 (.A(\soc_inst.cpu_core.id_imm[9] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold3002 (.A(\soc_inst.cpu_core.id_rs1_data[5] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold3003 (.A(\soc_inst.mem_ctrl.spi_addr[13] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold3004 (.A(_00562_),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold3005 (.A(\soc_inst.mem_ctrl.spi_data_out[8] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold3006 (.A(\soc_inst.cpu_core.alu.op[2] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold3007 (.A(\soc_inst.cpu_core.id_imm[5] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold3008 (.A(\soc_inst.mem_ctrl.spi_data_out[14] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold3009 (.A(\soc_inst.cpu_core.alu.a[5] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold3010 (.A(\soc_inst.cpu_core.id_rs1_data[11] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold3011 (.A(\soc_inst.core_mem_wdata[1] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold3012 (.A(\soc_inst.cpu_core.csr_file.mtval[0] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold3013 (.A(\soc_inst.core_instr_addr[17] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold3014 (.A(\soc_inst.cpu_core.ex_branch_target[27] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold3015 (.A(_02369_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold3016 (.A(\soc_inst.cpu_core.ex_alu_result[29] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold3017 (.A(\soc_inst.mem_ctrl.spi_addr[20] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold3018 (.A(_00569_),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold3019 (.A(\soc_inst.cpu_core.id_imm[1] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold3020 (.A(\soc_inst.cpu_core.id_imm[2] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold3021 (.A(\soc_inst.cpu_core.id_rs2_data[22] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold3022 (.A(\soc_inst.cpu_core.csr_file.mtval[3] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold3023 (.A(_00086_),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold3024 (.A(\soc_inst.cpu_core.id_imm[19] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold3025 (.A(\soc_inst.core_mem_addr[7] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold3026 (.A(\soc_inst.core_mem_addr[16] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold3027 (.A(\soc_inst.cpu_core.id_pc[10] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold3028 (.A(\soc_inst.cpu_core.csr_file.mtval[25] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold3029 (.A(\soc_inst.cpu_core.csr_file.mtval[30] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold3030 (.A(_07407_),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold3031 (.A(\soc_inst.cpu_core.ex_alu_result[4] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold3032 (.A(_01350_),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold3033 (.A(\soc_inst.cpu_core.id_rs2_data[21] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold3034 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.fsm_state[1] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold3035 (.A(\soc_inst.mem_ctrl.spi_data_out[7] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold3036 (.A(\soc_inst.cpu_core.id_rs2_data[24] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold3037 (.A(\soc_inst.cpu_core.csr_file.mcause[3] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold3038 (.A(\soc_inst.cpu_core.csr_file.mtval[22] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold3039 (.A(\soc_inst.cpu_core.csr_file.mtval[28] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold3040 (.A(\soc_inst.cpu_core.id_funct3[1] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold3041 (.A(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold3042 (.A(\soc_inst.i2c_inst.bit_cnt[0] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold3043 (.A(_00401_),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold3044 (.A(\soc_inst.cpu_core.id_rs1_data[28] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold3045 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[1] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold3046 (.A(\soc_inst.mem_ctrl.spi_addr[6] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold3047 (.A(\soc_inst.cpu_core.id_imm[18] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold3048 (.A(\soc_inst.mem_ctrl.spi_data_out[3] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold3049 (.A(\soc_inst.cpu_core.csr_file.mcause[1] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold3050 (.A(\soc_inst.core_instr_addr[20] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold3051 (.A(\soc_inst.mem_ctrl.spi_data_out[15] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold3052 (.A(\soc_inst.mem_ctrl.spi_data_out[1] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold3053 (.A(\soc_inst.cpu_core.id_rs2_data[27] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold3054 (.A(\soc_inst.core_instr_addr[19] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold3055 (.A(\soc_inst.cpu_core.id_rs2_data[26] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold3056 (.A(\soc_inst.cpu_core.id_rs1_data[16] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold3057 (.A(\soc_inst.cpu_core.alu.a[0] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold3058 (.A(\soc_inst.cpu_core.id_pc[17] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold3059 (.A(\soc_inst.core_instr_addr[16] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold3060 (.A(_00537_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold3061 (.A(\soc_inst.mem_ctrl.spi_addr[11] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold3062 (.A(_00560_),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold3063 (.A(\soc_inst.mem_ctrl.spi_data_out[5] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold3064 (.A(\soc_inst.pwm_inst.channel_counter[0][9] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold3065 (.A(\soc_inst.cpu_core.id_imm[29] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold3066 (.A(\soc_inst.cpu_core.alu.a[7] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold3067 (.A(\soc_inst.cpu_core.id_pc[14] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold3068 (.A(\soc_inst.mem_ctrl.spi_data_out[4] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold3069 (.A(\soc_inst.mem_ctrl.instr_ready_reg ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold3070 (.A(\soc_inst.cpu_core.csr_file.mepc[1] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold3071 (.A(\soc_inst.mem_ctrl.next_instr_ready_reg ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold3072 (.A(_00639_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold3073 (.A(\soc_inst.cpu_core.ex_alu_result[17] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold3074 (.A(\soc_inst.cpu_core.csr_file.mtval[29] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold3075 (.A(_07400_),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold3076 (.A(\soc_inst.cpu_core.id_funct3[0] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold3077 (.A(\soc_inst.cpu_core.alu.b[18] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold3078 (.A(_01175_),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold3079 (.A(\soc_inst.spi_inst.cpha ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold3080 (.A(\soc_inst.cpu_core.if_funct7[3] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold3081 (.A(\soc_inst.cpu_core.ex_alu_result[9] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold3082 (.A(_01355_),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold3083 (.A(\soc_inst.cpu_core.alu.b[29] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold3084 (.A(\soc_inst.cpu_core.id_rs1_data[29] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold3085 (.A(\soc_inst.cpu_core.csr_file.mtime[8] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold3086 (.A(_00219_),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold3087 (.A(\soc_inst.mem_ctrl.spi_addr[7] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold3088 (.A(\soc_inst.cpu_core.csr_file.mtval[23] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold3089 (.A(_07358_),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold3090 (.A(\soc_inst.cpu_core.id_imm[24] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold3091 (.A(\soc_inst.cpu_core.id_rs1_data[8] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold3092 (.A(\soc_inst.cpu_core.alu.b[26] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold3093 (.A(\soc_inst.cpu_core.csr_file.mtval[1] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold3094 (.A(\soc_inst.core_instr_addr[23] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold3095 (.A(\soc_inst.cpu_core.if_instr[5] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold3096 (.A(\soc_inst.spi_ena ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold3097 (.A(\soc_inst.cpu_core.id_pc[22] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold3098 (.A(\soc_inst.mem_ctrl.spi_addr[16] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold3099 (.A(\soc_inst.cpu_core.alu.b[9] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold3100 (.A(_04421_),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold3101 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[1] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold3102 (.A(\soc_inst.mem_ctrl.spi_addr[18] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold3103 (.A(\soc_inst.cpu_core.id_instr[5] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold3104 (.A(\soc_inst.cpu_core.id_imm[14] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold3105 (.A(\soc_inst.cpu_core.id_pc[15] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold3106 (.A(\soc_inst.spi_inst.cpol ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold3107 (.A(\soc_inst.i2c_inst.bit_cnt[3] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold3108 (.A(_09464_),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold3109 (.A(\soc_inst.pwm_inst.channel_counter[0][14] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold3110 (.A(\soc_inst.cpu_core.id_rs1_data[1] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold3111 (.A(\soc_inst.mem_ctrl.spi_mem_inst.write_enable ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold3112 (.A(_08656_),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold3113 (.A(_00015_),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold3114 (.A(\soc_inst.cpu_core.csr_file.mtval[24] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold3115 (.A(_07364_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold3116 (.A(\soc_inst.cpu_core.csr_file.mcause[0] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold3117 (.A(\soc_inst.cpu_core.ex_instr[7] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold3118 (.A(_01189_),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold3119 (.A(\soc_inst.cpu_core.csr_file.mtval[26] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold3120 (.A(_07379_),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold3121 (.A(\soc_inst.cpu_core.id_imm[12] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold3122 (.A(\soc_inst.cpu_core.id_imm[20] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold3123 (.A(\soc_inst.cpu_core.id_imm[23] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold3124 (.A(\soc_inst.cpu_core.alu.b[15] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold3125 (.A(\soc_inst.cpu_core.ex_alu_result[27] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold3126 (.A(\soc_inst.cpu_core.ex_alu_result[1] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold3127 (.A(_01347_),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold3128 (.A(\soc_inst.core_mem_addr[1] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold3129 (.A(\soc_inst.cpu_core.ex_alu_result[10] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold3130 (.A(\soc_inst.cpu_core.if_funct7[1] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold3131 (.A(\soc_inst.cpu_core.ex_alu_result[11] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold3132 (.A(_01357_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold3133 (.A(\soc_inst.cpu_core.ex_alu_result[15] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold3134 (.A(\soc_inst.cpu_core.csr_file.mcause[2] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold3135 (.A(\soc_inst.cpu_core.id_rs1_data[15] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold3136 (.A(\soc_inst.cpu_core.ex_alu_result[8] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold3137 (.A(_01354_),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold3138 (.A(\soc_inst.i2c_inst.state[0] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold3139 (.A(_00545_),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold3140 (.A(\soc_inst.cpu_core.id_rs1_data[19] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold3141 (.A(_00315_),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold3142 (.A(\soc_inst.cpu_core.id_pc[12] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold3143 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[0] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold3144 (.A(\soc_inst.cpu_core.csr_file.mtval[21] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold3145 (.A(\soc_inst.cpu_core.csr_file.mtval[16] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold3146 (.A(\soc_inst.cpu_core.csr_file.mepc[11] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold3147 (.A(_00532_),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold3148 (.A(\soc_inst.cpu_core.csr_file.mtval[27] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold3149 (.A(_07386_),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold3150 (.A(\soc_inst.cpu_core.csr_file.mtime[33] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold3151 (.A(_00200_),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold3152 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[4] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold3153 (.A(\soc_inst.cpu_core.csr_file.mtval[14] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold3154 (.A(_07284_),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold3155 (.A(\soc_inst.cpu_core.id_imm[17] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold3156 (.A(\soc_inst.cpu_core.ex_alu_result[24] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold3157 (.A(\soc_inst.cpu_core.if_instr[6] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold3158 (.A(\soc_inst.cpu_core.id_rs2_data[23] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold3159 (.A(\soc_inst.cpu_core.csr_file.mtval[15] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold3160 (.A(_07291_),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold3161 (.A(\soc_inst.i2c_inst.state[3] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold3162 (.A(\soc_inst.cpu_core.id_imm[15] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold3163 (.A(\soc_inst.cpu_core.alu.b[31] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold3164 (.A(_04467_),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold3165 (.A(\soc_inst.cpu_core.ex_alu_result[19] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold3166 (.A(\soc_inst.cpu_core.csr_file.mepc[3] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold3167 (.A(\soc_inst.cpu_core.csr_file.mepc[2] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold3168 (.A(\soc_inst.core_instr_addr[12] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold3169 (.A(\soc_inst.cpu_core._unused_mem_rd_addr[1] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold3170 (.A(\soc_inst.cpu_core.id_imm[26] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold3171 (.A(\soc_inst.cpu_core.id_rs1_data[26] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold3172 (.A(_01022_),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold3173 (.A(\soc_inst.cpu_core.csr_file.mtval[13] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold3174 (.A(_07277_),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold3175 (.A(\soc_inst.cpu_core.alu.b[14] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold3176 (.A(\soc_inst.cpu_core.csr_file.mtime[4] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold3177 (.A(_00215_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold3178 (.A(\soc_inst.cpu_core.id_imm[27] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold3179 (.A(_04310_),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold3180 (.A(\soc_inst.cpu_core.alu.a[31] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold3181 (.A(\soc_inst.cpu_core.csr_file.mtval[2] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold3182 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[4] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold3183 (.A(_11363_),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold3184 (.A(\soc_inst.core_mem_addr[14] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold3185 (.A(_01296_),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold3186 (.A(\soc_inst.mem_ctrl.spi_addr[17] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold3187 (.A(\soc_inst.cpu_core.ex_alu_result[2] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold3188 (.A(_01284_),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold3189 (.A(\soc_inst.cpu_core.csr_file.mtval[17] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold3190 (.A(_07307_),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold3191 (.A(\soc_inst.cpu_core.csr_file.mstatus[3] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold3192 (.A(\soc_inst.cpu_core.alu.a[2] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold3193 (.A(\soc_inst.cpu_core.alu.b[8] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold3194 (.A(\soc_inst.cpu_core.ex_alu_result[25] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold3195 (.A(\soc_inst.cpu_core.id_imm[11] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold3196 (.A(_04263_),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold3197 (.A(\soc_inst.cpu_core.id_rs1_data[21] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold3198 (.A(\soc_inst.cpu_core.id_imm[21] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold3199 (.A(\soc_inst.cpu_core.csr_file.mtval[20] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold3200 (.A(\soc_inst.cpu_core.ex_alu_result[3] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold3201 (.A(_01349_),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold3202 (.A(\soc_inst.mem_ctrl.spi_done ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold3203 (.A(_00007_),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold3204 (.A(\soc_inst.cpu_core.id_rs1_data[2] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold3205 (.A(\soc_inst.mem_ctrl.spi_data_out[0] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold3206 (.A(\soc_inst.cpu_core.alu.b[13] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold3207 (.A(_04427_),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold3208 (.A(\soc_inst.cpu_core.ex_alu_result[13] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold3209 (.A(_01295_),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold3210 (.A(\soc_inst.cpu_core.ex_alu_result[14] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold3211 (.A(\soc_inst.cpu_core.alu.a[12] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold3212 (.A(_05207_),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold3213 (.A(_01359_),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold3214 (.A(\soc_inst.cpu_core.id_imm[16] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold3215 (.A(\soc_inst.cpu_core.alu.a[30] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold3216 (.A(_00317_),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold3217 (.A(\soc_inst.cpu_core.mem_reg_we ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold3218 (.A(\soc_inst.core_mem_addr[0] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold3219 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[1] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold3220 (.A(\soc_inst.core_instr_addr[14] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold3221 (.A(\soc_inst.cpu_core.csr_file.mtval[19] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold3222 (.A(_07326_),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold3223 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.data_to_send[7] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold3224 (.A(_07638_),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold3225 (.A(_00316_),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold3226 (.A(\soc_inst.cpu_core.id_pc[16] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold3227 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[8] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold3228 (.A(\soc_inst.core_instr_data[8] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold3229 (.A(\soc_inst.uart_instances[0].uart_inst.uart_transmitter.cycle_counter[0] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold3230 (.A(\soc_inst.cpu_core.alu.a[10] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold3231 (.A(\soc_inst.mem_ctrl.spi_addr[5] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold3232 (.A(\soc_inst.core_instr_addr[13] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold3233 (.A(\soc_inst.cpu_core.alu.op[1] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold3234 (.A(\soc_inst.mem_ctrl.spi_mem_inst.init_cnt[9] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold3235 (.A(\soc_inst.cpu_core.id_pc[20] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold3236 (.A(\soc_inst.core_instr_addr[22] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold3237 (.A(\soc_inst.cpu_core.alu.b[17] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold3238 (.A(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold3239 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold3240 (.A(\soc_inst.cpu_core.alu.a[21] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold3241 (.A(\soc_inst.cpu_core.alu.b[19] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold3242 (.A(\soc_inst.mem_ctrl.spi_addr[9] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold3243 (.A(\soc_inst.cpu_core.alu.op[0] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold3244 (.A(\soc_inst.core_instr_data[11] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold3245 (.A(\soc_inst.cpu_core.alu.b[3] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold3246 (.A(\soc_inst.cpu_core.if_funct7[6] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold3247 (.A(\soc_inst.cpu_core.alu.a[26] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold3248 (.A(\soc_inst.mem_ctrl.spi_is_instr ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold3249 (.A(\soc_inst.cpu_core.alu.a[27] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold3250 (.A(\soc_inst.cpu_core.ex_alu_result[30] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold3251 (.A(\soc_inst.cpu_core.alu.a[28] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold3252 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[4] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold3253 (.A(\soc_inst.cpu_core.alu.a[9] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold3254 (.A(\soc_inst.cpu_core.csr_file.mtime[15] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold3255 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[5] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold3256 (.A(\soc_inst.cpu_core.csr_file.mtime[5] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold3257 (.A(\soc_inst.cpu_core.alu.a[24] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold3258 (.A(\soc_inst.uart_instances[0].uart_inst.uart_divider_reg[7] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold3259 (.A(\soc_inst.cpu_core.ex_alu_result[26] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold3260 (.A(\soc_inst.gpio_inst.int_pend_reg[4] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold3261 (.A(_08297_),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold3262 (.A(\soc_inst.core_instr_data[5] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold3263 (.A(\soc_inst.cpu_core.alu.a[11] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold3264 (.A(\soc_inst.core_instr_data[4] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold3265 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[12] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold3266 (.A(_11332_),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold3267 (.A(_02375_),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold3268 (.A(\soc_inst.core_instr_data[15] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold3269 (.A(\soc_inst.core_mem_wdata[2] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold3270 (.A(\soc_inst.core_instr_data[0] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold3271 (.A(\soc_inst.cpu_core.alu.a[25] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold3272 (.A(\soc_inst.cpu_core.alu.b[16] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold3273 (.A(\soc_inst.i2c_inst.state[2] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold3274 (.A(\soc_inst.cpu_core.alu.op[3] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold3275 (.A(\soc_inst.cpu_core.alu.a[15] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold3276 (.A(\soc_inst.spi_inst.len_sel[1] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold3277 (.A(\soc_inst.spi_inst.bit_counter[2] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold3278 (.A(_09246_),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold3279 (.A(\soc_inst.core_instr_data[9] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold3280 (.A(\soc_inst.cpu_core.id_rs2_data[20] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold3281 (.A(\soc_inst.cpu_core.id_rs2_data[30] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold3282 (.A(\soc_inst.cpu_core.alu.a[13] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold3283 (.A(\soc_inst.cpu_core.id_rs2_data[25] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold3284 (.A(\soc_inst.cpu_core.alu.a[8] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold3285 (.A(\soc_inst.core_instr_data[7] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold3286 (.A(\soc_inst.core_instr_data[10] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold3287 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[2] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold3288 (.A(_08634_),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold3289 (.A(_00010_),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold3290 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[0] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold3291 (.A(_02374_),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold3292 (.A(\soc_inst.cpu_core.csr_file.mtime[30] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold3293 (.A(\soc_inst.mem_ctrl.access_state[3] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold3294 (.A(\soc_inst.core_instr_data[6] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold3295 (.A(\soc_inst.cpu_core.alu.a[16] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold3296 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[3] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold3297 (.A(_00832_),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold3298 (.A(\soc_inst.cpu_core.csr_file.mtime[40] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold3299 (.A(\soc_inst.cpu_core.alu.a[17] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold3300 (.A(\soc_inst.cpu_core.csr_file.mtime[2] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold3301 (.A(\soc_inst.cpu_core.csr_file.mtime[17] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold3302 (.A(\soc_inst.core_instr_data[14] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold3303 (.A(uio_oe[5]),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold3304 (.A(_11247_),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold3305 (.A(\soc_inst.i2c_inst.state[1] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold3306 (.A(\soc_inst.cpu_core.alu.a[22] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold3307 (.A(\soc_inst.cpu_core.alu.a[20] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold3308 (.A(\soc_inst.cpu_core.alu.a[23] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold3309 (.A(\soc_inst.core_mem_addr[13] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold3310 (.A(\soc_inst.cpu_core.alu.a[14] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold3311 (.A(\soc_inst.cpu_core.alu.b[2] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold3312 (.A(_01159_),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold3313 (.A(\soc_inst.mem_ctrl.spi_mem_inst.bit_counter[2] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold3314 (.A(\soc_inst.cpu_core.alu.a[18] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold3315 (.A(\soc_inst.core_instr_data[13] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold3316 (.A(\soc_inst.cpu_core.alu.a[19] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold3317 (.A(\soc_inst.cpu_core.if_imm12[0] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold3318 (.A(\soc_inst.cpu_core.alu.b[4] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold3319 (.A(\soc_inst.cpu_core.csr_file.mtime[39] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold3320 (.A(\soc_inst.mem_ctrl.spi_mem_inst.fsm_state[14] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold3321 (.A(\soc_inst.cpu_core.alu.op[3] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold3322 (.A(\soc_inst.cpu_core.ex_alu_result[1] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold3323 (.A(_00266_),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold3324 (.A(\soc_inst.cpu_core.id_rs1_data[22] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold3325 (.A(_07094_),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold3326 (.A(\soc_inst.core_instr_addr[22] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold3327 (.A(\soc_inst.cpu_core.csr_file.mtime[9] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold3328 (.A(\soc_inst.i2c_inst.clk_cnt[1] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold3329 (.A(\soc_inst.cpu_core.if_funct7[3] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold3330 (.A(\soc_inst.cpu_core.ex_exception_pc[11] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold3331 (.A(\soc_inst.cpu_core.id_pc[22] ),
    .X(net3410));
 sg13g2_antennanp ANTENNA_1 (.A(_09707_));
 sg13g2_antennanp ANTENNA_2 (.A(net6433));
 sg13g2_antennanp ANTENNA_3 (.A(net6433));
 sg13g2_antennanp ANTENNA_4 (.A(net6433));
 sg13g2_antennanp ANTENNA_5 (.A(net6433));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_46 ();
 sg13g2_fill_1 FILLER_0_61 ();
 sg13g2_fill_1 FILLER_0_66 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_fill_1 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_fill_2 FILLER_0_164 ();
 sg13g2_fill_1 FILLER_0_166 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_4 FILLER_0_221 ();
 sg13g2_fill_2 FILLER_0_225 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_fill_2 FILLER_0_277 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_fill_1 FILLER_0_289 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_314 ();
 sg13g2_fill_1 FILLER_0_316 ();
 sg13g2_fill_2 FILLER_0_347 ();
 sg13g2_fill_1 FILLER_0_349 ();
 sg13g2_fill_2 FILLER_0_379 ();
 sg13g2_fill_1 FILLER_0_381 ();
 sg13g2_fill_2 FILLER_0_391 ();
 sg13g2_fill_1 FILLER_0_425 ();
 sg13g2_fill_2 FILLER_0_471 ();
 sg13g2_fill_1 FILLER_0_473 ();
 sg13g2_fill_2 FILLER_0_479 ();
 sg13g2_fill_1 FILLER_0_481 ();
 sg13g2_fill_2 FILLER_0_496 ();
 sg13g2_fill_2 FILLER_0_517 ();
 sg13g2_fill_1 FILLER_0_519 ();
 sg13g2_fill_1 FILLER_0_642 ();
 sg13g2_fill_1 FILLER_0_708 ();
 sg13g2_fill_2 FILLER_0_728 ();
 sg13g2_fill_1 FILLER_0_730 ();
 sg13g2_fill_1 FILLER_0_773 ();
 sg13g2_fill_1 FILLER_0_805 ();
 sg13g2_fill_1 FILLER_0_946 ();
 sg13g2_fill_2 FILLER_0_975 ();
 sg13g2_fill_1 FILLER_0_977 ();
 sg13g2_fill_2 FILLER_0_996 ();
 sg13g2_fill_2 FILLER_0_1024 ();
 sg13g2_fill_1 FILLER_0_1080 ();
 sg13g2_fill_2 FILLER_0_1107 ();
 sg13g2_decap_8 FILLER_0_1143 ();
 sg13g2_decap_8 FILLER_0_1150 ();
 sg13g2_fill_1 FILLER_0_1157 ();
 sg13g2_fill_1 FILLER_0_1185 ();
 sg13g2_fill_2 FILLER_0_1227 ();
 sg13g2_fill_1 FILLER_0_1247 ();
 sg13g2_fill_2 FILLER_0_1258 ();
 sg13g2_decap_4 FILLER_0_1341 ();
 sg13g2_fill_2 FILLER_0_1345 ();
 sg13g2_fill_2 FILLER_0_1372 ();
 sg13g2_fill_1 FILLER_0_1374 ();
 sg13g2_decap_4 FILLER_0_1394 ();
 sg13g2_fill_1 FILLER_0_1398 ();
 sg13g2_decap_8 FILLER_0_1439 ();
 sg13g2_decap_8 FILLER_0_1446 ();
 sg13g2_decap_8 FILLER_0_1453 ();
 sg13g2_decap_4 FILLER_0_1469 ();
 sg13g2_fill_2 FILLER_0_1473 ();
 sg13g2_decap_4 FILLER_0_1480 ();
 sg13g2_decap_4 FILLER_0_1494 ();
 sg13g2_decap_4 FILLER_0_1504 ();
 sg13g2_decap_8 FILLER_0_1513 ();
 sg13g2_decap_8 FILLER_0_1520 ();
 sg13g2_decap_8 FILLER_0_1527 ();
 sg13g2_decap_8 FILLER_0_1534 ();
 sg13g2_decap_4 FILLER_0_1541 ();
 sg13g2_fill_1 FILLER_0_1545 ();
 sg13g2_fill_2 FILLER_0_1565 ();
 sg13g2_fill_2 FILLER_0_1608 ();
 sg13g2_fill_2 FILLER_0_1678 ();
 sg13g2_fill_1 FILLER_0_1680 ();
 sg13g2_decap_4 FILLER_0_1709 ();
 sg13g2_fill_2 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_8 FILLER_0_1762 ();
 sg13g2_decap_8 FILLER_0_1769 ();
 sg13g2_fill_1 FILLER_0_1798 ();
 sg13g2_decap_8 FILLER_0_1803 ();
 sg13g2_decap_8 FILLER_0_1810 ();
 sg13g2_fill_2 FILLER_0_1817 ();
 sg13g2_decap_8 FILLER_0_1888 ();
 sg13g2_fill_1 FILLER_0_1895 ();
 sg13g2_fill_2 FILLER_0_1900 ();
 sg13g2_fill_1 FILLER_0_1902 ();
 sg13g2_fill_1 FILLER_0_1908 ();
 sg13g2_fill_2 FILLER_0_1913 ();
 sg13g2_decap_4 FILLER_0_1919 ();
 sg13g2_fill_1 FILLER_0_1951 ();
 sg13g2_decap_8 FILLER_0_1974 ();
 sg13g2_fill_2 FILLER_0_1981 ();
 sg13g2_fill_1 FILLER_0_1992 ();
 sg13g2_fill_2 FILLER_0_2006 ();
 sg13g2_fill_1 FILLER_0_2008 ();
 sg13g2_fill_2 FILLER_0_2040 ();
 sg13g2_fill_1 FILLER_0_2042 ();
 sg13g2_fill_2 FILLER_0_2052 ();
 sg13g2_fill_1 FILLER_0_2054 ();
 sg13g2_decap_8 FILLER_0_2068 ();
 sg13g2_decap_8 FILLER_0_2075 ();
 sg13g2_fill_2 FILLER_0_2082 ();
 sg13g2_fill_2 FILLER_0_2088 ();
 sg13g2_decap_8 FILLER_0_2122 ();
 sg13g2_decap_8 FILLER_0_2129 ();
 sg13g2_decap_4 FILLER_0_2136 ();
 sg13g2_decap_8 FILLER_0_2153 ();
 sg13g2_fill_2 FILLER_0_2160 ();
 sg13g2_decap_4 FILLER_0_2167 ();
 sg13g2_decap_8 FILLER_0_2175 ();
 sg13g2_decap_8 FILLER_0_2182 ();
 sg13g2_decap_8 FILLER_0_2189 ();
 sg13g2_fill_2 FILLER_0_2205 ();
 sg13g2_decap_8 FILLER_0_2216 ();
 sg13g2_decap_4 FILLER_0_2223 ();
 sg13g2_fill_1 FILLER_0_2231 ();
 sg13g2_fill_2 FILLER_0_2315 ();
 sg13g2_decap_8 FILLER_0_2322 ();
 sg13g2_fill_1 FILLER_0_2329 ();
 sg13g2_fill_1 FILLER_0_2334 ();
 sg13g2_decap_4 FILLER_0_2340 ();
 sg13g2_fill_2 FILLER_0_2344 ();
 sg13g2_decap_8 FILLER_0_2355 ();
 sg13g2_decap_8 FILLER_0_2362 ();
 sg13g2_fill_1 FILLER_0_2369 ();
 sg13g2_decap_4 FILLER_0_2397 ();
 sg13g2_fill_1 FILLER_0_2446 ();
 sg13g2_decap_8 FILLER_0_2468 ();
 sg13g2_decap_8 FILLER_0_2475 ();
 sg13g2_fill_1 FILLER_0_2482 ();
 sg13g2_decap_8 FILLER_0_2523 ();
 sg13g2_decap_4 FILLER_0_2530 ();
 sg13g2_fill_2 FILLER_0_2539 ();
 sg13g2_fill_1 FILLER_0_2607 ();
 sg13g2_fill_2 FILLER_0_2616 ();
 sg13g2_fill_1 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2640 ();
 sg13g2_decap_8 FILLER_0_2647 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_decap_4 FILLER_0_2668 ();
 sg13g2_fill_2 FILLER_0_2672 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_54 ();
 sg13g2_fill_1 FILLER_1_56 ();
 sg13g2_fill_1 FILLER_1_122 ();
 sg13g2_fill_2 FILLER_1_183 ();
 sg13g2_fill_1 FILLER_1_185 ();
 sg13g2_fill_2 FILLER_1_230 ();
 sg13g2_fill_1 FILLER_1_232 ();
 sg13g2_fill_1 FILLER_1_369 ();
 sg13g2_fill_1 FILLER_1_469 ();
 sg13g2_fill_2 FILLER_1_507 ();
 sg13g2_fill_2 FILLER_1_524 ();
 sg13g2_fill_2 FILLER_1_645 ();
 sg13g2_fill_1 FILLER_1_702 ();
 sg13g2_fill_1 FILLER_1_793 ();
 sg13g2_fill_2 FILLER_1_832 ();
 sg13g2_fill_1 FILLER_1_834 ();
 sg13g2_fill_1 FILLER_1_872 ();
 sg13g2_fill_2 FILLER_1_1286 ();
 sg13g2_fill_1 FILLER_1_1385 ();
 sg13g2_fill_2 FILLER_1_1444 ();
 sg13g2_fill_2 FILLER_1_1495 ();
 sg13g2_decap_8 FILLER_1_1532 ();
 sg13g2_decap_4 FILLER_1_1539 ();
 sg13g2_fill_2 FILLER_1_1543 ();
 sg13g2_fill_2 FILLER_1_1564 ();
 sg13g2_fill_2 FILLER_1_1643 ();
 sg13g2_fill_1 FILLER_1_1645 ();
 sg13g2_fill_1 FILLER_1_1660 ();
 sg13g2_decap_8 FILLER_1_1722 ();
 sg13g2_fill_2 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1758 ();
 sg13g2_fill_1 FILLER_1_1765 ();
 sg13g2_fill_1 FILLER_1_1850 ();
 sg13g2_fill_2 FILLER_1_1869 ();
 sg13g2_fill_1 FILLER_1_1871 ();
 sg13g2_decap_4 FILLER_1_1973 ();
 sg13g2_fill_2 FILLER_1_1977 ();
 sg13g2_fill_1 FILLER_1_2037 ();
 sg13g2_decap_8 FILLER_1_2066 ();
 sg13g2_fill_2 FILLER_1_2073 ();
 sg13g2_fill_2 FILLER_1_2138 ();
 sg13g2_fill_1 FILLER_1_2168 ();
 sg13g2_fill_1 FILLER_1_2178 ();
 sg13g2_fill_2 FILLER_1_2235 ();
 sg13g2_fill_2 FILLER_1_2250 ();
 sg13g2_fill_1 FILLER_1_2280 ();
 sg13g2_fill_2 FILLER_1_2330 ();
 sg13g2_fill_2 FILLER_1_2359 ();
 sg13g2_fill_2 FILLER_1_2365 ();
 sg13g2_fill_1 FILLER_1_2367 ();
 sg13g2_fill_2 FILLER_1_2373 ();
 sg13g2_fill_1 FILLER_1_2448 ();
 sg13g2_fill_2 FILLER_1_2477 ();
 sg13g2_fill_2 FILLER_1_2588 ();
 sg13g2_fill_1 FILLER_1_2590 ();
 sg13g2_fill_2 FILLER_1_2624 ();
 sg13g2_decap_8 FILLER_1_2654 ();
 sg13g2_decap_8 FILLER_1_2661 ();
 sg13g2_decap_4 FILLER_1_2668 ();
 sg13g2_fill_2 FILLER_1_2672 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_fill_2 FILLER_2_169 ();
 sg13g2_fill_1 FILLER_2_171 ();
 sg13g2_fill_1 FILLER_2_226 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_304 ();
 sg13g2_fill_2 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_348 ();
 sg13g2_fill_1 FILLER_2_417 ();
 sg13g2_fill_2 FILLER_2_529 ();
 sg13g2_fill_1 FILLER_2_569 ();
 sg13g2_fill_1 FILLER_2_603 ();
 sg13g2_fill_1 FILLER_2_646 ();
 sg13g2_fill_2 FILLER_2_680 ();
 sg13g2_fill_2 FILLER_2_720 ();
 sg13g2_fill_1 FILLER_2_722 ();
 sg13g2_fill_1 FILLER_2_756 ();
 sg13g2_fill_2 FILLER_2_878 ();
 sg13g2_fill_1 FILLER_2_880 ();
 sg13g2_fill_2 FILLER_2_935 ();
 sg13g2_fill_1 FILLER_2_937 ();
 sg13g2_fill_2 FILLER_2_1051 ();
 sg13g2_fill_1 FILLER_2_1118 ();
 sg13g2_fill_1 FILLER_2_1141 ();
 sg13g2_fill_2 FILLER_2_1202 ();
 sg13g2_fill_1 FILLER_2_1204 ();
 sg13g2_fill_2 FILLER_2_1294 ();
 sg13g2_fill_1 FILLER_2_1315 ();
 sg13g2_fill_2 FILLER_2_1467 ();
 sg13g2_fill_2 FILLER_2_1582 ();
 sg13g2_fill_1 FILLER_2_1584 ();
 sg13g2_fill_2 FILLER_2_1603 ();
 sg13g2_fill_2 FILLER_2_1680 ();
 sg13g2_fill_1 FILLER_2_1682 ();
 sg13g2_fill_2 FILLER_2_1798 ();
 sg13g2_fill_1 FILLER_2_1800 ();
 sg13g2_fill_1 FILLER_2_1829 ();
 sg13g2_fill_1 FILLER_2_1839 ();
 sg13g2_fill_2 FILLER_2_1896 ();
 sg13g2_fill_1 FILLER_2_1898 ();
 sg13g2_decap_4 FILLER_2_2064 ();
 sg13g2_fill_2 FILLER_2_2068 ();
 sg13g2_fill_2 FILLER_2_2203 ();
 sg13g2_fill_2 FILLER_2_2233 ();
 sg13g2_fill_1 FILLER_2_2268 ();
 sg13g2_fill_2 FILLER_2_2291 ();
 sg13g2_fill_1 FILLER_2_2302 ();
 sg13g2_fill_2 FILLER_2_2424 ();
 sg13g2_fill_1 FILLER_2_2435 ();
 sg13g2_fill_1 FILLER_2_2500 ();
 sg13g2_fill_2 FILLER_2_2519 ();
 sg13g2_fill_1 FILLER_2_2521 ();
 sg13g2_decap_8 FILLER_2_2654 ();
 sg13g2_decap_8 FILLER_2_2661 ();
 sg13g2_decap_4 FILLER_2_2668 ();
 sg13g2_fill_2 FILLER_2_2672 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_11 ();
 sg13g2_fill_2 FILLER_3_56 ();
 sg13g2_fill_1 FILLER_3_173 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_300 ();
 sg13g2_fill_1 FILLER_3_302 ();
 sg13g2_fill_2 FILLER_3_339 ();
 sg13g2_fill_1 FILLER_3_392 ();
 sg13g2_fill_2 FILLER_3_429 ();
 sg13g2_fill_1 FILLER_3_455 ();
 sg13g2_fill_2 FILLER_3_474 ();
 sg13g2_fill_2 FILLER_3_600 ();
 sg13g2_fill_2 FILLER_3_666 ();
 sg13g2_fill_1 FILLER_3_668 ();
 sg13g2_fill_1 FILLER_3_761 ();
 sg13g2_fill_2 FILLER_3_798 ();
 sg13g2_fill_1 FILLER_3_800 ();
 sg13g2_fill_2 FILLER_3_828 ();
 sg13g2_fill_1 FILLER_3_830 ();
 sg13g2_fill_2 FILLER_3_867 ();
 sg13g2_fill_1 FILLER_3_869 ();
 sg13g2_fill_1 FILLER_3_984 ();
 sg13g2_fill_2 FILLER_3_1091 ();
 sg13g2_fill_1 FILLER_3_1111 ();
 sg13g2_fill_2 FILLER_3_1130 ();
 sg13g2_fill_2 FILLER_3_1222 ();
 sg13g2_fill_1 FILLER_3_1233 ();
 sg13g2_fill_1 FILLER_3_1244 ();
 sg13g2_fill_2 FILLER_3_1283 ();
 sg13g2_fill_1 FILLER_3_1304 ();
 sg13g2_fill_2 FILLER_3_1353 ();
 sg13g2_fill_1 FILLER_3_1405 ();
 sg13g2_fill_1 FILLER_3_1420 ();
 sg13g2_fill_2 FILLER_3_1459 ();
 sg13g2_fill_1 FILLER_3_1477 ();
 sg13g2_fill_2 FILLER_3_1484 ();
 sg13g2_fill_1 FILLER_3_1519 ();
 sg13g2_decap_4 FILLER_3_1593 ();
 sg13g2_fill_2 FILLER_3_1597 ();
 sg13g2_fill_2 FILLER_3_1645 ();
 sg13g2_fill_2 FILLER_3_1674 ();
 sg13g2_fill_1 FILLER_3_1676 ();
 sg13g2_fill_2 FILLER_3_1684 ();
 sg13g2_fill_2 FILLER_3_1714 ();
 sg13g2_fill_1 FILLER_3_1716 ();
 sg13g2_fill_2 FILLER_3_1757 ();
 sg13g2_fill_1 FILLER_3_1759 ();
 sg13g2_fill_2 FILLER_3_1801 ();
 sg13g2_fill_1 FILLER_3_1803 ();
 sg13g2_fill_1 FILLER_3_1845 ();
 sg13g2_fill_1 FILLER_3_1855 ();
 sg13g2_fill_2 FILLER_3_1874 ();
 sg13g2_fill_1 FILLER_3_1876 ();
 sg13g2_fill_1 FILLER_3_1923 ();
 sg13g2_fill_2 FILLER_3_2022 ();
 sg13g2_fill_1 FILLER_3_2069 ();
 sg13g2_decap_4 FILLER_3_2120 ();
 sg13g2_fill_1 FILLER_3_2137 ();
 sg13g2_fill_1 FILLER_3_2143 ();
 sg13g2_fill_1 FILLER_3_2181 ();
 sg13g2_fill_1 FILLER_3_2303 ();
 sg13g2_fill_1 FILLER_3_2359 ();
 sg13g2_fill_2 FILLER_3_2400 ();
 sg13g2_fill_1 FILLER_3_2434 ();
 sg13g2_fill_2 FILLER_3_2467 ();
 sg13g2_fill_1 FILLER_3_2469 ();
 sg13g2_fill_2 FILLER_3_2501 ();
 sg13g2_fill_2 FILLER_3_2530 ();
 sg13g2_fill_1 FILLER_3_2588 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_59 ();
 sg13g2_fill_2 FILLER_4_115 ();
 sg13g2_fill_2 FILLER_4_141 ();
 sg13g2_fill_1 FILLER_4_143 ();
 sg13g2_fill_2 FILLER_4_201 ();
 sg13g2_fill_1 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_300 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_fill_2 FILLER_4_386 ();
 sg13g2_fill_1 FILLER_4_410 ();
 sg13g2_fill_1 FILLER_4_475 ();
 sg13g2_fill_1 FILLER_4_513 ();
 sg13g2_fill_2 FILLER_4_523 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_fill_1 FILLER_4_591 ();
 sg13g2_fill_1 FILLER_4_634 ();
 sg13g2_fill_2 FILLER_4_658 ();
 sg13g2_fill_2 FILLER_4_670 ();
 sg13g2_fill_2 FILLER_4_699 ();
 sg13g2_fill_1 FILLER_4_701 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_fill_1 FILLER_4_755 ();
 sg13g2_fill_2 FILLER_4_799 ();
 sg13g2_fill_2 FILLER_4_810 ();
 sg13g2_fill_2 FILLER_4_878 ();
 sg13g2_fill_1 FILLER_4_880 ();
 sg13g2_fill_1 FILLER_4_899 ();
 sg13g2_fill_1 FILLER_4_971 ();
 sg13g2_fill_2 FILLER_4_1079 ();
 sg13g2_fill_1 FILLER_4_1151 ();
 sg13g2_fill_1 FILLER_4_1317 ();
 sg13g2_fill_1 FILLER_4_1352 ();
 sg13g2_fill_1 FILLER_4_1362 ();
 sg13g2_fill_2 FILLER_4_1396 ();
 sg13g2_fill_2 FILLER_4_1435 ();
 sg13g2_fill_2 FILLER_4_1464 ();
 sg13g2_fill_2 FILLER_4_1484 ();
 sg13g2_fill_2 FILLER_4_1500 ();
 sg13g2_fill_1 FILLER_4_1512 ();
 sg13g2_decap_4 FILLER_4_1545 ();
 sg13g2_fill_2 FILLER_4_1562 ();
 sg13g2_fill_2 FILLER_4_1586 ();
 sg13g2_fill_2 FILLER_4_1602 ();
 sg13g2_fill_1 FILLER_4_1604 ();
 sg13g2_decap_8 FILLER_4_1642 ();
 sg13g2_fill_2 FILLER_4_1724 ();
 sg13g2_fill_1 FILLER_4_1726 ();
 sg13g2_fill_2 FILLER_4_1740 ();
 sg13g2_fill_1 FILLER_4_1742 ();
 sg13g2_fill_2 FILLER_4_1785 ();
 sg13g2_fill_1 FILLER_4_1787 ();
 sg13g2_fill_1 FILLER_4_1816 ();
 sg13g2_fill_2 FILLER_4_1911 ();
 sg13g2_fill_2 FILLER_4_1935 ();
 sg13g2_fill_1 FILLER_4_1959 ();
 sg13g2_fill_1 FILLER_4_1973 ();
 sg13g2_fill_2 FILLER_4_2023 ();
 sg13g2_fill_1 FILLER_4_2025 ();
 sg13g2_fill_1 FILLER_4_2129 ();
 sg13g2_fill_1 FILLER_4_2138 ();
 sg13g2_decap_8 FILLER_4_2180 ();
 sg13g2_fill_1 FILLER_4_2187 ();
 sg13g2_fill_2 FILLER_4_2197 ();
 sg13g2_fill_1 FILLER_4_2199 ();
 sg13g2_fill_2 FILLER_4_2213 ();
 sg13g2_fill_1 FILLER_4_2251 ();
 sg13g2_fill_1 FILLER_4_2288 ();
 sg13g2_fill_2 FILLER_4_2325 ();
 sg13g2_fill_1 FILLER_4_2327 ();
 sg13g2_fill_2 FILLER_4_2337 ();
 sg13g2_fill_2 FILLER_4_2352 ();
 sg13g2_fill_1 FILLER_4_2354 ();
 sg13g2_fill_1 FILLER_4_2399 ();
 sg13g2_fill_1 FILLER_4_2441 ();
 sg13g2_fill_2 FILLER_4_2470 ();
 sg13g2_fill_1 FILLER_4_2472 ();
 sg13g2_fill_2 FILLER_4_2495 ();
 sg13g2_fill_1 FILLER_4_2524 ();
 sg13g2_fill_2 FILLER_4_2557 ();
 sg13g2_fill_2 FILLER_4_2604 ();
 sg13g2_fill_1 FILLER_4_2606 ();
 sg13g2_fill_2 FILLER_4_2630 ();
 sg13g2_fill_1 FILLER_4_2632 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_decap_4 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_fill_2 FILLER_5_393 ();
 sg13g2_fill_1 FILLER_5_395 ();
 sg13g2_fill_1 FILLER_5_479 ();
 sg13g2_fill_2 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_500 ();
 sg13g2_fill_2 FILLER_5_556 ();
 sg13g2_fill_1 FILLER_5_558 ();
 sg13g2_fill_1 FILLER_5_605 ();
 sg13g2_fill_2 FILLER_5_628 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_fill_2 FILLER_5_654 ();
 sg13g2_fill_2 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_693 ();
 sg13g2_fill_1 FILLER_5_704 ();
 sg13g2_fill_2 FILLER_5_723 ();
 sg13g2_fill_1 FILLER_5_725 ();
 sg13g2_fill_2 FILLER_5_740 ();
 sg13g2_fill_2 FILLER_5_789 ();
 sg13g2_fill_1 FILLER_5_791 ();
 sg13g2_fill_1 FILLER_5_818 ();
 sg13g2_fill_2 FILLER_5_840 ();
 sg13g2_fill_1 FILLER_5_863 ();
 sg13g2_fill_1 FILLER_5_914 ();
 sg13g2_fill_2 FILLER_5_924 ();
 sg13g2_fill_2 FILLER_5_948 ();
 sg13g2_fill_1 FILLER_5_950 ();
 sg13g2_fill_2 FILLER_5_1024 ();
 sg13g2_fill_1 FILLER_5_1115 ();
 sg13g2_fill_2 FILLER_5_1189 ();
 sg13g2_fill_1 FILLER_5_1242 ();
 sg13g2_fill_1 FILLER_5_1310 ();
 sg13g2_fill_1 FILLER_5_1320 ();
 sg13g2_fill_1 FILLER_5_1346 ();
 sg13g2_fill_2 FILLER_5_1406 ();
 sg13g2_fill_1 FILLER_5_1408 ();
 sg13g2_fill_2 FILLER_5_1448 ();
 sg13g2_fill_1 FILLER_5_1455 ();
 sg13g2_decap_8 FILLER_5_1492 ();
 sg13g2_decap_4 FILLER_5_1499 ();
 sg13g2_decap_8 FILLER_5_1507 ();
 sg13g2_decap_8 FILLER_5_1542 ();
 sg13g2_fill_2 FILLER_5_1549 ();
 sg13g2_fill_1 FILLER_5_1551 ();
 sg13g2_fill_1 FILLER_5_1574 ();
 sg13g2_decap_4 FILLER_5_1588 ();
 sg13g2_fill_1 FILLER_5_1592 ();
 sg13g2_decap_8 FILLER_5_1630 ();
 sg13g2_decap_8 FILLER_5_1637 ();
 sg13g2_decap_4 FILLER_5_1644 ();
 sg13g2_decap_4 FILLER_5_1676 ();
 sg13g2_fill_1 FILLER_5_1693 ();
 sg13g2_fill_2 FILLER_5_1744 ();
 sg13g2_fill_1 FILLER_5_1786 ();
 sg13g2_fill_2 FILLER_5_1810 ();
 sg13g2_fill_1 FILLER_5_1812 ();
 sg13g2_fill_1 FILLER_5_1822 ();
 sg13g2_fill_2 FILLER_5_1851 ();
 sg13g2_fill_1 FILLER_5_1853 ();
 sg13g2_fill_2 FILLER_5_1884 ();
 sg13g2_fill_2 FILLER_5_1939 ();
 sg13g2_fill_1 FILLER_5_1941 ();
 sg13g2_fill_1 FILLER_5_2029 ();
 sg13g2_fill_2 FILLER_5_2084 ();
 sg13g2_fill_1 FILLER_5_2086 ();
 sg13g2_decap_8 FILLER_5_2132 ();
 sg13g2_decap_8 FILLER_5_2180 ();
 sg13g2_fill_1 FILLER_5_2187 ();
 sg13g2_fill_2 FILLER_5_2248 ();
 sg13g2_fill_1 FILLER_5_2250 ();
 sg13g2_fill_1 FILLER_5_2278 ();
 sg13g2_fill_1 FILLER_5_2339 ();
 sg13g2_fill_2 FILLER_5_2362 ();
 sg13g2_fill_1 FILLER_5_2364 ();
 sg13g2_fill_2 FILLER_5_2391 ();
 sg13g2_fill_2 FILLER_5_2429 ();
 sg13g2_fill_1 FILLER_5_2431 ();
 sg13g2_fill_1 FILLER_5_2441 ();
 sg13g2_fill_2 FILLER_5_2474 ();
 sg13g2_fill_1 FILLER_5_2476 ();
 sg13g2_fill_2 FILLER_5_2486 ();
 sg13g2_fill_2 FILLER_5_2506 ();
 sg13g2_fill_1 FILLER_5_2508 ();
 sg13g2_fill_1 FILLER_5_2518 ();
 sg13g2_fill_1 FILLER_5_2584 ();
 sg13g2_fill_1 FILLER_5_2594 ();
 sg13g2_fill_1 FILLER_5_2673 ();
 sg13g2_fill_2 FILLER_6_75 ();
 sg13g2_fill_1 FILLER_6_113 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_4 FILLER_6_166 ();
 sg13g2_fill_2 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_decap_8 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_fill_2 FILLER_6_204 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_1 FILLER_6_234 ();
 sg13g2_fill_2 FILLER_6_323 ();
 sg13g2_fill_2 FILLER_6_353 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_425 ();
 sg13g2_fill_2 FILLER_6_461 ();
 sg13g2_fill_1 FILLER_6_463 ();
 sg13g2_fill_2 FILLER_6_483 ();
 sg13g2_fill_2 FILLER_6_608 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_fill_1 FILLER_6_638 ();
 sg13g2_fill_1 FILLER_6_739 ();
 sg13g2_fill_2 FILLER_6_815 ();
 sg13g2_fill_1 FILLER_6_932 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1038 ();
 sg13g2_fill_2 FILLER_6_1062 ();
 sg13g2_fill_1 FILLER_6_1142 ();
 sg13g2_fill_2 FILLER_6_1266 ();
 sg13g2_fill_2 FILLER_6_1321 ();
 sg13g2_fill_2 FILLER_6_1336 ();
 sg13g2_fill_2 FILLER_6_1381 ();
 sg13g2_fill_1 FILLER_6_1383 ();
 sg13g2_fill_2 FILLER_6_1482 ();
 sg13g2_decap_8 FILLER_6_1487 ();
 sg13g2_fill_1 FILLER_6_1494 ();
 sg13g2_decap_8 FILLER_6_1504 ();
 sg13g2_fill_1 FILLER_6_1541 ();
 sg13g2_decap_8 FILLER_6_1551 ();
 sg13g2_fill_1 FILLER_6_1558 ();
 sg13g2_decap_4 FILLER_6_1623 ();
 sg13g2_fill_2 FILLER_6_1627 ();
 sg13g2_decap_8 FILLER_6_1695 ();
 sg13g2_decap_8 FILLER_6_1702 ();
 sg13g2_fill_1 FILLER_6_1709 ();
 sg13g2_decap_8 FILLER_6_1717 ();
 sg13g2_fill_1 FILLER_6_1724 ();
 sg13g2_fill_2 FILLER_6_1821 ();
 sg13g2_fill_2 FILLER_6_1867 ();
 sg13g2_fill_1 FILLER_6_1869 ();
 sg13g2_fill_2 FILLER_6_1902 ();
 sg13g2_fill_1 FILLER_6_1904 ();
 sg13g2_fill_2 FILLER_6_1972 ();
 sg13g2_fill_1 FILLER_6_1974 ();
 sg13g2_fill_2 FILLER_6_1985 ();
 sg13g2_fill_1 FILLER_6_1987 ();
 sg13g2_fill_2 FILLER_6_2042 ();
 sg13g2_fill_2 FILLER_6_2049 ();
 sg13g2_fill_1 FILLER_6_2051 ();
 sg13g2_fill_2 FILLER_6_2078 ();
 sg13g2_fill_2 FILLER_6_2089 ();
 sg13g2_fill_1 FILLER_6_2091 ();
 sg13g2_fill_1 FILLER_6_2127 ();
 sg13g2_fill_1 FILLER_6_2132 ();
 sg13g2_fill_1 FILLER_6_2143 ();
 sg13g2_decap_8 FILLER_6_2181 ();
 sg13g2_fill_1 FILLER_6_2188 ();
 sg13g2_fill_2 FILLER_6_2217 ();
 sg13g2_fill_1 FILLER_6_2219 ();
 sg13g2_fill_2 FILLER_6_2224 ();
 sg13g2_fill_1 FILLER_6_2226 ();
 sg13g2_fill_2 FILLER_6_2236 ();
 sg13g2_fill_1 FILLER_6_2259 ();
 sg13g2_fill_2 FILLER_6_2274 ();
 sg13g2_fill_1 FILLER_6_2276 ();
 sg13g2_fill_2 FILLER_6_2317 ();
 sg13g2_fill_2 FILLER_6_2332 ();
 sg13g2_fill_1 FILLER_6_2334 ();
 sg13g2_fill_1 FILLER_6_2453 ();
 sg13g2_decap_8 FILLER_6_2502 ();
 sg13g2_decap_4 FILLER_6_2509 ();
 sg13g2_fill_2 FILLER_6_2635 ();
 sg13g2_fill_1 FILLER_6_2637 ();
 sg13g2_fill_1 FILLER_7_126 ();
 sg13g2_decap_4 FILLER_7_130 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_decap_4 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_2 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_decap_4 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_276 ();
 sg13g2_fill_2 FILLER_7_325 ();
 sg13g2_fill_1 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_459 ();
 sg13g2_fill_2 FILLER_7_601 ();
 sg13g2_fill_1 FILLER_7_623 ();
 sg13g2_fill_2 FILLER_7_680 ();
 sg13g2_fill_2 FILLER_7_729 ();
 sg13g2_fill_1 FILLER_7_731 ();
 sg13g2_fill_1 FILLER_7_799 ();
 sg13g2_fill_1 FILLER_7_806 ();
 sg13g2_fill_2 FILLER_7_961 ();
 sg13g2_fill_1 FILLER_7_963 ();
 sg13g2_fill_2 FILLER_7_1018 ();
 sg13g2_fill_1 FILLER_7_1020 ();
 sg13g2_fill_1 FILLER_7_1107 ();
 sg13g2_fill_1 FILLER_7_1117 ();
 sg13g2_fill_1 FILLER_7_1217 ();
 sg13g2_fill_1 FILLER_7_1263 ();
 sg13g2_fill_1 FILLER_7_1370 ();
 sg13g2_fill_1 FILLER_7_1411 ();
 sg13g2_fill_2 FILLER_7_1429 ();
 sg13g2_fill_1 FILLER_7_1431 ();
 sg13g2_fill_2 FILLER_7_1436 ();
 sg13g2_fill_1 FILLER_7_1438 ();
 sg13g2_fill_2 FILLER_7_1466 ();
 sg13g2_fill_1 FILLER_7_1468 ();
 sg13g2_fill_2 FILLER_7_1496 ();
 sg13g2_fill_1 FILLER_7_1498 ();
 sg13g2_fill_2 FILLER_7_1598 ();
 sg13g2_decap_4 FILLER_7_1609 ();
 sg13g2_fill_1 FILLER_7_1613 ();
 sg13g2_fill_2 FILLER_7_1634 ();
 sg13g2_fill_2 FILLER_7_1777 ();
 sg13g2_fill_1 FILLER_7_1779 ();
 sg13g2_fill_2 FILLER_7_1817 ();
 sg13g2_fill_1 FILLER_7_1819 ();
 sg13g2_fill_2 FILLER_7_1838 ();
 sg13g2_fill_2 FILLER_7_1894 ();
 sg13g2_fill_2 FILLER_7_1940 ();
 sg13g2_fill_2 FILLER_7_1978 ();
 sg13g2_fill_2 FILLER_7_2021 ();
 sg13g2_fill_2 FILLER_7_2050 ();
 sg13g2_fill_1 FILLER_7_2052 ();
 sg13g2_fill_1 FILLER_7_2079 ();
 sg13g2_fill_2 FILLER_7_2139 ();
 sg13g2_fill_2 FILLER_7_2181 ();
 sg13g2_fill_1 FILLER_7_2260 ();
 sg13g2_fill_2 FILLER_7_2275 ();
 sg13g2_fill_2 FILLER_7_2304 ();
 sg13g2_fill_1 FILLER_7_2306 ();
 sg13g2_fill_2 FILLER_7_2334 ();
 sg13g2_fill_2 FILLER_7_2363 ();
 sg13g2_fill_2 FILLER_7_2414 ();
 sg13g2_fill_1 FILLER_7_2416 ();
 sg13g2_fill_2 FILLER_7_2458 ();
 sg13g2_fill_1 FILLER_7_2460 ();
 sg13g2_fill_1 FILLER_7_2497 ();
 sg13g2_fill_2 FILLER_7_2543 ();
 sg13g2_fill_2 FILLER_7_2559 ();
 sg13g2_fill_2 FILLER_7_2570 ();
 sg13g2_fill_2 FILLER_7_2581 ();
 sg13g2_fill_1 FILLER_7_2583 ();
 sg13g2_fill_1 FILLER_7_2673 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_decap_8 FILLER_8_134 ();
 sg13g2_decap_4 FILLER_8_141 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_fill_2 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_240 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_fill_1 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_fill_2 FILLER_8_369 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_fill_2 FILLER_8_395 ();
 sg13g2_fill_2 FILLER_8_402 ();
 sg13g2_fill_1 FILLER_8_404 ();
 sg13g2_fill_2 FILLER_8_547 ();
 sg13g2_fill_1 FILLER_8_567 ();
 sg13g2_fill_1 FILLER_8_622 ();
 sg13g2_fill_2 FILLER_8_728 ();
 sg13g2_fill_2 FILLER_8_771 ();
 sg13g2_fill_2 FILLER_8_846 ();
 sg13g2_fill_1 FILLER_8_865 ();
 sg13g2_fill_1 FILLER_8_973 ();
 sg13g2_fill_2 FILLER_8_1001 ();
 sg13g2_fill_1 FILLER_8_1017 ();
 sg13g2_fill_2 FILLER_8_1035 ();
 sg13g2_fill_1 FILLER_8_1068 ();
 sg13g2_fill_1 FILLER_8_1136 ();
 sg13g2_fill_1 FILLER_8_1283 ();
 sg13g2_fill_2 FILLER_8_1339 ();
 sg13g2_fill_1 FILLER_8_1341 ();
 sg13g2_fill_1 FILLER_8_1364 ();
 sg13g2_fill_1 FILLER_8_1408 ();
 sg13g2_decap_8 FILLER_8_1431 ();
 sg13g2_decap_8 FILLER_8_1438 ();
 sg13g2_fill_2 FILLER_8_1450 ();
 sg13g2_fill_1 FILLER_8_1461 ();
 sg13g2_fill_2 FILLER_8_1495 ();
 sg13g2_fill_1 FILLER_8_1574 ();
 sg13g2_fill_2 FILLER_8_1583 ();
 sg13g2_fill_1 FILLER_8_1585 ();
 sg13g2_fill_1 FILLER_8_1706 ();
 sg13g2_fill_2 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1749 ();
 sg13g2_decap_8 FILLER_8_1756 ();
 sg13g2_fill_1 FILLER_8_1843 ();
 sg13g2_fill_1 FILLER_8_1910 ();
 sg13g2_fill_2 FILLER_8_1929 ();
 sg13g2_fill_1 FILLER_8_1975 ();
 sg13g2_fill_1 FILLER_8_2024 ();
 sg13g2_fill_1 FILLER_8_2039 ();
 sg13g2_fill_2 FILLER_8_2094 ();
 sg13g2_fill_2 FILLER_8_2130 ();
 sg13g2_fill_1 FILLER_8_2164 ();
 sg13g2_fill_2 FILLER_8_2222 ();
 sg13g2_fill_1 FILLER_8_2224 ();
 sg13g2_fill_1 FILLER_8_2293 ();
 sg13g2_fill_2 FILLER_8_2321 ();
 sg13g2_fill_1 FILLER_8_2323 ();
 sg13g2_fill_1 FILLER_8_2373 ();
 sg13g2_fill_2 FILLER_8_2384 ();
 sg13g2_fill_1 FILLER_8_2386 ();
 sg13g2_fill_1 FILLER_8_2450 ();
 sg13g2_fill_1 FILLER_8_2487 ();
 sg13g2_fill_1 FILLER_8_2515 ();
 sg13g2_fill_2 FILLER_8_2596 ();
 sg13g2_fill_2 FILLER_8_2620 ();
 sg13g2_fill_1 FILLER_8_2622 ();
 sg13g2_fill_2 FILLER_8_2628 ();
 sg13g2_fill_1 FILLER_8_2635 ();
 sg13g2_fill_1 FILLER_8_2662 ();
 sg13g2_fill_2 FILLER_8_2672 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_1 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_fill_2 FILLER_9_126 ();
 sg13g2_fill_1 FILLER_9_128 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_fill_1 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_9_504 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_fill_2 FILLER_9_539 ();
 sg13g2_fill_2 FILLER_9_569 ();
 sg13g2_fill_2 FILLER_9_602 ();
 sg13g2_fill_1 FILLER_9_604 ();
 sg13g2_fill_2 FILLER_9_618 ();
 sg13g2_fill_2 FILLER_9_637 ();
 sg13g2_fill_1 FILLER_9_639 ();
 sg13g2_fill_1 FILLER_9_731 ();
 sg13g2_fill_1 FILLER_9_762 ();
 sg13g2_fill_1 FILLER_9_802 ();
 sg13g2_fill_2 FILLER_9_816 ();
 sg13g2_fill_1 FILLER_9_818 ();
 sg13g2_fill_2 FILLER_9_973 ();
 sg13g2_fill_1 FILLER_9_975 ();
 sg13g2_fill_2 FILLER_9_989 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_9_1070 ();
 sg13g2_fill_1 FILLER_9_1081 ();
 sg13g2_fill_2 FILLER_9_1117 ();
 sg13g2_fill_1 FILLER_9_1170 ();
 sg13g2_fill_1 FILLER_9_1248 ();
 sg13g2_fill_1 FILLER_9_1273 ();
 sg13g2_fill_1 FILLER_9_1329 ();
 sg13g2_fill_2 FILLER_9_1343 ();
 sg13g2_decap_4 FILLER_9_1381 ();
 sg13g2_fill_2 FILLER_9_1385 ();
 sg13g2_fill_2 FILLER_9_1392 ();
 sg13g2_fill_1 FILLER_9_1394 ();
 sg13g2_decap_8 FILLER_9_1423 ();
 sg13g2_decap_8 FILLER_9_1430 ();
 sg13g2_decap_8 FILLER_9_1437 ();
 sg13g2_decap_8 FILLER_9_1444 ();
 sg13g2_fill_2 FILLER_9_1451 ();
 sg13g2_fill_2 FILLER_9_1544 ();
 sg13g2_fill_2 FILLER_9_1556 ();
 sg13g2_fill_2 FILLER_9_1574 ();
 sg13g2_fill_1 FILLER_9_1589 ();
 sg13g2_fill_1 FILLER_9_1603 ();
 sg13g2_decap_4 FILLER_9_1632 ();
 sg13g2_fill_2 FILLER_9_1654 ();
 sg13g2_fill_1 FILLER_9_1656 ();
 sg13g2_fill_1 FILLER_9_1663 ();
 sg13g2_fill_1 FILLER_9_1708 ();
 sg13g2_fill_2 FILLER_9_1737 ();
 sg13g2_fill_2 FILLER_9_1743 ();
 sg13g2_fill_1 FILLER_9_1745 ();
 sg13g2_decap_4 FILLER_9_1755 ();
 sg13g2_fill_1 FILLER_9_1759 ();
 sg13g2_fill_1 FILLER_9_1806 ();
 sg13g2_fill_1 FILLER_9_1919 ();
 sg13g2_fill_2 FILLER_9_1943 ();
 sg13g2_fill_1 FILLER_9_1945 ();
 sg13g2_decap_8 FILLER_9_1973 ();
 sg13g2_decap_8 FILLER_9_1980 ();
 sg13g2_decap_8 FILLER_9_1987 ();
 sg13g2_decap_8 FILLER_9_1998 ();
 sg13g2_fill_1 FILLER_9_2005 ();
 sg13g2_fill_2 FILLER_9_2010 ();
 sg13g2_decap_4 FILLER_9_2028 ();
 sg13g2_fill_1 FILLER_9_2032 ();
 sg13g2_fill_2 FILLER_9_2037 ();
 sg13g2_fill_1 FILLER_9_2039 ();
 sg13g2_decap_4 FILLER_9_2081 ();
 sg13g2_fill_2 FILLER_9_2098 ();
 sg13g2_fill_1 FILLER_9_2124 ();
 sg13g2_fill_2 FILLER_9_2218 ();
 sg13g2_fill_1 FILLER_9_2220 ();
 sg13g2_fill_1 FILLER_9_2239 ();
 sg13g2_fill_2 FILLER_9_2276 ();
 sg13g2_fill_2 FILLER_9_2287 ();
 sg13g2_fill_1 FILLER_9_2289 ();
 sg13g2_fill_2 FILLER_9_2305 ();
 sg13g2_fill_2 FILLER_9_2319 ();
 sg13g2_fill_1 FILLER_9_2321 ();
 sg13g2_fill_1 FILLER_9_2331 ();
 sg13g2_fill_2 FILLER_9_2461 ();
 sg13g2_fill_1 FILLER_9_2673 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_5 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_fill_2 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_358 ();
 sg13g2_fill_2 FILLER_10_375 ();
 sg13g2_fill_2 FILLER_10_405 ();
 sg13g2_fill_2 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_464 ();
 sg13g2_fill_2 FILLER_10_583 ();
 sg13g2_fill_1 FILLER_10_585 ();
 sg13g2_fill_1 FILLER_10_611 ();
 sg13g2_fill_2 FILLER_10_696 ();
 sg13g2_fill_1 FILLER_10_698 ();
 sg13g2_fill_1 FILLER_10_737 ();
 sg13g2_fill_1 FILLER_10_747 ();
 sg13g2_fill_1 FILLER_10_870 ();
 sg13g2_fill_2 FILLER_10_928 ();
 sg13g2_fill_2 FILLER_10_1039 ();
 sg13g2_fill_1 FILLER_10_1051 ();
 sg13g2_fill_1 FILLER_10_1097 ();
 sg13g2_fill_1 FILLER_10_1220 ();
 sg13g2_fill_1 FILLER_10_1274 ();
 sg13g2_fill_1 FILLER_10_1343 ();
 sg13g2_fill_2 FILLER_10_1385 ();
 sg13g2_fill_2 FILLER_10_1405 ();
 sg13g2_fill_1 FILLER_10_1416 ();
 sg13g2_fill_2 FILLER_10_1429 ();
 sg13g2_fill_1 FILLER_10_1431 ();
 sg13g2_decap_8 FILLER_10_1447 ();
 sg13g2_fill_2 FILLER_10_1454 ();
 sg13g2_fill_1 FILLER_10_1456 ();
 sg13g2_fill_2 FILLER_10_1466 ();
 sg13g2_fill_2 FILLER_10_1491 ();
 sg13g2_fill_1 FILLER_10_1498 ();
 sg13g2_fill_1 FILLER_10_1511 ();
 sg13g2_fill_2 FILLER_10_1520 ();
 sg13g2_fill_1 FILLER_10_1522 ();
 sg13g2_fill_1 FILLER_10_1528 ();
 sg13g2_fill_1 FILLER_10_1568 ();
 sg13g2_fill_2 FILLER_10_1689 ();
 sg13g2_fill_1 FILLER_10_1708 ();
 sg13g2_fill_2 FILLER_10_1765 ();
 sg13g2_fill_2 FILLER_10_1772 ();
 sg13g2_fill_1 FILLER_10_1796 ();
 sg13g2_fill_1 FILLER_10_1811 ();
 sg13g2_decap_4 FILLER_10_1847 ();
 sg13g2_fill_1 FILLER_10_1851 ();
 sg13g2_fill_2 FILLER_10_1857 ();
 sg13g2_fill_1 FILLER_10_1859 ();
 sg13g2_decap_4 FILLER_10_1869 ();
 sg13g2_fill_2 FILLER_10_1919 ();
 sg13g2_fill_1 FILLER_10_1921 ();
 sg13g2_fill_2 FILLER_10_1932 ();
 sg13g2_fill_1 FILLER_10_1934 ();
 sg13g2_fill_2 FILLER_10_1943 ();
 sg13g2_decap_8 FILLER_10_1982 ();
 sg13g2_decap_8 FILLER_10_1989 ();
 sg13g2_decap_8 FILLER_10_1996 ();
 sg13g2_fill_2 FILLER_10_2003 ();
 sg13g2_fill_1 FILLER_10_2005 ();
 sg13g2_fill_1 FILLER_10_2047 ();
 sg13g2_fill_2 FILLER_10_2059 ();
 sg13g2_fill_1 FILLER_10_2061 ();
 sg13g2_fill_1 FILLER_10_2093 ();
 sg13g2_fill_2 FILLER_10_2183 ();
 sg13g2_fill_2 FILLER_10_2212 ();
 sg13g2_fill_2 FILLER_10_2275 ();
 sg13g2_fill_1 FILLER_10_2286 ();
 sg13g2_fill_1 FILLER_10_2299 ();
 sg13g2_decap_8 FILLER_10_2332 ();
 sg13g2_fill_2 FILLER_10_2339 ();
 sg13g2_fill_2 FILLER_10_2346 ();
 sg13g2_decap_8 FILLER_10_2380 ();
 sg13g2_fill_1 FILLER_10_2387 ();
 sg13g2_fill_1 FILLER_10_2409 ();
 sg13g2_fill_2 FILLER_10_2431 ();
 sg13g2_fill_1 FILLER_10_2433 ();
 sg13g2_fill_2 FILLER_10_2523 ();
 sg13g2_fill_2 FILLER_10_2534 ();
 sg13g2_fill_1 FILLER_10_2536 ();
 sg13g2_fill_2 FILLER_10_2585 ();
 sg13g2_fill_1 FILLER_10_2596 ();
 sg13g2_fill_2 FILLER_10_2610 ();
 sg13g2_fill_1 FILLER_10_2645 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_fill_2 FILLER_11_124 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_fill_2 FILLER_11_194 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_2 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_208 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_2 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_411 ();
 sg13g2_fill_2 FILLER_11_517 ();
 sg13g2_fill_1 FILLER_11_533 ();
 sg13g2_fill_2 FILLER_11_548 ();
 sg13g2_fill_1 FILLER_11_550 ();
 sg13g2_fill_1 FILLER_11_597 ();
 sg13g2_fill_1 FILLER_11_645 ();
 sg13g2_fill_2 FILLER_11_755 ();
 sg13g2_fill_2 FILLER_11_793 ();
 sg13g2_fill_2 FILLER_11_808 ();
 sg13g2_fill_1 FILLER_11_837 ();
 sg13g2_fill_2 FILLER_11_966 ();
 sg13g2_fill_1 FILLER_11_968 ();
 sg13g2_fill_2 FILLER_11_982 ();
 sg13g2_fill_1 FILLER_11_984 ();
 sg13g2_fill_1 FILLER_11_994 ();
 sg13g2_fill_1 FILLER_11_1013 ();
 sg13g2_fill_2 FILLER_11_1122 ();
 sg13g2_fill_1 FILLER_11_1124 ();
 sg13g2_fill_1 FILLER_11_1135 ();
 sg13g2_fill_1 FILLER_11_1222 ();
 sg13g2_fill_2 FILLER_11_1293 ();
 sg13g2_fill_1 FILLER_11_1295 ();
 sg13g2_decap_4 FILLER_11_1329 ();
 sg13g2_fill_1 FILLER_11_1333 ();
 sg13g2_fill_1 FILLER_11_1382 ();
 sg13g2_fill_2 FILLER_11_1406 ();
 sg13g2_fill_2 FILLER_11_1428 ();
 sg13g2_fill_2 FILLER_11_1438 ();
 sg13g2_decap_4 FILLER_11_1457 ();
 sg13g2_fill_1 FILLER_11_1461 ();
 sg13g2_fill_2 FILLER_11_1472 ();
 sg13g2_fill_2 FILLER_11_1482 ();
 sg13g2_fill_2 FILLER_11_1499 ();
 sg13g2_fill_2 FILLER_11_1509 ();
 sg13g2_fill_1 FILLER_11_1511 ();
 sg13g2_fill_2 FILLER_11_1527 ();
 sg13g2_fill_1 FILLER_11_1553 ();
 sg13g2_fill_2 FILLER_11_1563 ();
 sg13g2_fill_1 FILLER_11_1585 ();
 sg13g2_fill_2 FILLER_11_1678 ();
 sg13g2_decap_4 FILLER_11_1717 ();
 sg13g2_fill_1 FILLER_11_1721 ();
 sg13g2_decap_4 FILLER_11_1732 ();
 sg13g2_fill_1 FILLER_11_1736 ();
 sg13g2_decap_4 FILLER_11_1746 ();
 sg13g2_fill_2 FILLER_11_1812 ();
 sg13g2_decap_4 FILLER_11_1851 ();
 sg13g2_fill_2 FILLER_11_1855 ();
 sg13g2_decap_8 FILLER_11_1861 ();
 sg13g2_fill_1 FILLER_11_1868 ();
 sg13g2_fill_2 FILLER_11_1925 ();
 sg13g2_fill_1 FILLER_11_1927 ();
 sg13g2_fill_1 FILLER_11_1981 ();
 sg13g2_decap_4 FILLER_11_1991 ();
 sg13g2_fill_2 FILLER_11_1995 ();
 sg13g2_decap_4 FILLER_11_2014 ();
 sg13g2_decap_4 FILLER_11_2062 ();
 sg13g2_fill_2 FILLER_11_2066 ();
 sg13g2_decap_4 FILLER_11_2097 ();
 sg13g2_fill_1 FILLER_11_2101 ();
 sg13g2_decap_4 FILLER_11_2110 ();
 sg13g2_fill_1 FILLER_11_2114 ();
 sg13g2_fill_1 FILLER_11_2186 ();
 sg13g2_fill_2 FILLER_11_2255 ();
 sg13g2_fill_2 FILLER_11_2336 ();
 sg13g2_decap_4 FILLER_11_2343 ();
 sg13g2_fill_1 FILLER_11_2347 ();
 sg13g2_decap_8 FILLER_11_2364 ();
 sg13g2_decap_8 FILLER_11_2380 ();
 sg13g2_decap_4 FILLER_11_2387 ();
 sg13g2_fill_2 FILLER_11_2397 ();
 sg13g2_fill_1 FILLER_11_2417 ();
 sg13g2_fill_2 FILLER_11_2445 ();
 sg13g2_fill_2 FILLER_11_2459 ();
 sg13g2_fill_1 FILLER_11_2461 ();
 sg13g2_fill_1 FILLER_11_2546 ();
 sg13g2_fill_2 FILLER_11_2575 ();
 sg13g2_fill_1 FILLER_11_2577 ();
 sg13g2_fill_1 FILLER_11_2601 ();
 sg13g2_fill_2 FILLER_11_2638 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_36 ();
 sg13g2_fill_1 FILLER_12_38 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_110 ();
 sg13g2_decap_4 FILLER_12_114 ();
 sg13g2_decap_4 FILLER_12_125 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_decap_8 FILLER_12_145 ();
 sg13g2_decap_4 FILLER_12_157 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_decap_4 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_178 ();
 sg13g2_decap_4 FILLER_12_200 ();
 sg13g2_decap_4 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_369 ();
 sg13g2_fill_1 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_514 ();
 sg13g2_fill_2 FILLER_12_703 ();
 sg13g2_fill_1 FILLER_12_705 ();
 sg13g2_fill_1 FILLER_12_749 ();
 sg13g2_fill_2 FILLER_12_807 ();
 sg13g2_fill_1 FILLER_12_809 ();
 sg13g2_fill_1 FILLER_12_883 ();
 sg13g2_fill_1 FILLER_12_927 ();
 sg13g2_fill_2 FILLER_12_965 ();
 sg13g2_fill_2 FILLER_12_1076 ();
 sg13g2_fill_1 FILLER_12_1245 ();
 sg13g2_fill_1 FILLER_12_1286 ();
 sg13g2_fill_2 FILLER_12_1335 ();
 sg13g2_fill_1 FILLER_12_1337 ();
 sg13g2_fill_1 FILLER_12_1395 ();
 sg13g2_fill_1 FILLER_12_1420 ();
 sg13g2_fill_2 FILLER_12_1468 ();
 sg13g2_fill_1 FILLER_12_1470 ();
 sg13g2_fill_1 FILLER_12_1484 ();
 sg13g2_fill_2 FILLER_12_1550 ();
 sg13g2_fill_1 FILLER_12_1570 ();
 sg13g2_decap_4 FILLER_12_1579 ();
 sg13g2_fill_2 FILLER_12_1583 ();
 sg13g2_fill_2 FILLER_12_1647 ();
 sg13g2_fill_1 FILLER_12_1694 ();
 sg13g2_decap_4 FILLER_12_1730 ();
 sg13g2_fill_1 FILLER_12_1756 ();
 sg13g2_fill_1 FILLER_12_1770 ();
 sg13g2_fill_2 FILLER_12_1803 ();
 sg13g2_fill_1 FILLER_12_1805 ();
 sg13g2_fill_2 FILLER_12_1833 ();
 sg13g2_fill_1 FILLER_12_1835 ();
 sg13g2_decap_8 FILLER_12_1862 ();
 sg13g2_fill_1 FILLER_12_1869 ();
 sg13g2_fill_1 FILLER_12_1947 ();
 sg13g2_fill_2 FILLER_12_1960 ();
 sg13g2_fill_2 FILLER_12_2022 ();
 sg13g2_fill_1 FILLER_12_2024 ();
 sg13g2_fill_2 FILLER_12_2074 ();
 sg13g2_fill_1 FILLER_12_2076 ();
 sg13g2_fill_1 FILLER_12_2105 ();
 sg13g2_fill_1 FILLER_12_2115 ();
 sg13g2_decap_8 FILLER_12_2186 ();
 sg13g2_fill_1 FILLER_12_2193 ();
 sg13g2_fill_1 FILLER_12_2274 ();
 sg13g2_fill_1 FILLER_12_2304 ();
 sg13g2_fill_2 FILLER_12_2337 ();
 sg13g2_decap_8 FILLER_12_2372 ();
 sg13g2_decap_4 FILLER_12_2379 ();
 sg13g2_fill_1 FILLER_12_2383 ();
 sg13g2_fill_2 FILLER_12_2537 ();
 sg13g2_fill_2 FILLER_12_2560 ();
 sg13g2_fill_2 FILLER_12_2620 ();
 sg13g2_fill_1 FILLER_12_2622 ();
 sg13g2_fill_1 FILLER_12_2632 ();
 sg13g2_fill_2 FILLER_12_2651 ();
 sg13g2_fill_2 FILLER_12_2671 ();
 sg13g2_fill_1 FILLER_12_2673 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_fill_2 FILLER_13_173 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_fill_2 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_423 ();
 sg13g2_fill_2 FILLER_13_465 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_481 ();
 sg13g2_fill_2 FILLER_13_495 ();
 sg13g2_fill_2 FILLER_13_552 ();
 sg13g2_fill_2 FILLER_13_573 ();
 sg13g2_fill_1 FILLER_13_597 ();
 sg13g2_fill_2 FILLER_13_737 ();
 sg13g2_fill_1 FILLER_13_739 ();
 sg13g2_fill_2 FILLER_13_753 ();
 sg13g2_fill_2 FILLER_13_807 ();
 sg13g2_fill_1 FILLER_13_809 ();
 sg13g2_fill_2 FILLER_13_834 ();
 sg13g2_fill_2 FILLER_13_886 ();
 sg13g2_fill_2 FILLER_13_895 ();
 sg13g2_fill_2 FILLER_13_1000 ();
 sg13g2_fill_1 FILLER_13_1002 ();
 sg13g2_fill_1 FILLER_13_1026 ();
 sg13g2_fill_2 FILLER_13_1059 ();
 sg13g2_fill_1 FILLER_13_1065 ();
 sg13g2_fill_2 FILLER_13_1093 ();
 sg13g2_fill_1 FILLER_13_1136 ();
 sg13g2_fill_1 FILLER_13_1235 ();
 sg13g2_fill_2 FILLER_13_1295 ();
 sg13g2_fill_2 FILLER_13_1324 ();
 sg13g2_decap_4 FILLER_13_1342 ();
 sg13g2_fill_2 FILLER_13_1374 ();
 sg13g2_fill_1 FILLER_13_1376 ();
 sg13g2_fill_2 FILLER_13_1381 ();
 sg13g2_fill_1 FILLER_13_1396 ();
 sg13g2_fill_2 FILLER_13_1413 ();
 sg13g2_fill_1 FILLER_13_1415 ();
 sg13g2_fill_2 FILLER_13_1436 ();
 sg13g2_fill_1 FILLER_13_1438 ();
 sg13g2_decap_4 FILLER_13_1474 ();
 sg13g2_fill_2 FILLER_13_1485 ();
 sg13g2_fill_2 FILLER_13_1501 ();
 sg13g2_fill_1 FILLER_13_1503 ();
 sg13g2_fill_1 FILLER_13_1589 ();
 sg13g2_fill_2 FILLER_13_1627 ();
 sg13g2_decap_4 FILLER_13_1693 ();
 sg13g2_fill_2 FILLER_13_1697 ();
 sg13g2_fill_2 FILLER_13_1717 ();
 sg13g2_fill_1 FILLER_13_1747 ();
 sg13g2_decap_4 FILLER_13_1766 ();
 sg13g2_fill_1 FILLER_13_1770 ();
 sg13g2_fill_2 FILLER_13_1815 ();
 sg13g2_fill_2 FILLER_13_1822 ();
 sg13g2_fill_1 FILLER_13_1838 ();
 sg13g2_fill_1 FILLER_13_1875 ();
 sg13g2_fill_1 FILLER_13_1913 ();
 sg13g2_fill_2 FILLER_13_1925 ();
 sg13g2_fill_2 FILLER_13_1956 ();
 sg13g2_fill_2 FILLER_13_1964 ();
 sg13g2_fill_1 FILLER_13_1966 ();
 sg13g2_decap_4 FILLER_13_1993 ();
 sg13g2_fill_1 FILLER_13_2011 ();
 sg13g2_decap_4 FILLER_13_2024 ();
 sg13g2_fill_2 FILLER_13_2071 ();
 sg13g2_fill_1 FILLER_13_2073 ();
 sg13g2_decap_8 FILLER_13_2078 ();
 sg13g2_fill_1 FILLER_13_2118 ();
 sg13g2_decap_4 FILLER_13_2125 ();
 sg13g2_fill_1 FILLER_13_2129 ();
 sg13g2_fill_2 FILLER_13_2144 ();
 sg13g2_decap_4 FILLER_13_2186 ();
 sg13g2_fill_2 FILLER_13_2190 ();
 sg13g2_fill_1 FILLER_13_2259 ();
 sg13g2_fill_2 FILLER_13_2269 ();
 sg13g2_fill_1 FILLER_13_2271 ();
 sg13g2_fill_2 FILLER_13_2289 ();
 sg13g2_fill_1 FILLER_13_2291 ();
 sg13g2_fill_1 FILLER_13_2300 ();
 sg13g2_fill_1 FILLER_13_2352 ();
 sg13g2_decap_8 FILLER_13_2380 ();
 sg13g2_fill_1 FILLER_13_2387 ();
 sg13g2_fill_1 FILLER_13_2452 ();
 sg13g2_fill_2 FILLER_13_2509 ();
 sg13g2_fill_2 FILLER_13_2550 ();
 sg13g2_fill_2 FILLER_13_2588 ();
 sg13g2_fill_1 FILLER_13_2590 ();
 sg13g2_fill_2 FILLER_13_2671 ();
 sg13g2_fill_1 FILLER_13_2673 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_33 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_decap_4 FILLER_14_148 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_4 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_193 ();
 sg13g2_fill_2 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_4 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_388 ();
 sg13g2_fill_1 FILLER_14_426 ();
 sg13g2_fill_1 FILLER_14_473 ();
 sg13g2_fill_2 FILLER_14_524 ();
 sg13g2_fill_1 FILLER_14_526 ();
 sg13g2_fill_1 FILLER_14_544 ();
 sg13g2_fill_2 FILLER_14_675 ();
 sg13g2_fill_1 FILLER_14_737 ();
 sg13g2_fill_2 FILLER_14_756 ();
 sg13g2_fill_1 FILLER_14_758 ();
 sg13g2_fill_2 FILLER_14_914 ();
 sg13g2_fill_1 FILLER_14_916 ();
 sg13g2_fill_1 FILLER_14_984 ();
 sg13g2_fill_1 FILLER_14_1031 ();
 sg13g2_fill_2 FILLER_14_1075 ();
 sg13g2_fill_2 FILLER_14_1086 ();
 sg13g2_fill_2 FILLER_14_1098 ();
 sg13g2_fill_1 FILLER_14_1100 ();
 sg13g2_decap_4 FILLER_14_1119 ();
 sg13g2_fill_2 FILLER_14_1128 ();
 sg13g2_fill_2 FILLER_14_1156 ();
 sg13g2_fill_1 FILLER_14_1192 ();
 sg13g2_fill_1 FILLER_14_1256 ();
 sg13g2_fill_1 FILLER_14_1263 ();
 sg13g2_decap_4 FILLER_14_1302 ();
 sg13g2_fill_1 FILLER_14_1355 ();
 sg13g2_fill_2 FILLER_14_1434 ();
 sg13g2_fill_1 FILLER_14_1451 ();
 sg13g2_decap_4 FILLER_14_1462 ();
 sg13g2_decap_8 FILLER_14_1475 ();
 sg13g2_fill_2 FILLER_14_1482 ();
 sg13g2_decap_8 FILLER_14_1490 ();
 sg13g2_fill_2 FILLER_14_1497 ();
 sg13g2_fill_1 FILLER_14_1499 ();
 sg13g2_fill_2 FILLER_14_1504 ();
 sg13g2_fill_2 FILLER_14_1593 ();
 sg13g2_fill_2 FILLER_14_1614 ();
 sg13g2_fill_1 FILLER_14_1669 ();
 sg13g2_fill_1 FILLER_14_1679 ();
 sg13g2_fill_2 FILLER_14_1734 ();
 sg13g2_fill_1 FILLER_14_1736 ();
 sg13g2_decap_4 FILLER_14_1746 ();
 sg13g2_decap_8 FILLER_14_1778 ();
 sg13g2_fill_1 FILLER_14_1785 ();
 sg13g2_fill_1 FILLER_14_1817 ();
 sg13g2_fill_1 FILLER_14_1826 ();
 sg13g2_fill_1 FILLER_14_1835 ();
 sg13g2_decap_8 FILLER_14_1863 ();
 sg13g2_fill_1 FILLER_14_1870 ();
 sg13g2_fill_1 FILLER_14_1900 ();
 sg13g2_fill_2 FILLER_14_1925 ();
 sg13g2_fill_2 FILLER_14_1956 ();
 sg13g2_fill_2 FILLER_14_2012 ();
 sg13g2_fill_1 FILLER_14_2014 ();
 sg13g2_fill_1 FILLER_14_2053 ();
 sg13g2_fill_1 FILLER_14_2060 ();
 sg13g2_fill_2 FILLER_14_2083 ();
 sg13g2_fill_1 FILLER_14_2085 ();
 sg13g2_fill_2 FILLER_14_2090 ();
 sg13g2_fill_2 FILLER_14_2108 ();
 sg13g2_decap_4 FILLER_14_2129 ();
 sg13g2_fill_1 FILLER_14_2133 ();
 sg13g2_fill_2 FILLER_14_2138 ();
 sg13g2_fill_1 FILLER_14_2140 ();
 sg13g2_fill_1 FILLER_14_2177 ();
 sg13g2_fill_2 FILLER_14_2240 ();
 sg13g2_fill_2 FILLER_14_2252 ();
 sg13g2_fill_1 FILLER_14_2254 ();
 sg13g2_decap_4 FILLER_14_2268 ();
 sg13g2_fill_1 FILLER_14_2272 ();
 sg13g2_fill_2 FILLER_14_2333 ();
 sg13g2_fill_1 FILLER_14_2335 ();
 sg13g2_fill_2 FILLER_14_2340 ();
 sg13g2_fill_1 FILLER_14_2348 ();
 sg13g2_decap_8 FILLER_14_2367 ();
 sg13g2_fill_2 FILLER_14_2374 ();
 sg13g2_fill_1 FILLER_14_2376 ();
 sg13g2_fill_2 FILLER_14_2439 ();
 sg13g2_fill_1 FILLER_14_2441 ();
 sg13g2_fill_1 FILLER_14_2459 ();
 sg13g2_decap_8 FILLER_14_2504 ();
 sg13g2_decap_4 FILLER_14_2511 ();
 sg13g2_fill_1 FILLER_14_2515 ();
 sg13g2_fill_1 FILLER_14_2525 ();
 sg13g2_fill_2 FILLER_14_2581 ();
 sg13g2_fill_1 FILLER_14_2583 ();
 sg13g2_fill_2 FILLER_14_2620 ();
 sg13g2_fill_2 FILLER_14_2671 ();
 sg13g2_fill_1 FILLER_14_2673 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_432 ();
 sg13g2_fill_2 FILLER_15_538 ();
 sg13g2_fill_1 FILLER_15_567 ();
 sg13g2_fill_1 FILLER_15_574 ();
 sg13g2_fill_2 FILLER_15_589 ();
 sg13g2_fill_1 FILLER_15_591 ();
 sg13g2_fill_2 FILLER_15_714 ();
 sg13g2_fill_2 FILLER_15_734 ();
 sg13g2_fill_2 FILLER_15_763 ();
 sg13g2_fill_1 FILLER_15_806 ();
 sg13g2_fill_2 FILLER_15_833 ();
 sg13g2_fill_1 FILLER_15_884 ();
 sg13g2_fill_1 FILLER_15_1022 ();
 sg13g2_fill_2 FILLER_15_1035 ();
 sg13g2_fill_1 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1102 ();
 sg13g2_fill_2 FILLER_15_1109 ();
 sg13g2_fill_1 FILLER_15_1111 ();
 sg13g2_fill_2 FILLER_15_1125 ();
 sg13g2_fill_1 FILLER_15_1127 ();
 sg13g2_fill_2 FILLER_15_1143 ();
 sg13g2_decap_4 FILLER_15_1159 ();
 sg13g2_fill_2 FILLER_15_1163 ();
 sg13g2_fill_1 FILLER_15_1207 ();
 sg13g2_fill_2 FILLER_15_1215 ();
 sg13g2_fill_1 FILLER_15_1256 ();
 sg13g2_fill_1 FILLER_15_1266 ();
 sg13g2_decap_4 FILLER_15_1312 ();
 sg13g2_fill_1 FILLER_15_1316 ();
 sg13g2_fill_1 FILLER_15_1320 ();
 sg13g2_fill_2 FILLER_15_1327 ();
 sg13g2_fill_1 FILLER_15_1329 ();
 sg13g2_fill_2 FILLER_15_1339 ();
 sg13g2_fill_1 FILLER_15_1341 ();
 sg13g2_decap_4 FILLER_15_1348 ();
 sg13g2_fill_2 FILLER_15_1366 ();
 sg13g2_fill_2 FILLER_15_1448 ();
 sg13g2_fill_2 FILLER_15_1506 ();
 sg13g2_decap_8 FILLER_15_1518 ();
 sg13g2_fill_2 FILLER_15_1525 ();
 sg13g2_fill_1 FILLER_15_1527 ();
 sg13g2_fill_1 FILLER_15_1541 ();
 sg13g2_fill_1 FILLER_15_1566 ();
 sg13g2_fill_2 FILLER_15_1586 ();
 sg13g2_fill_1 FILLER_15_1597 ();
 sg13g2_fill_1 FILLER_15_1611 ();
 sg13g2_fill_1 FILLER_15_1628 ();
 sg13g2_fill_2 FILLER_15_1653 ();
 sg13g2_decap_4 FILLER_15_1688 ();
 sg13g2_fill_1 FILLER_15_1692 ();
 sg13g2_fill_2 FILLER_15_1721 ();
 sg13g2_fill_1 FILLER_15_1723 ();
 sg13g2_decap_4 FILLER_15_1759 ();
 sg13g2_fill_1 FILLER_15_1818 ();
 sg13g2_fill_2 FILLER_15_1842 ();
 sg13g2_fill_1 FILLER_15_1844 ();
 sg13g2_fill_2 FILLER_15_1850 ();
 sg13g2_fill_2 FILLER_15_1870 ();
 sg13g2_fill_1 FILLER_15_1872 ();
 sg13g2_fill_1 FILLER_15_1915 ();
 sg13g2_decap_4 FILLER_15_1930 ();
 sg13g2_fill_1 FILLER_15_1934 ();
 sg13g2_fill_2 FILLER_15_1976 ();
 sg13g2_decap_8 FILLER_15_2023 ();
 sg13g2_fill_1 FILLER_15_2030 ();
 sg13g2_decap_4 FILLER_15_2071 ();
 sg13g2_fill_2 FILLER_15_2111 ();
 sg13g2_fill_2 FILLER_15_2119 ();
 sg13g2_fill_1 FILLER_15_2121 ();
 sg13g2_decap_4 FILLER_15_2181 ();
 sg13g2_decap_8 FILLER_15_2244 ();
 sg13g2_fill_1 FILLER_15_2251 ();
 sg13g2_fill_2 FILLER_15_2261 ();
 sg13g2_decap_4 FILLER_15_2267 ();
 sg13g2_fill_1 FILLER_15_2271 ();
 sg13g2_decap_4 FILLER_15_2276 ();
 sg13g2_fill_2 FILLER_15_2280 ();
 sg13g2_decap_4 FILLER_15_2293 ();
 sg13g2_fill_2 FILLER_15_2360 ();
 sg13g2_fill_2 FILLER_15_2372 ();
 sg13g2_fill_1 FILLER_15_2379 ();
 sg13g2_fill_1 FILLER_15_2406 ();
 sg13g2_fill_1 FILLER_15_2456 ();
 sg13g2_fill_2 FILLER_15_2484 ();
 sg13g2_decap_8 FILLER_15_2499 ();
 sg13g2_fill_1 FILLER_15_2524 ();
 sg13g2_fill_1 FILLER_15_2571 ();
 sg13g2_fill_1 FILLER_15_2673 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_27 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_decap_8 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_171 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_decap_8 FILLER_16_192 ();
 sg13g2_fill_2 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_303 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_372 ();
 sg13g2_fill_1 FILLER_16_444 ();
 sg13g2_fill_2 FILLER_16_458 ();
 sg13g2_fill_1 FILLER_16_534 ();
 sg13g2_fill_1 FILLER_16_544 ();
 sg13g2_fill_2 FILLER_16_561 ();
 sg13g2_fill_1 FILLER_16_627 ();
 sg13g2_fill_2 FILLER_16_686 ();
 sg13g2_fill_2 FILLER_16_702 ();
 sg13g2_fill_2 FILLER_16_732 ();
 sg13g2_fill_2 FILLER_16_793 ();
 sg13g2_fill_2 FILLER_16_810 ();
 sg13g2_fill_1 FILLER_16_812 ();
 sg13g2_fill_1 FILLER_16_849 ();
 sg13g2_fill_2 FILLER_16_873 ();
 sg13g2_fill_2 FILLER_16_903 ();
 sg13g2_fill_1 FILLER_16_905 ();
 sg13g2_fill_2 FILLER_16_919 ();
 sg13g2_fill_2 FILLER_16_934 ();
 sg13g2_fill_1 FILLER_16_1006 ();
 sg13g2_fill_2 FILLER_16_1025 ();
 sg13g2_fill_2 FILLER_16_1097 ();
 sg13g2_fill_1 FILLER_16_1099 ();
 sg13g2_fill_2 FILLER_16_1142 ();
 sg13g2_fill_1 FILLER_16_1144 ();
 sg13g2_fill_1 FILLER_16_1159 ();
 sg13g2_fill_1 FILLER_16_1216 ();
 sg13g2_fill_2 FILLER_16_1227 ();
 sg13g2_fill_2 FILLER_16_1239 ();
 sg13g2_fill_1 FILLER_16_1272 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_fill_2 FILLER_16_1326 ();
 sg13g2_fill_1 FILLER_16_1328 ();
 sg13g2_decap_8 FILLER_16_1361 ();
 sg13g2_decap_8 FILLER_16_1368 ();
 sg13g2_fill_1 FILLER_16_1375 ();
 sg13g2_fill_2 FILLER_16_1380 ();
 sg13g2_fill_1 FILLER_16_1382 ();
 sg13g2_decap_4 FILLER_16_1388 ();
 sg13g2_fill_1 FILLER_16_1392 ();
 sg13g2_decap_4 FILLER_16_1407 ();
 sg13g2_decap_8 FILLER_16_1432 ();
 sg13g2_decap_8 FILLER_16_1439 ();
 sg13g2_decap_4 FILLER_16_1446 ();
 sg13g2_fill_2 FILLER_16_1450 ();
 sg13g2_decap_8 FILLER_16_1469 ();
 sg13g2_fill_2 FILLER_16_1494 ();
 sg13g2_decap_4 FILLER_16_1531 ();
 sg13g2_fill_1 FILLER_16_1560 ();
 sg13g2_fill_1 FILLER_16_1634 ();
 sg13g2_fill_2 FILLER_16_1678 ();
 sg13g2_decap_8 FILLER_16_1684 ();
 sg13g2_decap_8 FILLER_16_1691 ();
 sg13g2_decap_4 FILLER_16_1698 ();
 sg13g2_fill_2 FILLER_16_1707 ();
 sg13g2_fill_2 FILLER_16_1759 ();
 sg13g2_fill_1 FILLER_16_1805 ();
 sg13g2_decap_4 FILLER_16_1864 ();
 sg13g2_fill_1 FILLER_16_1868 ();
 sg13g2_decap_4 FILLER_16_1873 ();
 sg13g2_decap_4 FILLER_16_1917 ();
 sg13g2_fill_2 FILLER_16_1952 ();
 sg13g2_fill_1 FILLER_16_1954 ();
 sg13g2_fill_2 FILLER_16_1995 ();
 sg13g2_fill_1 FILLER_16_1997 ();
 sg13g2_fill_2 FILLER_16_2007 ();
 sg13g2_decap_4 FILLER_16_2099 ();
 sg13g2_fill_2 FILLER_16_2103 ();
 sg13g2_fill_2 FILLER_16_2128 ();
 sg13g2_fill_2 FILLER_16_2166 ();
 sg13g2_fill_1 FILLER_16_2168 ();
 sg13g2_decap_4 FILLER_16_2178 ();
 sg13g2_decap_4 FILLER_16_2190 ();
 sg13g2_fill_2 FILLER_16_2229 ();
 sg13g2_fill_1 FILLER_16_2275 ();
 sg13g2_fill_1 FILLER_16_2285 ();
 sg13g2_fill_2 FILLER_16_2295 ();
 sg13g2_fill_1 FILLER_16_2309 ();
 sg13g2_fill_2 FILLER_16_2315 ();
 sg13g2_fill_1 FILLER_16_2317 ();
 sg13g2_fill_2 FILLER_16_2336 ();
 sg13g2_fill_1 FILLER_16_2338 ();
 sg13g2_fill_2 FILLER_16_2406 ();
 sg13g2_fill_1 FILLER_16_2408 ();
 sg13g2_fill_1 FILLER_16_2431 ();
 sg13g2_fill_2 FILLER_16_2481 ();
 sg13g2_fill_1 FILLER_16_2483 ();
 sg13g2_decap_4 FILLER_16_2497 ();
 sg13g2_fill_2 FILLER_16_2528 ();
 sg13g2_fill_2 FILLER_16_2565 ();
 sg13g2_fill_2 FILLER_16_2603 ();
 sg13g2_fill_1 FILLER_16_2673 ();
 sg13g2_fill_2 FILLER_17_46 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_160 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_fill_2 FILLER_17_196 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_476 ();
 sg13g2_fill_1 FILLER_17_521 ();
 sg13g2_fill_2 FILLER_17_552 ();
 sg13g2_fill_2 FILLER_17_567 ();
 sg13g2_fill_1 FILLER_17_569 ();
 sg13g2_fill_2 FILLER_17_575 ();
 sg13g2_fill_1 FILLER_17_577 ();
 sg13g2_fill_2 FILLER_17_596 ();
 sg13g2_fill_1 FILLER_17_598 ();
 sg13g2_fill_1 FILLER_17_603 ();
 sg13g2_fill_2 FILLER_17_620 ();
 sg13g2_fill_2 FILLER_17_635 ();
 sg13g2_fill_2 FILLER_17_772 ();
 sg13g2_fill_2 FILLER_17_789 ();
 sg13g2_fill_1 FILLER_17_791 ();
 sg13g2_fill_2 FILLER_17_803 ();
 sg13g2_fill_1 FILLER_17_805 ();
 sg13g2_fill_2 FILLER_17_836 ();
 sg13g2_fill_2 FILLER_17_923 ();
 sg13g2_fill_2 FILLER_17_958 ();
 sg13g2_fill_1 FILLER_17_1018 ();
 sg13g2_fill_2 FILLER_17_1037 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_fill_2 FILLER_17_1145 ();
 sg13g2_fill_1 FILLER_17_1166 ();
 sg13g2_fill_2 FILLER_17_1194 ();
 sg13g2_fill_1 FILLER_17_1210 ();
 sg13g2_fill_2 FILLER_17_1224 ();
 sg13g2_fill_2 FILLER_17_1265 ();
 sg13g2_fill_2 FILLER_17_1305 ();
 sg13g2_decap_8 FILLER_17_1363 ();
 sg13g2_fill_2 FILLER_17_1370 ();
 sg13g2_decap_4 FILLER_17_1385 ();
 sg13g2_decap_8 FILLER_17_1440 ();
 sg13g2_fill_2 FILLER_17_1447 ();
 sg13g2_fill_1 FILLER_17_1449 ();
 sg13g2_fill_1 FILLER_17_1455 ();
 sg13g2_fill_2 FILLER_17_1484 ();
 sg13g2_fill_1 FILLER_17_1486 ();
 sg13g2_fill_2 FILLER_17_1500 ();
 sg13g2_fill_2 FILLER_17_1521 ();
 sg13g2_fill_1 FILLER_17_1523 ();
 sg13g2_fill_1 FILLER_17_1540 ();
 sg13g2_decap_4 FILLER_17_1588 ();
 sg13g2_fill_2 FILLER_17_1714 ();
 sg13g2_fill_1 FILLER_17_1716 ();
 sg13g2_fill_2 FILLER_17_1734 ();
 sg13g2_fill_1 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_fill_2 FILLER_17_1764 ();
 sg13g2_fill_1 FILLER_17_1798 ();
 sg13g2_fill_2 FILLER_17_1812 ();
 sg13g2_fill_1 FILLER_17_1814 ();
 sg13g2_decap_8 FILLER_17_1855 ();
 sg13g2_decap_4 FILLER_17_1862 ();
 sg13g2_fill_2 FILLER_17_1866 ();
 sg13g2_fill_2 FILLER_17_1903 ();
 sg13g2_fill_1 FILLER_17_1905 ();
 sg13g2_fill_2 FILLER_17_1933 ();
 sg13g2_fill_1 FILLER_17_1935 ();
 sg13g2_fill_2 FILLER_17_1968 ();
 sg13g2_fill_1 FILLER_17_1970 ();
 sg13g2_fill_1 FILLER_17_1992 ();
 sg13g2_decap_4 FILLER_17_2002 ();
 sg13g2_fill_2 FILLER_17_2038 ();
 sg13g2_fill_1 FILLER_17_2040 ();
 sg13g2_decap_8 FILLER_17_2068 ();
 sg13g2_fill_1 FILLER_17_2111 ();
 sg13g2_decap_8 FILLER_17_2144 ();
 sg13g2_decap_8 FILLER_17_2151 ();
 sg13g2_decap_8 FILLER_17_2158 ();
 sg13g2_decap_8 FILLER_17_2165 ();
 sg13g2_decap_8 FILLER_17_2172 ();
 sg13g2_fill_1 FILLER_17_2179 ();
 sg13g2_decap_8 FILLER_17_2184 ();
 sg13g2_decap_8 FILLER_17_2191 ();
 sg13g2_fill_2 FILLER_17_2198 ();
 sg13g2_fill_2 FILLER_17_2209 ();
 sg13g2_fill_1 FILLER_17_2216 ();
 sg13g2_fill_2 FILLER_17_2227 ();
 sg13g2_fill_2 FILLER_17_2319 ();
 sg13g2_fill_2 FILLER_17_2325 ();
 sg13g2_fill_2 FILLER_17_2349 ();
 sg13g2_fill_2 FILLER_17_2422 ();
 sg13g2_fill_1 FILLER_17_2424 ();
 sg13g2_decap_8 FILLER_17_2477 ();
 sg13g2_fill_2 FILLER_17_2484 ();
 sg13g2_fill_2 FILLER_17_2491 ();
 sg13g2_fill_2 FILLER_17_2523 ();
 sg13g2_fill_1 FILLER_17_2540 ();
 sg13g2_fill_2 FILLER_17_2567 ();
 sg13g2_fill_1 FILLER_17_2569 ();
 sg13g2_fill_2 FILLER_17_2596 ();
 sg13g2_fill_1 FILLER_17_2598 ();
 sg13g2_fill_2 FILLER_17_2613 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_426 ();
 sg13g2_fill_1 FILLER_18_475 ();
 sg13g2_fill_1 FILLER_18_507 ();
 sg13g2_fill_1 FILLER_18_565 ();
 sg13g2_fill_2 FILLER_18_570 ();
 sg13g2_fill_1 FILLER_18_588 ();
 sg13g2_fill_2 FILLER_18_607 ();
 sg13g2_fill_1 FILLER_18_637 ();
 sg13g2_fill_2 FILLER_18_647 ();
 sg13g2_fill_2 FILLER_18_667 ();
 sg13g2_fill_1 FILLER_18_700 ();
 sg13g2_fill_2 FILLER_18_826 ();
 sg13g2_fill_1 FILLER_18_944 ();
 sg13g2_fill_2 FILLER_18_963 ();
 sg13g2_fill_2 FILLER_18_975 ();
 sg13g2_fill_2 FILLER_18_1033 ();
 sg13g2_fill_2 FILLER_18_1053 ();
 sg13g2_fill_1 FILLER_18_1063 ();
 sg13g2_fill_2 FILLER_18_1080 ();
 sg13g2_fill_1 FILLER_18_1082 ();
 sg13g2_fill_2 FILLER_18_1153 ();
 sg13g2_fill_1 FILLER_18_1192 ();
 sg13g2_fill_1 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_fill_1 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1313 ();
 sg13g2_fill_1 FILLER_18_1335 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_4 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1473 ();
 sg13g2_fill_1 FILLER_18_1542 ();
 sg13g2_decap_4 FILLER_18_1607 ();
 sg13g2_fill_2 FILLER_18_1656 ();
 sg13g2_fill_2 FILLER_18_1671 ();
 sg13g2_fill_2 FILLER_18_1718 ();
 sg13g2_fill_1 FILLER_18_1720 ();
 sg13g2_decap_4 FILLER_18_1730 ();
 sg13g2_fill_2 FILLER_18_1734 ();
 sg13g2_decap_4 FILLER_18_1745 ();
 sg13g2_fill_1 FILLER_18_1749 ();
 sg13g2_fill_2 FILLER_18_1808 ();
 sg13g2_fill_2 FILLER_18_1860 ();
 sg13g2_fill_2 FILLER_18_1921 ();
 sg13g2_fill_1 FILLER_18_1969 ();
 sg13g2_fill_2 FILLER_18_2020 ();
 sg13g2_fill_2 FILLER_18_2036 ();
 sg13g2_fill_2 FILLER_18_2051 ();
 sg13g2_fill_1 FILLER_18_2072 ();
 sg13g2_fill_2 FILLER_18_2090 ();
 sg13g2_fill_2 FILLER_18_2128 ();
 sg13g2_fill_1 FILLER_18_2130 ();
 sg13g2_decap_8 FILLER_18_2135 ();
 sg13g2_decap_8 FILLER_18_2142 ();
 sg13g2_decap_8 FILLER_18_2149 ();
 sg13g2_fill_2 FILLER_18_2156 ();
 sg13g2_fill_1 FILLER_18_2158 ();
 sg13g2_fill_2 FILLER_18_2204 ();
 sg13g2_fill_2 FILLER_18_2225 ();
 sg13g2_fill_1 FILLER_18_2227 ();
 sg13g2_fill_2 FILLER_18_2256 ();
 sg13g2_fill_1 FILLER_18_2271 ();
 sg13g2_fill_2 FILLER_18_2335 ();
 sg13g2_fill_1 FILLER_18_2337 ();
 sg13g2_fill_1 FILLER_18_2416 ();
 sg13g2_fill_1 FILLER_18_2434 ();
 sg13g2_decap_8 FILLER_18_2510 ();
 sg13g2_decap_8 FILLER_18_2517 ();
 sg13g2_fill_1 FILLER_18_2524 ();
 sg13g2_decap_8 FILLER_18_2529 ();
 sg13g2_fill_2 FILLER_18_2577 ();
 sg13g2_fill_1 FILLER_18_2579 ();
 sg13g2_fill_2 FILLER_18_2638 ();
 sg13g2_fill_1 FILLER_18_2645 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_357 ();
 sg13g2_fill_1 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_411 ();
 sg13g2_fill_1 FILLER_19_460 ();
 sg13g2_fill_2 FILLER_19_593 ();
 sg13g2_fill_1 FILLER_19_595 ();
 sg13g2_fill_2 FILLER_19_633 ();
 sg13g2_fill_1 FILLER_19_651 ();
 sg13g2_fill_1 FILLER_19_740 ();
 sg13g2_fill_1 FILLER_19_815 ();
 sg13g2_fill_2 FILLER_19_895 ();
 sg13g2_fill_2 FILLER_19_968 ();
 sg13g2_fill_2 FILLER_19_983 ();
 sg13g2_fill_2 FILLER_19_1013 ();
 sg13g2_fill_1 FILLER_19_1015 ();
 sg13g2_fill_1 FILLER_19_1062 ();
 sg13g2_fill_2 FILLER_19_1097 ();
 sg13g2_fill_1 FILLER_19_1114 ();
 sg13g2_fill_1 FILLER_19_1125 ();
 sg13g2_fill_1 FILLER_19_1140 ();
 sg13g2_fill_1 FILLER_19_1213 ();
 sg13g2_fill_2 FILLER_19_1259 ();
 sg13g2_fill_1 FILLER_19_1261 ();
 sg13g2_fill_2 FILLER_19_1265 ();
 sg13g2_fill_2 FILLER_19_1285 ();
 sg13g2_decap_8 FILLER_19_1297 ();
 sg13g2_decap_4 FILLER_19_1304 ();
 sg13g2_fill_1 FILLER_19_1308 ();
 sg13g2_fill_2 FILLER_19_1374 ();
 sg13g2_fill_1 FILLER_19_1393 ();
 sg13g2_fill_1 FILLER_19_1400 ();
 sg13g2_fill_2 FILLER_19_1439 ();
 sg13g2_fill_2 FILLER_19_1493 ();
 sg13g2_fill_1 FILLER_19_1495 ();
 sg13g2_fill_2 FILLER_19_1508 ();
 sg13g2_fill_2 FILLER_19_1532 ();
 sg13g2_fill_1 FILLER_19_1534 ();
 sg13g2_fill_2 FILLER_19_1563 ();
 sg13g2_fill_1 FILLER_19_1565 ();
 sg13g2_decap_4 FILLER_19_1598 ();
 sg13g2_fill_2 FILLER_19_1602 ();
 sg13g2_fill_2 FILLER_19_1677 ();
 sg13g2_fill_2 FILLER_19_1731 ();
 sg13g2_fill_1 FILLER_19_1733 ();
 sg13g2_decap_4 FILLER_19_1741 ();
 sg13g2_fill_1 FILLER_19_1745 ();
 sg13g2_decap_8 FILLER_19_1764 ();
 sg13g2_decap_4 FILLER_19_1771 ();
 sg13g2_fill_1 FILLER_19_1797 ();
 sg13g2_decap_4 FILLER_19_1802 ();
 sg13g2_fill_1 FILLER_19_1806 ();
 sg13g2_fill_2 FILLER_19_1852 ();
 sg13g2_fill_1 FILLER_19_1875 ();
 sg13g2_fill_2 FILLER_19_1888 ();
 sg13g2_decap_4 FILLER_19_1913 ();
 sg13g2_fill_1 FILLER_19_1917 ();
 sg13g2_fill_2 FILLER_19_2013 ();
 sg13g2_fill_2 FILLER_19_2086 ();
 sg13g2_fill_1 FILLER_19_2112 ();
 sg13g2_fill_1 FILLER_19_2157 ();
 sg13g2_fill_2 FILLER_19_2394 ();
 sg13g2_fill_1 FILLER_19_2396 ();
 sg13g2_decap_8 FILLER_19_2419 ();
 sg13g2_fill_2 FILLER_19_2430 ();
 sg13g2_fill_1 FILLER_19_2432 ();
 sg13g2_fill_2 FILLER_19_2446 ();
 sg13g2_fill_1 FILLER_19_2452 ();
 sg13g2_fill_1 FILLER_19_2502 ();
 sg13g2_decap_8 FILLER_19_2516 ();
 sg13g2_decap_8 FILLER_19_2523 ();
 sg13g2_decap_4 FILLER_19_2530 ();
 sg13g2_fill_1 FILLER_19_2534 ();
 sg13g2_fill_2 FILLER_19_2581 ();
 sg13g2_fill_1 FILLER_19_2583 ();
 sg13g2_fill_2 FILLER_19_2624 ();
 sg13g2_fill_1 FILLER_19_2626 ();
 sg13g2_fill_1 FILLER_19_2673 ();
 sg13g2_fill_1 FILLER_20_17 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_decap_8 FILLER_20_178 ();
 sg13g2_decap_4 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_fill_2 FILLER_20_343 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_493 ();
 sg13g2_fill_2 FILLER_20_521 ();
 sg13g2_fill_2 FILLER_20_582 ();
 sg13g2_fill_2 FILLER_20_643 ();
 sg13g2_fill_1 FILLER_20_673 ();
 sg13g2_fill_1 FILLER_20_710 ();
 sg13g2_fill_2 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_783 ();
 sg13g2_fill_2 FILLER_20_932 ();
 sg13g2_fill_2 FILLER_20_1009 ();
 sg13g2_fill_2 FILLER_20_1017 ();
 sg13g2_fill_1 FILLER_20_1019 ();
 sg13g2_fill_1 FILLER_20_1061 ();
 sg13g2_fill_1 FILLER_20_1159 ();
 sg13g2_fill_2 FILLER_20_1182 ();
 sg13g2_fill_1 FILLER_20_1217 ();
 sg13g2_decap_4 FILLER_20_1282 ();
 sg13g2_decap_8 FILLER_20_1295 ();
 sg13g2_fill_1 FILLER_20_1334 ();
 sg13g2_fill_2 FILLER_20_1361 ();
 sg13g2_fill_1 FILLER_20_1363 ();
 sg13g2_fill_2 FILLER_20_1414 ();
 sg13g2_fill_1 FILLER_20_1416 ();
 sg13g2_fill_1 FILLER_20_1481 ();
 sg13g2_fill_2 FILLER_20_1491 ();
 sg13g2_fill_1 FILLER_20_1493 ();
 sg13g2_fill_2 FILLER_20_1551 ();
 sg13g2_fill_1 FILLER_20_1583 ();
 sg13g2_fill_1 FILLER_20_1612 ();
 sg13g2_fill_1 FILLER_20_1618 ();
 sg13g2_fill_2 FILLER_20_1625 ();
 sg13g2_fill_2 FILLER_20_1635 ();
 sg13g2_fill_1 FILLER_20_1637 ();
 sg13g2_fill_2 FILLER_20_1649 ();
 sg13g2_fill_1 FILLER_20_1651 ();
 sg13g2_fill_2 FILLER_20_1665 ();
 sg13g2_fill_2 FILLER_20_1700 ();
 sg13g2_fill_1 FILLER_20_1702 ();
 sg13g2_decap_4 FILLER_20_1755 ();
 sg13g2_decap_8 FILLER_20_1908 ();
 sg13g2_decap_4 FILLER_20_1915 ();
 sg13g2_fill_2 FILLER_20_1946 ();
 sg13g2_fill_1 FILLER_20_1948 ();
 sg13g2_fill_2 FILLER_20_1980 ();
 sg13g2_decap_4 FILLER_20_2018 ();
 sg13g2_fill_1 FILLER_20_2030 ();
 sg13g2_fill_2 FILLER_20_2057 ();
 sg13g2_fill_1 FILLER_20_2059 ();
 sg13g2_fill_2 FILLER_20_2257 ();
 sg13g2_fill_1 FILLER_20_2259 ();
 sg13g2_fill_2 FILLER_20_2268 ();
 sg13g2_fill_2 FILLER_20_2283 ();
 sg13g2_fill_1 FILLER_20_2285 ();
 sg13g2_fill_2 FILLER_20_2317 ();
 sg13g2_fill_2 FILLER_20_2363 ();
 sg13g2_fill_1 FILLER_20_2418 ();
 sg13g2_fill_2 FILLER_20_2468 ();
 sg13g2_fill_1 FILLER_20_2470 ();
 sg13g2_decap_8 FILLER_20_2512 ();
 sg13g2_decap_8 FILLER_20_2519 ();
 sg13g2_decap_8 FILLER_20_2526 ();
 sg13g2_decap_4 FILLER_20_2533 ();
 sg13g2_fill_2 FILLER_20_2564 ();
 sg13g2_fill_1 FILLER_20_2566 ();
 sg13g2_fill_1 FILLER_20_2603 ();
 sg13g2_fill_1 FILLER_20_2640 ();
 sg13g2_fill_1 FILLER_20_2673 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_fill_2 FILLER_21_418 ();
 sg13g2_fill_1 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_541 ();
 sg13g2_fill_1 FILLER_21_543 ();
 sg13g2_fill_2 FILLER_21_637 ();
 sg13g2_fill_1 FILLER_21_779 ();
 sg13g2_fill_2 FILLER_21_799 ();
 sg13g2_fill_1 FILLER_21_801 ();
 sg13g2_fill_1 FILLER_21_816 ();
 sg13g2_fill_2 FILLER_21_827 ();
 sg13g2_fill_2 FILLER_21_868 ();
 sg13g2_fill_2 FILLER_21_879 ();
 sg13g2_fill_1 FILLER_21_913 ();
 sg13g2_fill_2 FILLER_21_969 ();
 sg13g2_fill_2 FILLER_21_1006 ();
 sg13g2_fill_1 FILLER_21_1030 ();
 sg13g2_decap_4 FILLER_21_1051 ();
 sg13g2_fill_1 FILLER_21_1055 ();
 sg13g2_fill_2 FILLER_21_1064 ();
 sg13g2_fill_2 FILLER_21_1088 ();
 sg13g2_fill_2 FILLER_21_1104 ();
 sg13g2_fill_2 FILLER_21_1164 ();
 sg13g2_fill_1 FILLER_21_1193 ();
 sg13g2_fill_1 FILLER_21_1200 ();
 sg13g2_decap_4 FILLER_21_1291 ();
 sg13g2_fill_1 FILLER_21_1295 ();
 sg13g2_fill_2 FILLER_21_1341 ();
 sg13g2_fill_1 FILLER_21_1343 ();
 sg13g2_fill_2 FILLER_21_1391 ();
 sg13g2_fill_1 FILLER_21_1393 ();
 sg13g2_fill_1 FILLER_21_1456 ();
 sg13g2_fill_2 FILLER_21_1490 ();
 sg13g2_fill_2 FILLER_21_1526 ();
 sg13g2_fill_1 FILLER_21_1528 ();
 sg13g2_decap_4 FILLER_21_1612 ();
 sg13g2_fill_2 FILLER_21_1616 ();
 sg13g2_fill_2 FILLER_21_1632 ();
 sg13g2_decap_4 FILLER_21_1678 ();
 sg13g2_fill_1 FILLER_21_1682 ();
 sg13g2_fill_1 FILLER_21_1754 ();
 sg13g2_fill_1 FILLER_21_1764 ();
 sg13g2_fill_1 FILLER_21_1884 ();
 sg13g2_fill_2 FILLER_21_1906 ();
 sg13g2_fill_1 FILLER_21_1908 ();
 sg13g2_fill_1 FILLER_21_1930 ();
 sg13g2_fill_1 FILLER_21_2018 ();
 sg13g2_fill_1 FILLER_21_2033 ();
 sg13g2_fill_2 FILLER_21_2056 ();
 sg13g2_decap_8 FILLER_21_2071 ();
 sg13g2_fill_2 FILLER_21_2217 ();
 sg13g2_fill_2 FILLER_21_2232 ();
 sg13g2_fill_2 FILLER_21_2270 ();
 sg13g2_fill_2 FILLER_21_2304 ();
 sg13g2_fill_1 FILLER_21_2306 ();
 sg13g2_fill_2 FILLER_21_2348 ();
 sg13g2_fill_1 FILLER_21_2350 ();
 sg13g2_fill_1 FILLER_21_2368 ();
 sg13g2_fill_2 FILLER_21_2382 ();
 sg13g2_fill_1 FILLER_21_2384 ();
 sg13g2_fill_2 FILLER_21_2505 ();
 sg13g2_fill_1 FILLER_21_2533 ();
 sg13g2_fill_2 FILLER_21_2597 ();
 sg13g2_fill_2 FILLER_21_2613 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_fill_2 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_290 ();
 sg13g2_fill_2 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_625 ();
 sg13g2_fill_2 FILLER_22_738 ();
 sg13g2_fill_1 FILLER_22_750 ();
 sg13g2_fill_2 FILLER_22_769 ();
 sg13g2_fill_2 FILLER_22_808 ();
 sg13g2_fill_1 FILLER_22_831 ();
 sg13g2_fill_2 FILLER_22_841 ();
 sg13g2_fill_1 FILLER_22_843 ();
 sg13g2_fill_2 FILLER_22_977 ();
 sg13g2_fill_1 FILLER_22_979 ();
 sg13g2_fill_2 FILLER_22_989 ();
 sg13g2_fill_1 FILLER_22_991 ();
 sg13g2_fill_1 FILLER_22_1031 ();
 sg13g2_decap_8 FILLER_22_1047 ();
 sg13g2_decap_8 FILLER_22_1054 ();
 sg13g2_decap_4 FILLER_22_1061 ();
 sg13g2_fill_2 FILLER_22_1069 ();
 sg13g2_fill_1 FILLER_22_1071 ();
 sg13g2_fill_2 FILLER_22_1076 ();
 sg13g2_fill_1 FILLER_22_1214 ();
 sg13g2_fill_2 FILLER_22_1276 ();
 sg13g2_fill_1 FILLER_22_1306 ();
 sg13g2_fill_2 FILLER_22_1367 ();
 sg13g2_fill_1 FILLER_22_1369 ();
 sg13g2_decap_4 FILLER_22_1384 ();
 sg13g2_fill_2 FILLER_22_1442 ();
 sg13g2_fill_1 FILLER_22_1444 ();
 sg13g2_fill_1 FILLER_22_1550 ();
 sg13g2_fill_2 FILLER_22_1596 ();
 sg13g2_fill_2 FILLER_22_1610 ();
 sg13g2_fill_1 FILLER_22_1612 ();
 sg13g2_fill_1 FILLER_22_1623 ();
 sg13g2_decap_4 FILLER_22_1627 ();
 sg13g2_fill_2 FILLER_22_1637 ();
 sg13g2_fill_1 FILLER_22_1639 ();
 sg13g2_fill_2 FILLER_22_1645 ();
 sg13g2_fill_1 FILLER_22_1647 ();
 sg13g2_fill_2 FILLER_22_1689 ();
 sg13g2_fill_2 FILLER_22_1740 ();
 sg13g2_fill_1 FILLER_22_1742 ();
 sg13g2_fill_2 FILLER_22_1779 ();
 sg13g2_fill_1 FILLER_22_1781 ();
 sg13g2_fill_1 FILLER_22_1822 ();
 sg13g2_fill_2 FILLER_22_1882 ();
 sg13g2_fill_2 FILLER_22_1941 ();
 sg13g2_fill_1 FILLER_22_1959 ();
 sg13g2_fill_2 FILLER_22_2006 ();
 sg13g2_fill_1 FILLER_22_2008 ();
 sg13g2_decap_8 FILLER_22_2062 ();
 sg13g2_fill_2 FILLER_22_2077 ();
 sg13g2_fill_1 FILLER_22_2079 ();
 sg13g2_fill_1 FILLER_22_2099 ();
 sg13g2_fill_1 FILLER_22_2106 ();
 sg13g2_fill_2 FILLER_22_2157 ();
 sg13g2_fill_1 FILLER_22_2159 ();
 sg13g2_fill_1 FILLER_22_2195 ();
 sg13g2_fill_2 FILLER_22_2217 ();
 sg13g2_fill_2 FILLER_22_2268 ();
 sg13g2_fill_2 FILLER_22_2297 ();
 sg13g2_fill_1 FILLER_22_2299 ();
 sg13g2_fill_2 FILLER_22_2364 ();
 sg13g2_fill_1 FILLER_22_2441 ();
 sg13g2_fill_2 FILLER_22_2545 ();
 sg13g2_decap_4 FILLER_22_2584 ();
 sg13g2_fill_2 FILLER_22_2601 ();
 sg13g2_fill_1 FILLER_22_2603 ();
 sg13g2_fill_2 FILLER_22_2672 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_4 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_453 ();
 sg13g2_fill_2 FILLER_23_481 ();
 sg13g2_fill_1 FILLER_23_498 ();
 sg13g2_fill_1 FILLER_23_638 ();
 sg13g2_fill_1 FILLER_23_672 ();
 sg13g2_fill_2 FILLER_23_696 ();
 sg13g2_fill_1 FILLER_23_706 ();
 sg13g2_fill_2 FILLER_23_712 ();
 sg13g2_fill_2 FILLER_23_990 ();
 sg13g2_fill_1 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_1047 ();
 sg13g2_fill_1 FILLER_23_1054 ();
 sg13g2_decap_8 FILLER_23_1072 ();
 sg13g2_fill_1 FILLER_23_1079 ();
 sg13g2_fill_1 FILLER_23_1083 ();
 sg13g2_fill_1 FILLER_23_1112 ();
 sg13g2_fill_2 FILLER_23_1260 ();
 sg13g2_fill_1 FILLER_23_1330 ();
 sg13g2_fill_2 FILLER_23_1345 ();
 sg13g2_fill_2 FILLER_23_1372 ();
 sg13g2_fill_1 FILLER_23_1374 ();
 sg13g2_fill_2 FILLER_23_1384 ();
 sg13g2_fill_1 FILLER_23_1386 ();
 sg13g2_fill_1 FILLER_23_1402 ();
 sg13g2_fill_1 FILLER_23_1408 ();
 sg13g2_fill_2 FILLER_23_1479 ();
 sg13g2_fill_2 FILLER_23_1588 ();
 sg13g2_fill_1 FILLER_23_1620 ();
 sg13g2_decap_8 FILLER_23_1632 ();
 sg13g2_decap_8 FILLER_23_1681 ();
 sg13g2_decap_8 FILLER_23_1688 ();
 sg13g2_decap_4 FILLER_23_1695 ();
 sg13g2_fill_1 FILLER_23_1699 ();
 sg13g2_decap_8 FILLER_23_1730 ();
 sg13g2_fill_2 FILLER_23_1737 ();
 sg13g2_fill_1 FILLER_23_1739 ();
 sg13g2_fill_1 FILLER_23_1749 ();
 sg13g2_fill_2 FILLER_23_1755 ();
 sg13g2_fill_1 FILLER_23_1788 ();
 sg13g2_fill_1 FILLER_23_1802 ();
 sg13g2_fill_1 FILLER_23_1847 ();
 sg13g2_fill_2 FILLER_23_1871 ();
 sg13g2_fill_1 FILLER_23_1873 ();
 sg13g2_fill_1 FILLER_23_1916 ();
 sg13g2_fill_2 FILLER_23_1929 ();
 sg13g2_fill_1 FILLER_23_1931 ();
 sg13g2_fill_1 FILLER_23_1968 ();
 sg13g2_decap_4 FILLER_23_1995 ();
 sg13g2_fill_2 FILLER_23_1999 ();
 sg13g2_fill_1 FILLER_23_2098 ();
 sg13g2_fill_2 FILLER_23_2105 ();
 sg13g2_fill_1 FILLER_23_2107 ();
 sg13g2_fill_1 FILLER_23_2120 ();
 sg13g2_fill_2 FILLER_23_2138 ();
 sg13g2_fill_2 FILLER_23_2161 ();
 sg13g2_fill_1 FILLER_23_2181 ();
 sg13g2_fill_1 FILLER_23_2288 ();
 sg13g2_fill_1 FILLER_23_2302 ();
 sg13g2_fill_2 FILLER_23_2317 ();
 sg13g2_fill_1 FILLER_23_2358 ();
 sg13g2_fill_1 FILLER_23_2390 ();
 sg13g2_fill_2 FILLER_23_2452 ();
 sg13g2_fill_1 FILLER_23_2454 ();
 sg13g2_fill_2 FILLER_23_2507 ();
 sg13g2_fill_1 FILLER_23_2509 ();
 sg13g2_decap_8 FILLER_23_2579 ();
 sg13g2_fill_2 FILLER_23_2586 ();
 sg13g2_fill_1 FILLER_23_2628 ();
 sg13g2_fill_2 FILLER_23_2642 ();
 sg13g2_fill_1 FILLER_23_2644 ();
 sg13g2_fill_1 FILLER_23_2673 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_419 ();
 sg13g2_fill_2 FILLER_24_487 ();
 sg13g2_fill_1 FILLER_24_581 ();
 sg13g2_fill_1 FILLER_24_610 ();
 sg13g2_fill_1 FILLER_24_704 ();
 sg13g2_fill_2 FILLER_24_790 ();
 sg13g2_fill_1 FILLER_24_792 ();
 sg13g2_fill_2 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_834 ();
 sg13g2_fill_2 FILLER_24_862 ();
 sg13g2_fill_2 FILLER_24_977 ();
 sg13g2_fill_1 FILLER_24_979 ();
 sg13g2_fill_1 FILLER_24_998 ();
 sg13g2_fill_1 FILLER_24_1071 ();
 sg13g2_fill_1 FILLER_24_1178 ();
 sg13g2_fill_1 FILLER_24_1197 ();
 sg13g2_fill_2 FILLER_24_1226 ();
 sg13g2_decap_8 FILLER_24_1327 ();
 sg13g2_fill_2 FILLER_24_1338 ();
 sg13g2_fill_2 FILLER_24_1350 ();
 sg13g2_fill_2 FILLER_24_1373 ();
 sg13g2_fill_1 FILLER_24_1375 ();
 sg13g2_decap_8 FILLER_24_1393 ();
 sg13g2_fill_2 FILLER_24_1414 ();
 sg13g2_fill_2 FILLER_24_1425 ();
 sg13g2_fill_1 FILLER_24_1427 ();
 sg13g2_fill_2 FILLER_24_1446 ();
 sg13g2_fill_2 FILLER_24_1582 ();
 sg13g2_fill_1 FILLER_24_1584 ();
 sg13g2_fill_2 FILLER_24_1596 ();
 sg13g2_fill_2 FILLER_24_1612 ();
 sg13g2_decap_8 FILLER_24_1622 ();
 sg13g2_decap_8 FILLER_24_1629 ();
 sg13g2_fill_1 FILLER_24_1636 ();
 sg13g2_decap_8 FILLER_24_1688 ();
 sg13g2_fill_2 FILLER_24_1695 ();
 sg13g2_fill_2 FILLER_24_1702 ();
 sg13g2_decap_8 FILLER_24_1711 ();
 sg13g2_fill_2 FILLER_24_1718 ();
 sg13g2_fill_2 FILLER_24_1742 ();
 sg13g2_fill_1 FILLER_24_1744 ();
 sg13g2_fill_1 FILLER_24_1772 ();
 sg13g2_fill_1 FILLER_24_1808 ();
 sg13g2_fill_1 FILLER_24_1836 ();
 sg13g2_fill_2 FILLER_24_1882 ();
 sg13g2_fill_1 FILLER_24_1884 ();
 sg13g2_fill_1 FILLER_24_1903 ();
 sg13g2_fill_2 FILLER_24_1916 ();
 sg13g2_fill_2 FILLER_24_1930 ();
 sg13g2_fill_2 FILLER_24_1978 ();
 sg13g2_decap_4 FILLER_24_1989 ();
 sg13g2_decap_4 FILLER_24_2002 ();
 sg13g2_fill_1 FILLER_24_2006 ();
 sg13g2_fill_2 FILLER_24_2018 ();
 sg13g2_decap_8 FILLER_24_2047 ();
 sg13g2_fill_1 FILLER_24_2108 ();
 sg13g2_fill_2 FILLER_24_2235 ();
 sg13g2_fill_2 FILLER_24_2242 ();
 sg13g2_fill_1 FILLER_24_2244 ();
 sg13g2_fill_1 FILLER_24_2311 ();
 sg13g2_fill_1 FILLER_24_2338 ();
 sg13g2_fill_2 FILLER_24_2352 ();
 sg13g2_fill_1 FILLER_24_2354 ();
 sg13g2_fill_2 FILLER_24_2386 ();
 sg13g2_fill_1 FILLER_24_2388 ();
 sg13g2_fill_2 FILLER_24_2460 ();
 sg13g2_fill_1 FILLER_24_2475 ();
 sg13g2_fill_1 FILLER_24_2514 ();
 sg13g2_decap_8 FILLER_24_2571 ();
 sg13g2_fill_1 FILLER_24_2582 ();
 sg13g2_fill_1 FILLER_24_2587 ();
 sg13g2_fill_1 FILLER_24_2606 ();
 sg13g2_fill_1 FILLER_24_2616 ();
 sg13g2_fill_2 FILLER_24_2672 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_424 ();
 sg13g2_fill_1 FILLER_25_491 ();
 sg13g2_fill_2 FILLER_25_576 ();
 sg13g2_fill_1 FILLER_25_587 ();
 sg13g2_fill_2 FILLER_25_594 ();
 sg13g2_fill_1 FILLER_25_596 ();
 sg13g2_fill_1 FILLER_25_686 ();
 sg13g2_fill_2 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_fill_2 FILLER_25_717 ();
 sg13g2_fill_1 FILLER_25_719 ();
 sg13g2_fill_2 FILLER_25_782 ();
 sg13g2_fill_1 FILLER_25_784 ();
 sg13g2_fill_2 FILLER_25_825 ();
 sg13g2_fill_1 FILLER_25_837 ();
 sg13g2_fill_2 FILLER_25_844 ();
 sg13g2_fill_1 FILLER_25_846 ();
 sg13g2_fill_2 FILLER_25_1001 ();
 sg13g2_fill_1 FILLER_25_1026 ();
 sg13g2_fill_2 FILLER_25_1046 ();
 sg13g2_fill_2 FILLER_25_1063 ();
 sg13g2_decap_4 FILLER_25_1088 ();
 sg13g2_fill_2 FILLER_25_1092 ();
 sg13g2_fill_1 FILLER_25_1103 ();
 sg13g2_fill_2 FILLER_25_1107 ();
 sg13g2_fill_1 FILLER_25_1117 ();
 sg13g2_fill_2 FILLER_25_1128 ();
 sg13g2_fill_1 FILLER_25_1130 ();
 sg13g2_fill_2 FILLER_25_1163 ();
 sg13g2_fill_1 FILLER_25_1182 ();
 sg13g2_fill_1 FILLER_25_1344 ();
 sg13g2_decap_8 FILLER_25_1369 ();
 sg13g2_fill_1 FILLER_25_1376 ();
 sg13g2_fill_2 FILLER_25_1384 ();
 sg13g2_decap_8 FILLER_25_1395 ();
 sg13g2_fill_2 FILLER_25_1434 ();
 sg13g2_decap_8 FILLER_25_1442 ();
 sg13g2_decap_4 FILLER_25_1449 ();
 sg13g2_fill_1 FILLER_25_1453 ();
 sg13g2_fill_2 FILLER_25_1501 ();
 sg13g2_fill_2 FILLER_25_1574 ();
 sg13g2_fill_1 FILLER_25_1604 ();
 sg13g2_fill_1 FILLER_25_1615 ();
 sg13g2_fill_1 FILLER_25_1631 ();
 sg13g2_fill_2 FILLER_25_1645 ();
 sg13g2_fill_1 FILLER_25_1647 ();
 sg13g2_fill_1 FILLER_25_1661 ();
 sg13g2_decap_4 FILLER_25_1688 ();
 sg13g2_fill_2 FILLER_25_1692 ();
 sg13g2_decap_4 FILLER_25_1710 ();
 sg13g2_fill_2 FILLER_25_1714 ();
 sg13g2_fill_1 FILLER_25_1785 ();
 sg13g2_decap_8 FILLER_25_1790 ();
 sg13g2_decap_8 FILLER_25_1797 ();
 sg13g2_fill_1 FILLER_25_1841 ();
 sg13g2_fill_1 FILLER_25_1910 ();
 sg13g2_fill_2 FILLER_25_1916 ();
 sg13g2_fill_2 FILLER_25_1958 ();
 sg13g2_decap_8 FILLER_25_2001 ();
 sg13g2_decap_4 FILLER_25_2008 ();
 sg13g2_fill_1 FILLER_25_2012 ();
 sg13g2_fill_2 FILLER_25_2040 ();
 sg13g2_fill_1 FILLER_25_2042 ();
 sg13g2_decap_8 FILLER_25_2052 ();
 sg13g2_fill_2 FILLER_25_2059 ();
 sg13g2_fill_1 FILLER_25_2061 ();
 sg13g2_fill_2 FILLER_25_2072 ();
 sg13g2_fill_2 FILLER_25_2121 ();
 sg13g2_fill_2 FILLER_25_2202 ();
 sg13g2_fill_2 FILLER_25_2257 ();
 sg13g2_fill_1 FILLER_25_2259 ();
 sg13g2_fill_2 FILLER_25_2279 ();
 sg13g2_fill_1 FILLER_25_2281 ();
 sg13g2_fill_2 FILLER_25_2294 ();
 sg13g2_fill_1 FILLER_25_2296 ();
 sg13g2_fill_2 FILLER_25_2341 ();
 sg13g2_fill_1 FILLER_25_2366 ();
 sg13g2_fill_1 FILLER_25_2380 ();
 sg13g2_fill_1 FILLER_25_2417 ();
 sg13g2_fill_2 FILLER_25_2422 ();
 sg13g2_fill_1 FILLER_25_2424 ();
 sg13g2_fill_2 FILLER_25_2470 ();
 sg13g2_fill_1 FILLER_25_2472 ();
 sg13g2_decap_4 FILLER_25_2515 ();
 sg13g2_decap_8 FILLER_25_2528 ();
 sg13g2_decap_8 FILLER_25_2535 ();
 sg13g2_fill_1 FILLER_25_2542 ();
 sg13g2_decap_4 FILLER_25_2565 ();
 sg13g2_fill_1 FILLER_25_2569 ();
 sg13g2_fill_2 FILLER_25_2588 ();
 sg13g2_fill_1 FILLER_25_2590 ();
 sg13g2_fill_2 FILLER_25_2638 ();
 sg13g2_fill_1 FILLER_25_2640 ();
 sg13g2_fill_2 FILLER_25_2672 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_47 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_61 ();
 sg13g2_fill_2 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_576 ();
 sg13g2_fill_1 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_653 ();
 sg13g2_fill_1 FILLER_26_655 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_fill_2 FILLER_26_686 ();
 sg13g2_fill_1 FILLER_26_688 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_fill_1 FILLER_26_724 ();
 sg13g2_fill_1 FILLER_26_789 ();
 sg13g2_fill_2 FILLER_26_803 ();
 sg13g2_fill_1 FILLER_26_805 ();
 sg13g2_fill_2 FILLER_26_839 ();
 sg13g2_fill_2 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_856 ();
 sg13g2_fill_1 FILLER_26_929 ();
 sg13g2_fill_2 FILLER_26_966 ();
 sg13g2_fill_1 FILLER_26_968 ();
 sg13g2_fill_1 FILLER_26_1006 ();
 sg13g2_fill_2 FILLER_26_1035 ();
 sg13g2_fill_1 FILLER_26_1037 ();
 sg13g2_fill_1 FILLER_26_1043 ();
 sg13g2_fill_1 FILLER_26_1062 ();
 sg13g2_decap_8 FILLER_26_1073 ();
 sg13g2_decap_8 FILLER_26_1096 ();
 sg13g2_fill_2 FILLER_26_1103 ();
 sg13g2_fill_2 FILLER_26_1114 ();
 sg13g2_fill_1 FILLER_26_1116 ();
 sg13g2_fill_2 FILLER_26_1130 ();
 sg13g2_fill_2 FILLER_26_1208 ();
 sg13g2_fill_2 FILLER_26_1220 ();
 sg13g2_fill_1 FILLER_26_1254 ();
 sg13g2_fill_2 FILLER_26_1290 ();
 sg13g2_decap_4 FILLER_26_1329 ();
 sg13g2_fill_2 FILLER_26_1333 ();
 sg13g2_fill_2 FILLER_26_1368 ();
 sg13g2_fill_1 FILLER_26_1370 ();
 sg13g2_decap_8 FILLER_26_1445 ();
 sg13g2_decap_8 FILLER_26_1452 ();
 sg13g2_decap_8 FILLER_26_1459 ();
 sg13g2_fill_2 FILLER_26_1498 ();
 sg13g2_fill_2 FILLER_26_1513 ();
 sg13g2_decap_4 FILLER_26_1528 ();
 sg13g2_decap_8 FILLER_26_1573 ();
 sg13g2_decap_8 FILLER_26_1580 ();
 sg13g2_decap_8 FILLER_26_1587 ();
 sg13g2_decap_4 FILLER_26_1594 ();
 sg13g2_fill_2 FILLER_26_1626 ();
 sg13g2_fill_2 FILLER_26_1633 ();
 sg13g2_fill_1 FILLER_26_1635 ();
 sg13g2_fill_1 FILLER_26_1644 ();
 sg13g2_fill_2 FILLER_26_1650 ();
 sg13g2_fill_2 FILLER_26_1657 ();
 sg13g2_decap_8 FILLER_26_1694 ();
 sg13g2_fill_2 FILLER_26_1733 ();
 sg13g2_fill_2 FILLER_26_1787 ();
 sg13g2_fill_1 FILLER_26_1789 ();
 sg13g2_decap_8 FILLER_26_1795 ();
 sg13g2_fill_2 FILLER_26_1899 ();
 sg13g2_fill_1 FILLER_26_1901 ();
 sg13g2_fill_2 FILLER_26_1913 ();
 sg13g2_fill_1 FILLER_26_1915 ();
 sg13g2_decap_8 FILLER_26_1969 ();
 sg13g2_decap_8 FILLER_26_1976 ();
 sg13g2_decap_8 FILLER_26_1983 ();
 sg13g2_decap_8 FILLER_26_1990 ();
 sg13g2_decap_4 FILLER_26_1997 ();
 sg13g2_fill_1 FILLER_26_2001 ();
 sg13g2_decap_4 FILLER_26_2029 ();
 sg13g2_fill_2 FILLER_26_2050 ();
 sg13g2_fill_1 FILLER_26_2052 ();
 sg13g2_fill_1 FILLER_26_2163 ();
 sg13g2_fill_1 FILLER_26_2227 ();
 sg13g2_fill_2 FILLER_26_2273 ();
 sg13g2_fill_2 FILLER_26_2387 ();
 sg13g2_fill_2 FILLER_26_2416 ();
 sg13g2_fill_2 FILLER_26_2454 ();
 sg13g2_fill_1 FILLER_26_2456 ();
 sg13g2_fill_1 FILLER_26_2465 ();
 sg13g2_fill_2 FILLER_26_2490 ();
 sg13g2_decap_8 FILLER_26_2522 ();
 sg13g2_fill_2 FILLER_26_2569 ();
 sg13g2_fill_2 FILLER_26_2626 ();
 sg13g2_fill_1 FILLER_26_2643 ();
 sg13g2_fill_2 FILLER_26_2672 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_430 ();
 sg13g2_fill_2 FILLER_27_559 ();
 sg13g2_fill_2 FILLER_27_576 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_fill_1 FILLER_27_704 ();
 sg13g2_fill_2 FILLER_27_713 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_fill_2 FILLER_27_754 ();
 sg13g2_fill_1 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_792 ();
 sg13g2_fill_2 FILLER_27_820 ();
 sg13g2_fill_1 FILLER_27_822 ();
 sg13g2_fill_1 FILLER_27_857 ();
 sg13g2_fill_2 FILLER_27_884 ();
 sg13g2_fill_2 FILLER_27_929 ();
 sg13g2_fill_1 FILLER_27_931 ();
 sg13g2_fill_2 FILLER_27_950 ();
 sg13g2_fill_2 FILLER_27_1045 ();
 sg13g2_decap_4 FILLER_27_1059 ();
 sg13g2_fill_2 FILLER_27_1063 ();
 sg13g2_fill_2 FILLER_27_1070 ();
 sg13g2_fill_1 FILLER_27_1131 ();
 sg13g2_fill_1 FILLER_27_1137 ();
 sg13g2_fill_1 FILLER_27_1170 ();
 sg13g2_decap_8 FILLER_27_1320 ();
 sg13g2_decap_4 FILLER_27_1327 ();
 sg13g2_fill_1 FILLER_27_1331 ();
 sg13g2_decap_4 FILLER_27_1366 ();
 sg13g2_fill_2 FILLER_27_1388 ();
 sg13g2_fill_1 FILLER_27_1390 ();
 sg13g2_fill_2 FILLER_27_1397 ();
 sg13g2_fill_1 FILLER_27_1425 ();
 sg13g2_decap_8 FILLER_27_1448 ();
 sg13g2_decap_8 FILLER_27_1455 ();
 sg13g2_decap_4 FILLER_27_1462 ();
 sg13g2_fill_2 FILLER_27_1489 ();
 sg13g2_fill_1 FILLER_27_1491 ();
 sg13g2_fill_1 FILLER_27_1510 ();
 sg13g2_fill_1 FILLER_27_1527 ();
 sg13g2_decap_4 FILLER_27_1533 ();
 sg13g2_decap_8 FILLER_27_1566 ();
 sg13g2_fill_2 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1584 ();
 sg13g2_decap_8 FILLER_27_1591 ();
 sg13g2_fill_2 FILLER_27_1647 ();
 sg13g2_fill_1 FILLER_27_1649 ();
 sg13g2_decap_8 FILLER_27_1685 ();
 sg13g2_decap_8 FILLER_27_1692 ();
 sg13g2_fill_1 FILLER_27_1699 ();
 sg13g2_decap_8 FILLER_27_1713 ();
 sg13g2_decap_4 FILLER_27_1720 ();
 sg13g2_fill_1 FILLER_27_1737 ();
 sg13g2_fill_2 FILLER_27_1770 ();
 sg13g2_fill_1 FILLER_27_1772 ();
 sg13g2_fill_2 FILLER_27_1809 ();
 sg13g2_fill_1 FILLER_27_1811 ();
 sg13g2_fill_2 FILLER_27_1839 ();
 sg13g2_decap_8 FILLER_27_1850 ();
 sg13g2_fill_2 FILLER_27_1897 ();
 sg13g2_fill_1 FILLER_27_1899 ();
 sg13g2_fill_1 FILLER_27_1973 ();
 sg13g2_fill_2 FILLER_27_1979 ();
 sg13g2_fill_1 FILLER_27_1981 ();
 sg13g2_fill_2 FILLER_27_1986 ();
 sg13g2_fill_1 FILLER_27_1988 ();
 sg13g2_fill_1 FILLER_27_2008 ();
 sg13g2_decap_8 FILLER_27_2045 ();
 sg13g2_decap_4 FILLER_27_2052 ();
 sg13g2_fill_2 FILLER_27_2056 ();
 sg13g2_fill_1 FILLER_27_2130 ();
 sg13g2_fill_1 FILLER_27_2190 ();
 sg13g2_fill_2 FILLER_27_2226 ();
 sg13g2_fill_1 FILLER_27_2228 ();
 sg13g2_fill_2 FILLER_27_2325 ();
 sg13g2_fill_2 FILLER_27_2369 ();
 sg13g2_fill_1 FILLER_27_2371 ();
 sg13g2_fill_2 FILLER_27_2403 ();
 sg13g2_fill_2 FILLER_27_2432 ();
 sg13g2_fill_1 FILLER_27_2434 ();
 sg13g2_fill_2 FILLER_27_2450 ();
 sg13g2_fill_1 FILLER_27_2452 ();
 sg13g2_fill_2 FILLER_27_2462 ();
 sg13g2_fill_1 FILLER_27_2464 ();
 sg13g2_fill_2 FILLER_27_2483 ();
 sg13g2_fill_2 FILLER_27_2536 ();
 sg13g2_fill_1 FILLER_27_2544 ();
 sg13g2_fill_2 FILLER_27_2576 ();
 sg13g2_fill_2 FILLER_27_2619 ();
 sg13g2_fill_2 FILLER_27_2671 ();
 sg13g2_fill_1 FILLER_27_2673 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_512 ();
 sg13g2_fill_1 FILLER_28_629 ();
 sg13g2_fill_1 FILLER_28_658 ();
 sg13g2_decap_4 FILLER_28_695 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_4 FILLER_28_732 ();
 sg13g2_fill_1 FILLER_28_736 ();
 sg13g2_fill_2 FILLER_28_741 ();
 sg13g2_fill_1 FILLER_28_743 ();
 sg13g2_fill_2 FILLER_28_774 ();
 sg13g2_fill_1 FILLER_28_776 ();
 sg13g2_fill_2 FILLER_28_794 ();
 sg13g2_fill_1 FILLER_28_796 ();
 sg13g2_fill_2 FILLER_28_801 ();
 sg13g2_fill_2 FILLER_28_810 ();
 sg13g2_fill_1 FILLER_28_812 ();
 sg13g2_fill_1 FILLER_28_928 ();
 sg13g2_fill_2 FILLER_28_950 ();
 sg13g2_fill_1 FILLER_28_952 ();
 sg13g2_fill_2 FILLER_28_998 ();
 sg13g2_fill_1 FILLER_28_1000 ();
 sg13g2_fill_2 FILLER_28_1014 ();
 sg13g2_fill_1 FILLER_28_1016 ();
 sg13g2_fill_2 FILLER_28_1022 ();
 sg13g2_fill_2 FILLER_28_1029 ();
 sg13g2_fill_1 FILLER_28_1031 ();
 sg13g2_fill_1 FILLER_28_1045 ();
 sg13g2_fill_1 FILLER_28_1101 ();
 sg13g2_fill_2 FILLER_28_1161 ();
 sg13g2_fill_2 FILLER_28_1182 ();
 sg13g2_fill_2 FILLER_28_1221 ();
 sg13g2_fill_2 FILLER_28_1291 ();
 sg13g2_decap_8 FILLER_28_1330 ();
 sg13g2_decap_4 FILLER_28_1337 ();
 sg13g2_fill_2 FILLER_28_1341 ();
 sg13g2_decap_4 FILLER_28_1367 ();
 sg13g2_fill_1 FILLER_28_1381 ();
 sg13g2_fill_1 FILLER_28_1396 ();
 sg13g2_fill_1 FILLER_28_1419 ();
 sg13g2_decap_4 FILLER_28_1461 ();
 sg13g2_fill_1 FILLER_28_1465 ();
 sg13g2_fill_2 FILLER_28_1511 ();
 sg13g2_decap_4 FILLER_28_1568 ();
 sg13g2_decap_8 FILLER_28_1585 ();
 sg13g2_decap_4 FILLER_28_1592 ();
 sg13g2_fill_2 FILLER_28_1596 ();
 sg13g2_fill_2 FILLER_28_1617 ();
 sg13g2_fill_1 FILLER_28_1619 ();
 sg13g2_decap_4 FILLER_28_1634 ();
 sg13g2_fill_1 FILLER_28_1638 ();
 sg13g2_fill_1 FILLER_28_1652 ();
 sg13g2_decap_4 FILLER_28_1666 ();
 sg13g2_fill_2 FILLER_28_1684 ();
 sg13g2_decap_4 FILLER_28_1691 ();
 sg13g2_fill_2 FILLER_28_1699 ();
 sg13g2_fill_1 FILLER_28_1701 ();
 sg13g2_fill_2 FILLER_28_1706 ();
 sg13g2_fill_1 FILLER_28_1713 ();
 sg13g2_fill_2 FILLER_28_1718 ();
 sg13g2_fill_1 FILLER_28_1720 ();
 sg13g2_fill_2 FILLER_28_1725 ();
 sg13g2_fill_1 FILLER_28_1727 ();
 sg13g2_fill_2 FILLER_28_1736 ();
 sg13g2_fill_2 FILLER_28_1751 ();
 sg13g2_decap_8 FILLER_28_1814 ();
 sg13g2_fill_1 FILLER_28_1821 ();
 sg13g2_fill_1 FILLER_28_1832 ();
 sg13g2_fill_2 FILLER_28_1837 ();
 sg13g2_decap_4 FILLER_28_1848 ();
 sg13g2_fill_2 FILLER_28_1852 ();
 sg13g2_fill_2 FILLER_28_1885 ();
 sg13g2_fill_1 FILLER_28_1887 ();
 sg13g2_fill_2 FILLER_28_1915 ();
 sg13g2_fill_1 FILLER_28_1917 ();
 sg13g2_fill_2 FILLER_28_1954 ();
 sg13g2_fill_1 FILLER_28_1956 ();
 sg13g2_decap_4 FILLER_28_2024 ();
 sg13g2_fill_2 FILLER_28_2055 ();
 sg13g2_fill_1 FILLER_28_2057 ();
 sg13g2_fill_1 FILLER_28_2101 ();
 sg13g2_fill_1 FILLER_28_2126 ();
 sg13g2_fill_2 FILLER_28_2240 ();
 sg13g2_fill_1 FILLER_28_2269 ();
 sg13g2_fill_1 FILLER_28_2330 ();
 sg13g2_fill_2 FILLER_28_2362 ();
 sg13g2_fill_1 FILLER_28_2364 ();
 sg13g2_fill_2 FILLER_28_2371 ();
 sg13g2_fill_2 FILLER_28_2395 ();
 sg13g2_fill_2 FILLER_28_2463 ();
 sg13g2_fill_2 FILLER_28_2471 ();
 sg13g2_fill_2 FILLER_28_2488 ();
 sg13g2_fill_2 FILLER_28_2627 ();
 sg13g2_fill_1 FILLER_28_2629 ();
 sg13g2_fill_2 FILLER_28_2671 ();
 sg13g2_fill_1 FILLER_28_2673 ();
 sg13g2_fill_1 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_decap_4 FILLER_29_417 ();
 sg13g2_fill_1 FILLER_29_479 ();
 sg13g2_fill_2 FILLER_29_511 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_fill_2 FILLER_29_573 ();
 sg13g2_fill_1 FILLER_29_575 ();
 sg13g2_fill_1 FILLER_29_686 ();
 sg13g2_fill_2 FILLER_29_692 ();
 sg13g2_fill_1 FILLER_29_694 ();
 sg13g2_decap_8 FILLER_29_705 ();
 sg13g2_decap_8 FILLER_29_712 ();
 sg13g2_decap_8 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_decap_8 FILLER_29_733 ();
 sg13g2_decap_8 FILLER_29_740 ();
 sg13g2_decap_4 FILLER_29_747 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_fill_2 FILLER_29_825 ();
 sg13g2_fill_1 FILLER_29_827 ();
 sg13g2_fill_2 FILLER_29_914 ();
 sg13g2_fill_1 FILLER_29_916 ();
 sg13g2_fill_2 FILLER_29_937 ();
 sg13g2_fill_1 FILLER_29_962 ();
 sg13g2_fill_1 FILLER_29_968 ();
 sg13g2_fill_1 FILLER_29_1021 ();
 sg13g2_fill_2 FILLER_29_1045 ();
 sg13g2_decap_8 FILLER_29_1102 ();
 sg13g2_fill_2 FILLER_29_1109 ();
 sg13g2_fill_1 FILLER_29_1139 ();
 sg13g2_fill_1 FILLER_29_1283 ();
 sg13g2_fill_2 FILLER_29_1293 ();
 sg13g2_fill_1 FILLER_29_1311 ();
 sg13g2_fill_2 FILLER_29_1396 ();
 sg13g2_fill_1 FILLER_29_1398 ();
 sg13g2_fill_2 FILLER_29_1405 ();
 sg13g2_fill_1 FILLER_29_1446 ();
 sg13g2_decap_4 FILLER_29_1505 ();
 sg13g2_decap_8 FILLER_29_1537 ();
 sg13g2_decap_8 FILLER_29_1544 ();
 sg13g2_decap_8 FILLER_29_1551 ();
 sg13g2_fill_2 FILLER_29_1558 ();
 sg13g2_fill_1 FILLER_29_1569 ();
 sg13g2_fill_2 FILLER_29_1577 ();
 sg13g2_fill_1 FILLER_29_1579 ();
 sg13g2_decap_4 FILLER_29_1593 ();
 sg13g2_fill_1 FILLER_29_1597 ();
 sg13g2_fill_2 FILLER_29_1640 ();
 sg13g2_fill_1 FILLER_29_1647 ();
 sg13g2_fill_2 FILLER_29_1653 ();
 sg13g2_decap_8 FILLER_29_1659 ();
 sg13g2_fill_2 FILLER_29_1692 ();
 sg13g2_fill_1 FILLER_29_1694 ();
 sg13g2_fill_1 FILLER_29_1708 ();
 sg13g2_decap_8 FILLER_29_1724 ();
 sg13g2_decap_4 FILLER_29_1731 ();
 sg13g2_decap_8 FILLER_29_1753 ();
 sg13g2_fill_1 FILLER_29_1760 ();
 sg13g2_decap_4 FILLER_29_1846 ();
 sg13g2_fill_1 FILLER_29_1877 ();
 sg13g2_fill_1 FILLER_29_1897 ();
 sg13g2_fill_2 FILLER_29_1955 ();
 sg13g2_fill_1 FILLER_29_1957 ();
 sg13g2_fill_1 FILLER_29_1971 ();
 sg13g2_decap_8 FILLER_29_1999 ();
 sg13g2_fill_2 FILLER_29_2047 ();
 sg13g2_fill_2 FILLER_29_2110 ();
 sg13g2_fill_1 FILLER_29_2112 ();
 sg13g2_fill_1 FILLER_29_2242 ();
 sg13g2_fill_2 FILLER_29_2270 ();
 sg13g2_fill_1 FILLER_29_2272 ();
 sg13g2_decap_4 FILLER_29_2324 ();
 sg13g2_fill_2 FILLER_29_2380 ();
 sg13g2_fill_2 FILLER_29_2415 ();
 sg13g2_fill_1 FILLER_29_2417 ();
 sg13g2_fill_2 FILLER_29_2453 ();
 sg13g2_fill_1 FILLER_29_2482 ();
 sg13g2_fill_1 FILLER_29_2495 ();
 sg13g2_fill_2 FILLER_29_2616 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_decap_4 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_decap_4 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_285 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_fill_2 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_fill_1 FILLER_30_430 ();
 sg13g2_fill_1 FILLER_30_522 ();
 sg13g2_fill_2 FILLER_30_544 ();
 sg13g2_fill_1 FILLER_30_624 ();
 sg13g2_decap_4 FILLER_30_635 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_fill_1 FILLER_30_668 ();
 sg13g2_fill_2 FILLER_30_682 ();
 sg13g2_fill_1 FILLER_30_684 ();
 sg13g2_decap_8 FILLER_30_696 ();
 sg13g2_decap_8 FILLER_30_703 ();
 sg13g2_decap_8 FILLER_30_710 ();
 sg13g2_decap_4 FILLER_30_717 ();
 sg13g2_fill_2 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_748 ();
 sg13g2_decap_8 FILLER_30_755 ();
 sg13g2_fill_1 FILLER_30_784 ();
 sg13g2_fill_2 FILLER_30_794 ();
 sg13g2_fill_1 FILLER_30_805 ();
 sg13g2_fill_1 FILLER_30_879 ();
 sg13g2_fill_2 FILLER_30_930 ();
 sg13g2_fill_2 FILLER_30_942 ();
 sg13g2_fill_1 FILLER_30_951 ();
 sg13g2_fill_2 FILLER_30_965 ();
 sg13g2_fill_1 FILLER_30_967 ();
 sg13g2_fill_2 FILLER_30_1010 ();
 sg13g2_fill_1 FILLER_30_1012 ();
 sg13g2_fill_1 FILLER_30_1060 ();
 sg13g2_decap_8 FILLER_30_1096 ();
 sg13g2_decap_8 FILLER_30_1103 ();
 sg13g2_fill_2 FILLER_30_1145 ();
 sg13g2_fill_1 FILLER_30_1262 ();
 sg13g2_decap_8 FILLER_30_1349 ();
 sg13g2_decap_8 FILLER_30_1356 ();
 sg13g2_decap_8 FILLER_30_1363 ();
 sg13g2_decap_8 FILLER_30_1370 ();
 sg13g2_fill_1 FILLER_30_1377 ();
 sg13g2_fill_2 FILLER_30_1415 ();
 sg13g2_fill_1 FILLER_30_1417 ();
 sg13g2_fill_1 FILLER_30_1495 ();
 sg13g2_decap_4 FILLER_30_1535 ();
 sg13g2_fill_1 FILLER_30_1539 ();
 sg13g2_fill_1 FILLER_30_1544 ();
 sg13g2_fill_2 FILLER_30_1571 ();
 sg13g2_fill_1 FILLER_30_1594 ();
 sg13g2_fill_1 FILLER_30_1609 ();
 sg13g2_fill_2 FILLER_30_1627 ();
 sg13g2_decap_8 FILLER_30_1640 ();
 sg13g2_decap_8 FILLER_30_1647 ();
 sg13g2_decap_8 FILLER_30_1654 ();
 sg13g2_decap_8 FILLER_30_1661 ();
 sg13g2_fill_2 FILLER_30_1689 ();
 sg13g2_fill_2 FILLER_30_1722 ();
 sg13g2_fill_1 FILLER_30_1724 ();
 sg13g2_decap_8 FILLER_30_1733 ();
 sg13g2_fill_2 FILLER_30_1740 ();
 sg13g2_fill_1 FILLER_30_1742 ();
 sg13g2_fill_2 FILLER_30_1789 ();
 sg13g2_fill_1 FILLER_30_1791 ();
 sg13g2_fill_1 FILLER_30_1851 ();
 sg13g2_fill_2 FILLER_30_1916 ();
 sg13g2_fill_1 FILLER_30_1918 ();
 sg13g2_fill_1 FILLER_30_1941 ();
 sg13g2_fill_1 FILLER_30_1968 ();
 sg13g2_fill_1 FILLER_30_2001 ();
 sg13g2_fill_2 FILLER_30_2023 ();
 sg13g2_fill_1 FILLER_30_2025 ();
 sg13g2_fill_1 FILLER_30_2143 ();
 sg13g2_fill_1 FILLER_30_2171 ();
 sg13g2_fill_2 FILLER_30_2207 ();
 sg13g2_fill_1 FILLER_30_2209 ();
 sg13g2_fill_1 FILLER_30_2250 ();
 sg13g2_fill_2 FILLER_30_2260 ();
 sg13g2_fill_1 FILLER_30_2276 ();
 sg13g2_fill_2 FILLER_30_2283 ();
 sg13g2_decap_4 FILLER_30_2324 ();
 sg13g2_fill_2 FILLER_30_2328 ();
 sg13g2_fill_2 FILLER_30_2334 ();
 sg13g2_fill_1 FILLER_30_2336 ();
 sg13g2_fill_1 FILLER_30_2346 ();
 sg13g2_fill_2 FILLER_30_2397 ();
 sg13g2_fill_2 FILLER_30_2430 ();
 sg13g2_fill_1 FILLER_30_2432 ();
 sg13g2_fill_1 FILLER_30_2455 ();
 sg13g2_fill_1 FILLER_30_2461 ();
 sg13g2_fill_2 FILLER_30_2489 ();
 sg13g2_fill_1 FILLER_30_2491 ();
 sg13g2_fill_1 FILLER_30_2501 ();
 sg13g2_fill_1 FILLER_30_2568 ();
 sg13g2_fill_2 FILLER_30_2615 ();
 sg13g2_fill_1 FILLER_30_2645 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_20 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_decap_8 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_decap_4 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_1 FILLER_31_433 ();
 sg13g2_fill_1 FILLER_31_521 ();
 sg13g2_fill_2 FILLER_31_535 ();
 sg13g2_decap_4 FILLER_31_614 ();
 sg13g2_fill_1 FILLER_31_618 ();
 sg13g2_decap_8 FILLER_31_647 ();
 sg13g2_fill_2 FILLER_31_654 ();
 sg13g2_fill_2 FILLER_31_669 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_fill_2 FILLER_31_721 ();
 sg13g2_fill_1 FILLER_31_723 ();
 sg13g2_fill_2 FILLER_31_728 ();
 sg13g2_fill_1 FILLER_31_730 ();
 sg13g2_decap_8 FILLER_31_744 ();
 sg13g2_decap_8 FILLER_31_751 ();
 sg13g2_decap_8 FILLER_31_758 ();
 sg13g2_fill_2 FILLER_31_765 ();
 sg13g2_fill_1 FILLER_31_767 ();
 sg13g2_fill_1 FILLER_31_796 ();
 sg13g2_fill_2 FILLER_31_842 ();
 sg13g2_fill_2 FILLER_31_984 ();
 sg13g2_fill_1 FILLER_31_1078 ();
 sg13g2_fill_2 FILLER_31_1092 ();
 sg13g2_fill_1 FILLER_31_1094 ();
 sg13g2_fill_1 FILLER_31_1130 ();
 sg13g2_fill_2 FILLER_31_1180 ();
 sg13g2_fill_1 FILLER_31_1191 ();
 sg13g2_fill_2 FILLER_31_1211 ();
 sg13g2_fill_1 FILLER_31_1213 ();
 sg13g2_fill_1 FILLER_31_1269 ();
 sg13g2_fill_1 FILLER_31_1335 ();
 sg13g2_decap_8 FILLER_31_1368 ();
 sg13g2_decap_8 FILLER_31_1375 ();
 sg13g2_fill_1 FILLER_31_1441 ();
 sg13g2_fill_2 FILLER_31_1470 ();
 sg13g2_fill_1 FILLER_31_1472 ();
 sg13g2_fill_1 FILLER_31_1497 ();
 sg13g2_decap_8 FILLER_31_1507 ();
 sg13g2_decap_8 FILLER_31_1514 ();
 sg13g2_fill_1 FILLER_31_1521 ();
 sg13g2_decap_8 FILLER_31_1527 ();
 sg13g2_fill_1 FILLER_31_1534 ();
 sg13g2_fill_1 FILLER_31_1572 ();
 sg13g2_fill_2 FILLER_31_1577 ();
 sg13g2_fill_2 FILLER_31_1588 ();
 sg13g2_fill_1 FILLER_31_1590 ();
 sg13g2_decap_8 FILLER_31_1637 ();
 sg13g2_decap_4 FILLER_31_1644 ();
 sg13g2_fill_1 FILLER_31_1648 ();
 sg13g2_fill_1 FILLER_31_1655 ();
 sg13g2_fill_1 FILLER_31_1661 ();
 sg13g2_fill_1 FILLER_31_1667 ();
 sg13g2_fill_2 FILLER_31_1677 ();
 sg13g2_fill_1 FILLER_31_1717 ();
 sg13g2_decap_4 FILLER_31_1741 ();
 sg13g2_fill_2 FILLER_31_1745 ();
 sg13g2_fill_2 FILLER_31_1751 ();
 sg13g2_fill_1 FILLER_31_1794 ();
 sg13g2_fill_2 FILLER_31_1907 ();
 sg13g2_fill_1 FILLER_31_1909 ();
 sg13g2_fill_2 FILLER_31_1946 ();
 sg13g2_fill_1 FILLER_31_1965 ();
 sg13g2_fill_2 FILLER_31_1971 ();
 sg13g2_fill_1 FILLER_31_1973 ();
 sg13g2_fill_2 FILLER_31_1983 ();
 sg13g2_fill_1 FILLER_31_1993 ();
 sg13g2_fill_1 FILLER_31_2017 ();
 sg13g2_fill_1 FILLER_31_2046 ();
 sg13g2_fill_2 FILLER_31_2060 ();
 sg13g2_fill_2 FILLER_31_2089 ();
 sg13g2_fill_1 FILLER_31_2091 ();
 sg13g2_fill_1 FILLER_31_2155 ();
 sg13g2_fill_2 FILLER_31_2183 ();
 sg13g2_fill_2 FILLER_31_2236 ();
 sg13g2_fill_1 FILLER_31_2238 ();
 sg13g2_fill_2 FILLER_31_2271 ();
 sg13g2_fill_1 FILLER_31_2273 ();
 sg13g2_decap_8 FILLER_31_2313 ();
 sg13g2_fill_2 FILLER_31_2320 ();
 sg13g2_fill_1 FILLER_31_2322 ();
 sg13g2_fill_2 FILLER_31_2336 ();
 sg13g2_fill_1 FILLER_31_2338 ();
 sg13g2_fill_2 FILLER_31_2348 ();
 sg13g2_fill_1 FILLER_31_2350 ();
 sg13g2_fill_2 FILLER_31_2433 ();
 sg13g2_fill_2 FILLER_31_2440 ();
 sg13g2_fill_2 FILLER_31_2531 ();
 sg13g2_fill_1 FILLER_31_2607 ();
 sg13g2_fill_1 FILLER_31_2625 ();
 sg13g2_fill_2 FILLER_31_2635 ();
 sg13g2_fill_2 FILLER_31_2672 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_448 ();
 sg13g2_fill_1 FILLER_32_450 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_fill_2 FILLER_32_532 ();
 sg13g2_fill_1 FILLER_32_534 ();
 sg13g2_fill_1 FILLER_32_557 ();
 sg13g2_fill_2 FILLER_32_571 ();
 sg13g2_fill_1 FILLER_32_573 ();
 sg13g2_fill_2 FILLER_32_587 ();
 sg13g2_fill_2 FILLER_32_598 ();
 sg13g2_fill_2 FILLER_32_609 ();
 sg13g2_fill_1 FILLER_32_611 ();
 sg13g2_fill_2 FILLER_32_693 ();
 sg13g2_fill_1 FILLER_32_695 ();
 sg13g2_decap_8 FILLER_32_727 ();
 sg13g2_decap_8 FILLER_32_734 ();
 sg13g2_decap_4 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_751 ();
 sg13g2_decap_8 FILLER_32_758 ();
 sg13g2_fill_2 FILLER_32_765 ();
 sg13g2_fill_2 FILLER_32_812 ();
 sg13g2_fill_1 FILLER_32_814 ();
 sg13g2_fill_2 FILLER_32_834 ();
 sg13g2_fill_1 FILLER_32_918 ();
 sg13g2_fill_2 FILLER_32_948 ();
 sg13g2_fill_1 FILLER_32_1018 ();
 sg13g2_fill_1 FILLER_32_1037 ();
 sg13g2_fill_1 FILLER_32_1079 ();
 sg13g2_decap_4 FILLER_32_1089 ();
 sg13g2_fill_1 FILLER_32_1093 ();
 sg13g2_fill_2 FILLER_32_1130 ();
 sg13g2_fill_2 FILLER_32_1178 ();
 sg13g2_fill_1 FILLER_32_1228 ();
 sg13g2_fill_1 FILLER_32_1340 ();
 sg13g2_fill_1 FILLER_32_1358 ();
 sg13g2_fill_2 FILLER_32_1367 ();
 sg13g2_fill_1 FILLER_32_1369 ();
 sg13g2_fill_1 FILLER_32_1398 ();
 sg13g2_fill_2 FILLER_32_1425 ();
 sg13g2_fill_2 FILLER_32_1437 ();
 sg13g2_fill_1 FILLER_32_1439 ();
 sg13g2_fill_2 FILLER_32_1446 ();
 sg13g2_decap_4 FILLER_32_1495 ();
 sg13g2_fill_2 FILLER_32_1512 ();
 sg13g2_fill_2 FILLER_32_1520 ();
 sg13g2_fill_1 FILLER_32_1529 ();
 sg13g2_fill_1 FILLER_32_1535 ();
 sg13g2_fill_2 FILLER_32_1579 ();
 sg13g2_decap_8 FILLER_32_1627 ();
 sg13g2_decap_8 FILLER_32_1634 ();
 sg13g2_decap_4 FILLER_32_1641 ();
 sg13g2_fill_2 FILLER_32_1667 ();
 sg13g2_fill_1 FILLER_32_1669 ();
 sg13g2_fill_2 FILLER_32_1702 ();
 sg13g2_fill_1 FILLER_32_1716 ();
 sg13g2_decap_8 FILLER_32_1736 ();
 sg13g2_decap_4 FILLER_32_1743 ();
 sg13g2_decap_4 FILLER_32_1760 ();
 sg13g2_fill_1 FILLER_32_1764 ();
 sg13g2_fill_2 FILLER_32_1787 ();
 sg13g2_fill_1 FILLER_32_1811 ();
 sg13g2_fill_2 FILLER_32_1825 ();
 sg13g2_fill_1 FILLER_32_1842 ();
 sg13g2_fill_1 FILLER_32_1883 ();
 sg13g2_decap_4 FILLER_32_1953 ();
 sg13g2_fill_1 FILLER_32_2024 ();
 sg13g2_fill_2 FILLER_32_2069 ();
 sg13g2_fill_1 FILLER_32_2071 ();
 sg13g2_fill_2 FILLER_32_2126 ();
 sg13g2_fill_2 FILLER_32_2229 ();
 sg13g2_fill_1 FILLER_32_2231 ();
 sg13g2_fill_2 FILLER_32_2263 ();
 sg13g2_fill_1 FILLER_32_2265 ();
 sg13g2_decap_4 FILLER_32_2305 ();
 sg13g2_fill_2 FILLER_32_2309 ();
 sg13g2_fill_2 FILLER_32_2370 ();
 sg13g2_fill_2 FILLER_32_2465 ();
 sg13g2_fill_1 FILLER_32_2467 ();
 sg13g2_fill_1 FILLER_32_2473 ();
 sg13g2_fill_2 FILLER_32_2492 ();
 sg13g2_fill_1 FILLER_32_2568 ();
 sg13g2_fill_2 FILLER_32_2592 ();
 sg13g2_fill_2 FILLER_32_2624 ();
 sg13g2_fill_2 FILLER_32_2671 ();
 sg13g2_fill_1 FILLER_32_2673 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_366 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_fill_2 FILLER_33_450 ();
 sg13g2_fill_1 FILLER_33_452 ();
 sg13g2_fill_1 FILLER_33_506 ();
 sg13g2_fill_2 FILLER_33_515 ();
 sg13g2_fill_2 FILLER_33_529 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_fill_1 FILLER_33_548 ();
 sg13g2_fill_1 FILLER_33_594 ();
 sg13g2_fill_1 FILLER_33_604 ();
 sg13g2_fill_1 FILLER_33_642 ();
 sg13g2_decap_4 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_677 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_4 FILLER_33_690 ();
 sg13g2_fill_1 FILLER_33_710 ();
 sg13g2_decap_8 FILLER_33_719 ();
 sg13g2_fill_2 FILLER_33_726 ();
 sg13g2_fill_1 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_734 ();
 sg13g2_fill_2 FILLER_33_741 ();
 sg13g2_fill_1 FILLER_33_815 ();
 sg13g2_fill_1 FILLER_33_924 ();
 sg13g2_fill_1 FILLER_33_1053 ();
 sg13g2_fill_2 FILLER_33_1081 ();
 sg13g2_fill_1 FILLER_33_1083 ();
 sg13g2_fill_2 FILLER_33_1101 ();
 sg13g2_fill_2 FILLER_33_1154 ();
 sg13g2_fill_1 FILLER_33_1156 ();
 sg13g2_fill_2 FILLER_33_1167 ();
 sg13g2_fill_2 FILLER_33_1178 ();
 sg13g2_fill_2 FILLER_33_1238 ();
 sg13g2_fill_1 FILLER_33_1267 ();
 sg13g2_fill_2 FILLER_33_1322 ();
 sg13g2_fill_2 FILLER_33_1371 ();
 sg13g2_decap_4 FILLER_33_1395 ();
 sg13g2_fill_1 FILLER_33_1399 ();
 sg13g2_fill_1 FILLER_33_1424 ();
 sg13g2_fill_1 FILLER_33_1442 ();
 sg13g2_fill_2 FILLER_33_1452 ();
 sg13g2_fill_2 FILLER_33_1485 ();
 sg13g2_fill_1 FILLER_33_1524 ();
 sg13g2_fill_1 FILLER_33_1562 ();
 sg13g2_decap_8 FILLER_33_1580 ();
 sg13g2_decap_4 FILLER_33_1587 ();
 sg13g2_decap_8 FILLER_33_1620 ();
 sg13g2_decap_8 FILLER_33_1627 ();
 sg13g2_decap_8 FILLER_33_1634 ();
 sg13g2_fill_2 FILLER_33_1641 ();
 sg13g2_fill_1 FILLER_33_1643 ();
 sg13g2_decap_8 FILLER_33_1667 ();
 sg13g2_decap_4 FILLER_33_1674 ();
 sg13g2_decap_8 FILLER_33_1727 ();
 sg13g2_decap_8 FILLER_33_1734 ();
 sg13g2_decap_8 FILLER_33_1741 ();
 sg13g2_decap_4 FILLER_33_1748 ();
 sg13g2_fill_2 FILLER_33_1773 ();
 sg13g2_fill_2 FILLER_33_1823 ();
 sg13g2_fill_1 FILLER_33_1825 ();
 sg13g2_fill_2 FILLER_33_1888 ();
 sg13g2_decap_8 FILLER_33_1948 ();
 sg13g2_decap_4 FILLER_33_1955 ();
 sg13g2_fill_2 FILLER_33_1995 ();
 sg13g2_fill_2 FILLER_33_2003 ();
 sg13g2_fill_1 FILLER_33_2005 ();
 sg13g2_fill_1 FILLER_33_2012 ();
 sg13g2_fill_2 FILLER_33_2046 ();
 sg13g2_fill_1 FILLER_33_2048 ();
 sg13g2_fill_1 FILLER_33_2208 ();
 sg13g2_fill_2 FILLER_33_2306 ();
 sg13g2_fill_1 FILLER_33_2308 ();
 sg13g2_fill_2 FILLER_33_2349 ();
 sg13g2_fill_1 FILLER_33_2351 ();
 sg13g2_fill_2 FILLER_33_2437 ();
 sg13g2_fill_1 FILLER_33_2439 ();
 sg13g2_fill_2 FILLER_33_2457 ();
 sg13g2_fill_2 FILLER_33_2500 ();
 sg13g2_fill_2 FILLER_33_2538 ();
 sg13g2_fill_2 FILLER_33_2567 ();
 sg13g2_fill_1 FILLER_33_2569 ();
 sg13g2_fill_2 FILLER_33_2603 ();
 sg13g2_fill_2 FILLER_33_2671 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_decap_4 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_480 ();
 sg13g2_fill_1 FILLER_34_482 ();
 sg13g2_fill_2 FILLER_34_526 ();
 sg13g2_fill_1 FILLER_34_528 ();
 sg13g2_fill_1 FILLER_34_550 ();
 sg13g2_fill_2 FILLER_34_569 ();
 sg13g2_fill_1 FILLER_34_580 ();
 sg13g2_fill_2 FILLER_34_634 ();
 sg13g2_decap_8 FILLER_34_639 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_fill_1 FILLER_34_693 ();
 sg13g2_decap_4 FILLER_34_702 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_4 FILLER_34_726 ();
 sg13g2_fill_1 FILLER_34_730 ();
 sg13g2_decap_8 FILLER_34_737 ();
 sg13g2_decap_8 FILLER_34_744 ();
 sg13g2_decap_8 FILLER_34_751 ();
 sg13g2_decap_8 FILLER_34_758 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_fill_2 FILLER_34_772 ();
 sg13g2_decap_4 FILLER_34_783 ();
 sg13g2_fill_2 FILLER_34_787 ();
 sg13g2_decap_4 FILLER_34_802 ();
 sg13g2_decap_4 FILLER_34_842 ();
 sg13g2_fill_1 FILLER_34_879 ();
 sg13g2_fill_1 FILLER_34_894 ();
 sg13g2_fill_2 FILLER_34_1025 ();
 sg13g2_fill_1 FILLER_34_1027 ();
 sg13g2_fill_2 FILLER_34_1057 ();
 sg13g2_fill_2 FILLER_34_1096 ();
 sg13g2_fill_2 FILLER_34_1195 ();
 sg13g2_fill_2 FILLER_34_1229 ();
 sg13g2_fill_1 FILLER_34_1231 ();
 sg13g2_fill_2 FILLER_34_1246 ();
 sg13g2_fill_1 FILLER_34_1303 ();
 sg13g2_decap_8 FILLER_34_1353 ();
 sg13g2_fill_2 FILLER_34_1384 ();
 sg13g2_fill_2 FILLER_34_1393 ();
 sg13g2_fill_1 FILLER_34_1395 ();
 sg13g2_fill_2 FILLER_34_1404 ();
 sg13g2_fill_2 FILLER_34_1411 ();
 sg13g2_fill_1 FILLER_34_1428 ();
 sg13g2_fill_2 FILLER_34_1461 ();
 sg13g2_fill_1 FILLER_34_1463 ();
 sg13g2_fill_2 FILLER_34_1470 ();
 sg13g2_fill_1 FILLER_34_1472 ();
 sg13g2_fill_1 FILLER_34_1501 ();
 sg13g2_fill_2 FILLER_34_1555 ();
 sg13g2_decap_8 FILLER_34_1584 ();
 sg13g2_decap_4 FILLER_34_1591 ();
 sg13g2_fill_2 FILLER_34_1595 ();
 sg13g2_decap_8 FILLER_34_1624 ();
 sg13g2_decap_8 FILLER_34_1631 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_fill_1 FILLER_34_1640 ();
 sg13g2_fill_2 FILLER_34_1670 ();
 sg13g2_fill_1 FILLER_34_1672 ();
 sg13g2_decap_4 FILLER_34_1686 ();
 sg13g2_decap_8 FILLER_34_1708 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_4 FILLER_34_1729 ();
 sg13g2_fill_2 FILLER_34_1792 ();
 sg13g2_fill_1 FILLER_34_1794 ();
 sg13g2_decap_8 FILLER_34_1821 ();
 sg13g2_decap_8 FILLER_34_1828 ();
 sg13g2_fill_2 FILLER_34_1835 ();
 sg13g2_fill_1 FILLER_34_1837 ();
 sg13g2_fill_2 FILLER_34_1887 ();
 sg13g2_fill_1 FILLER_34_1895 ();
 sg13g2_fill_2 FILLER_34_1952 ();
 sg13g2_fill_1 FILLER_34_1954 ();
 sg13g2_fill_2 FILLER_34_1973 ();
 sg13g2_fill_1 FILLER_34_1975 ();
 sg13g2_fill_1 FILLER_34_1990 ();
 sg13g2_fill_2 FILLER_34_2004 ();
 sg13g2_fill_1 FILLER_34_2062 ();
 sg13g2_fill_1 FILLER_34_2094 ();
 sg13g2_fill_2 FILLER_34_2108 ();
 sg13g2_fill_1 FILLER_34_2110 ();
 sg13g2_fill_1 FILLER_34_2163 ();
 sg13g2_fill_2 FILLER_34_2226 ();
 sg13g2_fill_2 FILLER_34_2250 ();
 sg13g2_fill_1 FILLER_34_2252 ();
 sg13g2_fill_2 FILLER_34_2280 ();
 sg13g2_fill_1 FILLER_34_2282 ();
 sg13g2_fill_1 FILLER_34_2305 ();
 sg13g2_fill_2 FILLER_34_2319 ();
 sg13g2_fill_1 FILLER_34_2321 ();
 sg13g2_fill_2 FILLER_34_2349 ();
 sg13g2_fill_1 FILLER_34_2351 ();
 sg13g2_fill_1 FILLER_34_2379 ();
 sg13g2_fill_1 FILLER_34_2393 ();
 sg13g2_fill_1 FILLER_34_2460 ();
 sg13g2_fill_2 FILLER_34_2523 ();
 sg13g2_fill_2 FILLER_34_2566 ();
 sg13g2_fill_1 FILLER_34_2568 ();
 sg13g2_fill_2 FILLER_34_2614 ();
 sg13g2_fill_1 FILLER_34_2616 ();
 sg13g2_fill_2 FILLER_34_2649 ();
 sg13g2_fill_1 FILLER_34_2651 ();
 sg13g2_fill_1 FILLER_34_2673 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_40 ();
 sg13g2_fill_1 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_434 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_516 ();
 sg13g2_fill_2 FILLER_35_580 ();
 sg13g2_fill_1 FILLER_35_586 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_fill_1 FILLER_35_598 ();
 sg13g2_fill_2 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_639 ();
 sg13g2_decap_8 FILLER_35_646 ();
 sg13g2_decap_8 FILLER_35_653 ();
 sg13g2_decap_8 FILLER_35_660 ();
 sg13g2_decap_8 FILLER_35_667 ();
 sg13g2_fill_1 FILLER_35_674 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_fill_1 FILLER_35_728 ();
 sg13g2_fill_1 FILLER_35_734 ();
 sg13g2_decap_8 FILLER_35_747 ();
 sg13g2_decap_8 FILLER_35_754 ();
 sg13g2_decap_8 FILLER_35_761 ();
 sg13g2_decap_8 FILLER_35_768 ();
 sg13g2_decap_8 FILLER_35_775 ();
 sg13g2_decap_8 FILLER_35_782 ();
 sg13g2_fill_1 FILLER_35_789 ();
 sg13g2_fill_1 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_4 FILLER_35_812 ();
 sg13g2_fill_1 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_fill_1 FILLER_35_853 ();
 sg13g2_fill_2 FILLER_35_881 ();
 sg13g2_fill_1 FILLER_35_883 ();
 sg13g2_fill_1 FILLER_35_933 ();
 sg13g2_fill_2 FILLER_35_943 ();
 sg13g2_fill_1 FILLER_35_960 ();
 sg13g2_fill_2 FILLER_35_1012 ();
 sg13g2_fill_2 FILLER_35_1154 ();
 sg13g2_fill_1 FILLER_35_1156 ();
 sg13g2_fill_2 FILLER_35_1319 ();
 sg13g2_fill_2 FILLER_35_1343 ();
 sg13g2_decap_4 FILLER_35_1355 ();
 sg13g2_fill_2 FILLER_35_1369 ();
 sg13g2_fill_1 FILLER_35_1371 ();
 sg13g2_decap_8 FILLER_35_1378 ();
 sg13g2_decap_8 FILLER_35_1385 ();
 sg13g2_fill_1 FILLER_35_1392 ();
 sg13g2_fill_2 FILLER_35_1424 ();
 sg13g2_decap_8 FILLER_35_1464 ();
 sg13g2_fill_1 FILLER_35_1471 ();
 sg13g2_fill_1 FILLER_35_1505 ();
 sg13g2_fill_2 FILLER_35_1535 ();
 sg13g2_fill_1 FILLER_35_1542 ();
 sg13g2_fill_2 FILLER_35_1561 ();
 sg13g2_decap_8 FILLER_35_1567 ();
 sg13g2_decap_8 FILLER_35_1574 ();
 sg13g2_decap_4 FILLER_35_1594 ();
 sg13g2_decap_8 FILLER_35_1619 ();
 sg13g2_decap_4 FILLER_35_1626 ();
 sg13g2_decap_8 FILLER_35_1672 ();
 sg13g2_decap_8 FILLER_35_1679 ();
 sg13g2_fill_2 FILLER_35_1686 ();
 sg13g2_fill_1 FILLER_35_1688 ();
 sg13g2_decap_8 FILLER_35_1695 ();
 sg13g2_fill_2 FILLER_35_1702 ();
 sg13g2_decap_8 FILLER_35_1788 ();
 sg13g2_fill_2 FILLER_35_1795 ();
 sg13g2_fill_1 FILLER_35_1797 ();
 sg13g2_fill_2 FILLER_35_1816 ();
 sg13g2_decap_8 FILLER_35_1826 ();
 sg13g2_fill_2 FILLER_35_1874 ();
 sg13g2_fill_1 FILLER_35_1889 ();
 sg13g2_fill_2 FILLER_35_1896 ();
 sg13g2_fill_1 FILLER_35_1898 ();
 sg13g2_fill_2 FILLER_35_1923 ();
 sg13g2_fill_2 FILLER_35_1938 ();
 sg13g2_fill_2 FILLER_35_1997 ();
 sg13g2_fill_1 FILLER_35_1999 ();
 sg13g2_fill_2 FILLER_35_2012 ();
 sg13g2_fill_2 FILLER_35_2047 ();
 sg13g2_fill_1 FILLER_35_2049 ();
 sg13g2_fill_2 FILLER_35_2077 ();
 sg13g2_decap_4 FILLER_35_2149 ();
 sg13g2_fill_2 FILLER_35_2153 ();
 sg13g2_fill_2 FILLER_35_2256 ();
 sg13g2_fill_2 FILLER_35_2280 ();
 sg13g2_fill_1 FILLER_35_2417 ();
 sg13g2_fill_2 FILLER_35_2436 ();
 sg13g2_fill_2 FILLER_35_2464 ();
 sg13g2_fill_1 FILLER_35_2507 ();
 sg13g2_fill_2 FILLER_35_2548 ();
 sg13g2_fill_1 FILLER_35_2550 ();
 sg13g2_fill_1 FILLER_35_2587 ();
 sg13g2_fill_2 FILLER_35_2634 ();
 sg13g2_fill_1 FILLER_35_2636 ();
 sg13g2_fill_1 FILLER_35_2664 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_decap_4 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_2 FILLER_36_520 ();
 sg13g2_fill_1 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_537 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_decap_4 FILLER_36_586 ();
 sg13g2_fill_1 FILLER_36_590 ();
 sg13g2_fill_1 FILLER_36_607 ();
 sg13g2_fill_2 FILLER_36_663 ();
 sg13g2_fill_1 FILLER_36_665 ();
 sg13g2_fill_2 FILLER_36_683 ();
 sg13g2_fill_1 FILLER_36_685 ();
 sg13g2_decap_8 FILLER_36_696 ();
 sg13g2_decap_8 FILLER_36_703 ();
 sg13g2_decap_8 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_717 ();
 sg13g2_decap_8 FILLER_36_737 ();
 sg13g2_decap_8 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_760 ();
 sg13g2_decap_4 FILLER_36_769 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_fill_1 FILLER_36_847 ();
 sg13g2_decap_4 FILLER_36_875 ();
 sg13g2_fill_2 FILLER_36_923 ();
 sg13g2_fill_1 FILLER_36_933 ();
 sg13g2_fill_1 FILLER_36_1042 ();
 sg13g2_fill_2 FILLER_36_1091 ();
 sg13g2_fill_1 FILLER_36_1143 ();
 sg13g2_fill_2 FILLER_36_1180 ();
 sg13g2_fill_1 FILLER_36_1217 ();
 sg13g2_fill_2 FILLER_36_1231 ();
 sg13g2_fill_2 FILLER_36_1301 ();
 sg13g2_fill_2 FILLER_36_1330 ();
 sg13g2_decap_4 FILLER_36_1390 ();
 sg13g2_fill_2 FILLER_36_1394 ();
 sg13g2_decap_8 FILLER_36_1428 ();
 sg13g2_fill_2 FILLER_36_1435 ();
 sg13g2_decap_8 FILLER_36_1446 ();
 sg13g2_decap_4 FILLER_36_1462 ();
 sg13g2_fill_1 FILLER_36_1466 ();
 sg13g2_decap_8 FILLER_36_1508 ();
 sg13g2_fill_2 FILLER_36_1537 ();
 sg13g2_decap_8 FILLER_36_1561 ();
 sg13g2_decap_8 FILLER_36_1568 ();
 sg13g2_decap_8 FILLER_36_1575 ();
 sg13g2_decap_8 FILLER_36_1582 ();
 sg13g2_fill_2 FILLER_36_1589 ();
 sg13g2_fill_1 FILLER_36_1596 ();
 sg13g2_fill_2 FILLER_36_1602 ();
 sg13g2_fill_1 FILLER_36_1604 ();
 sg13g2_decap_8 FILLER_36_1626 ();
 sg13g2_fill_2 FILLER_36_1633 ();
 sg13g2_fill_2 FILLER_36_1658 ();
 sg13g2_decap_8 FILLER_36_1665 ();
 sg13g2_decap_8 FILLER_36_1676 ();
 sg13g2_decap_8 FILLER_36_1683 ();
 sg13g2_decap_8 FILLER_36_1690 ();
 sg13g2_decap_8 FILLER_36_1739 ();
 sg13g2_decap_8 FILLER_36_1780 ();
 sg13g2_fill_2 FILLER_36_1787 ();
 sg13g2_fill_1 FILLER_36_1789 ();
 sg13g2_fill_2 FILLER_36_1827 ();
 sg13g2_fill_1 FILLER_36_1829 ();
 sg13g2_fill_1 FILLER_36_1913 ();
 sg13g2_fill_2 FILLER_36_1955 ();
 sg13g2_fill_1 FILLER_36_1957 ();
 sg13g2_decap_4 FILLER_36_1963 ();
 sg13g2_fill_2 FILLER_36_2083 ();
 sg13g2_decap_4 FILLER_36_2155 ();
 sg13g2_fill_1 FILLER_36_2172 ();
 sg13g2_fill_2 FILLER_36_2231 ();
 sg13g2_fill_1 FILLER_36_2233 ();
 sg13g2_fill_2 FILLER_36_2284 ();
 sg13g2_fill_2 FILLER_36_2313 ();
 sg13g2_decap_4 FILLER_36_2341 ();
 sg13g2_fill_1 FILLER_36_2345 ();
 sg13g2_fill_1 FILLER_36_2378 ();
 sg13g2_fill_2 FILLER_36_2410 ();
 sg13g2_fill_1 FILLER_36_2448 ();
 sg13g2_fill_2 FILLER_36_2482 ();
 sg13g2_fill_1 FILLER_36_2484 ();
 sg13g2_fill_2 FILLER_36_2498 ();
 sg13g2_fill_1 FILLER_36_2500 ();
 sg13g2_fill_2 FILLER_36_2518 ();
 sg13g2_fill_2 FILLER_36_2552 ();
 sg13g2_fill_1 FILLER_36_2554 ();
 sg13g2_fill_2 FILLER_36_2569 ();
 sg13g2_fill_1 FILLER_36_2589 ();
 sg13g2_fill_1 FILLER_36_2644 ();
 sg13g2_fill_1 FILLER_36_2673 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_62 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_425 ();
 sg13g2_fill_2 FILLER_37_452 ();
 sg13g2_fill_1 FILLER_37_454 ();
 sg13g2_fill_2 FILLER_37_484 ();
 sg13g2_fill_2 FILLER_37_516 ();
 sg13g2_decap_4 FILLER_37_563 ();
 sg13g2_fill_2 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_578 ();
 sg13g2_fill_1 FILLER_37_582 ();
 sg13g2_fill_1 FILLER_37_596 ();
 sg13g2_fill_2 FILLER_37_610 ();
 sg13g2_fill_1 FILLER_37_612 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_4 FILLER_37_657 ();
 sg13g2_fill_2 FILLER_37_677 ();
 sg13g2_fill_1 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_704 ();
 sg13g2_fill_2 FILLER_37_711 ();
 sg13g2_decap_8 FILLER_37_736 ();
 sg13g2_decap_8 FILLER_37_743 ();
 sg13g2_fill_2 FILLER_37_750 ();
 sg13g2_decap_4 FILLER_37_757 ();
 sg13g2_fill_2 FILLER_37_761 ();
 sg13g2_fill_1 FILLER_37_794 ();
 sg13g2_fill_2 FILLER_37_862 ();
 sg13g2_fill_2 FILLER_37_880 ();
 sg13g2_fill_2 FILLER_37_924 ();
 sg13g2_fill_1 FILLER_37_940 ();
 sg13g2_fill_2 FILLER_37_961 ();
 sg13g2_fill_2 FILLER_37_977 ();
 sg13g2_fill_2 FILLER_37_1022 ();
 sg13g2_fill_2 FILLER_37_1035 ();
 sg13g2_fill_1 FILLER_37_1075 ();
 sg13g2_fill_2 FILLER_37_1143 ();
 sg13g2_decap_8 FILLER_37_1186 ();
 sg13g2_decap_8 FILLER_37_1193 ();
 sg13g2_fill_1 FILLER_37_1301 ();
 sg13g2_fill_1 FILLER_37_1397 ();
 sg13g2_fill_2 FILLER_37_1426 ();
 sg13g2_fill_2 FILLER_37_1469 ();
 sg13g2_fill_1 FILLER_37_1471 ();
 sg13g2_decap_4 FILLER_37_1514 ();
 sg13g2_fill_2 FILLER_37_1518 ();
 sg13g2_fill_1 FILLER_37_1524 ();
 sg13g2_fill_2 FILLER_37_1535 ();
 sg13g2_decap_4 FILLER_37_1545 ();
 sg13g2_decap_4 FILLER_37_1555 ();
 sg13g2_decap_4 FILLER_37_1565 ();
 sg13g2_fill_2 FILLER_37_1569 ();
 sg13g2_fill_1 FILLER_37_1583 ();
 sg13g2_fill_1 FILLER_37_1599 ();
 sg13g2_fill_1 FILLER_37_1634 ();
 sg13g2_fill_1 FILLER_37_1662 ();
 sg13g2_fill_1 FILLER_37_1676 ();
 sg13g2_decap_8 FILLER_37_1682 ();
 sg13g2_decap_4 FILLER_37_1689 ();
 sg13g2_fill_1 FILLER_37_1693 ();
 sg13g2_fill_2 FILLER_37_1707 ();
 sg13g2_decap_8 FILLER_37_1719 ();
 sg13g2_decap_8 FILLER_37_1726 ();
 sg13g2_decap_8 FILLER_37_1733 ();
 sg13g2_decap_4 FILLER_37_1753 ();
 sg13g2_decap_8 FILLER_37_1775 ();
 sg13g2_fill_2 FILLER_37_1782 ();
 sg13g2_fill_1 FILLER_37_1882 ();
 sg13g2_decap_8 FILLER_37_1929 ();
 sg13g2_fill_2 FILLER_37_1936 ();
 sg13g2_fill_1 FILLER_37_1996 ();
 sg13g2_fill_1 FILLER_37_2010 ();
 sg13g2_fill_1 FILLER_37_2039 ();
 sg13g2_fill_1 FILLER_37_2059 ();
 sg13g2_decap_4 FILLER_37_2077 ();
 sg13g2_decap_4 FILLER_37_2200 ();
 sg13g2_fill_2 FILLER_37_2255 ();
 sg13g2_fill_1 FILLER_37_2257 ();
 sg13g2_fill_1 FILLER_37_2267 ();
 sg13g2_fill_2 FILLER_37_2273 ();
 sg13g2_fill_2 FILLER_37_2297 ();
 sg13g2_fill_1 FILLER_37_2299 ();
 sg13g2_fill_2 FILLER_37_2365 ();
 sg13g2_fill_1 FILLER_37_2367 ();
 sg13g2_fill_2 FILLER_37_2413 ();
 sg13g2_fill_1 FILLER_37_2415 ();
 sg13g2_fill_2 FILLER_37_2464 ();
 sg13g2_fill_1 FILLER_37_2494 ();
 sg13g2_fill_1 FILLER_37_2565 ();
 sg13g2_fill_2 FILLER_37_2588 ();
 sg13g2_fill_2 FILLER_37_2618 ();
 sg13g2_fill_1 FILLER_37_2620 ();
 sg13g2_fill_2 FILLER_37_2671 ();
 sg13g2_fill_1 FILLER_37_2673 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_decap_4 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_492 ();
 sg13g2_fill_1 FILLER_38_534 ();
 sg13g2_fill_2 FILLER_38_548 ();
 sg13g2_decap_8 FILLER_38_566 ();
 sg13g2_decap_8 FILLER_38_573 ();
 sg13g2_decap_8 FILLER_38_580 ();
 sg13g2_fill_1 FILLER_38_587 ();
 sg13g2_fill_1 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_decap_8 FILLER_38_659 ();
 sg13g2_fill_2 FILLER_38_666 ();
 sg13g2_fill_1 FILLER_38_668 ();
 sg13g2_fill_1 FILLER_38_688 ();
 sg13g2_decap_4 FILLER_38_694 ();
 sg13g2_fill_2 FILLER_38_698 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_715 ();
 sg13g2_fill_2 FILLER_38_722 ();
 sg13g2_decap_4 FILLER_38_729 ();
 sg13g2_fill_2 FILLER_38_733 ();
 sg13g2_decap_4 FILLER_38_741 ();
 sg13g2_fill_2 FILLER_38_745 ();
 sg13g2_fill_2 FILLER_38_763 ();
 sg13g2_fill_1 FILLER_38_765 ();
 sg13g2_fill_1 FILLER_38_790 ();
 sg13g2_fill_2 FILLER_38_819 ();
 sg13g2_fill_1 FILLER_38_821 ();
 sg13g2_fill_2 FILLER_38_832 ();
 sg13g2_fill_1 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_38_844 ();
 sg13g2_fill_2 FILLER_38_863 ();
 sg13g2_fill_2 FILLER_38_899 ();
 sg13g2_fill_1 FILLER_38_901 ();
 sg13g2_fill_1 FILLER_38_927 ();
 sg13g2_fill_2 FILLER_38_976 ();
 sg13g2_fill_2 FILLER_38_1018 ();
 sg13g2_fill_1 FILLER_38_1020 ();
 sg13g2_fill_1 FILLER_38_1062 ();
 sg13g2_fill_1 FILLER_38_1097 ();
 sg13g2_fill_1 FILLER_38_1131 ();
 sg13g2_decap_4 FILLER_38_1182 ();
 sg13g2_fill_1 FILLER_38_1186 ();
 sg13g2_fill_2 FILLER_38_1213 ();
 sg13g2_fill_1 FILLER_38_1215 ();
 sg13g2_fill_2 FILLER_38_1241 ();
 sg13g2_fill_2 FILLER_38_1278 ();
 sg13g2_decap_8 FILLER_38_1289 ();
 sg13g2_fill_2 FILLER_38_1296 ();
 sg13g2_fill_1 FILLER_38_1298 ();
 sg13g2_fill_2 FILLER_38_1325 ();
 sg13g2_decap_4 FILLER_38_1409 ();
 sg13g2_fill_2 FILLER_38_1413 ();
 sg13g2_fill_2 FILLER_38_1449 ();
 sg13g2_fill_2 FILLER_38_1498 ();
 sg13g2_fill_1 FILLER_38_1500 ();
 sg13g2_decap_8 FILLER_38_1518 ();
 sg13g2_fill_2 FILLER_38_1525 ();
 sg13g2_fill_1 FILLER_38_1527 ();
 sg13g2_fill_2 FILLER_38_1541 ();
 sg13g2_fill_2 FILLER_38_1576 ();
 sg13g2_fill_1 FILLER_38_1589 ();
 sg13g2_fill_2 FILLER_38_1605 ();
 sg13g2_fill_1 FILLER_38_1607 ();
 sg13g2_fill_2 FILLER_38_1629 ();
 sg13g2_fill_1 FILLER_38_1631 ();
 sg13g2_fill_2 FILLER_38_1667 ();
 sg13g2_fill_1 FILLER_38_1669 ();
 sg13g2_decap_8 FILLER_38_1690 ();
 sg13g2_fill_1 FILLER_38_1697 ();
 sg13g2_fill_2 FILLER_38_1718 ();
 sg13g2_decap_8 FILLER_38_1730 ();
 sg13g2_decap_8 FILLER_38_1737 ();
 sg13g2_fill_2 FILLER_38_1744 ();
 sg13g2_decap_8 FILLER_38_1774 ();
 sg13g2_decap_8 FILLER_38_1781 ();
 sg13g2_fill_2 FILLER_38_1788 ();
 sg13g2_fill_1 FILLER_38_1790 ();
 sg13g2_fill_2 FILLER_38_1801 ();
 sg13g2_fill_1 FILLER_38_1803 ();
 sg13g2_fill_1 FILLER_38_1866 ();
 sg13g2_fill_2 FILLER_38_1889 ();
 sg13g2_fill_1 FILLER_38_1891 ();
 sg13g2_fill_2 FILLER_38_1922 ();
 sg13g2_decap_8 FILLER_38_1929 ();
 sg13g2_decap_8 FILLER_38_1936 ();
 sg13g2_decap_4 FILLER_38_1943 ();
 sg13g2_decap_8 FILLER_38_1998 ();
 sg13g2_decap_4 FILLER_38_2005 ();
 sg13g2_fill_2 FILLER_38_2021 ();
 sg13g2_decap_8 FILLER_38_2069 ();
 sg13g2_decap_8 FILLER_38_2076 ();
 sg13g2_decap_4 FILLER_38_2083 ();
 sg13g2_fill_1 FILLER_38_2087 ();
 sg13g2_fill_2 FILLER_38_2101 ();
 sg13g2_fill_1 FILLER_38_2103 ();
 sg13g2_fill_2 FILLER_38_2182 ();
 sg13g2_fill_1 FILLER_38_2184 ();
 sg13g2_fill_2 FILLER_38_2204 ();
 sg13g2_fill_1 FILLER_38_2230 ();
 sg13g2_decap_4 FILLER_38_2318 ();
 sg13g2_fill_2 FILLER_38_2322 ();
 sg13g2_fill_1 FILLER_38_2337 ();
 sg13g2_fill_1 FILLER_38_2351 ();
 sg13g2_fill_2 FILLER_38_2378 ();
 sg13g2_fill_1 FILLER_38_2380 ();
 sg13g2_fill_2 FILLER_38_2395 ();
 sg13g2_fill_1 FILLER_38_2397 ();
 sg13g2_fill_2 FILLER_38_2435 ();
 sg13g2_fill_2 FILLER_38_2465 ();
 sg13g2_fill_1 FILLER_38_2467 ();
 sg13g2_fill_1 FILLER_38_2512 ();
 sg13g2_fill_2 FILLER_38_2526 ();
 sg13g2_fill_1 FILLER_38_2604 ();
 sg13g2_fill_2 FILLER_38_2633 ();
 sg13g2_fill_1 FILLER_38_2635 ();
 sg13g2_fill_1 FILLER_38_2673 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_50 ();
 sg13g2_decap_8 FILLER_39_87 ();
 sg13g2_fill_2 FILLER_39_94 ();
 sg13g2_decap_8 FILLER_39_146 ();
 sg13g2_decap_8 FILLER_39_153 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_248 ();
 sg13g2_fill_1 FILLER_39_250 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_379 ();
 sg13g2_fill_2 FILLER_39_435 ();
 sg13g2_fill_1 FILLER_39_452 ();
 sg13g2_fill_2 FILLER_39_487 ();
 sg13g2_decap_8 FILLER_39_515 ();
 sg13g2_fill_2 FILLER_39_522 ();
 sg13g2_fill_1 FILLER_39_524 ();
 sg13g2_fill_2 FILLER_39_538 ();
 sg13g2_decap_4 FILLER_39_546 ();
 sg13g2_fill_1 FILLER_39_563 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_2 FILLER_39_606 ();
 sg13g2_fill_1 FILLER_39_608 ();
 sg13g2_decap_8 FILLER_39_636 ();
 sg13g2_decap_8 FILLER_39_643 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_decap_4 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_677 ();
 sg13g2_decap_8 FILLER_39_684 ();
 sg13g2_decap_4 FILLER_39_691 ();
 sg13g2_fill_2 FILLER_39_695 ();
 sg13g2_decap_8 FILLER_39_705 ();
 sg13g2_decap_8 FILLER_39_712 ();
 sg13g2_decap_8 FILLER_39_719 ();
 sg13g2_decap_8 FILLER_39_726 ();
 sg13g2_fill_2 FILLER_39_733 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_4 FILLER_39_779 ();
 sg13g2_fill_2 FILLER_39_783 ();
 sg13g2_decap_4 FILLER_39_878 ();
 sg13g2_fill_2 FILLER_39_897 ();
 sg13g2_fill_1 FILLER_39_899 ();
 sg13g2_fill_1 FILLER_39_946 ();
 sg13g2_fill_1 FILLER_39_1000 ();
 sg13g2_decap_4 FILLER_39_1103 ();
 sg13g2_fill_2 FILLER_39_1116 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_decap_4 FILLER_39_1147 ();
 sg13g2_fill_2 FILLER_39_1222 ();
 sg13g2_fill_1 FILLER_39_1224 ();
 sg13g2_fill_1 FILLER_39_1243 ();
 sg13g2_decap_8 FILLER_39_1293 ();
 sg13g2_fill_1 FILLER_39_1300 ();
 sg13g2_decap_8 FILLER_39_1304 ();
 sg13g2_fill_1 FILLER_39_1311 ();
 sg13g2_decap_4 FILLER_39_1318 ();
 sg13g2_fill_1 FILLER_39_1322 ();
 sg13g2_fill_1 FILLER_39_1326 ();
 sg13g2_decap_4 FILLER_39_1336 ();
 sg13g2_fill_1 FILLER_39_1362 ();
 sg13g2_fill_1 FILLER_39_1391 ();
 sg13g2_fill_2 FILLER_39_1412 ();
 sg13g2_fill_1 FILLER_39_1414 ();
 sg13g2_fill_2 FILLER_39_1452 ();
 sg13g2_fill_2 FILLER_39_1491 ();
 sg13g2_fill_2 FILLER_39_1522 ();
 sg13g2_decap_4 FILLER_39_1533 ();
 sg13g2_fill_2 FILLER_39_1537 ();
 sg13g2_fill_2 FILLER_39_1592 ();
 sg13g2_decap_8 FILLER_39_1610 ();
 sg13g2_decap_8 FILLER_39_1617 ();
 sg13g2_decap_8 FILLER_39_1624 ();
 sg13g2_decap_8 FILLER_39_1631 ();
 sg13g2_fill_2 FILLER_39_1638 ();
 sg13g2_fill_1 FILLER_39_1640 ();
 sg13g2_decap_4 FILLER_39_1659 ();
 sg13g2_decap_8 FILLER_39_1688 ();
 sg13g2_decap_8 FILLER_39_1695 ();
 sg13g2_decap_8 FILLER_39_1702 ();
 sg13g2_decap_4 FILLER_39_1709 ();
 sg13g2_fill_2 FILLER_39_1713 ();
 sg13g2_decap_4 FILLER_39_1735 ();
 sg13g2_fill_1 FILLER_39_1739 ();
 sg13g2_fill_2 FILLER_39_1760 ();
 sg13g2_decap_4 FILLER_39_1780 ();
 sg13g2_fill_2 FILLER_39_1784 ();
 sg13g2_fill_2 FILLER_39_1857 ();
 sg13g2_fill_1 FILLER_39_1886 ();
 sg13g2_decap_8 FILLER_39_1896 ();
 sg13g2_fill_2 FILLER_39_1957 ();
 sg13g2_fill_1 FILLER_39_1959 ();
 sg13g2_fill_1 FILLER_39_2006 ();
 sg13g2_decap_8 FILLER_39_2016 ();
 sg13g2_decap_4 FILLER_39_2023 ();
 sg13g2_fill_1 FILLER_39_2027 ();
 sg13g2_fill_1 FILLER_39_2055 ();
 sg13g2_decap_4 FILLER_39_2060 ();
 sg13g2_fill_1 FILLER_39_2064 ();
 sg13g2_fill_2 FILLER_39_2069 ();
 sg13g2_fill_1 FILLER_39_2071 ();
 sg13g2_fill_1 FILLER_39_2098 ();
 sg13g2_fill_2 FILLER_39_2151 ();
 sg13g2_fill_1 FILLER_39_2153 ();
 sg13g2_fill_2 FILLER_39_2193 ();
 sg13g2_fill_1 FILLER_39_2195 ();
 sg13g2_fill_1 FILLER_39_2235 ();
 sg13g2_fill_2 FILLER_39_2257 ();
 sg13g2_fill_2 FILLER_39_2281 ();
 sg13g2_decap_8 FILLER_39_2315 ();
 sg13g2_fill_2 FILLER_39_2322 ();
 sg13g2_fill_2 FILLER_39_2337 ();
 sg13g2_decap_4 FILLER_39_2431 ();
 sg13g2_fill_1 FILLER_39_2435 ();
 sg13g2_fill_1 FILLER_39_2446 ();
 sg13g2_fill_2 FILLER_39_2480 ();
 sg13g2_fill_1 FILLER_39_2482 ();
 sg13g2_fill_1 FILLER_39_2523 ();
 sg13g2_fill_1 FILLER_39_2552 ();
 sg13g2_fill_2 FILLER_39_2581 ();
 sg13g2_decap_8 FILLER_39_2611 ();
 sg13g2_fill_2 FILLER_39_2636 ();
 sg13g2_fill_1 FILLER_39_2638 ();
 sg13g2_decap_8 FILLER_39_2667 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_21 ();
 sg13g2_fill_2 FILLER_40_41 ();
 sg13g2_fill_1 FILLER_40_83 ();
 sg13g2_fill_1 FILLER_40_93 ();
 sg13g2_decap_8 FILLER_40_146 ();
 sg13g2_decap_4 FILLER_40_153 ();
 sg13g2_fill_2 FILLER_40_183 ();
 sg13g2_fill_1 FILLER_40_185 ();
 sg13g2_decap_4 FILLER_40_206 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_decap_4 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_364 ();
 sg13g2_fill_1 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_505 ();
 sg13g2_decap_4 FILLER_40_525 ();
 sg13g2_fill_2 FILLER_40_529 ();
 sg13g2_fill_2 FILLER_40_547 ();
 sg13g2_fill_2 FILLER_40_559 ();
 sg13g2_decap_8 FILLER_40_566 ();
 sg13g2_decap_8 FILLER_40_573 ();
 sg13g2_fill_2 FILLER_40_580 ();
 sg13g2_fill_1 FILLER_40_587 ();
 sg13g2_decap_4 FILLER_40_596 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_decap_8 FILLER_40_645 ();
 sg13g2_fill_1 FILLER_40_652 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_4 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_703 ();
 sg13g2_decap_8 FILLER_40_710 ();
 sg13g2_fill_1 FILLER_40_731 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_4 FILLER_40_780 ();
 sg13g2_fill_1 FILLER_40_784 ();
 sg13g2_fill_2 FILLER_40_845 ();
 sg13g2_fill_1 FILLER_40_847 ();
 sg13g2_fill_2 FILLER_40_947 ();
 sg13g2_fill_2 FILLER_40_961 ();
 sg13g2_fill_1 FILLER_40_963 ();
 sg13g2_fill_2 FILLER_40_986 ();
 sg13g2_fill_1 FILLER_40_1068 ();
 sg13g2_decap_8 FILLER_40_1149 ();
 sg13g2_fill_2 FILLER_40_1156 ();
 sg13g2_fill_1 FILLER_40_1195 ();
 sg13g2_decap_8 FILLER_40_1223 ();
 sg13g2_fill_1 FILLER_40_1230 ();
 sg13g2_fill_1 FILLER_40_1259 ();
 sg13g2_decap_8 FILLER_40_1316 ();
 sg13g2_fill_1 FILLER_40_1323 ();
 sg13g2_fill_1 FILLER_40_1333 ();
 sg13g2_fill_1 FILLER_40_1343 ();
 sg13g2_fill_2 FILLER_40_1349 ();
 sg13g2_fill_1 FILLER_40_1351 ();
 sg13g2_decap_8 FILLER_40_1356 ();
 sg13g2_decap_4 FILLER_40_1363 ();
 sg13g2_fill_2 FILLER_40_1367 ();
 sg13g2_fill_1 FILLER_40_1381 ();
 sg13g2_fill_2 FILLER_40_1386 ();
 sg13g2_decap_8 FILLER_40_1409 ();
 sg13g2_decap_8 FILLER_40_1416 ();
 sg13g2_decap_8 FILLER_40_1423 ();
 sg13g2_decap_4 FILLER_40_1435 ();
 sg13g2_fill_1 FILLER_40_1439 ();
 sg13g2_fill_2 FILLER_40_1454 ();
 sg13g2_fill_1 FILLER_40_1456 ();
 sg13g2_decap_8 FILLER_40_1553 ();
 sg13g2_decap_4 FILLER_40_1560 ();
 sg13g2_decap_8 FILLER_40_1605 ();
 sg13g2_fill_2 FILLER_40_1612 ();
 sg13g2_fill_1 FILLER_40_1614 ();
 sg13g2_decap_8 FILLER_40_1620 ();
 sg13g2_decap_8 FILLER_40_1627 ();
 sg13g2_decap_8 FILLER_40_1634 ();
 sg13g2_decap_8 FILLER_40_1641 ();
 sg13g2_decap_4 FILLER_40_1648 ();
 sg13g2_fill_2 FILLER_40_1652 ();
 sg13g2_decap_4 FILLER_40_1659 ();
 sg13g2_fill_1 FILLER_40_1669 ();
 sg13g2_decap_8 FILLER_40_1674 ();
 sg13g2_decap_8 FILLER_40_1681 ();
 sg13g2_decap_8 FILLER_40_1688 ();
 sg13g2_decap_8 FILLER_40_1695 ();
 sg13g2_decap_8 FILLER_40_1702 ();
 sg13g2_decap_8 FILLER_40_1709 ();
 sg13g2_decap_8 FILLER_40_1716 ();
 sg13g2_fill_2 FILLER_40_1723 ();
 sg13g2_decap_4 FILLER_40_1735 ();
 sg13g2_fill_2 FILLER_40_1782 ();
 sg13g2_fill_1 FILLER_40_1784 ();
 sg13g2_fill_2 FILLER_40_1826 ();
 sg13g2_fill_1 FILLER_40_1828 ();
 sg13g2_decap_4 FILLER_40_1856 ();
 sg13g2_decap_8 FILLER_40_1887 ();
 sg13g2_fill_2 FILLER_40_1894 ();
 sg13g2_fill_1 FILLER_40_1896 ();
 sg13g2_fill_1 FILLER_40_1946 ();
 sg13g2_fill_2 FILLER_40_1983 ();
 sg13g2_fill_2 FILLER_40_2016 ();
 sg13g2_fill_1 FILLER_40_2018 ();
 sg13g2_fill_2 FILLER_40_2051 ();
 sg13g2_fill_1 FILLER_40_2058 ();
 sg13g2_decap_4 FILLER_40_2082 ();
 sg13g2_fill_1 FILLER_40_2086 ();
 sg13g2_fill_2 FILLER_40_2152 ();
 sg13g2_fill_1 FILLER_40_2154 ();
 sg13g2_fill_2 FILLER_40_2212 ();
 sg13g2_fill_1 FILLER_40_2285 ();
 sg13g2_decap_8 FILLER_40_2313 ();
 sg13g2_decap_4 FILLER_40_2346 ();
 sg13g2_fill_1 FILLER_40_2350 ();
 sg13g2_fill_2 FILLER_40_2377 ();
 sg13g2_fill_2 FILLER_40_2397 ();
 sg13g2_decap_8 FILLER_40_2426 ();
 sg13g2_fill_1 FILLER_40_2433 ();
 sg13g2_fill_2 FILLER_40_2475 ();
 sg13g2_fill_2 FILLER_40_2533 ();
 sg13g2_decap_4 FILLER_40_2540 ();
 sg13g2_fill_1 FILLER_40_2544 ();
 sg13g2_fill_2 FILLER_40_2554 ();
 sg13g2_fill_2 FILLER_40_2573 ();
 sg13g2_fill_1 FILLER_40_2596 ();
 sg13g2_decap_8 FILLER_40_2611 ();
 sg13g2_fill_2 FILLER_40_2618 ();
 sg13g2_fill_1 FILLER_40_2620 ();
 sg13g2_decap_8 FILLER_40_2665 ();
 sg13g2_fill_2 FILLER_40_2672 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_46 ();
 sg13g2_fill_1 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_1 FILLER_41_145 ();
 sg13g2_fill_2 FILLER_41_151 ();
 sg13g2_fill_1 FILLER_41_153 ();
 sg13g2_decap_4 FILLER_41_160 ();
 sg13g2_decap_8 FILLER_41_199 ();
 sg13g2_decap_4 FILLER_41_206 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_311 ();
 sg13g2_decap_4 FILLER_41_327 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_1 FILLER_41_381 ();
 sg13g2_fill_2 FILLER_41_403 ();
 sg13g2_fill_1 FILLER_41_405 ();
 sg13g2_fill_2 FILLER_41_439 ();
 sg13g2_fill_1 FILLER_41_525 ();
 sg13g2_fill_2 FILLER_41_569 ();
 sg13g2_fill_2 FILLER_41_577 ();
 sg13g2_fill_1 FILLER_41_579 ();
 sg13g2_fill_2 FILLER_41_601 ();
 sg13g2_decap_4 FILLER_41_650 ();
 sg13g2_fill_1 FILLER_41_690 ();
 sg13g2_decap_4 FILLER_41_704 ();
 sg13g2_fill_2 FILLER_41_708 ();
 sg13g2_fill_1 FILLER_41_751 ();
 sg13g2_fill_1 FILLER_41_802 ();
 sg13g2_fill_2 FILLER_41_824 ();
 sg13g2_fill_1 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_fill_2 FILLER_41_866 ();
 sg13g2_fill_2 FILLER_41_942 ();
 sg13g2_fill_1 FILLER_41_1016 ();
 sg13g2_fill_1 FILLER_41_1031 ();
 sg13g2_fill_2 FILLER_41_1049 ();
 sg13g2_fill_2 FILLER_41_1078 ();
 sg13g2_fill_2 FILLER_41_1123 ();
 sg13g2_fill_1 FILLER_41_1125 ();
 sg13g2_fill_2 FILLER_41_1134 ();
 sg13g2_fill_2 FILLER_41_1217 ();
 sg13g2_decap_8 FILLER_41_1223 ();
 sg13g2_fill_1 FILLER_41_1230 ();
 sg13g2_decap_8 FILLER_41_1244 ();
 sg13g2_fill_1 FILLER_41_1251 ();
 sg13g2_fill_2 FILLER_41_1258 ();
 sg13g2_fill_1 FILLER_41_1260 ();
 sg13g2_decap_8 FILLER_41_1274 ();
 sg13g2_decap_4 FILLER_41_1281 ();
 sg13g2_fill_1 FILLER_41_1313 ();
 sg13g2_fill_1 FILLER_41_1342 ();
 sg13g2_fill_2 FILLER_41_1370 ();
 sg13g2_fill_1 FILLER_41_1372 ();
 sg13g2_fill_2 FILLER_41_1389 ();
 sg13g2_decap_8 FILLER_41_1404 ();
 sg13g2_decap_4 FILLER_41_1411 ();
 sg13g2_fill_1 FILLER_41_1415 ();
 sg13g2_fill_1 FILLER_41_1455 ();
 sg13g2_fill_2 FILLER_41_1464 ();
 sg13g2_fill_2 FILLER_41_1471 ();
 sg13g2_fill_1 FILLER_41_1473 ();
 sg13g2_fill_1 FILLER_41_1491 ();
 sg13g2_fill_2 FILLER_41_1538 ();
 sg13g2_decap_8 FILLER_41_1557 ();
 sg13g2_fill_1 FILLER_41_1569 ();
 sg13g2_fill_1 FILLER_41_1575 ();
 sg13g2_decap_8 FILLER_41_1581 ();
 sg13g2_fill_1 FILLER_41_1588 ();
 sg13g2_decap_8 FILLER_41_1593 ();
 sg13g2_decap_4 FILLER_41_1600 ();
 sg13g2_decap_4 FILLER_41_1617 ();
 sg13g2_decap_8 FILLER_41_1626 ();
 sg13g2_decap_4 FILLER_41_1633 ();
 sg13g2_fill_1 FILLER_41_1637 ();
 sg13g2_decap_8 FILLER_41_1650 ();
 sg13g2_fill_1 FILLER_41_1657 ();
 sg13g2_decap_8 FILLER_41_1671 ();
 sg13g2_decap_8 FILLER_41_1678 ();
 sg13g2_decap_4 FILLER_41_1685 ();
 sg13g2_fill_1 FILLER_41_1698 ();
 sg13g2_fill_1 FILLER_41_1749 ();
 sg13g2_decap_8 FILLER_41_1774 ();
 sg13g2_decap_8 FILLER_41_1781 ();
 sg13g2_decap_8 FILLER_41_1788 ();
 sg13g2_decap_4 FILLER_41_1795 ();
 sg13g2_fill_2 FILLER_41_1799 ();
 sg13g2_decap_4 FILLER_41_1819 ();
 sg13g2_fill_2 FILLER_41_1823 ();
 sg13g2_decap_8 FILLER_41_1829 ();
 sg13g2_decap_8 FILLER_41_1836 ();
 sg13g2_decap_4 FILLER_41_1843 ();
 sg13g2_fill_2 FILLER_41_1870 ();
 sg13g2_fill_2 FILLER_41_1917 ();
 sg13g2_fill_1 FILLER_41_1919 ();
 sg13g2_decap_8 FILLER_41_1938 ();
 sg13g2_decap_8 FILLER_41_1945 ();
 sg13g2_fill_1 FILLER_41_1952 ();
 sg13g2_fill_2 FILLER_41_1980 ();
 sg13g2_fill_2 FILLER_41_2014 ();
 sg13g2_fill_1 FILLER_41_2078 ();
 sg13g2_fill_1 FILLER_41_2178 ();
 sg13g2_fill_2 FILLER_41_2244 ();
 sg13g2_decap_4 FILLER_41_2383 ();
 sg13g2_fill_2 FILLER_41_2439 ();
 sg13g2_fill_1 FILLER_41_2441 ();
 sg13g2_fill_2 FILLER_41_2470 ();
 sg13g2_fill_1 FILLER_41_2472 ();
 sg13g2_fill_2 FILLER_41_2482 ();
 sg13g2_decap_8 FILLER_41_2489 ();
 sg13g2_decap_4 FILLER_41_2501 ();
 sg13g2_fill_2 FILLER_41_2505 ();
 sg13g2_fill_2 FILLER_41_2538 ();
 sg13g2_decap_8 FILLER_41_2549 ();
 sg13g2_fill_1 FILLER_41_2556 ();
 sg13g2_decap_8 FILLER_41_2561 ();
 sg13g2_decap_4 FILLER_41_2568 ();
 sg13g2_fill_2 FILLER_41_2572 ();
 sg13g2_decap_4 FILLER_41_2587 ();
 sg13g2_fill_2 FILLER_41_2591 ();
 sg13g2_decap_8 FILLER_41_2597 ();
 sg13g2_fill_2 FILLER_41_2604 ();
 sg13g2_fill_1 FILLER_41_2606 ();
 sg13g2_fill_1 FILLER_41_2619 ();
 sg13g2_fill_2 FILLER_41_2634 ();
 sg13g2_fill_1 FILLER_41_2636 ();
 sg13g2_fill_1 FILLER_41_2673 ();
 sg13g2_fill_2 FILLER_42_16 ();
 sg13g2_fill_1 FILLER_42_18 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_114 ();
 sg13g2_decap_4 FILLER_42_157 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_201 ();
 sg13g2_decap_4 FILLER_42_227 ();
 sg13g2_fill_1 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_fill_2 FILLER_42_252 ();
 sg13g2_fill_1 FILLER_42_254 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_decap_4 FILLER_42_298 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_decap_4 FILLER_42_313 ();
 sg13g2_decap_4 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_359 ();
 sg13g2_fill_2 FILLER_42_378 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_1 FILLER_42_409 ();
 sg13g2_fill_2 FILLER_42_446 ();
 sg13g2_fill_2 FILLER_42_491 ();
 sg13g2_fill_1 FILLER_42_506 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_591 ();
 sg13g2_decap_8 FILLER_42_598 ();
 sg13g2_decap_4 FILLER_42_612 ();
 sg13g2_fill_2 FILLER_42_616 ();
 sg13g2_fill_2 FILLER_42_654 ();
 sg13g2_fill_2 FILLER_42_712 ();
 sg13g2_fill_1 FILLER_42_714 ();
 sg13g2_decap_4 FILLER_42_722 ();
 sg13g2_fill_1 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_fill_2 FILLER_42_813 ();
 sg13g2_fill_2 FILLER_42_843 ();
 sg13g2_fill_2 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_873 ();
 sg13g2_decap_8 FILLER_42_880 ();
 sg13g2_fill_2 FILLER_42_887 ();
 sg13g2_fill_1 FILLER_42_914 ();
 sg13g2_fill_1 FILLER_42_924 ();
 sg13g2_fill_2 FILLER_42_977 ();
 sg13g2_fill_2 FILLER_42_1049 ();
 sg13g2_decap_4 FILLER_42_1094 ();
 sg13g2_decap_8 FILLER_42_1103 ();
 sg13g2_fill_2 FILLER_42_1110 ();
 sg13g2_fill_2 FILLER_42_1145 ();
 sg13g2_fill_1 FILLER_42_1147 ();
 sg13g2_fill_2 FILLER_42_1161 ();
 sg13g2_fill_1 FILLER_42_1163 ();
 sg13g2_fill_1 FILLER_42_1187 ();
 sg13g2_fill_2 FILLER_42_1218 ();
 sg13g2_fill_1 FILLER_42_1233 ();
 sg13g2_fill_2 FILLER_42_1244 ();
 sg13g2_fill_2 FILLER_42_1347 ();
 sg13g2_decap_4 FILLER_42_1375 ();
 sg13g2_fill_2 FILLER_42_1385 ();
 sg13g2_fill_1 FILLER_42_1387 ();
 sg13g2_fill_1 FILLER_42_1396 ();
 sg13g2_fill_1 FILLER_42_1403 ();
 sg13g2_fill_2 FILLER_42_1432 ();
 sg13g2_fill_1 FILLER_42_1434 ();
 sg13g2_decap_8 FILLER_42_1477 ();
 sg13g2_fill_1 FILLER_42_1484 ();
 sg13g2_decap_8 FILLER_42_1518 ();
 sg13g2_decap_8 FILLER_42_1525 ();
 sg13g2_decap_8 FILLER_42_1532 ();
 sg13g2_fill_1 FILLER_42_1539 ();
 sg13g2_decap_8 FILLER_42_1553 ();
 sg13g2_decap_8 FILLER_42_1560 ();
 sg13g2_decap_4 FILLER_42_1567 ();
 sg13g2_decap_8 FILLER_42_1581 ();
 sg13g2_decap_8 FILLER_42_1614 ();
 sg13g2_fill_2 FILLER_42_1621 ();
 sg13g2_decap_8 FILLER_42_1628 ();
 sg13g2_fill_1 FILLER_42_1635 ();
 sg13g2_decap_8 FILLER_42_1640 ();
 sg13g2_decap_8 FILLER_42_1647 ();
 sg13g2_decap_4 FILLER_42_1654 ();
 sg13g2_fill_1 FILLER_42_1658 ();
 sg13g2_fill_2 FILLER_42_1686 ();
 sg13g2_fill_1 FILLER_42_1688 ();
 sg13g2_fill_2 FILLER_42_1699 ();
 sg13g2_fill_1 FILLER_42_1701 ();
 sg13g2_fill_1 FILLER_42_1707 ();
 sg13g2_decap_8 FILLER_42_1733 ();
 sg13g2_decap_8 FILLER_42_1740 ();
 sg13g2_decap_4 FILLER_42_1747 ();
 sg13g2_fill_1 FILLER_42_1751 ();
 sg13g2_decap_8 FILLER_42_1764 ();
 sg13g2_decap_8 FILLER_42_1771 ();
 sg13g2_fill_2 FILLER_42_1778 ();
 sg13g2_fill_2 FILLER_42_1793 ();
 sg13g2_fill_1 FILLER_42_1795 ();
 sg13g2_decap_8 FILLER_42_1828 ();
 sg13g2_decap_4 FILLER_42_1835 ();
 sg13g2_fill_2 FILLER_42_1839 ();
 sg13g2_decap_4 FILLER_42_1846 ();
 sg13g2_fill_1 FILLER_42_1850 ();
 sg13g2_fill_2 FILLER_42_1864 ();
 sg13g2_fill_2 FILLER_42_1883 ();
 sg13g2_fill_1 FILLER_42_1885 ();
 sg13g2_fill_1 FILLER_42_1913 ();
 sg13g2_decap_8 FILLER_42_1941 ();
 sg13g2_fill_2 FILLER_42_1979 ();
 sg13g2_fill_1 FILLER_42_2008 ();
 sg13g2_decap_4 FILLER_42_2049 ();
 sg13g2_decap_4 FILLER_42_2119 ();
 sg13g2_fill_2 FILLER_42_2213 ();
 sg13g2_fill_1 FILLER_42_2221 ();
 sg13g2_fill_1 FILLER_42_2300 ();
 sg13g2_fill_1 FILLER_42_2436 ();
 sg13g2_fill_2 FILLER_42_2450 ();
 sg13g2_fill_1 FILLER_42_2452 ();
 sg13g2_decap_4 FILLER_42_2466 ();
 sg13g2_decap_8 FILLER_42_2474 ();
 sg13g2_decap_8 FILLER_42_2481 ();
 sg13g2_decap_8 FILLER_42_2488 ();
 sg13g2_decap_8 FILLER_42_2495 ();
 sg13g2_decap_8 FILLER_42_2502 ();
 sg13g2_fill_2 FILLER_42_2509 ();
 sg13g2_decap_8 FILLER_42_2528 ();
 sg13g2_decap_8 FILLER_42_2535 ();
 sg13g2_decap_4 FILLER_42_2542 ();
 sg13g2_fill_2 FILLER_42_2546 ();
 sg13g2_decap_8 FILLER_42_2561 ();
 sg13g2_fill_2 FILLER_42_2573 ();
 sg13g2_fill_2 FILLER_42_2607 ();
 sg13g2_fill_1 FILLER_42_2609 ();
 sg13g2_decap_4 FILLER_42_2657 ();
 sg13g2_fill_1 FILLER_42_2661 ();
 sg13g2_decap_8 FILLER_42_2666 ();
 sg13g2_fill_1 FILLER_42_2673 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_38 ();
 sg13g2_fill_1 FILLER_43_40 ();
 sg13g2_decap_4 FILLER_43_77 ();
 sg13g2_fill_2 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_4 FILLER_43_166 ();
 sg13g2_fill_1 FILLER_43_180 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_decap_4 FILLER_43_212 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_235 ();
 sg13g2_fill_2 FILLER_43_241 ();
 sg13g2_fill_1 FILLER_43_243 ();
 sg13g2_decap_8 FILLER_43_250 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_fill_2 FILLER_43_264 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_fill_2 FILLER_43_367 ();
 sg13g2_fill_1 FILLER_43_425 ();
 sg13g2_fill_2 FILLER_43_533 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_4 FILLER_43_551 ();
 sg13g2_fill_2 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_594 ();
 sg13g2_decap_4 FILLER_43_601 ();
 sg13g2_fill_1 FILLER_43_605 ();
 sg13g2_fill_2 FILLER_43_616 ();
 sg13g2_decap_4 FILLER_43_623 ();
 sg13g2_fill_2 FILLER_43_627 ();
 sg13g2_fill_2 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_636 ();
 sg13g2_fill_2 FILLER_43_661 ();
 sg13g2_fill_1 FILLER_43_672 ();
 sg13g2_fill_1 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_714 ();
 sg13g2_fill_1 FILLER_43_741 ();
 sg13g2_fill_1 FILLER_43_767 ();
 sg13g2_fill_1 FILLER_43_831 ();
 sg13g2_fill_1 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_872 ();
 sg13g2_decap_4 FILLER_43_879 ();
 sg13g2_fill_2 FILLER_43_936 ();
 sg13g2_fill_1 FILLER_43_938 ();
 sg13g2_fill_1 FILLER_43_1000 ();
 sg13g2_fill_1 FILLER_43_1019 ();
 sg13g2_fill_2 FILLER_43_1059 ();
 sg13g2_decap_8 FILLER_43_1100 ();
 sg13g2_decap_8 FILLER_43_1107 ();
 sg13g2_decap_8 FILLER_43_1114 ();
 sg13g2_decap_4 FILLER_43_1121 ();
 sg13g2_fill_1 FILLER_43_1125 ();
 sg13g2_decap_8 FILLER_43_1149 ();
 sg13g2_fill_2 FILLER_43_1217 ();
 sg13g2_fill_1 FILLER_43_1219 ();
 sg13g2_fill_2 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1226 ();
 sg13g2_fill_2 FILLER_43_1277 ();
 sg13g2_fill_1 FILLER_43_1279 ();
 sg13g2_fill_2 FILLER_43_1355 ();
 sg13g2_fill_1 FILLER_43_1357 ();
 sg13g2_fill_2 FILLER_43_1374 ();
 sg13g2_decap_4 FILLER_43_1382 ();
 sg13g2_fill_1 FILLER_43_1386 ();
 sg13g2_fill_1 FILLER_43_1391 ();
 sg13g2_fill_1 FILLER_43_1420 ();
 sg13g2_decap_4 FILLER_43_1431 ();
 sg13g2_fill_2 FILLER_43_1435 ();
 sg13g2_fill_2 FILLER_43_1466 ();
 sg13g2_fill_1 FILLER_43_1468 ();
 sg13g2_fill_1 FILLER_43_1483 ();
 sg13g2_decap_4 FILLER_43_1512 ();
 sg13g2_fill_1 FILLER_43_1525 ();
 sg13g2_decap_8 FILLER_43_1529 ();
 sg13g2_fill_1 FILLER_43_1536 ();
 sg13g2_decap_8 FILLER_43_1546 ();
 sg13g2_decap_8 FILLER_43_1553 ();
 sg13g2_fill_2 FILLER_43_1560 ();
 sg13g2_fill_2 FILLER_43_1585 ();
 sg13g2_fill_1 FILLER_43_1587 ();
 sg13g2_fill_2 FILLER_43_1599 ();
 sg13g2_fill_1 FILLER_43_1601 ();
 sg13g2_fill_2 FILLER_43_1615 ();
 sg13g2_fill_2 FILLER_43_1622 ();
 sg13g2_fill_1 FILLER_43_1624 ();
 sg13g2_fill_1 FILLER_43_1630 ();
 sg13g2_decap_8 FILLER_43_1636 ();
 sg13g2_decap_8 FILLER_43_1643 ();
 sg13g2_fill_2 FILLER_43_1655 ();
 sg13g2_fill_1 FILLER_43_1657 ();
 sg13g2_decap_4 FILLER_43_1663 ();
 sg13g2_fill_2 FILLER_43_1667 ();
 sg13g2_decap_8 FILLER_43_1675 ();
 sg13g2_decap_8 FILLER_43_1682 ();
 sg13g2_decap_4 FILLER_43_1694 ();
 sg13g2_decap_8 FILLER_43_1721 ();
 sg13g2_decap_8 FILLER_43_1728 ();
 sg13g2_decap_8 FILLER_43_1735 ();
 sg13g2_decap_8 FILLER_43_1742 ();
 sg13g2_fill_1 FILLER_43_1753 ();
 sg13g2_decap_8 FILLER_43_1758 ();
 sg13g2_decap_4 FILLER_43_1765 ();
 sg13g2_fill_2 FILLER_43_1769 ();
 sg13g2_fill_2 FILLER_43_1834 ();
 sg13g2_decap_4 FILLER_43_1891 ();
 sg13g2_fill_2 FILLER_43_1895 ();
 sg13g2_fill_1 FILLER_43_1933 ();
 sg13g2_decap_8 FILLER_43_1947 ();
 sg13g2_fill_2 FILLER_43_1954 ();
 sg13g2_fill_1 FILLER_43_1956 ();
 sg13g2_decap_8 FILLER_43_1984 ();
 sg13g2_decap_8 FILLER_43_1991 ();
 sg13g2_fill_2 FILLER_43_1998 ();
 sg13g2_fill_1 FILLER_43_2013 ();
 sg13g2_decap_8 FILLER_43_2051 ();
 sg13g2_decap_8 FILLER_43_2058 ();
 sg13g2_fill_2 FILLER_43_2065 ();
 sg13g2_fill_2 FILLER_43_2093 ();
 sg13g2_decap_4 FILLER_43_2108 ();
 sg13g2_decap_4 FILLER_43_2202 ();
 sg13g2_fill_2 FILLER_43_2206 ();
 sg13g2_fill_2 FILLER_43_2226 ();
 sg13g2_decap_4 FILLER_43_2259 ();
 sg13g2_fill_2 FILLER_43_2263 ();
 sg13g2_fill_2 FILLER_43_2278 ();
 sg13g2_fill_1 FILLER_43_2280 ();
 sg13g2_fill_1 FILLER_43_2299 ();
 sg13g2_decap_4 FILLER_43_2327 ();
 sg13g2_fill_1 FILLER_43_2331 ();
 sg13g2_fill_1 FILLER_43_2345 ();
 sg13g2_fill_2 FILLER_43_2425 ();
 sg13g2_fill_1 FILLER_43_2427 ();
 sg13g2_decap_4 FILLER_43_2433 ();
 sg13g2_fill_1 FILLER_43_2437 ();
 sg13g2_fill_1 FILLER_43_2451 ();
 sg13g2_fill_2 FILLER_43_2460 ();
 sg13g2_decap_4 FILLER_43_2475 ();
 sg13g2_fill_2 FILLER_43_2479 ();
 sg13g2_decap_8 FILLER_43_2494 ();
 sg13g2_fill_2 FILLER_43_2501 ();
 sg13g2_fill_1 FILLER_43_2503 ();
 sg13g2_decap_4 FILLER_43_2535 ();
 sg13g2_fill_2 FILLER_43_2578 ();
 sg13g2_fill_1 FILLER_43_2580 ();
 sg13g2_fill_2 FILLER_43_2662 ();
 sg13g2_fill_1 FILLER_43_2664 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_38 ();
 sg13g2_fill_1 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_2 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_164 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_2 FILLER_44_178 ();
 sg13g2_fill_1 FILLER_44_217 ();
 sg13g2_fill_2 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_350 ();
 sg13g2_fill_2 FILLER_44_477 ();
 sg13g2_fill_1 FILLER_44_507 ();
 sg13g2_fill_2 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_541 ();
 sg13g2_fill_2 FILLER_44_552 ();
 sg13g2_decap_4 FILLER_44_591 ();
 sg13g2_fill_2 FILLER_44_618 ();
 sg13g2_decap_4 FILLER_44_648 ();
 sg13g2_fill_1 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_fill_1 FILLER_44_705 ();
 sg13g2_decap_4 FILLER_44_730 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_fill_2 FILLER_44_765 ();
 sg13g2_fill_1 FILLER_44_776 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_2 FILLER_44_870 ();
 sg13g2_fill_1 FILLER_44_872 ();
 sg13g2_fill_2 FILLER_44_878 ();
 sg13g2_decap_4 FILLER_44_886 ();
 sg13g2_fill_1 FILLER_44_890 ();
 sg13g2_fill_2 FILLER_44_958 ();
 sg13g2_fill_2 FILLER_44_978 ();
 sg13g2_fill_1 FILLER_44_980 ();
 sg13g2_fill_2 FILLER_44_1020 ();
 sg13g2_fill_1 FILLER_44_1022 ();
 sg13g2_fill_2 FILLER_44_1057 ();
 sg13g2_fill_1 FILLER_44_1085 ();
 sg13g2_fill_2 FILLER_44_1095 ();
 sg13g2_fill_1 FILLER_44_1107 ();
 sg13g2_fill_2 FILLER_44_1113 ();
 sg13g2_fill_1 FILLER_44_1119 ();
 sg13g2_fill_1 FILLER_44_1129 ();
 sg13g2_fill_2 FILLER_44_1175 ();
 sg13g2_fill_2 FILLER_44_1222 ();
 sg13g2_fill_1 FILLER_44_1224 ();
 sg13g2_fill_1 FILLER_44_1253 ();
 sg13g2_fill_1 FILLER_44_1288 ();
 sg13g2_fill_2 FILLER_44_1339 ();
 sg13g2_decap_4 FILLER_44_1370 ();
 sg13g2_fill_2 FILLER_44_1392 ();
 sg13g2_fill_1 FILLER_44_1532 ();
 sg13g2_decap_4 FILLER_44_1553 ();
 sg13g2_decap_4 FILLER_44_1572 ();
 sg13g2_fill_1 FILLER_44_1576 ();
 sg13g2_decap_4 FILLER_44_1582 ();
 sg13g2_fill_2 FILLER_44_1586 ();
 sg13g2_decap_4 FILLER_44_1594 ();
 sg13g2_fill_1 FILLER_44_1598 ();
 sg13g2_decap_8 FILLER_44_1610 ();
 sg13g2_fill_2 FILLER_44_1617 ();
 sg13g2_fill_1 FILLER_44_1619 ();
 sg13g2_decap_4 FILLER_44_1624 ();
 sg13g2_fill_2 FILLER_44_1628 ();
 sg13g2_fill_2 FILLER_44_1633 ();
 sg13g2_decap_8 FILLER_44_1639 ();
 sg13g2_decap_8 FILLER_44_1646 ();
 sg13g2_decap_8 FILLER_44_1653 ();
 sg13g2_decap_8 FILLER_44_1660 ();
 sg13g2_decap_8 FILLER_44_1667 ();
 sg13g2_decap_8 FILLER_44_1674 ();
 sg13g2_fill_2 FILLER_44_1681 ();
 sg13g2_fill_1 FILLER_44_1683 ();
 sg13g2_decap_8 FILLER_44_1689 ();
 sg13g2_fill_2 FILLER_44_1696 ();
 sg13g2_decap_4 FILLER_44_1702 ();
 sg13g2_fill_2 FILLER_44_1706 ();
 sg13g2_decap_8 FILLER_44_1712 ();
 sg13g2_fill_1 FILLER_44_1719 ();
 sg13g2_decap_4 FILLER_44_1748 ();
 sg13g2_fill_2 FILLER_44_1752 ();
 sg13g2_decap_4 FILLER_44_1767 ();
 sg13g2_fill_1 FILLER_44_1771 ();
 sg13g2_fill_2 FILLER_44_1807 ();
 sg13g2_decap_4 FILLER_44_1822 ();
 sg13g2_decap_8 FILLER_44_1836 ();
 sg13g2_fill_2 FILLER_44_1843 ();
 sg13g2_fill_2 FILLER_44_1849 ();
 sg13g2_fill_2 FILLER_44_1864 ();
 sg13g2_fill_1 FILLER_44_1866 ();
 sg13g2_fill_2 FILLER_44_1917 ();
 sg13g2_fill_1 FILLER_44_1919 ();
 sg13g2_decap_8 FILLER_44_1942 ();
 sg13g2_fill_2 FILLER_44_1949 ();
 sg13g2_fill_1 FILLER_44_1951 ();
 sg13g2_fill_1 FILLER_44_1965 ();
 sg13g2_fill_1 FILLER_44_1980 ();
 sg13g2_decap_8 FILLER_44_1998 ();
 sg13g2_decap_8 FILLER_44_2005 ();
 sg13g2_fill_2 FILLER_44_2012 ();
 sg13g2_fill_1 FILLER_44_2027 ();
 sg13g2_decap_4 FILLER_44_2058 ();
 sg13g2_fill_1 FILLER_44_2062 ();
 sg13g2_fill_1 FILLER_44_2083 ();
 sg13g2_fill_1 FILLER_44_2108 ();
 sg13g2_fill_2 FILLER_44_2113 ();
 sg13g2_fill_1 FILLER_44_2115 ();
 sg13g2_fill_2 FILLER_44_2185 ();
 sg13g2_fill_2 FILLER_44_2192 ();
 sg13g2_fill_2 FILLER_44_2259 ();
 sg13g2_fill_1 FILLER_44_2304 ();
 sg13g2_fill_2 FILLER_44_2309 ();
 sg13g2_fill_2 FILLER_44_2363 ();
 sg13g2_fill_2 FILLER_44_2387 ();
 sg13g2_fill_1 FILLER_44_2389 ();
 sg13g2_fill_2 FILLER_44_2417 ();
 sg13g2_fill_1 FILLER_44_2419 ();
 sg13g2_fill_1 FILLER_44_2452 ();
 sg13g2_fill_1 FILLER_44_2545 ();
 sg13g2_fill_1 FILLER_44_2596 ();
 sg13g2_fill_1 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2666 ();
 sg13g2_fill_1 FILLER_44_2673 ();
 sg13g2_decap_8 FILLER_45_83 ();
 sg13g2_decap_4 FILLER_45_90 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_135 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_338 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_2 FILLER_45_371 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_411 ();
 sg13g2_fill_1 FILLER_45_428 ();
 sg13g2_fill_1 FILLER_45_524 ();
 sg13g2_decap_4 FILLER_45_562 ();
 sg13g2_fill_2 FILLER_45_587 ();
 sg13g2_fill_1 FILLER_45_589 ();
 sg13g2_fill_2 FILLER_45_595 ();
 sg13g2_decap_4 FILLER_45_607 ();
 sg13g2_fill_1 FILLER_45_611 ();
 sg13g2_fill_2 FILLER_45_625 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_1 FILLER_45_665 ();
 sg13g2_decap_4 FILLER_45_697 ();
 sg13g2_fill_1 FILLER_45_701 ();
 sg13g2_fill_1 FILLER_45_750 ();
 sg13g2_fill_1 FILLER_45_778 ();
 sg13g2_fill_1 FILLER_45_786 ();
 sg13g2_fill_1 FILLER_45_805 ();
 sg13g2_fill_2 FILLER_45_821 ();
 sg13g2_fill_1 FILLER_45_823 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_873 ();
 sg13g2_decap_8 FILLER_45_880 ();
 sg13g2_fill_2 FILLER_45_942 ();
 sg13g2_fill_2 FILLER_45_1007 ();
 sg13g2_fill_1 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1025 ();
 sg13g2_fill_1 FILLER_45_1027 ();
 sg13g2_fill_2 FILLER_45_1056 ();
 sg13g2_fill_1 FILLER_45_1061 ();
 sg13g2_fill_1 FILLER_45_1066 ();
 sg13g2_fill_1 FILLER_45_1127 ();
 sg13g2_fill_1 FILLER_45_1179 ();
 sg13g2_fill_1 FILLER_45_1234 ();
 sg13g2_fill_2 FILLER_45_1290 ();
 sg13g2_fill_2 FILLER_45_1337 ();
 sg13g2_fill_2 FILLER_45_1347 ();
 sg13g2_fill_2 FILLER_45_1371 ();
 sg13g2_decap_8 FILLER_45_1420 ();
 sg13g2_decap_8 FILLER_45_1427 ();
 sg13g2_decap_8 FILLER_45_1434 ();
 sg13g2_decap_8 FILLER_45_1441 ();
 sg13g2_fill_1 FILLER_45_1481 ();
 sg13g2_fill_2 FILLER_45_1515 ();
 sg13g2_fill_1 FILLER_45_1517 ();
 sg13g2_fill_1 FILLER_45_1555 ();
 sg13g2_decap_8 FILLER_45_1581 ();
 sg13g2_decap_8 FILLER_45_1588 ();
 sg13g2_decap_8 FILLER_45_1595 ();
 sg13g2_fill_2 FILLER_45_1602 ();
 sg13g2_fill_2 FILLER_45_1614 ();
 sg13g2_decap_8 FILLER_45_1631 ();
 sg13g2_decap_8 FILLER_45_1638 ();
 sg13g2_decap_8 FILLER_45_1645 ();
 sg13g2_decap_8 FILLER_45_1652 ();
 sg13g2_decap_4 FILLER_45_1659 ();
 sg13g2_fill_2 FILLER_45_1663 ();
 sg13g2_fill_2 FILLER_45_1670 ();
 sg13g2_fill_2 FILLER_45_1680 ();
 sg13g2_fill_1 FILLER_45_1682 ();
 sg13g2_decap_8 FILLER_45_1697 ();
 sg13g2_decap_8 FILLER_45_1704 ();
 sg13g2_decap_4 FILLER_45_1711 ();
 sg13g2_fill_2 FILLER_45_1715 ();
 sg13g2_decap_8 FILLER_45_1764 ();
 sg13g2_fill_1 FILLER_45_1771 ();
 sg13g2_fill_2 FILLER_45_1825 ();
 sg13g2_decap_4 FILLER_45_1837 ();
 sg13g2_fill_2 FILLER_45_1841 ();
 sg13g2_fill_1 FILLER_45_1848 ();
 sg13g2_fill_2 FILLER_45_1853 ();
 sg13g2_fill_2 FILLER_45_1901 ();
 sg13g2_fill_1 FILLER_45_1916 ();
 sg13g2_fill_2 FILLER_45_1996 ();
 sg13g2_fill_1 FILLER_45_1998 ();
 sg13g2_fill_2 FILLER_45_2004 ();
 sg13g2_decap_4 FILLER_45_2010 ();
 sg13g2_fill_2 FILLER_45_2014 ();
 sg13g2_fill_2 FILLER_45_2055 ();
 sg13g2_fill_1 FILLER_45_2057 ();
 sg13g2_decap_4 FILLER_45_2071 ();
 sg13g2_fill_1 FILLER_45_2094 ();
 sg13g2_fill_1 FILLER_45_2114 ();
 sg13g2_fill_2 FILLER_45_2125 ();
 sg13g2_fill_1 FILLER_45_2179 ();
 sg13g2_fill_1 FILLER_45_2214 ();
 sg13g2_decap_4 FILLER_45_2270 ();
 sg13g2_fill_1 FILLER_45_2274 ();
 sg13g2_decap_8 FILLER_45_2288 ();
 sg13g2_decap_4 FILLER_45_2295 ();
 sg13g2_fill_1 FILLER_45_2299 ();
 sg13g2_fill_2 FILLER_45_2359 ();
 sg13g2_fill_1 FILLER_45_2361 ();
 sg13g2_fill_1 FILLER_45_2379 ();
 sg13g2_fill_2 FILLER_45_2399 ();
 sg13g2_fill_1 FILLER_45_2485 ();
 sg13g2_decap_4 FILLER_45_2504 ();
 sg13g2_fill_2 FILLER_45_2508 ();
 sg13g2_fill_1 FILLER_45_2581 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_29 ();
 sg13g2_fill_2 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_fill_1 FILLER_46_158 ();
 sg13g2_fill_2 FILLER_46_186 ();
 sg13g2_fill_1 FILLER_46_188 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_302 ();
 sg13g2_fill_1 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_563 ();
 sg13g2_fill_2 FILLER_46_605 ();
 sg13g2_decap_4 FILLER_46_665 ();
 sg13g2_fill_2 FILLER_46_682 ();
 sg13g2_fill_1 FILLER_46_749 ();
 sg13g2_fill_2 FILLER_46_759 ();
 sg13g2_fill_2 FILLER_46_770 ();
 sg13g2_fill_1 FILLER_46_786 ();
 sg13g2_fill_1 FILLER_46_796 ();
 sg13g2_fill_1 FILLER_46_823 ();
 sg13g2_fill_1 FILLER_46_883 ();
 sg13g2_decap_8 FILLER_46_890 ();
 sg13g2_fill_2 FILLER_46_897 ();
 sg13g2_fill_2 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_921 ();
 sg13g2_fill_2 FILLER_46_941 ();
 sg13g2_fill_2 FILLER_46_956 ();
 sg13g2_fill_2 FILLER_46_977 ();
 sg13g2_fill_1 FILLER_46_987 ();
 sg13g2_fill_2 FILLER_46_1022 ();
 sg13g2_decap_4 FILLER_46_1054 ();
 sg13g2_fill_1 FILLER_46_1085 ();
 sg13g2_decap_8 FILLER_46_1141 ();
 sg13g2_fill_2 FILLER_46_1148 ();
 sg13g2_fill_1 FILLER_46_1150 ();
 sg13g2_fill_2 FILLER_46_1174 ();
 sg13g2_fill_2 FILLER_46_1242 ();
 sg13g2_fill_1 FILLER_46_1244 ();
 sg13g2_fill_2 FILLER_46_1286 ();
 sg13g2_fill_1 FILLER_46_1346 ();
 sg13g2_fill_1 FILLER_46_1354 ();
 sg13g2_fill_2 FILLER_46_1370 ();
 sg13g2_fill_1 FILLER_46_1372 ();
 sg13g2_fill_2 FILLER_46_1389 ();
 sg13g2_fill_1 FILLER_46_1391 ();
 sg13g2_fill_2 FILLER_46_1421 ();
 sg13g2_fill_1 FILLER_46_1423 ();
 sg13g2_decap_8 FILLER_46_1427 ();
 sg13g2_decap_8 FILLER_46_1434 ();
 sg13g2_fill_2 FILLER_46_1520 ();
 sg13g2_fill_1 FILLER_46_1538 ();
 sg13g2_fill_2 FILLER_46_1552 ();
 sg13g2_fill_1 FILLER_46_1554 ();
 sg13g2_decap_8 FILLER_46_1563 ();
 sg13g2_decap_4 FILLER_46_1570 ();
 sg13g2_fill_1 FILLER_46_1574 ();
 sg13g2_decap_8 FILLER_46_1581 ();
 sg13g2_decap_4 FILLER_46_1588 ();
 sg13g2_fill_2 FILLER_46_1592 ();
 sg13g2_decap_8 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1605 ();
 sg13g2_fill_1 FILLER_46_1612 ();
 sg13g2_decap_4 FILLER_46_1618 ();
 sg13g2_fill_2 FILLER_46_1622 ();
 sg13g2_fill_1 FILLER_46_1629 ();
 sg13g2_decap_4 FILLER_46_1645 ();
 sg13g2_fill_2 FILLER_46_1649 ();
 sg13g2_fill_2 FILLER_46_1670 ();
 sg13g2_fill_2 FILLER_46_1677 ();
 sg13g2_decap_8 FILLER_46_1692 ();
 sg13g2_fill_1 FILLER_46_1699 ();
 sg13g2_decap_4 FILLER_46_1714 ();
 sg13g2_fill_1 FILLER_46_1718 ();
 sg13g2_fill_1 FILLER_46_1739 ();
 sg13g2_decap_8 FILLER_46_1765 ();
 sg13g2_decap_8 FILLER_46_1772 ();
 sg13g2_decap_4 FILLER_46_1779 ();
 sg13g2_fill_1 FILLER_46_1783 ();
 sg13g2_fill_1 FILLER_46_1807 ();
 sg13g2_decap_4 FILLER_46_1858 ();
 sg13g2_fill_2 FILLER_46_1875 ();
 sg13g2_fill_2 FILLER_46_1882 ();
 sg13g2_fill_2 FILLER_46_1898 ();
 sg13g2_fill_1 FILLER_46_1900 ();
 sg13g2_decap_8 FILLER_46_1941 ();
 sg13g2_fill_1 FILLER_46_1948 ();
 sg13g2_fill_2 FILLER_46_1990 ();
 sg13g2_fill_1 FILLER_46_1992 ();
 sg13g2_fill_1 FILLER_46_2043 ();
 sg13g2_fill_2 FILLER_46_2103 ();
 sg13g2_fill_1 FILLER_46_2105 ();
 sg13g2_fill_2 FILLER_46_2145 ();
 sg13g2_fill_2 FILLER_46_2211 ();
 sg13g2_fill_1 FILLER_46_2213 ();
 sg13g2_fill_2 FILLER_46_2241 ();
 sg13g2_fill_2 FILLER_46_2255 ();
 sg13g2_fill_1 FILLER_46_2257 ();
 sg13g2_fill_2 FILLER_46_2297 ();
 sg13g2_fill_1 FILLER_46_2299 ();
 sg13g2_fill_1 FILLER_46_2313 ();
 sg13g2_fill_1 FILLER_46_2327 ();
 sg13g2_fill_2 FILLER_46_2333 ();
 sg13g2_fill_1 FILLER_46_2384 ();
 sg13g2_fill_1 FILLER_46_2394 ();
 sg13g2_fill_2 FILLER_46_2452 ();
 sg13g2_fill_1 FILLER_46_2519 ();
 sg13g2_fill_1 FILLER_46_2528 ();
 sg13g2_fill_2 FILLER_46_2538 ();
 sg13g2_fill_2 FILLER_46_2652 ();
 sg13g2_fill_1 FILLER_46_2654 ();
 sg13g2_fill_1 FILLER_46_2673 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_fill_2 FILLER_47_48 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_136 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_decap_4 FILLER_47_184 ();
 sg13g2_fill_1 FILLER_47_188 ();
 sg13g2_fill_2 FILLER_47_193 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_fill_2 FILLER_47_226 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_fill_2 FILLER_47_501 ();
 sg13g2_fill_1 FILLER_47_555 ();
 sg13g2_fill_1 FILLER_47_581 ();
 sg13g2_fill_2 FILLER_47_588 ();
 sg13g2_fill_1 FILLER_47_618 ();
 sg13g2_fill_1 FILLER_47_669 ();
 sg13g2_fill_2 FILLER_47_675 ();
 sg13g2_fill_2 FILLER_47_691 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_fill_1 FILLER_47_699 ();
 sg13g2_fill_2 FILLER_47_709 ();
 sg13g2_fill_2 FILLER_47_783 ();
 sg13g2_fill_1 FILLER_47_804 ();
 sg13g2_decap_4 FILLER_47_906 ();
 sg13g2_fill_1 FILLER_47_910 ();
 sg13g2_fill_1 FILLER_47_938 ();
 sg13g2_fill_2 FILLER_47_985 ();
 sg13g2_fill_2 FILLER_47_1014 ();
 sg13g2_fill_1 FILLER_47_1016 ();
 sg13g2_fill_2 FILLER_47_1030 ();
 sg13g2_fill_1 FILLER_47_1032 ();
 sg13g2_fill_1 FILLER_47_1042 ();
 sg13g2_decap_4 FILLER_47_1057 ();
 sg13g2_fill_1 FILLER_47_1089 ();
 sg13g2_decap_4 FILLER_47_1102 ();
 sg13g2_fill_1 FILLER_47_1106 ();
 sg13g2_decap_4 FILLER_47_1125 ();
 sg13g2_decap_4 FILLER_47_1155 ();
 sg13g2_fill_2 FILLER_47_1224 ();
 sg13g2_decap_4 FILLER_47_1277 ();
 sg13g2_fill_1 FILLER_47_1394 ();
 sg13g2_fill_2 FILLER_47_1487 ();
 sg13g2_fill_1 FILLER_47_1489 ();
 sg13g2_fill_1 FILLER_47_1515 ();
 sg13g2_decap_8 FILLER_47_1549 ();
 sg13g2_decap_4 FILLER_47_1556 ();
 sg13g2_fill_1 FILLER_47_1560 ();
 sg13g2_decap_8 FILLER_47_1572 ();
 sg13g2_decap_4 FILLER_47_1579 ();
 sg13g2_decap_4 FILLER_47_1591 ();
 sg13g2_fill_2 FILLER_47_1605 ();
 sg13g2_fill_1 FILLER_47_1607 ();
 sg13g2_fill_2 FILLER_47_1618 ();
 sg13g2_fill_1 FILLER_47_1620 ();
 sg13g2_fill_2 FILLER_47_1625 ();
 sg13g2_fill_1 FILLER_47_1627 ();
 sg13g2_decap_8 FILLER_47_1633 ();
 sg13g2_decap_8 FILLER_47_1640 ();
 sg13g2_decap_8 FILLER_47_1647 ();
 sg13g2_fill_1 FILLER_47_1654 ();
 sg13g2_fill_1 FILLER_47_1660 ();
 sg13g2_decap_8 FILLER_47_1677 ();
 sg13g2_decap_4 FILLER_47_1684 ();
 sg13g2_fill_1 FILLER_47_1688 ();
 sg13g2_fill_1 FILLER_47_1699 ();
 sg13g2_decap_8 FILLER_47_1717 ();
 sg13g2_decap_8 FILLER_47_1724 ();
 sg13g2_decap_8 FILLER_47_1735 ();
 sg13g2_fill_1 FILLER_47_1742 ();
 sg13g2_decap_8 FILLER_47_1765 ();
 sg13g2_decap_8 FILLER_47_1772 ();
 sg13g2_fill_2 FILLER_47_1779 ();
 sg13g2_fill_1 FILLER_47_1781 ();
 sg13g2_fill_1 FILLER_47_1787 ();
 sg13g2_decap_4 FILLER_47_1798 ();
 sg13g2_fill_1 FILLER_47_1812 ();
 sg13g2_fill_1 FILLER_47_1826 ();
 sg13g2_decap_8 FILLER_47_1872 ();
 sg13g2_fill_2 FILLER_47_1879 ();
 sg13g2_decap_4 FILLER_47_1890 ();
 sg13g2_fill_2 FILLER_47_1948 ();
 sg13g2_fill_1 FILLER_47_1950 ();
 sg13g2_fill_1 FILLER_47_1996 ();
 sg13g2_fill_2 FILLER_47_2034 ();
 sg13g2_fill_1 FILLER_47_2036 ();
 sg13g2_fill_2 FILLER_47_2050 ();
 sg13g2_fill_2 FILLER_47_2082 ();
 sg13g2_fill_1 FILLER_47_2136 ();
 sg13g2_fill_1 FILLER_47_2206 ();
 sg13g2_fill_1 FILLER_47_2265 ();
 sg13g2_fill_2 FILLER_47_2453 ();
 sg13g2_fill_1 FILLER_47_2479 ();
 sg13g2_fill_1 FILLER_47_2512 ();
 sg13g2_decap_4 FILLER_47_2535 ();
 sg13g2_fill_1 FILLER_47_2539 ();
 sg13g2_fill_2 FILLER_47_2550 ();
 sg13g2_decap_4 FILLER_47_2563 ();
 sg13g2_fill_1 FILLER_47_2612 ();
 sg13g2_fill_2 FILLER_47_2618 ();
 sg13g2_decap_4 FILLER_47_2668 ();
 sg13g2_fill_2 FILLER_47_2672 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_1 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_fill_2 FILLER_48_174 ();
 sg13g2_decap_4 FILLER_48_184 ();
 sg13g2_fill_1 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_fill_2 FILLER_48_356 ();
 sg13g2_fill_1 FILLER_48_403 ();
 sg13g2_fill_1 FILLER_48_506 ();
 sg13g2_fill_1 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_550 ();
 sg13g2_fill_1 FILLER_48_557 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_583 ();
 sg13g2_fill_1 FILLER_48_585 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_decap_4 FILLER_48_607 ();
 sg13g2_decap_4 FILLER_48_624 ();
 sg13g2_fill_2 FILLER_48_638 ();
 sg13g2_fill_1 FILLER_48_640 ();
 sg13g2_fill_1 FILLER_48_647 ();
 sg13g2_decap_8 FILLER_48_657 ();
 sg13g2_decap_8 FILLER_48_664 ();
 sg13g2_decap_4 FILLER_48_671 ();
 sg13g2_decap_4 FILLER_48_679 ();
 sg13g2_fill_1 FILLER_48_683 ();
 sg13g2_fill_2 FILLER_48_715 ();
 sg13g2_decap_4 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_846 ();
 sg13g2_fill_2 FILLER_48_908 ();
 sg13g2_fill_1 FILLER_48_910 ();
 sg13g2_fill_2 FILLER_48_933 ();
 sg13g2_fill_1 FILLER_48_935 ();
 sg13g2_fill_2 FILLER_48_967 ();
 sg13g2_fill_1 FILLER_48_969 ();
 sg13g2_fill_1 FILLER_48_991 ();
 sg13g2_fill_2 FILLER_48_1016 ();
 sg13g2_fill_1 FILLER_48_1061 ();
 sg13g2_fill_2 FILLER_48_1074 ();
 sg13g2_decap_4 FILLER_48_1085 ();
 sg13g2_decap_4 FILLER_48_1099 ();
 sg13g2_fill_2 FILLER_48_1103 ();
 sg13g2_decap_8 FILLER_48_1122 ();
 sg13g2_decap_4 FILLER_48_1134 ();
 sg13g2_fill_1 FILLER_48_1138 ();
 sg13g2_decap_4 FILLER_48_1152 ();
 sg13g2_fill_2 FILLER_48_1224 ();
 sg13g2_fill_2 FILLER_48_1238 ();
 sg13g2_decap_8 FILLER_48_1243 ();
 sg13g2_decap_4 FILLER_48_1250 ();
 sg13g2_fill_1 FILLER_48_1254 ();
 sg13g2_fill_2 FILLER_48_1290 ();
 sg13g2_fill_2 FILLER_48_1359 ();
 sg13g2_fill_2 FILLER_48_1376 ();
 sg13g2_fill_1 FILLER_48_1413 ();
 sg13g2_fill_1 FILLER_48_1420 ();
 sg13g2_fill_2 FILLER_48_1460 ();
 sg13g2_fill_1 FILLER_48_1462 ();
 sg13g2_fill_2 FILLER_48_1469 ();
 sg13g2_fill_1 FILLER_48_1471 ();
 sg13g2_fill_2 FILLER_48_1509 ();
 sg13g2_fill_2 FILLER_48_1516 ();
 sg13g2_fill_2 FILLER_48_1527 ();
 sg13g2_decap_4 FILLER_48_1557 ();
 sg13g2_fill_2 FILLER_48_1572 ();
 sg13g2_fill_1 FILLER_48_1574 ();
 sg13g2_fill_1 FILLER_48_1589 ();
 sg13g2_decap_4 FILLER_48_1602 ();
 sg13g2_fill_2 FILLER_48_1606 ();
 sg13g2_decap_8 FILLER_48_1632 ();
 sg13g2_decap_8 FILLER_48_1639 ();
 sg13g2_fill_1 FILLER_48_1657 ();
 sg13g2_decap_8 FILLER_48_1671 ();
 sg13g2_decap_8 FILLER_48_1678 ();
 sg13g2_fill_2 FILLER_48_1693 ();
 sg13g2_fill_1 FILLER_48_1695 ();
 sg13g2_decap_8 FILLER_48_1710 ();
 sg13g2_fill_2 FILLER_48_1717 ();
 sg13g2_fill_1 FILLER_48_1719 ();
 sg13g2_fill_2 FILLER_48_1744 ();
 sg13g2_decap_8 FILLER_48_1755 ();
 sg13g2_decap_8 FILLER_48_1762 ();
 sg13g2_decap_8 FILLER_48_1769 ();
 sg13g2_fill_2 FILLER_48_1776 ();
 sg13g2_fill_1 FILLER_48_1778 ();
 sg13g2_fill_2 FILLER_48_1832 ();
 sg13g2_fill_2 FILLER_48_1847 ();
 sg13g2_fill_1 FILLER_48_1849 ();
 sg13g2_fill_1 FILLER_48_1863 ();
 sg13g2_decap_4 FILLER_48_1882 ();
 sg13g2_fill_2 FILLER_48_1905 ();
 sg13g2_fill_1 FILLER_48_1957 ();
 sg13g2_fill_2 FILLER_48_2170 ();
 sg13g2_fill_1 FILLER_48_2172 ();
 sg13g2_fill_1 FILLER_48_2245 ();
 sg13g2_fill_1 FILLER_48_2280 ();
 sg13g2_fill_1 FILLER_48_2379 ();
 sg13g2_fill_1 FILLER_48_2411 ();
 sg13g2_fill_1 FILLER_48_2433 ();
 sg13g2_fill_2 FILLER_48_2470 ();
 sg13g2_fill_1 FILLER_48_2472 ();
 sg13g2_fill_2 FILLER_48_2501 ();
 sg13g2_fill_1 FILLER_48_2539 ();
 sg13g2_decap_4 FILLER_48_2556 ();
 sg13g2_decap_4 FILLER_48_2587 ();
 sg13g2_fill_2 FILLER_48_2604 ();
 sg13g2_decap_4 FILLER_48_2669 ();
 sg13g2_fill_1 FILLER_48_2673 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_fill_2 FILLER_49_143 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_fill_2 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_445 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_decap_8 FILLER_49_547 ();
 sg13g2_decap_8 FILLER_49_554 ();
 sg13g2_decap_8 FILLER_49_566 ();
 sg13g2_decap_8 FILLER_49_573 ();
 sg13g2_fill_1 FILLER_49_580 ();
 sg13g2_fill_2 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_640 ();
 sg13g2_decap_8 FILLER_49_652 ();
 sg13g2_decap_8 FILLER_49_659 ();
 sg13g2_decap_8 FILLER_49_666 ();
 sg13g2_fill_2 FILLER_49_673 ();
 sg13g2_fill_2 FILLER_49_712 ();
 sg13g2_fill_1 FILLER_49_723 ();
 sg13g2_fill_1 FILLER_49_739 ();
 sg13g2_fill_1 FILLER_49_810 ();
 sg13g2_fill_1 FILLER_49_838 ();
 sg13g2_fill_2 FILLER_49_880 ();
 sg13g2_fill_2 FILLER_49_926 ();
 sg13g2_fill_2 FILLER_49_963 ();
 sg13g2_fill_1 FILLER_49_965 ();
 sg13g2_fill_1 FILLER_49_1030 ();
 sg13g2_fill_2 FILLER_49_1062 ();
 sg13g2_fill_1 FILLER_49_1064 ();
 sg13g2_fill_1 FILLER_49_1078 ();
 sg13g2_fill_2 FILLER_49_1110 ();
 sg13g2_fill_1 FILLER_49_1112 ();
 sg13g2_fill_1 FILLER_49_1129 ();
 sg13g2_fill_2 FILLER_49_1139 ();
 sg13g2_fill_2 FILLER_49_1168 ();
 sg13g2_fill_1 FILLER_49_1170 ();
 sg13g2_fill_2 FILLER_49_1179 ();
 sg13g2_fill_1 FILLER_49_1181 ();
 sg13g2_fill_2 FILLER_49_1236 ();
 sg13g2_decap_4 FILLER_49_1290 ();
 sg13g2_fill_1 FILLER_49_1294 ();
 sg13g2_fill_1 FILLER_49_1347 ();
 sg13g2_fill_2 FILLER_49_1366 ();
 sg13g2_fill_2 FILLER_49_1382 ();
 sg13g2_fill_1 FILLER_49_1401 ();
 sg13g2_fill_2 FILLER_49_1473 ();
 sg13g2_fill_2 FILLER_49_1481 ();
 sg13g2_fill_1 FILLER_49_1483 ();
 sg13g2_decap_8 FILLER_49_1512 ();
 sg13g2_decap_4 FILLER_49_1519 ();
 sg13g2_fill_1 FILLER_49_1531 ();
 sg13g2_fill_2 FILLER_49_1537 ();
 sg13g2_decap_4 FILLER_49_1549 ();
 sg13g2_fill_1 FILLER_49_1566 ();
 sg13g2_fill_2 FILLER_49_1573 ();
 sg13g2_decap_4 FILLER_49_1579 ();
 sg13g2_fill_1 FILLER_49_1586 ();
 sg13g2_decap_4 FILLER_49_1601 ();
 sg13g2_fill_2 FILLER_49_1623 ();
 sg13g2_decap_8 FILLER_49_1630 ();
 sg13g2_decap_8 FILLER_49_1637 ();
 sg13g2_decap_8 FILLER_49_1644 ();
 sg13g2_decap_8 FILLER_49_1651 ();
 sg13g2_decap_8 FILLER_49_1658 ();
 sg13g2_fill_1 FILLER_49_1665 ();
 sg13g2_decap_8 FILLER_49_1669 ();
 sg13g2_decap_8 FILLER_49_1676 ();
 sg13g2_fill_2 FILLER_49_1683 ();
 sg13g2_fill_2 FILLER_49_1721 ();
 sg13g2_decap_8 FILLER_49_1765 ();
 sg13g2_fill_1 FILLER_49_1772 ();
 sg13g2_fill_2 FILLER_49_1804 ();
 sg13g2_fill_1 FILLER_49_1806 ();
 sg13g2_decap_4 FILLER_49_1839 ();
 sg13g2_fill_2 FILLER_49_1936 ();
 sg13g2_fill_2 FILLER_49_1987 ();
 sg13g2_fill_1 FILLER_49_1989 ();
 sg13g2_fill_1 FILLER_49_2008 ();
 sg13g2_fill_2 FILLER_49_2037 ();
 sg13g2_fill_1 FILLER_49_2039 ();
 sg13g2_decap_8 FILLER_49_2066 ();
 sg13g2_fill_2 FILLER_49_2073 ();
 sg13g2_fill_1 FILLER_49_2075 ();
 sg13g2_fill_1 FILLER_49_2103 ();
 sg13g2_fill_2 FILLER_49_2163 ();
 sg13g2_fill_2 FILLER_49_2204 ();
 sg13g2_fill_2 FILLER_49_2225 ();
 sg13g2_fill_1 FILLER_49_2242 ();
 sg13g2_fill_2 FILLER_49_2397 ();
 sg13g2_fill_2 FILLER_49_2418 ();
 sg13g2_fill_1 FILLER_49_2447 ();
 sg13g2_fill_1 FILLER_49_2461 ();
 sg13g2_fill_1 FILLER_49_2480 ();
 sg13g2_fill_2 FILLER_49_2508 ();
 sg13g2_fill_1 FILLER_49_2510 ();
 sg13g2_fill_2 FILLER_49_2597 ();
 sg13g2_fill_1 FILLER_49_2599 ();
 sg13g2_decap_4 FILLER_49_2626 ();
 sg13g2_fill_2 FILLER_49_2630 ();
 sg13g2_decap_4 FILLER_49_2668 ();
 sg13g2_fill_2 FILLER_49_2672 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_61 ();
 sg13g2_fill_1 FILLER_50_68 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_fill_2 FILLER_50_257 ();
 sg13g2_fill_1 FILLER_50_259 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_379 ();
 sg13g2_fill_2 FILLER_50_399 ();
 sg13g2_fill_2 FILLER_50_484 ();
 sg13g2_fill_1 FILLER_50_499 ();
 sg13g2_fill_1 FILLER_50_537 ();
 sg13g2_fill_1 FILLER_50_579 ();
 sg13g2_fill_2 FILLER_50_606 ();
 sg13g2_fill_1 FILLER_50_608 ();
 sg13g2_decap_8 FILLER_50_632 ();
 sg13g2_decap_4 FILLER_50_639 ();
 sg13g2_decap_4 FILLER_50_659 ();
 sg13g2_fill_2 FILLER_50_741 ();
 sg13g2_fill_1 FILLER_50_756 ();
 sg13g2_fill_2 FILLER_50_845 ();
 sg13g2_fill_1 FILLER_50_939 ();
 sg13g2_fill_1 FILLER_50_955 ();
 sg13g2_fill_1 FILLER_50_1017 ();
 sg13g2_fill_2 FILLER_50_1036 ();
 sg13g2_fill_1 FILLER_50_1066 ();
 sg13g2_fill_2 FILLER_50_1139 ();
 sg13g2_fill_2 FILLER_50_1157 ();
 sg13g2_fill_1 FILLER_50_1159 ();
 sg13g2_fill_1 FILLER_50_1165 ();
 sg13g2_fill_2 FILLER_50_1182 ();
 sg13g2_fill_1 FILLER_50_1184 ();
 sg13g2_fill_1 FILLER_50_1190 ();
 sg13g2_fill_1 FILLER_50_1240 ();
 sg13g2_fill_1 FILLER_50_1289 ();
 sg13g2_decap_4 FILLER_50_1313 ();
 sg13g2_fill_2 FILLER_50_1344 ();
 sg13g2_fill_2 FILLER_50_1381 ();
 sg13g2_fill_1 FILLER_50_1383 ();
 sg13g2_fill_1 FILLER_50_1406 ();
 sg13g2_decap_8 FILLER_50_1513 ();
 sg13g2_fill_2 FILLER_50_1534 ();
 sg13g2_decap_4 FILLER_50_1559 ();
 sg13g2_fill_1 FILLER_50_1563 ();
 sg13g2_decap_4 FILLER_50_1591 ();
 sg13g2_fill_1 FILLER_50_1595 ();
 sg13g2_decap_8 FILLER_50_1601 ();
 sg13g2_decap_4 FILLER_50_1608 ();
 sg13g2_fill_2 FILLER_50_1612 ();
 sg13g2_decap_4 FILLER_50_1634 ();
 sg13g2_decap_8 FILLER_50_1643 ();
 sg13g2_decap_8 FILLER_50_1650 ();
 sg13g2_decap_4 FILLER_50_1657 ();
 sg13g2_decap_8 FILLER_50_1711 ();
 sg13g2_fill_2 FILLER_50_1718 ();
 sg13g2_fill_1 FILLER_50_1720 ();
 sg13g2_fill_2 FILLER_50_1739 ();
 sg13g2_fill_1 FILLER_50_1741 ();
 sg13g2_fill_2 FILLER_50_1772 ();
 sg13g2_fill_1 FILLER_50_1774 ();
 sg13g2_fill_1 FILLER_50_1785 ();
 sg13g2_fill_1 FILLER_50_1823 ();
 sg13g2_fill_2 FILLER_50_1909 ();
 sg13g2_fill_1 FILLER_50_1924 ();
 sg13g2_fill_1 FILLER_50_1983 ();
 sg13g2_fill_1 FILLER_50_1997 ();
 sg13g2_decap_8 FILLER_50_2033 ();
 sg13g2_fill_2 FILLER_50_2040 ();
 sg13g2_decap_8 FILLER_50_2063 ();
 sg13g2_fill_1 FILLER_50_2070 ();
 sg13g2_fill_2 FILLER_50_2084 ();
 sg13g2_fill_1 FILLER_50_2116 ();
 sg13g2_fill_1 FILLER_50_2193 ();
 sg13g2_fill_1 FILLER_50_2284 ();
 sg13g2_fill_1 FILLER_50_2345 ();
 sg13g2_fill_2 FILLER_50_2377 ();
 sg13g2_fill_1 FILLER_50_2392 ();
 sg13g2_fill_2 FILLER_50_2398 ();
 sg13g2_fill_1 FILLER_50_2400 ();
 sg13g2_fill_1 FILLER_50_2460 ();
 sg13g2_fill_2 FILLER_50_2564 ();
 sg13g2_fill_1 FILLER_50_2566 ();
 sg13g2_fill_2 FILLER_50_2579 ();
 sg13g2_fill_2 FILLER_50_2634 ();
 sg13g2_fill_1 FILLER_50_2650 ();
 sg13g2_fill_1 FILLER_50_2673 ();
 sg13g2_fill_1 FILLER_51_49 ();
 sg13g2_fill_2 FILLER_51_104 ();
 sg13g2_fill_1 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_125 ();
 sg13g2_fill_2 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_186 ();
 sg13g2_fill_2 FILLER_51_196 ();
 sg13g2_fill_1 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_212 ();
 sg13g2_fill_1 FILLER_51_264 ();
 sg13g2_fill_2 FILLER_51_371 ();
 sg13g2_fill_1 FILLER_51_405 ();
 sg13g2_fill_1 FILLER_51_411 ();
 sg13g2_fill_1 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_545 ();
 sg13g2_fill_1 FILLER_51_573 ();
 sg13g2_fill_2 FILLER_51_604 ();
 sg13g2_fill_1 FILLER_51_615 ();
 sg13g2_fill_1 FILLER_51_620 ();
 sg13g2_fill_1 FILLER_51_626 ();
 sg13g2_fill_1 FILLER_51_648 ();
 sg13g2_decap_8 FILLER_51_677 ();
 sg13g2_fill_2 FILLER_51_719 ();
 sg13g2_decap_4 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_894 ();
 sg13g2_decap_8 FILLER_51_901 ();
 sg13g2_decap_4 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_954 ();
 sg13g2_fill_2 FILLER_51_963 ();
 sg13g2_fill_2 FILLER_51_1016 ();
 sg13g2_fill_1 FILLER_51_1056 ();
 sg13g2_fill_1 FILLER_51_1088 ();
 sg13g2_fill_2 FILLER_51_1102 ();
 sg13g2_fill_1 FILLER_51_1104 ();
 sg13g2_decap_8 FILLER_51_1118 ();
 sg13g2_fill_2 FILLER_51_1125 ();
 sg13g2_fill_1 FILLER_51_1127 ();
 sg13g2_fill_2 FILLER_51_1167 ();
 sg13g2_fill_1 FILLER_51_1169 ();
 sg13g2_fill_1 FILLER_51_1211 ();
 sg13g2_fill_2 FILLER_51_1217 ();
 sg13g2_fill_2 FILLER_51_1225 ();
 sg13g2_decap_4 FILLER_51_1321 ();
 sg13g2_fill_1 FILLER_51_1325 ();
 sg13g2_fill_2 FILLER_51_1332 ();
 sg13g2_fill_2 FILLER_51_1389 ();
 sg13g2_fill_2 FILLER_51_1407 ();
 sg13g2_fill_2 FILLER_51_1451 ();
 sg13g2_fill_1 FILLER_51_1466 ();
 sg13g2_fill_2 FILLER_51_1482 ();
 sg13g2_decap_8 FILLER_51_1508 ();
 sg13g2_fill_2 FILLER_51_1515 ();
 sg13g2_fill_2 FILLER_51_1531 ();
 sg13g2_fill_1 FILLER_51_1533 ();
 sg13g2_decap_8 FILLER_51_1561 ();
 sg13g2_decap_8 FILLER_51_1568 ();
 sg13g2_decap_8 FILLER_51_1575 ();
 sg13g2_decap_4 FILLER_51_1582 ();
 sg13g2_fill_2 FILLER_51_1586 ();
 sg13g2_fill_2 FILLER_51_1597 ();
 sg13g2_fill_1 FILLER_51_1599 ();
 sg13g2_decap_8 FILLER_51_1650 ();
 sg13g2_fill_2 FILLER_51_1657 ();
 sg13g2_fill_1 FILLER_51_1659 ();
 sg13g2_decap_8 FILLER_51_1681 ();
 sg13g2_decap_8 FILLER_51_1692 ();
 sg13g2_decap_8 FILLER_51_1715 ();
 sg13g2_fill_2 FILLER_51_1722 ();
 sg13g2_fill_1 FILLER_51_1724 ();
 sg13g2_decap_8 FILLER_51_1766 ();
 sg13g2_fill_2 FILLER_51_1773 ();
 sg13g2_fill_2 FILLER_51_1815 ();
 sg13g2_fill_1 FILLER_51_1817 ();
 sg13g2_fill_1 FILLER_51_1849 ();
 sg13g2_decap_4 FILLER_51_1863 ();
 sg13g2_fill_2 FILLER_51_1909 ();
 sg13g2_fill_2 FILLER_51_1951 ();
 sg13g2_fill_1 FILLER_51_1993 ();
 sg13g2_decap_8 FILLER_51_2021 ();
 sg13g2_decap_8 FILLER_51_2028 ();
 sg13g2_decap_8 FILLER_51_2035 ();
 sg13g2_fill_1 FILLER_51_2042 ();
 sg13g2_fill_1 FILLER_51_2092 ();
 sg13g2_fill_2 FILLER_51_2120 ();
 sg13g2_fill_1 FILLER_51_2229 ();
 sg13g2_fill_1 FILLER_51_2253 ();
 sg13g2_fill_2 FILLER_51_2271 ();
 sg13g2_fill_2 FILLER_51_2326 ();
 sg13g2_fill_1 FILLER_51_2328 ();
 sg13g2_fill_1 FILLER_51_2349 ();
 sg13g2_fill_2 FILLER_51_2362 ();
 sg13g2_fill_2 FILLER_51_2382 ();
 sg13g2_fill_1 FILLER_51_2384 ();
 sg13g2_fill_2 FILLER_51_2403 ();
 sg13g2_fill_2 FILLER_51_2426 ();
 sg13g2_fill_2 FILLER_51_2447 ();
 sg13g2_fill_2 FILLER_51_2503 ();
 sg13g2_fill_1 FILLER_51_2505 ();
 sg13g2_fill_2 FILLER_51_2519 ();
 sg13g2_fill_1 FILLER_51_2521 ();
 sg13g2_fill_1 FILLER_51_2588 ();
 sg13g2_fill_2 FILLER_51_2671 ();
 sg13g2_fill_1 FILLER_51_2673 ();
 sg13g2_fill_2 FILLER_52_35 ();
 sg13g2_fill_1 FILLER_52_194 ();
 sg13g2_fill_2 FILLER_52_208 ();
 sg13g2_fill_1 FILLER_52_210 ();
 sg13g2_fill_2 FILLER_52_346 ();
 sg13g2_fill_1 FILLER_52_363 ();
 sg13g2_fill_2 FILLER_52_547 ();
 sg13g2_fill_1 FILLER_52_589 ();
 sg13g2_fill_2 FILLER_52_600 ();
 sg13g2_fill_1 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_fill_1 FILLER_52_653 ();
 sg13g2_fill_2 FILLER_52_658 ();
 sg13g2_fill_1 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_666 ();
 sg13g2_decap_8 FILLER_52_675 ();
 sg13g2_decap_4 FILLER_52_682 ();
 sg13g2_fill_2 FILLER_52_826 ();
 sg13g2_fill_1 FILLER_52_828 ();
 sg13g2_fill_1 FILLER_52_838 ();
 sg13g2_fill_1 FILLER_52_905 ();
 sg13g2_fill_1 FILLER_52_924 ();
 sg13g2_fill_2 FILLER_52_937 ();
 sg13g2_fill_2 FILLER_52_992 ();
 sg13g2_fill_2 FILLER_52_1011 ();
 sg13g2_fill_1 FILLER_52_1013 ();
 sg13g2_decap_4 FILLER_52_1022 ();
 sg13g2_fill_2 FILLER_52_1026 ();
 sg13g2_fill_1 FILLER_52_1033 ();
 sg13g2_fill_1 FILLER_52_1057 ();
 sg13g2_fill_1 FILLER_52_1089 ();
 sg13g2_fill_2 FILLER_52_1094 ();
 sg13g2_fill_1 FILLER_52_1096 ();
 sg13g2_decap_4 FILLER_52_1105 ();
 sg13g2_fill_2 FILLER_52_1109 ();
 sg13g2_decap_8 FILLER_52_1114 ();
 sg13g2_decap_8 FILLER_52_1121 ();
 sg13g2_fill_2 FILLER_52_1146 ();
 sg13g2_fill_2 FILLER_52_1173 ();
 sg13g2_fill_1 FILLER_52_1175 ();
 sg13g2_fill_1 FILLER_52_1193 ();
 sg13g2_fill_2 FILLER_52_1209 ();
 sg13g2_fill_1 FILLER_52_1224 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_decap_8 FILLER_52_1325 ();
 sg13g2_fill_2 FILLER_52_1332 ();
 sg13g2_fill_1 FILLER_52_1343 ();
 sg13g2_fill_2 FILLER_52_1362 ();
 sg13g2_fill_1 FILLER_52_1364 ();
 sg13g2_decap_4 FILLER_52_1383 ();
 sg13g2_fill_2 FILLER_52_1387 ();
 sg13g2_decap_4 FILLER_52_1398 ();
 sg13g2_fill_2 FILLER_52_1407 ();
 sg13g2_fill_2 FILLER_52_1427 ();
 sg13g2_fill_1 FILLER_52_1429 ();
 sg13g2_fill_2 FILLER_52_1504 ();
 sg13g2_fill_1 FILLER_52_1506 ();
 sg13g2_fill_1 FILLER_52_1515 ();
 sg13g2_fill_1 FILLER_52_1521 ();
 sg13g2_fill_1 FILLER_52_1535 ();
 sg13g2_decap_8 FILLER_52_1565 ();
 sg13g2_fill_2 FILLER_52_1572 ();
 sg13g2_decap_8 FILLER_52_1598 ();
 sg13g2_fill_1 FILLER_52_1605 ();
 sg13g2_decap_8 FILLER_52_1611 ();
 sg13g2_fill_2 FILLER_52_1618 ();
 sg13g2_fill_2 FILLER_52_1629 ();
 sg13g2_fill_1 FILLER_52_1631 ();
 sg13g2_decap_8 FILLER_52_1645 ();
 sg13g2_fill_2 FILLER_52_1652 ();
 sg13g2_fill_1 FILLER_52_1654 ();
 sg13g2_fill_1 FILLER_52_1659 ();
 sg13g2_decap_8 FILLER_52_1675 ();
 sg13g2_decap_8 FILLER_52_1682 ();
 sg13g2_decap_4 FILLER_52_1689 ();
 sg13g2_fill_1 FILLER_52_1693 ();
 sg13g2_decap_8 FILLER_52_1720 ();
 sg13g2_decap_8 FILLER_52_1727 ();
 sg13g2_fill_1 FILLER_52_1744 ();
 sg13g2_decap_8 FILLER_52_1768 ();
 sg13g2_fill_1 FILLER_52_1775 ();
 sg13g2_decap_8 FILLER_52_1780 ();
 sg13g2_fill_2 FILLER_52_1787 ();
 sg13g2_fill_1 FILLER_52_1789 ();
 sg13g2_fill_1 FILLER_52_1795 ();
 sg13g2_fill_1 FILLER_52_1810 ();
 sg13g2_fill_2 FILLER_52_1820 ();
 sg13g2_fill_1 FILLER_52_1822 ();
 sg13g2_decap_4 FILLER_52_1864 ();
 sg13g2_fill_1 FILLER_52_1881 ();
 sg13g2_fill_1 FILLER_52_1887 ();
 sg13g2_fill_1 FILLER_52_1901 ();
 sg13g2_fill_1 FILLER_52_1915 ();
 sg13g2_fill_2 FILLER_52_1938 ();
 sg13g2_fill_1 FILLER_52_1985 ();
 sg13g2_fill_2 FILLER_52_2027 ();
 sg13g2_fill_1 FILLER_52_2029 ();
 sg13g2_fill_2 FILLER_52_2034 ();
 sg13g2_fill_2 FILLER_52_2080 ();
 sg13g2_fill_2 FILLER_52_2117 ();
 sg13g2_fill_2 FILLER_52_2132 ();
 sg13g2_fill_1 FILLER_52_2134 ();
 sg13g2_fill_2 FILLER_52_2140 ();
 sg13g2_fill_1 FILLER_52_2173 ();
 sg13g2_fill_1 FILLER_52_2240 ();
 sg13g2_fill_2 FILLER_52_2254 ();
 sg13g2_fill_1 FILLER_52_2256 ();
 sg13g2_fill_1 FILLER_52_2288 ();
 sg13g2_fill_2 FILLER_52_2342 ();
 sg13g2_fill_2 FILLER_52_2370 ();
 sg13g2_fill_2 FILLER_52_2416 ();
 sg13g2_fill_1 FILLER_52_2428 ();
 sg13g2_fill_1 FILLER_52_2434 ();
 sg13g2_fill_2 FILLER_52_2457 ();
 sg13g2_fill_2 FILLER_52_2483 ();
 sg13g2_fill_2 FILLER_52_2523 ();
 sg13g2_fill_2 FILLER_52_2542 ();
 sg13g2_fill_1 FILLER_52_2544 ();
 sg13g2_decap_8 FILLER_52_2549 ();
 sg13g2_decap_4 FILLER_52_2556 ();
 sg13g2_fill_2 FILLER_52_2560 ();
 sg13g2_fill_1 FILLER_52_2587 ();
 sg13g2_fill_2 FILLER_52_2614 ();
 sg13g2_fill_1 FILLER_52_2616 ();
 sg13g2_fill_1 FILLER_52_2644 ();
 sg13g2_fill_1 FILLER_52_2673 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_fill_2 FILLER_53_64 ();
 sg13g2_fill_2 FILLER_53_94 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_175 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_fill_2 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_561 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_fill_1 FILLER_53_596 ();
 sg13g2_fill_2 FILLER_53_646 ();
 sg13g2_fill_2 FILLER_53_653 ();
 sg13g2_fill_2 FILLER_53_660 ();
 sg13g2_decap_4 FILLER_53_676 ();
 sg13g2_fill_2 FILLER_53_693 ();
 sg13g2_fill_1 FILLER_53_729 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_833 ();
 sg13g2_fill_1 FILLER_53_868 ();
 sg13g2_fill_2 FILLER_53_895 ();
 sg13g2_fill_1 FILLER_53_944 ();
 sg13g2_decap_4 FILLER_53_1001 ();
 sg13g2_fill_2 FILLER_53_1005 ();
 sg13g2_fill_1 FILLER_53_1016 ();
 sg13g2_fill_2 FILLER_53_1022 ();
 sg13g2_fill_2 FILLER_53_1043 ();
 sg13g2_fill_1 FILLER_53_1045 ();
 sg13g2_fill_1 FILLER_53_1084 ();
 sg13g2_fill_2 FILLER_53_1100 ();
 sg13g2_fill_1 FILLER_53_1116 ();
 sg13g2_fill_2 FILLER_53_1149 ();
 sg13g2_fill_1 FILLER_53_1165 ();
 sg13g2_fill_1 FILLER_53_1180 ();
 sg13g2_fill_1 FILLER_53_1216 ();
 sg13g2_fill_1 FILLER_53_1234 ();
 sg13g2_fill_2 FILLER_53_1362 ();
 sg13g2_fill_1 FILLER_53_1364 ();
 sg13g2_fill_2 FILLER_53_1370 ();
 sg13g2_fill_1 FILLER_53_1372 ();
 sg13g2_fill_2 FILLER_53_1408 ();
 sg13g2_fill_1 FILLER_53_1414 ();
 sg13g2_decap_4 FILLER_53_1424 ();
 sg13g2_fill_2 FILLER_53_1463 ();
 sg13g2_fill_1 FILLER_53_1465 ();
 sg13g2_fill_1 FILLER_53_1526 ();
 sg13g2_decap_8 FILLER_53_1562 ();
 sg13g2_decap_4 FILLER_53_1569 ();
 sg13g2_decap_8 FILLER_53_1603 ();
 sg13g2_fill_2 FILLER_53_1610 ();
 sg13g2_fill_1 FILLER_53_1612 ();
 sg13g2_fill_1 FILLER_53_1617 ();
 sg13g2_decap_8 FILLER_53_1638 ();
 sg13g2_decap_8 FILLER_53_1645 ();
 sg13g2_decap_8 FILLER_53_1663 ();
 sg13g2_decap_8 FILLER_53_1670 ();
 sg13g2_decap_4 FILLER_53_1677 ();
 sg13g2_fill_1 FILLER_53_1681 ();
 sg13g2_decap_4 FILLER_53_1686 ();
 sg13g2_fill_1 FILLER_53_1690 ();
 sg13g2_fill_2 FILLER_53_1696 ();
 sg13g2_fill_1 FILLER_53_1711 ();
 sg13g2_fill_2 FILLER_53_1726 ();
 sg13g2_fill_2 FILLER_53_1733 ();
 sg13g2_fill_1 FILLER_53_1735 ();
 sg13g2_decap_8 FILLER_53_1758 ();
 sg13g2_decap_8 FILLER_53_1765 ();
 sg13g2_decap_4 FILLER_53_1772 ();
 sg13g2_fill_2 FILLER_53_1776 ();
 sg13g2_fill_1 FILLER_53_1802 ();
 sg13g2_fill_2 FILLER_53_1816 ();
 sg13g2_fill_2 FILLER_53_1826 ();
 sg13g2_fill_2 FILLER_53_1860 ();
 sg13g2_fill_1 FILLER_53_1893 ();
 sg13g2_decap_8 FILLER_53_1903 ();
 sg13g2_decap_4 FILLER_53_1910 ();
 sg13g2_fill_1 FILLER_53_1914 ();
 sg13g2_fill_2 FILLER_53_1982 ();
 sg13g2_fill_1 FILLER_53_1993 ();
 sg13g2_fill_1 FILLER_53_2034 ();
 sg13g2_fill_2 FILLER_53_2085 ();
 sg13g2_fill_2 FILLER_53_2101 ();
 sg13g2_fill_1 FILLER_53_2103 ();
 sg13g2_fill_1 FILLER_53_2183 ();
 sg13g2_fill_2 FILLER_53_2218 ();
 sg13g2_fill_1 FILLER_53_2220 ();
 sg13g2_fill_1 FILLER_53_2231 ();
 sg13g2_fill_1 FILLER_53_2254 ();
 sg13g2_fill_1 FILLER_53_2266 ();
 sg13g2_fill_2 FILLER_53_2285 ();
 sg13g2_fill_2 FILLER_53_2354 ();
 sg13g2_fill_2 FILLER_53_2383 ();
 sg13g2_fill_1 FILLER_53_2385 ();
 sg13g2_fill_2 FILLER_53_2416 ();
 sg13g2_fill_2 FILLER_53_2450 ();
 sg13g2_fill_1 FILLER_53_2452 ();
 sg13g2_fill_1 FILLER_53_2466 ();
 sg13g2_fill_2 FILLER_53_2471 ();
 sg13g2_fill_2 FILLER_53_2552 ();
 sg13g2_fill_1 FILLER_53_2554 ();
 sg13g2_decap_4 FILLER_53_2561 ();
 sg13g2_fill_1 FILLER_53_2565 ();
 sg13g2_fill_2 FILLER_53_2582 ();
 sg13g2_fill_2 FILLER_53_2620 ();
 sg13g2_fill_1 FILLER_53_2622 ();
 sg13g2_fill_2 FILLER_53_2659 ();
 sg13g2_decap_4 FILLER_53_2670 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_115 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_228 ();
 sg13g2_fill_1 FILLER_54_271 ();
 sg13g2_fill_1 FILLER_54_344 ();
 sg13g2_fill_1 FILLER_54_452 ();
 sg13g2_fill_1 FILLER_54_488 ();
 sg13g2_fill_1 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_fill_2 FILLER_54_636 ();
 sg13g2_fill_1 FILLER_54_638 ();
 sg13g2_fill_1 FILLER_54_697 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_fill_1 FILLER_54_741 ();
 sg13g2_fill_2 FILLER_54_791 ();
 sg13g2_fill_1 FILLER_54_830 ();
 sg13g2_fill_2 FILLER_54_866 ();
 sg13g2_fill_1 FILLER_54_909 ();
 sg13g2_fill_2 FILLER_54_949 ();
 sg13g2_fill_1 FILLER_54_1022 ();
 sg13g2_fill_2 FILLER_54_1051 ();
 sg13g2_fill_1 FILLER_54_1053 ();
 sg13g2_fill_2 FILLER_54_1100 ();
 sg13g2_fill_2 FILLER_54_1135 ();
 sg13g2_fill_1 FILLER_54_1265 ();
 sg13g2_fill_1 FILLER_54_1354 ();
 sg13g2_decap_4 FILLER_54_1399 ();
 sg13g2_fill_1 FILLER_54_1403 ();
 sg13g2_fill_2 FILLER_54_1422 ();
 sg13g2_fill_1 FILLER_54_1424 ();
 sg13g2_decap_4 FILLER_54_1501 ();
 sg13g2_fill_1 FILLER_54_1505 ();
 sg13g2_fill_1 FILLER_54_1545 ();
 sg13g2_fill_1 FILLER_54_1558 ();
 sg13g2_decap_8 FILLER_54_1563 ();
 sg13g2_decap_4 FILLER_54_1570 ();
 sg13g2_fill_1 FILLER_54_1574 ();
 sg13g2_fill_2 FILLER_54_1583 ();
 sg13g2_fill_1 FILLER_54_1585 ();
 sg13g2_decap_8 FILLER_54_1606 ();
 sg13g2_fill_1 FILLER_54_1623 ();
 sg13g2_decap_8 FILLER_54_1634 ();
 sg13g2_fill_2 FILLER_54_1641 ();
 sg13g2_fill_1 FILLER_54_1666 ();
 sg13g2_decap_4 FILLER_54_1702 ();
 sg13g2_fill_2 FILLER_54_1706 ();
 sg13g2_fill_1 FILLER_54_1712 ();
 sg13g2_fill_2 FILLER_54_1718 ();
 sg13g2_fill_1 FILLER_54_1720 ();
 sg13g2_decap_8 FILLER_54_1731 ();
 sg13g2_fill_2 FILLER_54_1738 ();
 sg13g2_fill_1 FILLER_54_1740 ();
 sg13g2_decap_8 FILLER_54_1753 ();
 sg13g2_decap_8 FILLER_54_1760 ();
 sg13g2_decap_8 FILLER_54_1767 ();
 sg13g2_fill_2 FILLER_54_1783 ();
 sg13g2_fill_1 FILLER_54_1785 ();
 sg13g2_fill_2 FILLER_54_1810 ();
 sg13g2_fill_1 FILLER_54_1812 ();
 sg13g2_decap_8 FILLER_54_1831 ();
 sg13g2_fill_2 FILLER_54_1838 ();
 sg13g2_fill_1 FILLER_54_1840 ();
 sg13g2_fill_1 FILLER_54_1846 ();
 sg13g2_fill_1 FILLER_54_1920 ();
 sg13g2_fill_2 FILLER_54_1957 ();
 sg13g2_fill_1 FILLER_54_1959 ();
 sg13g2_fill_1 FILLER_54_1983 ();
 sg13g2_fill_1 FILLER_54_2020 ();
 sg13g2_fill_2 FILLER_54_2060 ();
 sg13g2_fill_1 FILLER_54_2062 ();
 sg13g2_fill_2 FILLER_54_2090 ();
 sg13g2_fill_2 FILLER_54_2188 ();
 sg13g2_fill_2 FILLER_54_2222 ();
 sg13g2_fill_1 FILLER_54_2298 ();
 sg13g2_fill_1 FILLER_54_2340 ();
 sg13g2_fill_2 FILLER_54_2394 ();
 sg13g2_fill_1 FILLER_54_2396 ();
 sg13g2_fill_2 FILLER_54_2536 ();
 sg13g2_fill_1 FILLER_54_2538 ();
 sg13g2_fill_2 FILLER_54_2612 ();
 sg13g2_fill_1 FILLER_54_2614 ();
 sg13g2_decap_4 FILLER_54_2668 ();
 sg13g2_fill_2 FILLER_54_2672 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_23 ();
 sg13g2_fill_1 FILLER_55_25 ();
 sg13g2_fill_1 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_fill_2 FILLER_55_62 ();
 sg13g2_fill_2 FILLER_55_69 ();
 sg13g2_fill_2 FILLER_55_181 ();
 sg13g2_fill_2 FILLER_55_240 ();
 sg13g2_fill_2 FILLER_55_270 ();
 sg13g2_fill_1 FILLER_55_272 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_314 ();
 sg13g2_fill_2 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_391 ();
 sg13g2_fill_2 FILLER_55_538 ();
 sg13g2_fill_1 FILLER_55_586 ();
 sg13g2_fill_2 FILLER_55_611 ();
 sg13g2_fill_2 FILLER_55_635 ();
 sg13g2_fill_2 FILLER_55_655 ();
 sg13g2_fill_1 FILLER_55_657 ();
 sg13g2_fill_1 FILLER_55_769 ();
 sg13g2_fill_2 FILLER_55_783 ();
 sg13g2_fill_2 FILLER_55_825 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_fill_1 FILLER_55_914 ();
 sg13g2_fill_1 FILLER_55_921 ();
 sg13g2_fill_2 FILLER_55_949 ();
 sg13g2_fill_1 FILLER_55_951 ();
 sg13g2_fill_1 FILLER_55_956 ();
 sg13g2_fill_1 FILLER_55_971 ();
 sg13g2_decap_8 FILLER_55_989 ();
 sg13g2_decap_4 FILLER_55_996 ();
 sg13g2_fill_1 FILLER_55_1000 ();
 sg13g2_fill_1 FILLER_55_1015 ();
 sg13g2_fill_1 FILLER_55_1040 ();
 sg13g2_fill_2 FILLER_55_1081 ();
 sg13g2_fill_1 FILLER_55_1125 ();
 sg13g2_fill_1 FILLER_55_1190 ();
 sg13g2_fill_2 FILLER_55_1227 ();
 sg13g2_decap_4 FILLER_55_1321 ();
 sg13g2_fill_1 FILLER_55_1325 ();
 sg13g2_fill_2 FILLER_55_1342 ();
 sg13g2_fill_1 FILLER_55_1377 ();
 sg13g2_decap_8 FILLER_55_1384 ();
 sg13g2_fill_2 FILLER_55_1391 ();
 sg13g2_fill_1 FILLER_55_1393 ();
 sg13g2_fill_2 FILLER_55_1419 ();
 sg13g2_fill_1 FILLER_55_1467 ();
 sg13g2_fill_2 FILLER_55_1481 ();
 sg13g2_fill_1 FILLER_55_1483 ();
 sg13g2_fill_2 FILLER_55_1521 ();
 sg13g2_fill_1 FILLER_55_1528 ();
 sg13g2_fill_1 FILLER_55_1534 ();
 sg13g2_decap_8 FILLER_55_1555 ();
 sg13g2_decap_8 FILLER_55_1562 ();
 sg13g2_decap_4 FILLER_55_1569 ();
 sg13g2_fill_1 FILLER_55_1573 ();
 sg13g2_fill_2 FILLER_55_1577 ();
 sg13g2_fill_1 FILLER_55_1584 ();
 sg13g2_fill_2 FILLER_55_1589 ();
 sg13g2_fill_1 FILLER_55_1591 ();
 sg13g2_fill_1 FILLER_55_1597 ();
 sg13g2_fill_1 FILLER_55_1603 ();
 sg13g2_fill_2 FILLER_55_1622 ();
 sg13g2_fill_1 FILLER_55_1624 ();
 sg13g2_decap_8 FILLER_55_1631 ();
 sg13g2_decap_8 FILLER_55_1638 ();
 sg13g2_decap_8 FILLER_55_1645 ();
 sg13g2_decap_4 FILLER_55_1692 ();
 sg13g2_fill_2 FILLER_55_1696 ();
 sg13g2_decap_8 FILLER_55_1725 ();
 sg13g2_decap_4 FILLER_55_1732 ();
 sg13g2_decap_8 FILLER_55_1760 ();
 sg13g2_fill_1 FILLER_55_1808 ();
 sg13g2_decap_4 FILLER_55_1835 ();
 sg13g2_fill_1 FILLER_55_1839 ();
 sg13g2_fill_2 FILLER_55_1862 ();
 sg13g2_fill_2 FILLER_55_1945 ();
 sg13g2_fill_1 FILLER_55_1953 ();
 sg13g2_fill_2 FILLER_55_1997 ();
 sg13g2_fill_2 FILLER_55_2045 ();
 sg13g2_fill_1 FILLER_55_2047 ();
 sg13g2_fill_2 FILLER_55_2063 ();
 sg13g2_fill_2 FILLER_55_2114 ();
 sg13g2_fill_1 FILLER_55_2116 ();
 sg13g2_fill_1 FILLER_55_2130 ();
 sg13g2_fill_2 FILLER_55_2144 ();
 sg13g2_fill_2 FILLER_55_2178 ();
 sg13g2_fill_1 FILLER_55_2180 ();
 sg13g2_fill_2 FILLER_55_2218 ();
 sg13g2_fill_1 FILLER_55_2220 ();
 sg13g2_fill_2 FILLER_55_2255 ();
 sg13g2_fill_1 FILLER_55_2257 ();
 sg13g2_fill_2 FILLER_55_2386 ();
 sg13g2_fill_1 FILLER_55_2426 ();
 sg13g2_fill_2 FILLER_55_2458 ();
 sg13g2_fill_2 FILLER_55_2497 ();
 sg13g2_fill_1 FILLER_55_2582 ();
 sg13g2_fill_2 FILLER_55_2610 ();
 sg13g2_fill_1 FILLER_55_2612 ();
 sg13g2_fill_2 FILLER_55_2639 ();
 sg13g2_fill_1 FILLER_55_2673 ();
 sg13g2_fill_2 FILLER_56_41 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_2 FILLER_56_71 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_fill_1 FILLER_56_331 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_2 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_437 ();
 sg13g2_fill_2 FILLER_56_568 ();
 sg13g2_fill_1 FILLER_56_570 ();
 sg13g2_fill_1 FILLER_56_605 ();
 sg13g2_fill_1 FILLER_56_631 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_2 FILLER_56_669 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_742 ();
 sg13g2_fill_2 FILLER_56_789 ();
 sg13g2_fill_2 FILLER_56_869 ();
 sg13g2_fill_1 FILLER_56_871 ();
 sg13g2_fill_2 FILLER_56_949 ();
 sg13g2_fill_1 FILLER_56_970 ();
 sg13g2_fill_1 FILLER_56_981 ();
 sg13g2_decap_4 FILLER_56_996 ();
 sg13g2_fill_2 FILLER_56_1000 ();
 sg13g2_fill_1 FILLER_56_1030 ();
 sg13g2_fill_1 FILLER_56_1040 ();
 sg13g2_fill_2 FILLER_56_1064 ();
 sg13g2_fill_1 FILLER_56_1066 ();
 sg13g2_decap_4 FILLER_56_1085 ();
 sg13g2_fill_2 FILLER_56_1157 ();
 sg13g2_fill_1 FILLER_56_1159 ();
 sg13g2_fill_2 FILLER_56_1197 ();
 sg13g2_fill_1 FILLER_56_1199 ();
 sg13g2_fill_2 FILLER_56_1226 ();
 sg13g2_fill_1 FILLER_56_1228 ();
 sg13g2_fill_1 FILLER_56_1262 ();
 sg13g2_fill_2 FILLER_56_1282 ();
 sg13g2_decap_8 FILLER_56_1322 ();
 sg13g2_fill_2 FILLER_56_1329 ();
 sg13g2_fill_1 FILLER_56_1344 ();
 sg13g2_fill_2 FILLER_56_1379 ();
 sg13g2_decap_8 FILLER_56_1385 ();
 sg13g2_decap_4 FILLER_56_1392 ();
 sg13g2_decap_8 FILLER_56_1429 ();
 sg13g2_fill_1 FILLER_56_1436 ();
 sg13g2_fill_2 FILLER_56_1490 ();
 sg13g2_fill_1 FILLER_56_1492 ();
 sg13g2_fill_1 FILLER_56_1529 ();
 sg13g2_fill_2 FILLER_56_1540 ();
 sg13g2_fill_1 FILLER_56_1574 ();
 sg13g2_fill_2 FILLER_56_1580 ();
 sg13g2_decap_8 FILLER_56_1590 ();
 sg13g2_decap_4 FILLER_56_1597 ();
 sg13g2_fill_2 FILLER_56_1606 ();
 sg13g2_decap_8 FILLER_56_1629 ();
 sg13g2_decap_8 FILLER_56_1636 ();
 sg13g2_decap_4 FILLER_56_1643 ();
 sg13g2_fill_1 FILLER_56_1647 ();
 sg13g2_fill_1 FILLER_56_1675 ();
 sg13g2_decap_8 FILLER_56_1682 ();
 sg13g2_fill_1 FILLER_56_1689 ();
 sg13g2_fill_2 FILLER_56_1695 ();
 sg13g2_fill_1 FILLER_56_1697 ();
 sg13g2_fill_2 FILLER_56_1701 ();
 sg13g2_decap_8 FILLER_56_1713 ();
 sg13g2_decap_8 FILLER_56_1720 ();
 sg13g2_fill_2 FILLER_56_1727 ();
 sg13g2_decap_8 FILLER_56_1753 ();
 sg13g2_decap_8 FILLER_56_1760 ();
 sg13g2_fill_1 FILLER_56_1767 ();
 sg13g2_fill_1 FILLER_56_1800 ();
 sg13g2_fill_2 FILLER_56_1810 ();
 sg13g2_decap_4 FILLER_56_1844 ();
 sg13g2_fill_2 FILLER_56_1848 ();
 sg13g2_fill_1 FILLER_56_1874 ();
 sg13g2_fill_2 FILLER_56_1899 ();
 sg13g2_fill_1 FILLER_56_1952 ();
 sg13g2_fill_1 FILLER_56_1959 ();
 sg13g2_fill_1 FILLER_56_1997 ();
 sg13g2_fill_1 FILLER_56_2012 ();
 sg13g2_fill_1 FILLER_56_2032 ();
 sg13g2_fill_2 FILLER_56_2108 ();
 sg13g2_fill_2 FILLER_56_2136 ();
 sg13g2_fill_1 FILLER_56_2138 ();
 sg13g2_fill_2 FILLER_56_2204 ();
 sg13g2_fill_1 FILLER_56_2206 ();
 sg13g2_fill_2 FILLER_56_2290 ();
 sg13g2_fill_2 FILLER_56_2338 ();
 sg13g2_fill_1 FILLER_56_2340 ();
 sg13g2_fill_2 FILLER_56_2354 ();
 sg13g2_fill_2 FILLER_56_2382 ();
 sg13g2_fill_1 FILLER_56_2384 ();
 sg13g2_fill_2 FILLER_56_2402 ();
 sg13g2_fill_1 FILLER_56_2404 ();
 sg13g2_fill_1 FILLER_56_2418 ();
 sg13g2_fill_1 FILLER_56_2432 ();
 sg13g2_fill_1 FILLER_56_2442 ();
 sg13g2_fill_2 FILLER_56_2456 ();
 sg13g2_fill_1 FILLER_56_2471 ();
 sg13g2_fill_1 FILLER_56_2481 ();
 sg13g2_fill_1 FILLER_56_2514 ();
 sg13g2_fill_2 FILLER_56_2547 ();
 sg13g2_fill_1 FILLER_56_2612 ();
 sg13g2_fill_1 FILLER_56_2673 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_2 FILLER_57_231 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_fill_2 FILLER_57_265 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_359 ();
 sg13g2_fill_1 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_548 ();
 sg13g2_fill_1 FILLER_57_566 ();
 sg13g2_fill_2 FILLER_57_584 ();
 sg13g2_fill_1 FILLER_57_586 ();
 sg13g2_fill_1 FILLER_57_713 ();
 sg13g2_fill_2 FILLER_57_719 ();
 sg13g2_fill_2 FILLER_57_767 ();
 sg13g2_fill_2 FILLER_57_782 ();
 sg13g2_fill_1 FILLER_57_784 ();
 sg13g2_fill_2 FILLER_57_801 ();
 sg13g2_decap_4 FILLER_57_808 ();
 sg13g2_fill_2 FILLER_57_838 ();
 sg13g2_fill_1 FILLER_57_840 ();
 sg13g2_fill_2 FILLER_57_863 ();
 sg13g2_fill_1 FILLER_57_865 ();
 sg13g2_fill_2 FILLER_57_899 ();
 sg13g2_fill_1 FILLER_57_901 ();
 sg13g2_fill_2 FILLER_57_911 ();
 sg13g2_fill_1 FILLER_57_913 ();
 sg13g2_fill_2 FILLER_57_923 ();
 sg13g2_fill_1 FILLER_57_1019 ();
 sg13g2_fill_1 FILLER_57_1089 ();
 sg13g2_fill_2 FILLER_57_1094 ();
 sg13g2_fill_1 FILLER_57_1186 ();
 sg13g2_fill_1 FILLER_57_1227 ();
 sg13g2_fill_2 FILLER_57_1325 ();
 sg13g2_fill_1 FILLER_57_1327 ();
 sg13g2_decap_4 FILLER_57_1346 ();
 sg13g2_fill_2 FILLER_57_1350 ();
 sg13g2_fill_1 FILLER_57_1365 ();
 sg13g2_fill_2 FILLER_57_1372 ();
 sg13g2_fill_2 FILLER_57_1449 ();
 sg13g2_fill_1 FILLER_57_1478 ();
 sg13g2_fill_1 FILLER_57_1561 ();
 sg13g2_fill_1 FILLER_57_1583 ();
 sg13g2_decap_4 FILLER_57_1599 ();
 sg13g2_fill_1 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1640 ();
 sg13g2_decap_8 FILLER_57_1651 ();
 sg13g2_fill_1 FILLER_57_1658 ();
 sg13g2_fill_2 FILLER_57_1664 ();
 sg13g2_decap_8 FILLER_57_1679 ();
 sg13g2_decap_8 FILLER_57_1686 ();
 sg13g2_decap_8 FILLER_57_1693 ();
 sg13g2_decap_8 FILLER_57_1700 ();
 sg13g2_decap_8 FILLER_57_1707 ();
 sg13g2_decap_4 FILLER_57_1718 ();
 sg13g2_fill_2 FILLER_57_1722 ();
 sg13g2_decap_8 FILLER_57_1750 ();
 sg13g2_fill_2 FILLER_57_1757 ();
 sg13g2_fill_1 FILLER_57_1799 ();
 sg13g2_decap_4 FILLER_57_1817 ();
 sg13g2_fill_2 FILLER_57_1838 ();
 sg13g2_fill_1 FILLER_57_1849 ();
 sg13g2_fill_2 FILLER_57_1854 ();
 sg13g2_fill_1 FILLER_57_1889 ();
 sg13g2_fill_1 FILLER_57_1899 ();
 sg13g2_decap_4 FILLER_57_1913 ();
 sg13g2_fill_2 FILLER_57_1930 ();
 sg13g2_fill_2 FILLER_57_1963 ();
 sg13g2_fill_1 FILLER_57_1965 ();
 sg13g2_fill_1 FILLER_57_1991 ();
 sg13g2_fill_2 FILLER_57_2019 ();
 sg13g2_fill_2 FILLER_57_2057 ();
 sg13g2_fill_1 FILLER_57_2135 ();
 sg13g2_fill_1 FILLER_57_2149 ();
 sg13g2_fill_2 FILLER_57_2183 ();
 sg13g2_fill_2 FILLER_57_2245 ();
 sg13g2_fill_1 FILLER_57_2247 ();
 sg13g2_fill_1 FILLER_57_2300 ();
 sg13g2_decap_8 FILLER_57_2332 ();
 sg13g2_fill_2 FILLER_57_2339 ();
 sg13g2_fill_2 FILLER_57_2367 ();
 sg13g2_fill_1 FILLER_57_2378 ();
 sg13g2_fill_2 FILLER_57_2430 ();
 sg13g2_decap_4 FILLER_57_2446 ();
 sg13g2_fill_2 FILLER_57_2468 ();
 sg13g2_fill_1 FILLER_57_2470 ();
 sg13g2_fill_2 FILLER_57_2477 ();
 sg13g2_fill_1 FILLER_57_2479 ();
 sg13g2_fill_2 FILLER_57_2507 ();
 sg13g2_fill_1 FILLER_57_2509 ();
 sg13g2_fill_1 FILLER_57_2561 ();
 sg13g2_fill_2 FILLER_57_2574 ();
 sg13g2_fill_1 FILLER_57_2581 ();
 sg13g2_fill_1 FILLER_57_2600 ();
 sg13g2_fill_1 FILLER_57_2632 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_118 ();
 sg13g2_fill_2 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_208 ();
 sg13g2_fill_1 FILLER_58_220 ();
 sg13g2_fill_2 FILLER_58_340 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_358 ();
 sg13g2_fill_2 FILLER_58_458 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_fill_2 FILLER_58_505 ();
 sg13g2_fill_1 FILLER_58_511 ();
 sg13g2_fill_1 FILLER_58_577 ();
 sg13g2_fill_2 FILLER_58_587 ();
 sg13g2_fill_1 FILLER_58_601 ();
 sg13g2_fill_2 FILLER_58_618 ();
 sg13g2_fill_2 FILLER_58_687 ();
 sg13g2_fill_2 FILLER_58_753 ();
 sg13g2_decap_4 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_961 ();
 sg13g2_decap_4 FILLER_58_998 ();
 sg13g2_fill_1 FILLER_58_1002 ();
 sg13g2_fill_2 FILLER_58_1012 ();
 sg13g2_fill_1 FILLER_58_1054 ();
 sg13g2_fill_1 FILLER_58_1062 ();
 sg13g2_decap_8 FILLER_58_1073 ();
 sg13g2_decap_4 FILLER_58_1080 ();
 sg13g2_fill_2 FILLER_58_1084 ();
 sg13g2_fill_1 FILLER_58_1126 ();
 sg13g2_fill_2 FILLER_58_1132 ();
 sg13g2_fill_1 FILLER_58_1160 ();
 sg13g2_decap_4 FILLER_58_1223 ();
 sg13g2_fill_2 FILLER_58_1227 ();
 sg13g2_decap_4 FILLER_58_1321 ();
 sg13g2_fill_2 FILLER_58_1325 ();
 sg13g2_decap_8 FILLER_58_1355 ();
 sg13g2_fill_1 FILLER_58_1362 ();
 sg13g2_fill_2 FILLER_58_1391 ();
 sg13g2_fill_2 FILLER_58_1434 ();
 sg13g2_decap_8 FILLER_58_1477 ();
 sg13g2_fill_2 FILLER_58_1484 ();
 sg13g2_fill_1 FILLER_58_1486 ();
 sg13g2_decap_8 FILLER_58_1490 ();
 sg13g2_decap_8 FILLER_58_1497 ();
 sg13g2_decap_8 FILLER_58_1504 ();
 sg13g2_fill_2 FILLER_58_1511 ();
 sg13g2_fill_2 FILLER_58_1526 ();
 sg13g2_fill_1 FILLER_58_1528 ();
 sg13g2_fill_2 FILLER_58_1547 ();
 sg13g2_fill_2 FILLER_58_1568 ();
 sg13g2_fill_1 FILLER_58_1585 ();
 sg13g2_fill_1 FILLER_58_1591 ();
 sg13g2_fill_2 FILLER_58_1600 ();
 sg13g2_fill_1 FILLER_58_1602 ();
 sg13g2_decap_4 FILLER_58_1628 ();
 sg13g2_fill_1 FILLER_58_1632 ();
 sg13g2_decap_8 FILLER_58_1642 ();
 sg13g2_decap_4 FILLER_58_1649 ();
 sg13g2_decap_8 FILLER_58_1656 ();
 sg13g2_decap_4 FILLER_58_1663 ();
 sg13g2_fill_1 FILLER_58_1667 ();
 sg13g2_decap_8 FILLER_58_1687 ();
 sg13g2_decap_8 FILLER_58_1694 ();
 sg13g2_decap_4 FILLER_58_1701 ();
 sg13g2_fill_1 FILLER_58_1705 ();
 sg13g2_decap_8 FILLER_58_1716 ();
 sg13g2_decap_4 FILLER_58_1723 ();
 sg13g2_fill_1 FILLER_58_1727 ();
 sg13g2_decap_8 FILLER_58_1732 ();
 sg13g2_decap_8 FILLER_58_1739 ();
 sg13g2_decap_8 FILLER_58_1746 ();
 sg13g2_decap_8 FILLER_58_1753 ();
 sg13g2_decap_8 FILLER_58_1760 ();
 sg13g2_decap_8 FILLER_58_1767 ();
 sg13g2_fill_1 FILLER_58_1774 ();
 sg13g2_decap_4 FILLER_58_1802 ();
 sg13g2_fill_2 FILLER_58_1806 ();
 sg13g2_decap_4 FILLER_58_1843 ();
 sg13g2_fill_2 FILLER_58_1847 ();
 sg13g2_fill_1 FILLER_58_1911 ();
 sg13g2_fill_1 FILLER_58_1939 ();
 sg13g2_fill_2 FILLER_58_1944 ();
 sg13g2_fill_1 FILLER_58_1946 ();
 sg13g2_fill_2 FILLER_58_1953 ();
 sg13g2_fill_1 FILLER_58_2032 ();
 sg13g2_fill_1 FILLER_58_2073 ();
 sg13g2_fill_2 FILLER_58_2196 ();
 sg13g2_fill_2 FILLER_58_2269 ();
 sg13g2_fill_2 FILLER_58_2323 ();
 sg13g2_decap_8 FILLER_58_2338 ();
 sg13g2_fill_2 FILLER_58_2345 ();
 sg13g2_fill_2 FILLER_58_2398 ();
 sg13g2_fill_1 FILLER_58_2400 ();
 sg13g2_decap_8 FILLER_58_2433 ();
 sg13g2_decap_4 FILLER_58_2440 ();
 sg13g2_fill_1 FILLER_58_2444 ();
 sg13g2_fill_2 FILLER_58_2485 ();
 sg13g2_fill_2 FILLER_58_2496 ();
 sg13g2_fill_1 FILLER_58_2498 ();
 sg13g2_fill_1 FILLER_58_2535 ();
 sg13g2_fill_1 FILLER_58_2590 ();
 sg13g2_fill_2 FILLER_58_2671 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_2 FILLER_59_47 ();
 sg13g2_fill_1 FILLER_59_81 ();
 sg13g2_fill_2 FILLER_59_103 ();
 sg13g2_fill_1 FILLER_59_105 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_1 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_fill_1 FILLER_59_302 ();
 sg13g2_fill_2 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_428 ();
 sg13g2_fill_2 FILLER_59_438 ();
 sg13g2_fill_1 FILLER_59_440 ();
 sg13g2_fill_1 FILLER_59_450 ();
 sg13g2_fill_1 FILLER_59_500 ();
 sg13g2_fill_1 FILLER_59_551 ();
 sg13g2_fill_1 FILLER_59_580 ();
 sg13g2_fill_1 FILLER_59_649 ();
 sg13g2_fill_1 FILLER_59_677 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_fill_1 FILLER_59_721 ();
 sg13g2_fill_2 FILLER_59_741 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_fill_1 FILLER_59_856 ();
 sg13g2_decap_4 FILLER_59_867 ();
 sg13g2_decap_8 FILLER_59_884 ();
 sg13g2_decap_4 FILLER_59_891 ();
 sg13g2_fill_1 FILLER_59_895 ();
 sg13g2_decap_4 FILLER_59_1009 ();
 sg13g2_fill_2 FILLER_59_1013 ();
 sg13g2_fill_2 FILLER_59_1048 ();
 sg13g2_fill_1 FILLER_59_1234 ();
 sg13g2_fill_2 FILLER_59_1301 ();
 sg13g2_decap_4 FILLER_59_1350 ();
 sg13g2_fill_2 FILLER_59_1354 ();
 sg13g2_fill_2 FILLER_59_1382 ();
 sg13g2_fill_1 FILLER_59_1384 ();
 sg13g2_decap_8 FILLER_59_1424 ();
 sg13g2_decap_4 FILLER_59_1431 ();
 sg13g2_fill_1 FILLER_59_1435 ();
 sg13g2_decap_4 FILLER_59_1441 ();
 sg13g2_fill_2 FILLER_59_1515 ();
 sg13g2_decap_8 FILLER_59_1552 ();
 sg13g2_decap_8 FILLER_59_1559 ();
 sg13g2_fill_2 FILLER_59_1566 ();
 sg13g2_fill_1 FILLER_59_1568 ();
 sg13g2_decap_4 FILLER_59_1579 ();
 sg13g2_fill_1 FILLER_59_1583 ();
 sg13g2_fill_1 FILLER_59_1588 ();
 sg13g2_decap_8 FILLER_59_1594 ();
 sg13g2_fill_2 FILLER_59_1601 ();
 sg13g2_fill_1 FILLER_59_1603 ();
 sg13g2_decap_4 FILLER_59_1610 ();
 sg13g2_fill_2 FILLER_59_1614 ();
 sg13g2_fill_1 FILLER_59_1621 ();
 sg13g2_fill_1 FILLER_59_1627 ();
 sg13g2_fill_2 FILLER_59_1634 ();
 sg13g2_decap_8 FILLER_59_1649 ();
 sg13g2_decap_4 FILLER_59_1656 ();
 sg13g2_fill_1 FILLER_59_1660 ();
 sg13g2_decap_4 FILLER_59_1683 ();
 sg13g2_decap_8 FILLER_59_1697 ();
 sg13g2_decap_8 FILLER_59_1728 ();
 sg13g2_decap_8 FILLER_59_1735 ();
 sg13g2_decap_8 FILLER_59_1742 ();
 sg13g2_decap_8 FILLER_59_1749 ();
 sg13g2_decap_8 FILLER_59_1756 ();
 sg13g2_fill_2 FILLER_59_1763 ();
 sg13g2_fill_2 FILLER_59_1796 ();
 sg13g2_fill_2 FILLER_59_1843 ();
 sg13g2_fill_2 FILLER_59_1873 ();
 sg13g2_fill_1 FILLER_59_1875 ();
 sg13g2_fill_1 FILLER_59_2015 ();
 sg13g2_fill_1 FILLER_59_2074 ();
 sg13g2_fill_2 FILLER_59_2170 ();
 sg13g2_fill_1 FILLER_59_2172 ();
 sg13g2_fill_1 FILLER_59_2210 ();
 sg13g2_fill_2 FILLER_59_2290 ();
 sg13g2_decap_8 FILLER_59_2332 ();
 sg13g2_decap_8 FILLER_59_2339 ();
 sg13g2_fill_2 FILLER_59_2391 ();
 sg13g2_fill_1 FILLER_59_2393 ();
 sg13g2_fill_2 FILLER_59_2436 ();
 sg13g2_fill_1 FILLER_59_2438 ();
 sg13g2_fill_1 FILLER_59_2481 ();
 sg13g2_fill_2 FILLER_59_2513 ();
 sg13g2_fill_2 FILLER_59_2575 ();
 sg13g2_fill_2 FILLER_59_2595 ();
 sg13g2_fill_1 FILLER_59_2597 ();
 sg13g2_fill_2 FILLER_59_2630 ();
 sg13g2_fill_1 FILLER_59_2673 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_71 ();
 sg13g2_fill_2 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_fill_2 FILLER_60_187 ();
 sg13g2_fill_2 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_fill_1 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_499 ();
 sg13g2_fill_1 FILLER_60_501 ();
 sg13g2_fill_2 FILLER_60_553 ();
 sg13g2_fill_2 FILLER_60_615 ();
 sg13g2_fill_1 FILLER_60_654 ();
 sg13g2_fill_1 FILLER_60_707 ();
 sg13g2_fill_1 FILLER_60_743 ();
 sg13g2_fill_2 FILLER_60_807 ();
 sg13g2_decap_4 FILLER_60_859 ();
 sg13g2_decap_8 FILLER_60_890 ();
 sg13g2_fill_2 FILLER_60_897 ();
 sg13g2_fill_1 FILLER_60_899 ();
 sg13g2_decap_4 FILLER_60_925 ();
 sg13g2_fill_2 FILLER_60_938 ();
 sg13g2_fill_1 FILLER_60_940 ();
 sg13g2_fill_2 FILLER_60_950 ();
 sg13g2_fill_1 FILLER_60_952 ();
 sg13g2_fill_1 FILLER_60_962 ();
 sg13g2_fill_1 FILLER_60_977 ();
 sg13g2_decap_8 FILLER_60_987 ();
 sg13g2_decap_8 FILLER_60_994 ();
 sg13g2_decap_8 FILLER_60_1001 ();
 sg13g2_fill_1 FILLER_60_1008 ();
 sg13g2_decap_8 FILLER_60_1019 ();
 sg13g2_decap_8 FILLER_60_1026 ();
 sg13g2_decap_4 FILLER_60_1033 ();
 sg13g2_fill_2 FILLER_60_1037 ();
 sg13g2_fill_2 FILLER_60_1100 ();
 sg13g2_fill_2 FILLER_60_1115 ();
 sg13g2_fill_2 FILLER_60_1296 ();
 sg13g2_fill_2 FILLER_60_1307 ();
 sg13g2_fill_2 FILLER_60_1349 ();
 sg13g2_fill_1 FILLER_60_1351 ();
 sg13g2_fill_1 FILLER_60_1380 ();
 sg13g2_fill_2 FILLER_60_1389 ();
 sg13g2_fill_1 FILLER_60_1391 ();
 sg13g2_fill_2 FILLER_60_1412 ();
 sg13g2_decap_8 FILLER_60_1419 ();
 sg13g2_fill_1 FILLER_60_1426 ();
 sg13g2_fill_1 FILLER_60_1489 ();
 sg13g2_fill_2 FILLER_60_1504 ();
 sg13g2_decap_4 FILLER_60_1515 ();
 sg13g2_fill_2 FILLER_60_1519 ();
 sg13g2_fill_2 FILLER_60_1530 ();
 sg13g2_decap_8 FILLER_60_1547 ();
 sg13g2_fill_2 FILLER_60_1554 ();
 sg13g2_decap_8 FILLER_60_1562 ();
 sg13g2_decap_4 FILLER_60_1569 ();
 sg13g2_fill_2 FILLER_60_1573 ();
 sg13g2_decap_4 FILLER_60_1579 ();
 sg13g2_fill_2 FILLER_60_1583 ();
 sg13g2_decap_8 FILLER_60_1597 ();
 sg13g2_decap_4 FILLER_60_1604 ();
 sg13g2_fill_1 FILLER_60_1608 ();
 sg13g2_fill_2 FILLER_60_1622 ();
 sg13g2_fill_1 FILLER_60_1624 ();
 sg13g2_decap_8 FILLER_60_1633 ();
 sg13g2_decap_8 FILLER_60_1640 ();
 sg13g2_decap_4 FILLER_60_1647 ();
 sg13g2_fill_2 FILLER_60_1651 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_decap_4 FILLER_60_1693 ();
 sg13g2_fill_2 FILLER_60_1697 ();
 sg13g2_decap_8 FILLER_60_1730 ();
 sg13g2_fill_2 FILLER_60_1810 ();
 sg13g2_fill_1 FILLER_60_1812 ();
 sg13g2_fill_1 FILLER_60_1840 ();
 sg13g2_fill_2 FILLER_60_1880 ();
 sg13g2_fill_1 FILLER_60_1924 ();
 sg13g2_fill_2 FILLER_60_1929 ();
 sg13g2_fill_1 FILLER_60_2011 ();
 sg13g2_fill_1 FILLER_60_2038 ();
 sg13g2_fill_1 FILLER_60_2066 ();
 sg13g2_fill_2 FILLER_60_2093 ();
 sg13g2_fill_2 FILLER_60_2131 ();
 sg13g2_fill_2 FILLER_60_2290 ();
 sg13g2_fill_1 FILLER_60_2292 ();
 sg13g2_decap_4 FILLER_60_2329 ();
 sg13g2_fill_1 FILLER_60_2360 ();
 sg13g2_fill_1 FILLER_60_2407 ();
 sg13g2_fill_1 FILLER_60_2422 ();
 sg13g2_fill_2 FILLER_60_2440 ();
 sg13g2_fill_1 FILLER_60_2473 ();
 sg13g2_fill_2 FILLER_60_2483 ();
 sg13g2_fill_1 FILLER_60_2485 ();
 sg13g2_fill_1 FILLER_60_2504 ();
 sg13g2_decap_8 FILLER_60_2527 ();
 sg13g2_fill_1 FILLER_60_2534 ();
 sg13g2_decap_8 FILLER_60_2539 ();
 sg13g2_fill_2 FILLER_60_2546 ();
 sg13g2_fill_1 FILLER_60_2594 ();
 sg13g2_fill_2 FILLER_60_2641 ();
 sg13g2_fill_2 FILLER_60_2671 ();
 sg13g2_fill_1 FILLER_60_2673 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_72 ();
 sg13g2_fill_2 FILLER_61_79 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_fill_1 FILLER_61_136 ();
 sg13g2_fill_1 FILLER_61_176 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_fill_2 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_262 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_300 ();
 sg13g2_fill_2 FILLER_61_307 ();
 sg13g2_fill_2 FILLER_61_379 ();
 sg13g2_fill_2 FILLER_61_451 ();
 sg13g2_fill_2 FILLER_61_462 ();
 sg13g2_fill_1 FILLER_61_464 ();
 sg13g2_fill_1 FILLER_61_476 ();
 sg13g2_fill_1 FILLER_61_513 ();
 sg13g2_fill_1 FILLER_61_519 ();
 sg13g2_fill_1 FILLER_61_548 ();
 sg13g2_fill_2 FILLER_61_621 ();
 sg13g2_fill_1 FILLER_61_724 ();
 sg13g2_decap_4 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_863 ();
 sg13g2_decap_8 FILLER_61_880 ();
 sg13g2_decap_4 FILLER_61_920 ();
 sg13g2_decap_8 FILLER_61_929 ();
 sg13g2_decap_8 FILLER_61_936 ();
 sg13g2_fill_2 FILLER_61_943 ();
 sg13g2_fill_1 FILLER_61_949 ();
 sg13g2_decap_8 FILLER_61_975 ();
 sg13g2_decap_8 FILLER_61_982 ();
 sg13g2_decap_8 FILLER_61_989 ();
 sg13g2_decap_8 FILLER_61_996 ();
 sg13g2_decap_8 FILLER_61_1031 ();
 sg13g2_fill_2 FILLER_61_1038 ();
 sg13g2_fill_1 FILLER_61_1081 ();
 sg13g2_fill_2 FILLER_61_1091 ();
 sg13g2_fill_2 FILLER_61_1179 ();
 sg13g2_fill_1 FILLER_61_1196 ();
 sg13g2_fill_1 FILLER_61_1259 ();
 sg13g2_fill_1 FILLER_61_1304 ();
 sg13g2_fill_2 FILLER_61_1343 ();
 sg13g2_fill_2 FILLER_61_1358 ();
 sg13g2_fill_1 FILLER_61_1360 ();
 sg13g2_decap_4 FILLER_61_1395 ();
 sg13g2_fill_1 FILLER_61_1399 ();
 sg13g2_fill_1 FILLER_61_1420 ();
 sg13g2_fill_2 FILLER_61_1429 ();
 sg13g2_fill_2 FILLER_61_1477 ();
 sg13g2_decap_8 FILLER_61_1522 ();
 sg13g2_fill_2 FILLER_61_1529 ();
 sg13g2_fill_1 FILLER_61_1538 ();
 sg13g2_decap_8 FILLER_61_1553 ();
 sg13g2_decap_8 FILLER_61_1560 ();
 sg13g2_decap_4 FILLER_61_1567 ();
 sg13g2_fill_2 FILLER_61_1597 ();
 sg13g2_fill_1 FILLER_61_1599 ();
 sg13g2_fill_2 FILLER_61_1614 ();
 sg13g2_fill_1 FILLER_61_1616 ();
 sg13g2_fill_2 FILLER_61_1635 ();
 sg13g2_fill_1 FILLER_61_1656 ();
 sg13g2_fill_1 FILLER_61_1663 ();
 sg13g2_fill_1 FILLER_61_1677 ();
 sg13g2_decap_8 FILLER_61_1688 ();
 sg13g2_decap_8 FILLER_61_1695 ();
 sg13g2_decap_4 FILLER_61_1702 ();
 sg13g2_fill_2 FILLER_61_1706 ();
 sg13g2_decap_8 FILLER_61_1718 ();
 sg13g2_decap_8 FILLER_61_1725 ();
 sg13g2_fill_2 FILLER_61_1732 ();
 sg13g2_fill_1 FILLER_61_1734 ();
 sg13g2_fill_1 FILLER_61_1789 ();
 sg13g2_fill_2 FILLER_61_1808 ();
 sg13g2_decap_4 FILLER_61_1837 ();
 sg13g2_fill_1 FILLER_61_1870 ();
 sg13g2_fill_2 FILLER_61_1877 ();
 sg13g2_fill_2 FILLER_61_1885 ();
 sg13g2_fill_2 FILLER_61_1912 ();
 sg13g2_fill_1 FILLER_61_1914 ();
 sg13g2_fill_1 FILLER_61_1933 ();
 sg13g2_fill_2 FILLER_61_1961 ();
 sg13g2_decap_4 FILLER_61_2022 ();
 sg13g2_fill_1 FILLER_61_2026 ();
 sg13g2_fill_2 FILLER_61_2137 ();
 sg13g2_fill_1 FILLER_61_2219 ();
 sg13g2_fill_1 FILLER_61_2285 ();
 sg13g2_fill_2 FILLER_61_2317 ();
 sg13g2_fill_1 FILLER_61_2319 ();
 sg13g2_fill_2 FILLER_61_2329 ();
 sg13g2_fill_1 FILLER_61_2331 ();
 sg13g2_fill_2 FILLER_61_2342 ();
 sg13g2_fill_1 FILLER_61_2344 ();
 sg13g2_fill_1 FILLER_61_2355 ();
 sg13g2_decap_4 FILLER_61_2365 ();
 sg13g2_fill_2 FILLER_61_2439 ();
 sg13g2_fill_1 FILLER_61_2441 ();
 sg13g2_fill_1 FILLER_61_2452 ();
 sg13g2_fill_2 FILLER_61_2468 ();
 sg13g2_fill_1 FILLER_61_2470 ();
 sg13g2_fill_2 FILLER_61_2477 ();
 sg13g2_fill_1 FILLER_61_2484 ();
 sg13g2_decap_8 FILLER_61_2517 ();
 sg13g2_decap_8 FILLER_61_2524 ();
 sg13g2_decap_8 FILLER_61_2531 ();
 sg13g2_decap_8 FILLER_61_2538 ();
 sg13g2_fill_2 FILLER_61_2545 ();
 sg13g2_fill_2 FILLER_61_2564 ();
 sg13g2_fill_2 FILLER_61_2590 ();
 sg13g2_fill_1 FILLER_61_2592 ();
 sg13g2_fill_1 FILLER_61_2602 ();
 sg13g2_fill_1 FILLER_61_2630 ();
 sg13g2_decap_4 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_61_2672 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_59 ();
 sg13g2_fill_2 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_276 ();
 sg13g2_fill_1 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_319 ();
 sg13g2_fill_1 FILLER_62_321 ();
 sg13g2_fill_2 FILLER_62_327 ();
 sg13g2_fill_2 FILLER_62_448 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_fill_2 FILLER_62_693 ();
 sg13g2_fill_2 FILLER_62_736 ();
 sg13g2_fill_1 FILLER_62_761 ();
 sg13g2_fill_1 FILLER_62_810 ();
 sg13g2_decap_4 FILLER_62_913 ();
 sg13g2_fill_2 FILLER_62_917 ();
 sg13g2_decap_4 FILLER_62_932 ();
 sg13g2_fill_2 FILLER_62_936 ();
 sg13g2_decap_8 FILLER_62_943 ();
 sg13g2_decap_8 FILLER_62_950 ();
 sg13g2_decap_8 FILLER_62_957 ();
 sg13g2_decap_8 FILLER_62_964 ();
 sg13g2_decap_8 FILLER_62_971 ();
 sg13g2_decap_8 FILLER_62_978 ();
 sg13g2_decap_4 FILLER_62_985 ();
 sg13g2_fill_2 FILLER_62_989 ();
 sg13g2_decap_8 FILLER_62_996 ();
 sg13g2_decap_4 FILLER_62_1003 ();
 sg13g2_fill_2 FILLER_62_1007 ();
 sg13g2_decap_8 FILLER_62_1018 ();
 sg13g2_decap_8 FILLER_62_1025 ();
 sg13g2_decap_8 FILLER_62_1032 ();
 sg13g2_decap_8 FILLER_62_1039 ();
 sg13g2_decap_8 FILLER_62_1046 ();
 sg13g2_decap_8 FILLER_62_1053 ();
 sg13g2_fill_1 FILLER_62_1060 ();
 sg13g2_fill_1 FILLER_62_1105 ();
 sg13g2_fill_2 FILLER_62_1133 ();
 sg13g2_fill_2 FILLER_62_1145 ();
 sg13g2_fill_1 FILLER_62_1147 ();
 sg13g2_fill_1 FILLER_62_1166 ();
 sg13g2_fill_2 FILLER_62_1195 ();
 sg13g2_fill_1 FILLER_62_1244 ();
 sg13g2_decap_4 FILLER_62_1268 ();
 sg13g2_fill_2 FILLER_62_1272 ();
 sg13g2_decap_4 FILLER_62_1277 ();
 sg13g2_fill_2 FILLER_62_1323 ();
 sg13g2_fill_2 FILLER_62_1392 ();
 sg13g2_fill_1 FILLER_62_1394 ();
 sg13g2_fill_1 FILLER_62_1417 ();
 sg13g2_fill_2 FILLER_62_1481 ();
 sg13g2_fill_1 FILLER_62_1483 ();
 sg13g2_fill_1 FILLER_62_1497 ();
 sg13g2_fill_2 FILLER_62_1526 ();
 sg13g2_fill_1 FILLER_62_1528 ();
 sg13g2_decap_8 FILLER_62_1559 ();
 sg13g2_fill_1 FILLER_62_1566 ();
 sg13g2_fill_1 FILLER_62_1571 ();
 sg13g2_fill_2 FILLER_62_1595 ();
 sg13g2_fill_1 FILLER_62_1597 ();
 sg13g2_fill_1 FILLER_62_1611 ();
 sg13g2_decap_8 FILLER_62_1629 ();
 sg13g2_fill_2 FILLER_62_1636 ();
 sg13g2_fill_1 FILLER_62_1638 ();
 sg13g2_fill_2 FILLER_62_1669 ();
 sg13g2_fill_1 FILLER_62_1671 ();
 sg13g2_decap_8 FILLER_62_1697 ();
 sg13g2_decap_8 FILLER_62_1714 ();
 sg13g2_decap_8 FILLER_62_1721 ();
 sg13g2_decap_8 FILLER_62_1728 ();
 sg13g2_fill_2 FILLER_62_1735 ();
 sg13g2_fill_2 FILLER_62_1747 ();
 sg13g2_fill_1 FILLER_62_1791 ();
 sg13g2_decap_8 FILLER_62_1841 ();
 sg13g2_decap_4 FILLER_62_1848 ();
 sg13g2_fill_1 FILLER_62_1852 ();
 sg13g2_fill_2 FILLER_62_1865 ();
 sg13g2_fill_1 FILLER_62_1867 ();
 sg13g2_decap_8 FILLER_62_1941 ();
 sg13g2_fill_1 FILLER_62_1948 ();
 sg13g2_decap_4 FILLER_62_2012 ();
 sg13g2_decap_8 FILLER_62_2029 ();
 sg13g2_fill_1 FILLER_62_2045 ();
 sg13g2_fill_1 FILLER_62_2069 ();
 sg13g2_fill_2 FILLER_62_2082 ();
 sg13g2_fill_2 FILLER_62_2106 ();
 sg13g2_decap_4 FILLER_62_2134 ();
 sg13g2_fill_1 FILLER_62_2138 ();
 sg13g2_fill_2 FILLER_62_2178 ();
 sg13g2_fill_1 FILLER_62_2180 ();
 sg13g2_fill_1 FILLER_62_2249 ();
 sg13g2_fill_2 FILLER_62_2304 ();
 sg13g2_fill_1 FILLER_62_2306 ();
 sg13g2_fill_1 FILLER_62_2321 ();
 sg13g2_fill_2 FILLER_62_2361 ();
 sg13g2_fill_1 FILLER_62_2363 ();
 sg13g2_fill_2 FILLER_62_2369 ();
 sg13g2_fill_1 FILLER_62_2371 ();
 sg13g2_decap_4 FILLER_62_2376 ();
 sg13g2_fill_1 FILLER_62_2380 ();
 sg13g2_fill_2 FILLER_62_2396 ();
 sg13g2_fill_1 FILLER_62_2398 ();
 sg13g2_fill_2 FILLER_62_2408 ();
 sg13g2_fill_1 FILLER_62_2436 ();
 sg13g2_decap_8 FILLER_62_2441 ();
 sg13g2_fill_2 FILLER_62_2448 ();
 sg13g2_fill_1 FILLER_62_2450 ();
 sg13g2_fill_2 FILLER_62_2481 ();
 sg13g2_fill_1 FILLER_62_2483 ();
 sg13g2_decap_8 FILLER_62_2530 ();
 sg13g2_decap_8 FILLER_62_2537 ();
 sg13g2_fill_1 FILLER_62_2557 ();
 sg13g2_fill_2 FILLER_62_2624 ();
 sg13g2_fill_2 FILLER_62_2631 ();
 sg13g2_fill_1 FILLER_62_2673 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_47 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_236 ();
 sg13g2_fill_2 FILLER_63_250 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_329 ();
 sg13g2_fill_1 FILLER_63_386 ();
 sg13g2_fill_1 FILLER_63_465 ();
 sg13g2_fill_2 FILLER_63_507 ();
 sg13g2_fill_1 FILLER_63_509 ();
 sg13g2_fill_2 FILLER_63_594 ();
 sg13g2_fill_1 FILLER_63_596 ();
 sg13g2_fill_2 FILLER_63_610 ();
 sg13g2_fill_1 FILLER_63_612 ();
 sg13g2_fill_1 FILLER_63_627 ();
 sg13g2_fill_1 FILLER_63_687 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_fill_1 FILLER_63_852 ();
 sg13g2_decap_8 FILLER_63_899 ();
 sg13g2_decap_4 FILLER_63_906 ();
 sg13g2_fill_2 FILLER_63_910 ();
 sg13g2_decap_8 FILLER_63_944 ();
 sg13g2_decap_4 FILLER_63_951 ();
 sg13g2_fill_1 FILLER_63_955 ();
 sg13g2_decap_8 FILLER_63_960 ();
 sg13g2_decap_8 FILLER_63_967 ();
 sg13g2_decap_4 FILLER_63_974 ();
 sg13g2_fill_2 FILLER_63_978 ();
 sg13g2_decap_8 FILLER_63_985 ();
 sg13g2_fill_1 FILLER_63_992 ();
 sg13g2_decap_8 FILLER_63_1000 ();
 sg13g2_decap_8 FILLER_63_1007 ();
 sg13g2_fill_2 FILLER_63_1014 ();
 sg13g2_fill_1 FILLER_63_1016 ();
 sg13g2_decap_8 FILLER_63_1022 ();
 sg13g2_decap_8 FILLER_63_1029 ();
 sg13g2_decap_8 FILLER_63_1036 ();
 sg13g2_decap_8 FILLER_63_1043 ();
 sg13g2_decap_8 FILLER_63_1050 ();
 sg13g2_decap_8 FILLER_63_1057 ();
 sg13g2_fill_1 FILLER_63_1064 ();
 sg13g2_fill_1 FILLER_63_1074 ();
 sg13g2_fill_1 FILLER_63_1090 ();
 sg13g2_fill_2 FILLER_63_1119 ();
 sg13g2_fill_2 FILLER_63_1134 ();
 sg13g2_fill_1 FILLER_63_1191 ();
 sg13g2_fill_2 FILLER_63_1233 ();
 sg13g2_fill_1 FILLER_63_1277 ();
 sg13g2_decap_4 FILLER_63_1282 ();
 sg13g2_fill_1 FILLER_63_1286 ();
 sg13g2_fill_1 FILLER_63_1315 ();
 sg13g2_decap_4 FILLER_63_1350 ();
 sg13g2_fill_2 FILLER_63_1354 ();
 sg13g2_decap_4 FILLER_63_1391 ();
 sg13g2_fill_2 FILLER_63_1395 ();
 sg13g2_decap_4 FILLER_63_1401 ();
 sg13g2_fill_1 FILLER_63_1409 ();
 sg13g2_decap_4 FILLER_63_1414 ();
 sg13g2_fill_1 FILLER_63_1418 ();
 sg13g2_fill_1 FILLER_63_1448 ();
 sg13g2_fill_2 FILLER_63_1468 ();
 sg13g2_decap_4 FILLER_63_1498 ();
 sg13g2_fill_2 FILLER_63_1524 ();
 sg13g2_fill_1 FILLER_63_1526 ();
 sg13g2_decap_4 FILLER_63_1565 ();
 sg13g2_fill_2 FILLER_63_1569 ();
 sg13g2_fill_2 FILLER_63_1576 ();
 sg13g2_fill_2 FILLER_63_1592 ();
 sg13g2_fill_2 FILLER_63_1615 ();
 sg13g2_fill_1 FILLER_63_1617 ();
 sg13g2_decap_8 FILLER_63_1636 ();
 sg13g2_fill_2 FILLER_63_1643 ();
 sg13g2_decap_4 FILLER_63_1660 ();
 sg13g2_fill_1 FILLER_63_1694 ();
 sg13g2_decap_8 FILLER_63_1721 ();
 sg13g2_decap_8 FILLER_63_1728 ();
 sg13g2_fill_2 FILLER_63_1808 ();
 sg13g2_fill_1 FILLER_63_1810 ();
 sg13g2_decap_8 FILLER_63_1815 ();
 sg13g2_decap_8 FILLER_63_1822 ();
 sg13g2_decap_8 FILLER_63_1829 ();
 sg13g2_decap_4 FILLER_63_1836 ();
 sg13g2_fill_1 FILLER_63_1840 ();
 sg13g2_fill_2 FILLER_63_1850 ();
 sg13g2_decap_4 FILLER_63_1856 ();
 sg13g2_decap_8 FILLER_63_1917 ();
 sg13g2_decap_8 FILLER_63_1937 ();
 sg13g2_decap_8 FILLER_63_1944 ();
 sg13g2_decap_4 FILLER_63_1951 ();
 sg13g2_fill_2 FILLER_63_1964 ();
 sg13g2_fill_2 FILLER_63_2042 ();
 sg13g2_fill_1 FILLER_63_2044 ();
 sg13g2_fill_2 FILLER_63_2081 ();
 sg13g2_fill_2 FILLER_63_2108 ();
 sg13g2_fill_1 FILLER_63_2110 ();
 sg13g2_fill_2 FILLER_63_2132 ();
 sg13g2_fill_2 FILLER_63_2173 ();
 sg13g2_fill_1 FILLER_63_2175 ();
 sg13g2_fill_2 FILLER_63_2189 ();
 sg13g2_fill_1 FILLER_63_2191 ();
 sg13g2_fill_2 FILLER_63_2202 ();
 sg13g2_fill_1 FILLER_63_2255 ();
 sg13g2_decap_4 FILLER_63_2295 ();
 sg13g2_fill_1 FILLER_63_2308 ();
 sg13g2_fill_1 FILLER_63_2315 ();
 sg13g2_fill_2 FILLER_63_2334 ();
 sg13g2_fill_1 FILLER_63_2336 ();
 sg13g2_decap_4 FILLER_63_2376 ();
 sg13g2_fill_2 FILLER_63_2380 ();
 sg13g2_fill_1 FILLER_63_2470 ();
 sg13g2_fill_1 FILLER_63_2498 ();
 sg13g2_fill_1 FILLER_63_2532 ();
 sg13g2_decap_4 FILLER_63_2538 ();
 sg13g2_fill_2 FILLER_63_2542 ();
 sg13g2_fill_2 FILLER_63_2550 ();
 sg13g2_fill_1 FILLER_63_2600 ();
 sg13g2_fill_2 FILLER_63_2628 ();
 sg13g2_fill_1 FILLER_63_2630 ();
 sg13g2_fill_2 FILLER_63_2635 ();
 sg13g2_fill_2 FILLER_63_2672 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_227 ();
 sg13g2_fill_2 FILLER_64_299 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_391 ();
 sg13g2_fill_2 FILLER_64_410 ();
 sg13g2_fill_1 FILLER_64_412 ();
 sg13g2_fill_2 FILLER_64_468 ();
 sg13g2_fill_1 FILLER_64_470 ();
 sg13g2_fill_1 FILLER_64_527 ();
 sg13g2_fill_2 FILLER_64_573 ();
 sg13g2_fill_1 FILLER_64_603 ();
 sg13g2_fill_2 FILLER_64_621 ();
 sg13g2_fill_1 FILLER_64_738 ();
 sg13g2_fill_2 FILLER_64_798 ();
 sg13g2_decap_8 FILLER_64_841 ();
 sg13g2_fill_1 FILLER_64_848 ();
 sg13g2_fill_2 FILLER_64_869 ();
 sg13g2_fill_1 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_64_904 ();
 sg13g2_decap_4 FILLER_64_911 ();
 sg13g2_fill_2 FILLER_64_920 ();
 sg13g2_fill_1 FILLER_64_922 ();
 sg13g2_decap_4 FILLER_64_936 ();
 sg13g2_fill_1 FILLER_64_940 ();
 sg13g2_decap_4 FILLER_64_951 ();
 sg13g2_fill_2 FILLER_64_955 ();
 sg13g2_fill_1 FILLER_64_961 ();
 sg13g2_decap_4 FILLER_64_970 ();
 sg13g2_fill_2 FILLER_64_974 ();
 sg13g2_decap_8 FILLER_64_995 ();
 sg13g2_decap_8 FILLER_64_1002 ();
 sg13g2_decap_4 FILLER_64_1009 ();
 sg13g2_fill_2 FILLER_64_1013 ();
 sg13g2_decap_8 FILLER_64_1033 ();
 sg13g2_decap_8 FILLER_64_1040 ();
 sg13g2_fill_2 FILLER_64_1047 ();
 sg13g2_fill_1 FILLER_64_1049 ();
 sg13g2_decap_8 FILLER_64_1058 ();
 sg13g2_decap_4 FILLER_64_1065 ();
 sg13g2_fill_1 FILLER_64_1069 ();
 sg13g2_fill_2 FILLER_64_1083 ();
 sg13g2_fill_1 FILLER_64_1094 ();
 sg13g2_fill_2 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1219 ();
 sg13g2_fill_1 FILLER_64_1278 ();
 sg13g2_decap_4 FILLER_64_1288 ();
 sg13g2_fill_1 FILLER_64_1292 ();
 sg13g2_decap_8 FILLER_64_1356 ();
 sg13g2_fill_1 FILLER_64_1363 ();
 sg13g2_decap_8 FILLER_64_1394 ();
 sg13g2_fill_1 FILLER_64_1401 ();
 sg13g2_fill_1 FILLER_64_1423 ();
 sg13g2_decap_8 FILLER_64_1449 ();
 sg13g2_fill_2 FILLER_64_1456 ();
 sg13g2_fill_1 FILLER_64_1458 ();
 sg13g2_decap_8 FILLER_64_1505 ();
 sg13g2_decap_8 FILLER_64_1512 ();
 sg13g2_fill_2 FILLER_64_1519 ();
 sg13g2_fill_1 FILLER_64_1521 ();
 sg13g2_fill_2 FILLER_64_1527 ();
 sg13g2_fill_1 FILLER_64_1529 ();
 sg13g2_decap_8 FILLER_64_1555 ();
 sg13g2_fill_2 FILLER_64_1566 ();
 sg13g2_fill_1 FILLER_64_1568 ();
 sg13g2_fill_1 FILLER_64_1574 ();
 sg13g2_fill_1 FILLER_64_1590 ();
 sg13g2_fill_2 FILLER_64_1605 ();
 sg13g2_fill_1 FILLER_64_1617 ();
 sg13g2_fill_2 FILLER_64_1629 ();
 sg13g2_fill_1 FILLER_64_1631 ();
 sg13g2_decap_8 FILLER_64_1641 ();
 sg13g2_fill_2 FILLER_64_1648 ();
 sg13g2_fill_2 FILLER_64_1654 ();
 sg13g2_decap_8 FILLER_64_1681 ();
 sg13g2_fill_1 FILLER_64_1688 ();
 sg13g2_decap_4 FILLER_64_1695 ();
 sg13g2_decap_8 FILLER_64_1706 ();
 sg13g2_decap_8 FILLER_64_1713 ();
 sg13g2_fill_2 FILLER_64_1725 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_decap_4 FILLER_64_1738 ();
 sg13g2_fill_2 FILLER_64_1742 ();
 sg13g2_fill_2 FILLER_64_1775 ();
 sg13g2_fill_2 FILLER_64_1791 ();
 sg13g2_fill_1 FILLER_64_1793 ();
 sg13g2_decap_8 FILLER_64_1821 ();
 sg13g2_fill_2 FILLER_64_1838 ();
 sg13g2_fill_1 FILLER_64_1840 ();
 sg13g2_fill_1 FILLER_64_1914 ();
 sg13g2_fill_1 FILLER_64_1928 ();
 sg13g2_fill_2 FILLER_64_1942 ();
 sg13g2_fill_1 FILLER_64_1944 ();
 sg13g2_fill_1 FILLER_64_1954 ();
 sg13g2_fill_2 FILLER_64_1959 ();
 sg13g2_fill_1 FILLER_64_1988 ();
 sg13g2_fill_1 FILLER_64_1998 ();
 sg13g2_fill_1 FILLER_64_2012 ();
 sg13g2_decap_8 FILLER_64_2044 ();
 sg13g2_fill_1 FILLER_64_2051 ();
 sg13g2_fill_1 FILLER_64_2056 ();
 sg13g2_fill_2 FILLER_64_2102 ();
 sg13g2_fill_1 FILLER_64_2104 ();
 sg13g2_decap_4 FILLER_64_2118 ();
 sg13g2_fill_1 FILLER_64_2131 ();
 sg13g2_fill_2 FILLER_64_2232 ();
 sg13g2_fill_2 FILLER_64_2271 ();
 sg13g2_fill_2 FILLER_64_2282 ();
 sg13g2_fill_1 FILLER_64_2284 ();
 sg13g2_fill_2 FILLER_64_2302 ();
 sg13g2_fill_1 FILLER_64_2350 ();
 sg13g2_decap_8 FILLER_64_2375 ();
 sg13g2_fill_2 FILLER_64_2422 ();
 sg13g2_fill_1 FILLER_64_2424 ();
 sg13g2_decap_4 FILLER_64_2452 ();
 sg13g2_fill_2 FILLER_64_2456 ();
 sg13g2_fill_1 FILLER_64_2476 ();
 sg13g2_fill_2 FILLER_64_2512 ();
 sg13g2_fill_1 FILLER_64_2514 ();
 sg13g2_fill_2 FILLER_64_2536 ();
 sg13g2_fill_1 FILLER_64_2550 ();
 sg13g2_fill_2 FILLER_64_2658 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_fill_1 FILLER_65_8 ();
 sg13g2_fill_2 FILLER_65_31 ();
 sg13g2_fill_1 FILLER_65_33 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_fill_2 FILLER_65_230 ();
 sg13g2_fill_2 FILLER_65_288 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_fill_2 FILLER_65_363 ();
 sg13g2_fill_2 FILLER_65_385 ();
 sg13g2_fill_1 FILLER_65_387 ();
 sg13g2_fill_2 FILLER_65_403 ();
 sg13g2_fill_1 FILLER_65_442 ();
 sg13g2_fill_2 FILLER_65_519 ();
 sg13g2_fill_1 FILLER_65_521 ();
 sg13g2_fill_2 FILLER_65_556 ();
 sg13g2_fill_1 FILLER_65_567 ();
 sg13g2_fill_1 FILLER_65_662 ();
 sg13g2_decap_4 FILLER_65_850 ();
 sg13g2_fill_2 FILLER_65_854 ();
 sg13g2_decap_8 FILLER_65_905 ();
 sg13g2_decap_8 FILLER_65_912 ();
 sg13g2_decap_8 FILLER_65_919 ();
 sg13g2_decap_8 FILLER_65_926 ();
 sg13g2_decap_8 FILLER_65_933 ();
 sg13g2_fill_2 FILLER_65_940 ();
 sg13g2_fill_1 FILLER_65_942 ();
 sg13g2_decap_8 FILLER_65_957 ();
 sg13g2_decap_8 FILLER_65_964 ();
 sg13g2_decap_4 FILLER_65_971 ();
 sg13g2_fill_2 FILLER_65_975 ();
 sg13g2_decap_8 FILLER_65_981 ();
 sg13g2_decap_8 FILLER_65_1001 ();
 sg13g2_fill_2 FILLER_65_1008 ();
 sg13g2_fill_1 FILLER_65_1010 ();
 sg13g2_decap_8 FILLER_65_1024 ();
 sg13g2_decap_8 FILLER_65_1031 ();
 sg13g2_fill_2 FILLER_65_1038 ();
 sg13g2_decap_8 FILLER_65_1049 ();
 sg13g2_decap_8 FILLER_65_1056 ();
 sg13g2_decap_8 FILLER_65_1063 ();
 sg13g2_decap_8 FILLER_65_1070 ();
 sg13g2_decap_4 FILLER_65_1077 ();
 sg13g2_fill_1 FILLER_65_1081 ();
 sg13g2_decap_4 FILLER_65_1097 ();
 sg13g2_fill_2 FILLER_65_1101 ();
 sg13g2_fill_1 FILLER_65_1177 ();
 sg13g2_fill_2 FILLER_65_1209 ();
 sg13g2_fill_1 FILLER_65_1211 ();
 sg13g2_fill_2 FILLER_65_1286 ();
 sg13g2_fill_2 FILLER_65_1297 ();
 sg13g2_fill_1 FILLER_65_1309 ();
 sg13g2_fill_2 FILLER_65_1315 ();
 sg13g2_decap_8 FILLER_65_1327 ();
 sg13g2_fill_1 FILLER_65_1334 ();
 sg13g2_decap_8 FILLER_65_1338 ();
 sg13g2_decap_8 FILLER_65_1345 ();
 sg13g2_decap_8 FILLER_65_1352 ();
 sg13g2_decap_8 FILLER_65_1359 ();
 sg13g2_decap_4 FILLER_65_1366 ();
 sg13g2_fill_1 FILLER_65_1370 ();
 sg13g2_decap_8 FILLER_65_1376 ();
 sg13g2_decap_8 FILLER_65_1383 ();
 sg13g2_fill_2 FILLER_65_1390 ();
 sg13g2_fill_2 FILLER_65_1432 ();
 sg13g2_fill_1 FILLER_65_1447 ();
 sg13g2_decap_4 FILLER_65_1452 ();
 sg13g2_decap_4 FILLER_65_1460 ();
 sg13g2_fill_1 FILLER_65_1521 ();
 sg13g2_decap_4 FILLER_65_1537 ();
 sg13g2_decap_4 FILLER_65_1595 ();
 sg13g2_fill_1 FILLER_65_1599 ();
 sg13g2_fill_2 FILLER_65_1614 ();
 sg13g2_decap_4 FILLER_65_1625 ();
 sg13g2_fill_1 FILLER_65_1629 ();
 sg13g2_fill_2 FILLER_65_1639 ();
 sg13g2_fill_1 FILLER_65_1641 ();
 sg13g2_fill_1 FILLER_65_1650 ();
 sg13g2_fill_2 FILLER_65_1665 ();
 sg13g2_fill_1 FILLER_65_1667 ();
 sg13g2_fill_2 FILLER_65_1707 ();
 sg13g2_fill_1 FILLER_65_1709 ();
 sg13g2_fill_2 FILLER_65_1745 ();
 sg13g2_fill_2 FILLER_65_1752 ();
 sg13g2_decap_4 FILLER_65_1767 ();
 sg13g2_fill_2 FILLER_65_1803 ();
 sg13g2_fill_1 FILLER_65_1805 ();
 sg13g2_fill_2 FILLER_65_1842 ();
 sg13g2_fill_1 FILLER_65_1854 ();
 sg13g2_fill_2 FILLER_65_1880 ();
 sg13g2_fill_1 FILLER_65_1882 ();
 sg13g2_decap_8 FILLER_65_1923 ();
 sg13g2_decap_8 FILLER_65_1930 ();
 sg13g2_fill_1 FILLER_65_1973 ();
 sg13g2_fill_2 FILLER_65_2023 ();
 sg13g2_fill_1 FILLER_65_2057 ();
 sg13g2_fill_2 FILLER_65_2083 ();
 sg13g2_fill_1 FILLER_65_2085 ();
 sg13g2_fill_1 FILLER_65_2130 ();
 sg13g2_fill_1 FILLER_65_2157 ();
 sg13g2_fill_2 FILLER_65_2207 ();
 sg13g2_fill_1 FILLER_65_2222 ();
 sg13g2_fill_2 FILLER_65_2236 ();
 sg13g2_fill_1 FILLER_65_2238 ();
 sg13g2_fill_1 FILLER_65_2244 ();
 sg13g2_fill_1 FILLER_65_2398 ();
 sg13g2_fill_2 FILLER_65_2417 ();
 sg13g2_fill_1 FILLER_65_2419 ();
 sg13g2_decap_8 FILLER_65_2460 ();
 sg13g2_decap_4 FILLER_65_2467 ();
 sg13g2_fill_2 FILLER_65_2503 ();
 sg13g2_fill_1 FILLER_65_2505 ();
 sg13g2_decap_4 FILLER_65_2530 ();
 sg13g2_fill_1 FILLER_65_2534 ();
 sg13g2_fill_2 FILLER_65_2563 ();
 sg13g2_fill_1 FILLER_65_2565 ();
 sg13g2_fill_2 FILLER_65_2606 ();
 sg13g2_fill_1 FILLER_65_2608 ();
 sg13g2_fill_2 FILLER_65_2622 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_43 ();
 sg13g2_fill_2 FILLER_66_68 ();
 sg13g2_fill_2 FILLER_66_75 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_fill_1 FILLER_66_106 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_fill_2 FILLER_66_334 ();
 sg13g2_fill_1 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_386 ();
 sg13g2_fill_1 FILLER_66_388 ();
 sg13g2_fill_2 FILLER_66_403 ();
 sg13g2_fill_2 FILLER_66_441 ();
 sg13g2_fill_1 FILLER_66_443 ();
 sg13g2_fill_2 FILLER_66_458 ();
 sg13g2_fill_1 FILLER_66_471 ();
 sg13g2_fill_1 FILLER_66_481 ();
 sg13g2_fill_2 FILLER_66_505 ();
 sg13g2_fill_1 FILLER_66_517 ();
 sg13g2_fill_2 FILLER_66_556 ();
 sg13g2_fill_1 FILLER_66_558 ();
 sg13g2_fill_1 FILLER_66_667 ();
 sg13g2_fill_2 FILLER_66_722 ();
 sg13g2_fill_2 FILLER_66_742 ();
 sg13g2_fill_1 FILLER_66_757 ();
 sg13g2_decap_4 FILLER_66_829 ();
 sg13g2_decap_4 FILLER_66_910 ();
 sg13g2_fill_1 FILLER_66_914 ();
 sg13g2_decap_4 FILLER_66_919 ();
 sg13g2_fill_1 FILLER_66_923 ();
 sg13g2_fill_2 FILLER_66_930 ();
 sg13g2_fill_1 FILLER_66_932 ();
 sg13g2_decap_4 FILLER_66_938 ();
 sg13g2_fill_2 FILLER_66_942 ();
 sg13g2_fill_2 FILLER_66_967 ();
 sg13g2_decap_8 FILLER_66_974 ();
 sg13g2_decap_8 FILLER_66_981 ();
 sg13g2_decap_4 FILLER_66_988 ();
 sg13g2_fill_1 FILLER_66_992 ();
 sg13g2_fill_2 FILLER_66_998 ();
 sg13g2_fill_1 FILLER_66_1000 ();
 sg13g2_decap_8 FILLER_66_1007 ();
 sg13g2_decap_4 FILLER_66_1014 ();
 sg13g2_fill_1 FILLER_66_1018 ();
 sg13g2_decap_8 FILLER_66_1026 ();
 sg13g2_decap_4 FILLER_66_1033 ();
 sg13g2_fill_1 FILLER_66_1037 ();
 sg13g2_decap_8 FILLER_66_1043 ();
 sg13g2_fill_1 FILLER_66_1050 ();
 sg13g2_decap_8 FILLER_66_1090 ();
 sg13g2_decap_8 FILLER_66_1097 ();
 sg13g2_decap_8 FILLER_66_1104 ();
 sg13g2_decap_8 FILLER_66_1116 ();
 sg13g2_decap_4 FILLER_66_1123 ();
 sg13g2_fill_1 FILLER_66_1127 ();
 sg13g2_fill_1 FILLER_66_1133 ();
 sg13g2_fill_2 FILLER_66_1160 ();
 sg13g2_fill_1 FILLER_66_1162 ();
 sg13g2_fill_1 FILLER_66_1226 ();
 sg13g2_fill_2 FILLER_66_1260 ();
 sg13g2_decap_4 FILLER_66_1300 ();
 sg13g2_fill_2 FILLER_66_1304 ();
 sg13g2_decap_8 FILLER_66_1340 ();
 sg13g2_decap_8 FILLER_66_1347 ();
 sg13g2_decap_4 FILLER_66_1354 ();
 sg13g2_fill_1 FILLER_66_1358 ();
 sg13g2_fill_1 FILLER_66_1384 ();
 sg13g2_fill_2 FILLER_66_1395 ();
 sg13g2_fill_1 FILLER_66_1397 ();
 sg13g2_decap_4 FILLER_66_1421 ();
 sg13g2_fill_1 FILLER_66_1425 ();
 sg13g2_fill_1 FILLER_66_1455 ();
 sg13g2_fill_2 FILLER_66_1466 ();
 sg13g2_fill_1 FILLER_66_1517 ();
 sg13g2_decap_8 FILLER_66_1561 ();
 sg13g2_fill_1 FILLER_66_1568 ();
 sg13g2_decap_8 FILLER_66_1589 ();
 sg13g2_fill_2 FILLER_66_1603 ();
 sg13g2_fill_2 FILLER_66_1609 ();
 sg13g2_fill_2 FILLER_66_1624 ();
 sg13g2_fill_1 FILLER_66_1626 ();
 sg13g2_fill_2 FILLER_66_1640 ();
 sg13g2_decap_8 FILLER_66_1678 ();
 sg13g2_fill_1 FILLER_66_1685 ();
 sg13g2_fill_1 FILLER_66_1691 ();
 sg13g2_fill_2 FILLER_66_1705 ();
 sg13g2_fill_1 FILLER_66_1707 ();
 sg13g2_fill_1 FILLER_66_1736 ();
 sg13g2_fill_2 FILLER_66_1840 ();
 sg13g2_fill_1 FILLER_66_1842 ();
 sg13g2_fill_2 FILLER_66_1882 ();
 sg13g2_fill_1 FILLER_66_1884 ();
 sg13g2_fill_1 FILLER_66_1936 ();
 sg13g2_fill_1 FILLER_66_1964 ();
 sg13g2_fill_2 FILLER_66_1984 ();
 sg13g2_fill_2 FILLER_66_2053 ();
 sg13g2_fill_2 FILLER_66_2189 ();
 sg13g2_fill_2 FILLER_66_2204 ();
 sg13g2_fill_2 FILLER_66_2219 ();
 sg13g2_fill_2 FILLER_66_2247 ();
 sg13g2_fill_1 FILLER_66_2249 ();
 sg13g2_fill_1 FILLER_66_2291 ();
 sg13g2_decap_8 FILLER_66_2305 ();
 sg13g2_decap_4 FILLER_66_2312 ();
 sg13g2_fill_2 FILLER_66_2316 ();
 sg13g2_fill_2 FILLER_66_2322 ();
 sg13g2_fill_2 FILLER_66_2339 ();
 sg13g2_fill_2 FILLER_66_2349 ();
 sg13g2_fill_1 FILLER_66_2351 ();
 sg13g2_fill_2 FILLER_66_2370 ();
 sg13g2_fill_2 FILLER_66_2403 ();
 sg13g2_fill_1 FILLER_66_2405 ();
 sg13g2_fill_1 FILLER_66_2464 ();
 sg13g2_fill_2 FILLER_66_2469 ();
 sg13g2_fill_1 FILLER_66_2471 ();
 sg13g2_fill_2 FILLER_66_2476 ();
 sg13g2_fill_1 FILLER_66_2478 ();
 sg13g2_fill_1 FILLER_66_2485 ();
 sg13g2_fill_2 FILLER_66_2492 ();
 sg13g2_fill_1 FILLER_66_2494 ();
 sg13g2_fill_2 FILLER_66_2504 ();
 sg13g2_fill_1 FILLER_66_2506 ();
 sg13g2_fill_1 FILLER_66_2541 ();
 sg13g2_fill_1 FILLER_66_2554 ();
 sg13g2_fill_2 FILLER_66_2589 ();
 sg13g2_fill_1 FILLER_66_2673 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_236 ();
 sg13g2_fill_2 FILLER_67_281 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_fill_2 FILLER_67_334 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_430 ();
 sg13g2_fill_1 FILLER_67_483 ();
 sg13g2_fill_1 FILLER_67_507 ();
 sg13g2_fill_2 FILLER_67_549 ();
 sg13g2_fill_1 FILLER_67_551 ();
 sg13g2_fill_2 FILLER_67_557 ();
 sg13g2_fill_1 FILLER_67_559 ();
 sg13g2_fill_2 FILLER_67_636 ();
 sg13g2_fill_2 FILLER_67_666 ();
 sg13g2_fill_2 FILLER_67_708 ();
 sg13g2_fill_1 FILLER_67_773 ();
 sg13g2_fill_2 FILLER_67_779 ();
 sg13g2_decap_4 FILLER_67_863 ();
 sg13g2_fill_2 FILLER_67_917 ();
 sg13g2_fill_2 FILLER_67_944 ();
 sg13g2_fill_2 FILLER_67_966 ();
 sg13g2_fill_2 FILLER_67_979 ();
 sg13g2_decap_8 FILLER_67_985 ();
 sg13g2_decap_4 FILLER_67_992 ();
 sg13g2_fill_1 FILLER_67_996 ();
 sg13g2_decap_4 FILLER_67_1005 ();
 sg13g2_fill_1 FILLER_67_1009 ();
 sg13g2_decap_8 FILLER_67_1021 ();
 sg13g2_decap_8 FILLER_67_1028 ();
 sg13g2_decap_8 FILLER_67_1035 ();
 sg13g2_fill_1 FILLER_67_1042 ();
 sg13g2_decap_4 FILLER_67_1056 ();
 sg13g2_fill_2 FILLER_67_1078 ();
 sg13g2_decap_8 FILLER_67_1109 ();
 sg13g2_decap_8 FILLER_67_1116 ();
 sg13g2_decap_8 FILLER_67_1123 ();
 sg13g2_fill_2 FILLER_67_1130 ();
 sg13g2_fill_2 FILLER_67_1145 ();
 sg13g2_fill_1 FILLER_67_1147 ();
 sg13g2_fill_1 FILLER_67_1171 ();
 sg13g2_fill_2 FILLER_67_1185 ();
 sg13g2_fill_2 FILLER_67_1205 ();
 sg13g2_fill_1 FILLER_67_1207 ();
 sg13g2_fill_2 FILLER_67_1217 ();
 sg13g2_fill_1 FILLER_67_1219 ();
 sg13g2_fill_2 FILLER_67_1248 ();
 sg13g2_fill_1 FILLER_67_1276 ();
 sg13g2_decap_4 FILLER_67_1352 ();
 sg13g2_fill_2 FILLER_67_1356 ();
 sg13g2_fill_2 FILLER_67_1409 ();
 sg13g2_fill_1 FILLER_67_1501 ();
 sg13g2_fill_2 FILLER_67_1539 ();
 sg13g2_decap_4 FILLER_67_1549 ();
 sg13g2_fill_2 FILLER_67_1558 ();
 sg13g2_decap_8 FILLER_67_1584 ();
 sg13g2_fill_2 FILLER_67_1591 ();
 sg13g2_fill_1 FILLER_67_1593 ();
 sg13g2_fill_1 FILLER_67_1617 ();
 sg13g2_fill_2 FILLER_67_1628 ();
 sg13g2_fill_1 FILLER_67_1630 ();
 sg13g2_fill_2 FILLER_67_1648 ();
 sg13g2_decap_8 FILLER_67_1691 ();
 sg13g2_fill_2 FILLER_67_1698 ();
 sg13g2_fill_1 FILLER_67_1700 ();
 sg13g2_fill_2 FILLER_67_1738 ();
 sg13g2_fill_1 FILLER_67_1740 ();
 sg13g2_fill_2 FILLER_67_1812 ();
 sg13g2_fill_2 FILLER_67_1893 ();
 sg13g2_fill_1 FILLER_67_1906 ();
 sg13g2_decap_8 FILLER_67_1934 ();
 sg13g2_fill_2 FILLER_67_1941 ();
 sg13g2_fill_1 FILLER_67_1943 ();
 sg13g2_fill_1 FILLER_67_1993 ();
 sg13g2_fill_1 FILLER_67_2044 ();
 sg13g2_fill_2 FILLER_67_2081 ();
 sg13g2_fill_1 FILLER_67_2098 ();
 sg13g2_fill_2 FILLER_67_2105 ();
 sg13g2_fill_1 FILLER_67_2134 ();
 sg13g2_fill_1 FILLER_67_2196 ();
 sg13g2_fill_2 FILLER_67_2202 ();
 sg13g2_fill_1 FILLER_67_2271 ();
 sg13g2_fill_2 FILLER_67_2295 ();
 sg13g2_fill_1 FILLER_67_2297 ();
 sg13g2_fill_1 FILLER_67_2315 ();
 sg13g2_fill_2 FILLER_67_2321 ();
 sg13g2_fill_1 FILLER_67_2323 ();
 sg13g2_fill_2 FILLER_67_2328 ();
 sg13g2_fill_2 FILLER_67_2343 ();
 sg13g2_fill_2 FILLER_67_2359 ();
 sg13g2_fill_1 FILLER_67_2425 ();
 sg13g2_fill_2 FILLER_67_2435 ();
 sg13g2_fill_1 FILLER_67_2437 ();
 sg13g2_fill_2 FILLER_67_2474 ();
 sg13g2_fill_1 FILLER_67_2481 ();
 sg13g2_fill_2 FILLER_67_2509 ();
 sg13g2_fill_2 FILLER_67_2547 ();
 sg13g2_fill_1 FILLER_67_2549 ();
 sg13g2_fill_2 FILLER_67_2643 ();
 sg13g2_fill_1 FILLER_67_2645 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_29 ();
 sg13g2_fill_1 FILLER_68_31 ();
 sg13g2_fill_2 FILLER_68_131 ();
 sg13g2_fill_2 FILLER_68_142 ();
 sg13g2_fill_2 FILLER_68_153 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_1 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_376 ();
 sg13g2_fill_1 FILLER_68_393 ();
 sg13g2_fill_2 FILLER_68_404 ();
 sg13g2_fill_1 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_417 ();
 sg13g2_fill_1 FILLER_68_598 ();
 sg13g2_fill_1 FILLER_68_773 ();
 sg13g2_fill_1 FILLER_68_871 ();
 sg13g2_decap_4 FILLER_68_890 ();
 sg13g2_decap_8 FILLER_68_907 ();
 sg13g2_decap_8 FILLER_68_914 ();
 sg13g2_decap_4 FILLER_68_921 ();
 sg13g2_fill_2 FILLER_68_925 ();
 sg13g2_fill_2 FILLER_68_945 ();
 sg13g2_fill_1 FILLER_68_961 ();
 sg13g2_fill_2 FILLER_68_972 ();
 sg13g2_fill_1 FILLER_68_980 ();
 sg13g2_fill_2 FILLER_68_994 ();
 sg13g2_fill_2 FILLER_68_1018 ();
 sg13g2_fill_1 FILLER_68_1020 ();
 sg13g2_decap_4 FILLER_68_1034 ();
 sg13g2_fill_1 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1070 ();
 sg13g2_fill_2 FILLER_68_1082 ();
 sg13g2_decap_4 FILLER_68_1090 ();
 sg13g2_decap_8 FILLER_68_1109 ();
 sg13g2_decap_8 FILLER_68_1116 ();
 sg13g2_decap_8 FILLER_68_1123 ();
 sg13g2_fill_1 FILLER_68_1130 ();
 sg13g2_fill_2 FILLER_68_1151 ();
 sg13g2_fill_1 FILLER_68_1153 ();
 sg13g2_fill_2 FILLER_68_1337 ();
 sg13g2_fill_2 FILLER_68_1394 ();
 sg13g2_fill_1 FILLER_68_1396 ();
 sg13g2_fill_2 FILLER_68_1471 ();
 sg13g2_fill_1 FILLER_68_1510 ();
 sg13g2_fill_2 FILLER_68_1544 ();
 sg13g2_fill_1 FILLER_68_1546 ();
 sg13g2_fill_1 FILLER_68_1552 ();
 sg13g2_fill_2 FILLER_68_1572 ();
 sg13g2_fill_1 FILLER_68_1574 ();
 sg13g2_fill_2 FILLER_68_1579 ();
 sg13g2_fill_1 FILLER_68_1585 ();
 sg13g2_fill_2 FILLER_68_1603 ();
 sg13g2_fill_2 FILLER_68_1622 ();
 sg13g2_fill_2 FILLER_68_1638 ();
 sg13g2_fill_1 FILLER_68_1645 ();
 sg13g2_fill_2 FILLER_68_1660 ();
 sg13g2_fill_2 FILLER_68_1666 ();
 sg13g2_fill_2 FILLER_68_1707 ();
 sg13g2_fill_2 FILLER_68_1746 ();
 sg13g2_fill_2 FILLER_68_1828 ();
 sg13g2_fill_1 FILLER_68_1830 ();
 sg13g2_decap_4 FILLER_68_1862 ();
 sg13g2_fill_2 FILLER_68_1866 ();
 sg13g2_decap_8 FILLER_68_1873 ();
 sg13g2_decap_4 FILLER_68_1880 ();
 sg13g2_fill_1 FILLER_68_1884 ();
 sg13g2_fill_2 FILLER_68_1895 ();
 sg13g2_fill_1 FILLER_68_1897 ();
 sg13g2_fill_1 FILLER_68_1910 ();
 sg13g2_decap_8 FILLER_68_1920 ();
 sg13g2_decap_8 FILLER_68_1927 ();
 sg13g2_fill_1 FILLER_68_1934 ();
 sg13g2_decap_4 FILLER_68_1986 ();
 sg13g2_decap_8 FILLER_68_1995 ();
 sg13g2_decap_8 FILLER_68_2002 ();
 sg13g2_decap_4 FILLER_68_2040 ();
 sg13g2_fill_2 FILLER_68_2044 ();
 sg13g2_fill_2 FILLER_68_2253 ();
 sg13g2_fill_1 FILLER_68_2268 ();
 sg13g2_fill_2 FILLER_68_2323 ();
 sg13g2_fill_2 FILLER_68_2379 ();
 sg13g2_fill_2 FILLER_68_2413 ();
 sg13g2_fill_1 FILLER_68_2415 ();
 sg13g2_fill_2 FILLER_68_2547 ();
 sg13g2_fill_1 FILLER_68_2549 ();
 sg13g2_fill_2 FILLER_68_2563 ();
 sg13g2_fill_2 FILLER_68_2584 ();
 sg13g2_fill_1 FILLER_68_2586 ();
 sg13g2_fill_1 FILLER_68_2616 ();
 sg13g2_fill_1 FILLER_68_2630 ();
 sg13g2_fill_2 FILLER_68_2672 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_73 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_166 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_304 ();
 sg13g2_fill_1 FILLER_69_318 ();
 sg13g2_fill_1 FILLER_69_333 ();
 sg13g2_fill_1 FILLER_69_437 ();
 sg13g2_fill_2 FILLER_69_443 ();
 sg13g2_fill_1 FILLER_69_476 ();
 sg13g2_fill_2 FILLER_69_528 ();
 sg13g2_fill_1 FILLER_69_572 ();
 sg13g2_fill_1 FILLER_69_586 ();
 sg13g2_fill_2 FILLER_69_666 ();
 sg13g2_fill_1 FILLER_69_682 ();
 sg13g2_fill_2 FILLER_69_720 ();
 sg13g2_fill_1 FILLER_69_746 ();
 sg13g2_fill_1 FILLER_69_756 ();
 sg13g2_fill_2 FILLER_69_817 ();
 sg13g2_fill_2 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_875 ();
 sg13g2_decap_8 FILLER_69_882 ();
 sg13g2_decap_8 FILLER_69_922 ();
 sg13g2_decap_4 FILLER_69_929 ();
 sg13g2_fill_2 FILLER_69_933 ();
 sg13g2_fill_2 FILLER_69_940 ();
 sg13g2_fill_1 FILLER_69_958 ();
 sg13g2_fill_1 FILLER_69_964 ();
 sg13g2_decap_8 FILLER_69_978 ();
 sg13g2_fill_1 FILLER_69_985 ();
 sg13g2_fill_2 FILLER_69_1002 ();
 sg13g2_decap_4 FILLER_69_1029 ();
 sg13g2_fill_2 FILLER_69_1055 ();
 sg13g2_decap_8 FILLER_69_1066 ();
 sg13g2_fill_1 FILLER_69_1073 ();
 sg13g2_decap_4 FILLER_69_1079 ();
 sg13g2_fill_1 FILLER_69_1097 ();
 sg13g2_decap_8 FILLER_69_1103 ();
 sg13g2_decap_8 FILLER_69_1110 ();
 sg13g2_decap_8 FILLER_69_1117 ();
 sg13g2_decap_8 FILLER_69_1124 ();
 sg13g2_fill_2 FILLER_69_1131 ();
 sg13g2_fill_2 FILLER_69_1141 ();
 sg13g2_fill_1 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1152 ();
 sg13g2_fill_2 FILLER_69_1159 ();
 sg13g2_fill_1 FILLER_69_1161 ();
 sg13g2_fill_1 FILLER_69_1213 ();
 sg13g2_fill_1 FILLER_69_1251 ();
 sg13g2_fill_2 FILLER_69_1304 ();
 sg13g2_fill_1 FILLER_69_1402 ();
 sg13g2_decap_8 FILLER_69_1446 ();
 sg13g2_decap_8 FILLER_69_1453 ();
 sg13g2_decap_8 FILLER_69_1460 ();
 sg13g2_fill_1 FILLER_69_1467 ();
 sg13g2_fill_2 FILLER_69_1499 ();
 sg13g2_fill_1 FILLER_69_1501 ();
 sg13g2_fill_2 FILLER_69_1540 ();
 sg13g2_fill_2 FILLER_69_1605 ();
 sg13g2_decap_8 FILLER_69_1634 ();
 sg13g2_decap_4 FILLER_69_1641 ();
 sg13g2_fill_1 FILLER_69_1645 ();
 sg13g2_fill_2 FILLER_69_1651 ();
 sg13g2_fill_1 FILLER_69_1653 ();
 sg13g2_fill_1 FILLER_69_1659 ();
 sg13g2_decap_8 FILLER_69_1677 ();
 sg13g2_fill_1 FILLER_69_1694 ();
 sg13g2_decap_8 FILLER_69_1699 ();
 sg13g2_decap_8 FILLER_69_1706 ();
 sg13g2_fill_2 FILLER_69_1713 ();
 sg13g2_fill_1 FILLER_69_1715 ();
 sg13g2_fill_1 FILLER_69_1743 ();
 sg13g2_fill_1 FILLER_69_1758 ();
 sg13g2_fill_2 FILLER_69_1764 ();
 sg13g2_fill_2 FILLER_69_1776 ();
 sg13g2_fill_1 FILLER_69_1778 ();
 sg13g2_decap_8 FILLER_69_1819 ();
 sg13g2_decap_8 FILLER_69_1826 ();
 sg13g2_decap_8 FILLER_69_1833 ();
 sg13g2_fill_2 FILLER_69_1844 ();
 sg13g2_fill_1 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1852 ();
 sg13g2_fill_1 FILLER_69_1854 ();
 sg13g2_fill_2 FILLER_69_1876 ();
 sg13g2_decap_8 FILLER_69_1882 ();
 sg13g2_fill_2 FILLER_69_1889 ();
 sg13g2_decap_8 FILLER_69_1928 ();
 sg13g2_decap_4 FILLER_69_1944 ();
 sg13g2_fill_2 FILLER_69_1948 ();
 sg13g2_decap_4 FILLER_69_1963 ();
 sg13g2_fill_2 FILLER_69_1985 ();
 sg13g2_fill_1 FILLER_69_2009 ();
 sg13g2_fill_1 FILLER_69_2016 ();
 sg13g2_fill_1 FILLER_69_2031 ();
 sg13g2_decap_8 FILLER_69_2041 ();
 sg13g2_decap_8 FILLER_69_2048 ();
 sg13g2_fill_1 FILLER_69_2055 ();
 sg13g2_fill_2 FILLER_69_2092 ();
 sg13g2_fill_2 FILLER_69_2105 ();
 sg13g2_fill_1 FILLER_69_2107 ();
 sg13g2_fill_1 FILLER_69_2176 ();
 sg13g2_fill_2 FILLER_69_2186 ();
 sg13g2_fill_2 FILLER_69_2198 ();
 sg13g2_fill_1 FILLER_69_2226 ();
 sg13g2_fill_2 FILLER_69_2267 ();
 sg13g2_fill_1 FILLER_69_2269 ();
 sg13g2_fill_1 FILLER_69_2288 ();
 sg13g2_fill_2 FILLER_69_2294 ();
 sg13g2_fill_1 FILLER_69_2296 ();
 sg13g2_fill_2 FILLER_69_2343 ();
 sg13g2_fill_1 FILLER_69_2345 ();
 sg13g2_fill_1 FILLER_69_2386 ();
 sg13g2_fill_2 FILLER_69_2392 ();
 sg13g2_fill_1 FILLER_69_2394 ();
 sg13g2_fill_2 FILLER_69_2431 ();
 sg13g2_fill_1 FILLER_69_2433 ();
 sg13g2_fill_2 FILLER_69_2447 ();
 sg13g2_fill_1 FILLER_69_2449 ();
 sg13g2_fill_2 FILLER_69_2463 ();
 sg13g2_fill_1 FILLER_69_2465 ();
 sg13g2_fill_1 FILLER_69_2484 ();
 sg13g2_fill_2 FILLER_69_2498 ();
 sg13g2_fill_2 FILLER_69_2540 ();
 sg13g2_fill_1 FILLER_69_2542 ();
 sg13g2_fill_2 FILLER_69_2556 ();
 sg13g2_fill_2 FILLER_69_2590 ();
 sg13g2_fill_1 FILLER_69_2625 ();
 sg13g2_fill_2 FILLER_69_2672 ();
 sg13g2_fill_1 FILLER_70_29 ();
 sg13g2_fill_2 FILLER_70_66 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_185 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_2 FILLER_70_259 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_295 ();
 sg13g2_fill_2 FILLER_70_311 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_340 ();
 sg13g2_fill_2 FILLER_70_408 ();
 sg13g2_fill_1 FILLER_70_410 ();
 sg13g2_fill_2 FILLER_70_474 ();
 sg13g2_fill_1 FILLER_70_476 ();
 sg13g2_fill_2 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_488 ();
 sg13g2_fill_1 FILLER_70_554 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_decap_8 FILLER_70_865 ();
 sg13g2_decap_8 FILLER_70_885 ();
 sg13g2_decap_4 FILLER_70_892 ();
 sg13g2_fill_1 FILLER_70_896 ();
 sg13g2_fill_1 FILLER_70_906 ();
 sg13g2_decap_8 FILLER_70_915 ();
 sg13g2_decap_4 FILLER_70_922 ();
 sg13g2_fill_2 FILLER_70_926 ();
 sg13g2_decap_8 FILLER_70_932 ();
 sg13g2_fill_2 FILLER_70_939 ();
 sg13g2_fill_1 FILLER_70_945 ();
 sg13g2_fill_2 FILLER_70_956 ();
 sg13g2_fill_2 FILLER_70_977 ();
 sg13g2_fill_1 FILLER_70_979 ();
 sg13g2_decap_4 FILLER_70_985 ();
 sg13g2_decap_4 FILLER_70_1015 ();
 sg13g2_fill_1 FILLER_70_1019 ();
 sg13g2_decap_4 FILLER_70_1048 ();
 sg13g2_decap_8 FILLER_70_1058 ();
 sg13g2_decap_8 FILLER_70_1065 ();
 sg13g2_decap_8 FILLER_70_1072 ();
 sg13g2_decap_8 FILLER_70_1079 ();
 sg13g2_decap_8 FILLER_70_1086 ();
 sg13g2_decap_8 FILLER_70_1093 ();
 sg13g2_decap_4 FILLER_70_1100 ();
 sg13g2_decap_8 FILLER_70_1109 ();
 sg13g2_decap_8 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_fill_2 FILLER_70_1137 ();
 sg13g2_fill_1 FILLER_70_1139 ();
 sg13g2_fill_2 FILLER_70_1147 ();
 sg13g2_fill_1 FILLER_70_1149 ();
 sg13g2_decap_4 FILLER_70_1159 ();
 sg13g2_fill_1 FILLER_70_1272 ();
 sg13g2_decap_8 FILLER_70_1360 ();
 sg13g2_fill_2 FILLER_70_1379 ();
 sg13g2_decap_4 FILLER_70_1436 ();
 sg13g2_fill_2 FILLER_70_1458 ();
 sg13g2_fill_1 FILLER_70_1460 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_fill_2 FILLER_70_1541 ();
 sg13g2_fill_2 FILLER_70_1567 ();
 sg13g2_fill_1 FILLER_70_1569 ();
 sg13g2_fill_2 FILLER_70_1588 ();
 sg13g2_decap_8 FILLER_70_1624 ();
 sg13g2_decap_8 FILLER_70_1631 ();
 sg13g2_fill_1 FILLER_70_1638 ();
 sg13g2_fill_1 FILLER_70_1654 ();
 sg13g2_fill_2 FILLER_70_1676 ();
 sg13g2_decap_4 FILLER_70_1714 ();
 sg13g2_fill_1 FILLER_70_1718 ();
 sg13g2_fill_1 FILLER_70_1747 ();
 sg13g2_fill_1 FILLER_70_1757 ();
 sg13g2_fill_1 FILLER_70_1834 ();
 sg13g2_fill_1 FILLER_70_1843 ();
 sg13g2_decap_4 FILLER_70_1884 ();
 sg13g2_fill_2 FILLER_70_1893 ();
 sg13g2_decap_8 FILLER_70_1946 ();
 sg13g2_fill_2 FILLER_70_1953 ();
 sg13g2_fill_2 FILLER_70_2003 ();
 sg13g2_fill_1 FILLER_70_2005 ();
 sg13g2_fill_2 FILLER_70_2012 ();
 sg13g2_fill_1 FILLER_70_2014 ();
 sg13g2_fill_2 FILLER_70_2021 ();
 sg13g2_fill_1 FILLER_70_2071 ();
 sg13g2_fill_1 FILLER_70_2077 ();
 sg13g2_fill_2 FILLER_70_2187 ();
 sg13g2_fill_1 FILLER_70_2189 ();
 sg13g2_fill_1 FILLER_70_2221 ();
 sg13g2_fill_2 FILLER_70_2227 ();
 sg13g2_fill_1 FILLER_70_2229 ();
 sg13g2_fill_1 FILLER_70_2252 ();
 sg13g2_fill_2 FILLER_70_2266 ();
 sg13g2_fill_1 FILLER_70_2268 ();
 sg13g2_fill_1 FILLER_70_2346 ();
 sg13g2_decap_4 FILLER_70_2360 ();
 sg13g2_fill_1 FILLER_70_2364 ();
 sg13g2_fill_1 FILLER_70_2404 ();
 sg13g2_fill_2 FILLER_70_2450 ();
 sg13g2_fill_1 FILLER_70_2452 ();
 sg13g2_fill_2 FILLER_70_2510 ();
 sg13g2_fill_1 FILLER_70_2512 ();
 sg13g2_fill_2 FILLER_70_2548 ();
 sg13g2_fill_2 FILLER_70_2559 ();
 sg13g2_fill_1 FILLER_70_2561 ();
 sg13g2_fill_1 FILLER_70_2639 ();
 sg13g2_fill_1 FILLER_70_2645 ();
 sg13g2_fill_2 FILLER_71_8 ();
 sg13g2_fill_1 FILLER_71_10 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_fill_2 FILLER_71_123 ();
 sg13g2_fill_2 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_fill_2 FILLER_71_326 ();
 sg13g2_fill_1 FILLER_71_328 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_fill_2 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_477 ();
 sg13g2_fill_1 FILLER_71_492 ();
 sg13g2_fill_2 FILLER_71_568 ();
 sg13g2_fill_1 FILLER_71_570 ();
 sg13g2_fill_2 FILLER_71_608 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_715 ();
 sg13g2_fill_2 FILLER_71_776 ();
 sg13g2_fill_1 FILLER_71_912 ();
 sg13g2_fill_2 FILLER_71_918 ();
 sg13g2_fill_1 FILLER_71_920 ();
 sg13g2_decap_8 FILLER_71_934 ();
 sg13g2_decap_8 FILLER_71_941 ();
 sg13g2_decap_4 FILLER_71_948 ();
 sg13g2_decap_4 FILLER_71_956 ();
 sg13g2_decap_4 FILLER_71_964 ();
 sg13g2_fill_1 FILLER_71_968 ();
 sg13g2_fill_1 FILLER_71_977 ();
 sg13g2_fill_2 FILLER_71_985 ();
 sg13g2_fill_1 FILLER_71_987 ();
 sg13g2_fill_2 FILLER_71_1003 ();
 sg13g2_fill_1 FILLER_71_1005 ();
 sg13g2_decap_8 FILLER_71_1052 ();
 sg13g2_decap_8 FILLER_71_1065 ();
 sg13g2_decap_8 FILLER_71_1072 ();
 sg13g2_decap_8 FILLER_71_1079 ();
 sg13g2_fill_1 FILLER_71_1086 ();
 sg13g2_decap_8 FILLER_71_1093 ();
 sg13g2_fill_2 FILLER_71_1100 ();
 sg13g2_decap_8 FILLER_71_1106 ();
 sg13g2_decap_8 FILLER_71_1113 ();
 sg13g2_decap_8 FILLER_71_1120 ();
 sg13g2_decap_4 FILLER_71_1127 ();
 sg13g2_fill_2 FILLER_71_1131 ();
 sg13g2_decap_8 FILLER_71_1138 ();
 sg13g2_decap_8 FILLER_71_1145 ();
 sg13g2_decap_8 FILLER_71_1152 ();
 sg13g2_decap_4 FILLER_71_1159 ();
 sg13g2_fill_2 FILLER_71_1168 ();
 sg13g2_fill_1 FILLER_71_1170 ();
 sg13g2_fill_1 FILLER_71_1252 ();
 sg13g2_fill_1 FILLER_71_1259 ();
 sg13g2_fill_1 FILLER_71_1310 ();
 sg13g2_fill_2 FILLER_71_1368 ();
 sg13g2_fill_1 FILLER_71_1407 ();
 sg13g2_decap_8 FILLER_71_1429 ();
 sg13g2_fill_1 FILLER_71_1436 ();
 sg13g2_fill_1 FILLER_71_1543 ();
 sg13g2_fill_1 FILLER_71_1613 ();
 sg13g2_fill_2 FILLER_71_1632 ();
 sg13g2_fill_1 FILLER_71_1634 ();
 sg13g2_fill_1 FILLER_71_1647 ();
 sg13g2_fill_2 FILLER_71_1666 ();
 sg13g2_fill_2 FILLER_71_1746 ();
 sg13g2_fill_2 FILLER_71_1767 ();
 sg13g2_fill_2 FILLER_71_1841 ();
 sg13g2_fill_2 FILLER_71_1885 ();
 sg13g2_fill_1 FILLER_71_1887 ();
 sg13g2_decap_8 FILLER_71_1938 ();
 sg13g2_decap_4 FILLER_71_1945 ();
 sg13g2_fill_1 FILLER_71_1984 ();
 sg13g2_decap_8 FILLER_71_2061 ();
 sg13g2_fill_2 FILLER_71_2068 ();
 sg13g2_decap_8 FILLER_71_2074 ();
 sg13g2_fill_1 FILLER_71_2081 ();
 sg13g2_fill_2 FILLER_71_2088 ();
 sg13g2_fill_1 FILLER_71_2090 ();
 sg13g2_fill_1 FILLER_71_2106 ();
 sg13g2_fill_2 FILLER_71_2165 ();
 sg13g2_fill_2 FILLER_71_2195 ();
 sg13g2_fill_2 FILLER_71_2261 ();
 sg13g2_fill_1 FILLER_71_2304 ();
 sg13g2_fill_1 FILLER_71_2318 ();
 sg13g2_fill_1 FILLER_71_2328 ();
 sg13g2_fill_1 FILLER_71_2364 ();
 sg13g2_fill_2 FILLER_71_2391 ();
 sg13g2_fill_1 FILLER_71_2406 ();
 sg13g2_fill_2 FILLER_71_2451 ();
 sg13g2_fill_1 FILLER_71_2453 ();
 sg13g2_fill_1 FILLER_71_2494 ();
 sg13g2_fill_1 FILLER_71_2513 ();
 sg13g2_fill_2 FILLER_71_2532 ();
 sg13g2_fill_2 FILLER_71_2551 ();
 sg13g2_fill_1 FILLER_71_2553 ();
 sg13g2_fill_2 FILLER_71_2581 ();
 sg13g2_fill_1 FILLER_71_2583 ();
 sg13g2_fill_2 FILLER_71_2620 ();
 sg13g2_fill_2 FILLER_71_2644 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_27 ();
 sg13g2_fill_2 FILLER_72_64 ();
 sg13g2_fill_2 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_102 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_2 FILLER_72_377 ();
 sg13g2_fill_2 FILLER_72_385 ();
 sg13g2_fill_1 FILLER_72_387 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_1 FILLER_72_436 ();
 sg13g2_fill_2 FILLER_72_457 ();
 sg13g2_fill_2 FILLER_72_464 ();
 sg13g2_fill_1 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_480 ();
 sg13g2_fill_2 FILLER_72_494 ();
 sg13g2_fill_1 FILLER_72_515 ();
 sg13g2_fill_2 FILLER_72_529 ();
 sg13g2_fill_1 FILLER_72_531 ();
 sg13g2_fill_1 FILLER_72_560 ();
 sg13g2_fill_2 FILLER_72_589 ();
 sg13g2_fill_2 FILLER_72_632 ();
 sg13g2_fill_1 FILLER_72_634 ();
 sg13g2_fill_1 FILLER_72_662 ();
 sg13g2_fill_1 FILLER_72_829 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_fill_2 FILLER_72_862 ();
 sg13g2_fill_1 FILLER_72_908 ();
 sg13g2_fill_2 FILLER_72_943 ();
 sg13g2_decap_4 FILLER_72_962 ();
 sg13g2_decap_8 FILLER_72_979 ();
 sg13g2_decap_4 FILLER_72_986 ();
 sg13g2_fill_2 FILLER_72_995 ();
 sg13g2_fill_1 FILLER_72_997 ();
 sg13g2_decap_4 FILLER_72_1008 ();
 sg13g2_fill_1 FILLER_72_1012 ();
 sg13g2_decap_4 FILLER_72_1022 ();
 sg13g2_fill_1 FILLER_72_1026 ();
 sg13g2_fill_2 FILLER_72_1047 ();
 sg13g2_fill_1 FILLER_72_1049 ();
 sg13g2_fill_2 FILLER_72_1054 ();
 sg13g2_fill_1 FILLER_72_1056 ();
 sg13g2_decap_8 FILLER_72_1071 ();
 sg13g2_fill_1 FILLER_72_1078 ();
 sg13g2_decap_8 FILLER_72_1084 ();
 sg13g2_decap_4 FILLER_72_1091 ();
 sg13g2_fill_2 FILLER_72_1095 ();
 sg13g2_fill_2 FILLER_72_1101 ();
 sg13g2_decap_8 FILLER_72_1116 ();
 sg13g2_decap_8 FILLER_72_1123 ();
 sg13g2_fill_2 FILLER_72_1130 ();
 sg13g2_fill_1 FILLER_72_1132 ();
 sg13g2_decap_4 FILLER_72_1138 ();
 sg13g2_decap_8 FILLER_72_1147 ();
 sg13g2_decap_8 FILLER_72_1154 ();
 sg13g2_decap_4 FILLER_72_1161 ();
 sg13g2_decap_8 FILLER_72_1170 ();
 sg13g2_fill_2 FILLER_72_1177 ();
 sg13g2_fill_2 FILLER_72_1241 ();
 sg13g2_fill_1 FILLER_72_1271 ();
 sg13g2_fill_2 FILLER_72_1407 ();
 sg13g2_fill_2 FILLER_72_1427 ();
 sg13g2_fill_1 FILLER_72_1433 ();
 sg13g2_fill_2 FILLER_72_1466 ();
 sg13g2_fill_1 FILLER_72_1468 ();
 sg13g2_fill_1 FILLER_72_1480 ();
 sg13g2_fill_2 FILLER_72_1534 ();
 sg13g2_fill_1 FILLER_72_1571 ();
 sg13g2_fill_2 FILLER_72_1582 ();
 sg13g2_fill_1 FILLER_72_1673 ();
 sg13g2_fill_1 FILLER_72_1741 ();
 sg13g2_fill_1 FILLER_72_1751 ();
 sg13g2_fill_1 FILLER_72_1792 ();
 sg13g2_fill_1 FILLER_72_1952 ();
 sg13g2_fill_2 FILLER_72_2061 ();
 sg13g2_fill_1 FILLER_72_2063 ();
 sg13g2_fill_2 FILLER_72_2077 ();
 sg13g2_fill_1 FILLER_72_2079 ();
 sg13g2_fill_2 FILLER_72_2125 ();
 sg13g2_fill_1 FILLER_72_2127 ();
 sg13g2_fill_2 FILLER_72_2169 ();
 sg13g2_fill_1 FILLER_72_2171 ();
 sg13g2_fill_1 FILLER_72_2194 ();
 sg13g2_fill_1 FILLER_72_2222 ();
 sg13g2_fill_2 FILLER_72_2227 ();
 sg13g2_fill_1 FILLER_72_2288 ();
 sg13g2_fill_1 FILLER_72_2326 ();
 sg13g2_fill_1 FILLER_72_2407 ();
 sg13g2_fill_2 FILLER_72_2449 ();
 sg13g2_fill_1 FILLER_72_2563 ();
 sg13g2_fill_1 FILLER_72_2645 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_56 ();
 sg13g2_fill_2 FILLER_73_152 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_318 ();
 sg13g2_fill_1 FILLER_73_320 ();
 sg13g2_fill_2 FILLER_73_359 ();
 sg13g2_fill_2 FILLER_73_380 ();
 sg13g2_fill_2 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_403 ();
 sg13g2_fill_1 FILLER_73_431 ();
 sg13g2_fill_1 FILLER_73_442 ();
 sg13g2_fill_2 FILLER_73_498 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_fill_2 FILLER_73_567 ();
 sg13g2_fill_1 FILLER_73_612 ();
 sg13g2_fill_1 FILLER_73_761 ();
 sg13g2_fill_2 FILLER_73_767 ();
 sg13g2_fill_1 FILLER_73_824 ();
 sg13g2_decap_8 FILLER_73_853 ();
 sg13g2_fill_1 FILLER_73_897 ();
 sg13g2_decap_4 FILLER_73_933 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_decap_8 FILLER_73_976 ();
 sg13g2_decap_8 FILLER_73_983 ();
 sg13g2_decap_8 FILLER_73_990 ();
 sg13g2_fill_2 FILLER_73_997 ();
 sg13g2_decap_8 FILLER_73_1028 ();
 sg13g2_decap_8 FILLER_73_1035 ();
 sg13g2_fill_1 FILLER_73_1042 ();
 sg13g2_decap_8 FILLER_73_1076 ();
 sg13g2_decap_8 FILLER_73_1083 ();
 sg13g2_fill_2 FILLER_73_1090 ();
 sg13g2_fill_1 FILLER_73_1102 ();
 sg13g2_fill_1 FILLER_73_1112 ();
 sg13g2_fill_1 FILLER_73_1127 ();
 sg13g2_fill_1 FILLER_73_1141 ();
 sg13g2_decap_4 FILLER_73_1153 ();
 sg13g2_decap_4 FILLER_73_1175 ();
 sg13g2_fill_2 FILLER_73_1179 ();
 sg13g2_fill_1 FILLER_73_1223 ();
 sg13g2_fill_1 FILLER_73_1247 ();
 sg13g2_fill_1 FILLER_73_1289 ();
 sg13g2_fill_1 FILLER_73_1318 ();
 sg13g2_fill_2 FILLER_73_1347 ();
 sg13g2_fill_2 FILLER_73_1358 ();
 sg13g2_fill_2 FILLER_73_1403 ();
 sg13g2_fill_1 FILLER_73_1405 ();
 sg13g2_fill_2 FILLER_73_1442 ();
 sg13g2_fill_1 FILLER_73_1444 ();
 sg13g2_fill_1 FILLER_73_1457 ();
 sg13g2_fill_1 FILLER_73_1472 ();
 sg13g2_fill_2 FILLER_73_1479 ();
 sg13g2_fill_2 FILLER_73_1494 ();
 sg13g2_fill_1 FILLER_73_1496 ();
 sg13g2_fill_1 FILLER_73_1539 ();
 sg13g2_fill_2 FILLER_73_1620 ();
 sg13g2_decap_4 FILLER_73_1632 ();
 sg13g2_fill_2 FILLER_73_1636 ();
 sg13g2_fill_2 FILLER_73_1691 ();
 sg13g2_fill_1 FILLER_73_1693 ();
 sg13g2_fill_1 FILLER_73_1735 ();
 sg13g2_fill_1 FILLER_73_1740 ();
 sg13g2_fill_1 FILLER_73_1745 ();
 sg13g2_fill_2 FILLER_73_1792 ();
 sg13g2_fill_1 FILLER_73_1794 ();
 sg13g2_fill_2 FILLER_73_1827 ();
 sg13g2_fill_1 FILLER_73_1829 ();
 sg13g2_fill_2 FILLER_73_1836 ();
 sg13g2_fill_2 FILLER_73_2014 ();
 sg13g2_fill_2 FILLER_73_2028 ();
 sg13g2_fill_1 FILLER_73_2030 ();
 sg13g2_fill_1 FILLER_73_2093 ();
 sg13g2_fill_2 FILLER_73_2145 ();
 sg13g2_fill_2 FILLER_73_2193 ();
 sg13g2_fill_1 FILLER_73_2325 ();
 sg13g2_fill_2 FILLER_73_2377 ();
 sg13g2_fill_1 FILLER_73_2379 ();
 sg13g2_fill_2 FILLER_73_2398 ();
 sg13g2_fill_2 FILLER_73_2450 ();
 sg13g2_fill_1 FILLER_73_2452 ();
 sg13g2_fill_2 FILLER_73_2503 ();
 sg13g2_fill_1 FILLER_73_2550 ();
 sg13g2_fill_2 FILLER_73_2583 ();
 sg13g2_fill_1 FILLER_73_2585 ();
 sg13g2_fill_2 FILLER_73_2608 ();
 sg13g2_fill_1 FILLER_74_31 ();
 sg13g2_fill_2 FILLER_74_45 ();
 sg13g2_fill_2 FILLER_74_158 ();
 sg13g2_fill_2 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_2 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_302 ();
 sg13g2_fill_2 FILLER_74_309 ();
 sg13g2_fill_1 FILLER_74_343 ();
 sg13g2_fill_2 FILLER_74_366 ();
 sg13g2_fill_1 FILLER_74_450 ();
 sg13g2_fill_1 FILLER_74_485 ();
 sg13g2_fill_2 FILLER_74_508 ();
 sg13g2_fill_1 FILLER_74_510 ();
 sg13g2_fill_2 FILLER_74_531 ();
 sg13g2_fill_1 FILLER_74_533 ();
 sg13g2_fill_1 FILLER_74_543 ();
 sg13g2_fill_2 FILLER_74_550 ();
 sg13g2_fill_1 FILLER_74_552 ();
 sg13g2_fill_2 FILLER_74_574 ();
 sg13g2_fill_1 FILLER_74_576 ();
 sg13g2_fill_2 FILLER_74_603 ();
 sg13g2_fill_1 FILLER_74_614 ();
 sg13g2_fill_1 FILLER_74_702 ();
 sg13g2_fill_2 FILLER_74_713 ();
 sg13g2_fill_1 FILLER_74_756 ();
 sg13g2_fill_1 FILLER_74_832 ();
 sg13g2_fill_2 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_74_881 ();
 sg13g2_fill_1 FILLER_74_883 ();
 sg13g2_decap_8 FILLER_74_900 ();
 sg13g2_decap_4 FILLER_74_907 ();
 sg13g2_fill_2 FILLER_74_931 ();
 sg13g2_decap_8 FILLER_74_937 ();
 sg13g2_fill_1 FILLER_74_944 ();
 sg13g2_decap_4 FILLER_74_964 ();
 sg13g2_decap_8 FILLER_74_976 ();
 sg13g2_decap_8 FILLER_74_983 ();
 sg13g2_decap_8 FILLER_74_990 ();
 sg13g2_fill_1 FILLER_74_997 ();
 sg13g2_decap_8 FILLER_74_1013 ();
 sg13g2_decap_8 FILLER_74_1020 ();
 sg13g2_decap_8 FILLER_74_1027 ();
 sg13g2_decap_8 FILLER_74_1034 ();
 sg13g2_decap_8 FILLER_74_1041 ();
 sg13g2_decap_8 FILLER_74_1048 ();
 sg13g2_decap_4 FILLER_74_1055 ();
 sg13g2_fill_1 FILLER_74_1059 ();
 sg13g2_decap_8 FILLER_74_1065 ();
 sg13g2_decap_8 FILLER_74_1072 ();
 sg13g2_decap_8 FILLER_74_1079 ();
 sg13g2_decap_4 FILLER_74_1086 ();
 sg13g2_decap_8 FILLER_74_1095 ();
 sg13g2_decap_8 FILLER_74_1102 ();
 sg13g2_decap_8 FILLER_74_1109 ();
 sg13g2_fill_2 FILLER_74_1120 ();
 sg13g2_fill_1 FILLER_74_1122 ();
 sg13g2_decap_8 FILLER_74_1138 ();
 sg13g2_fill_2 FILLER_74_1151 ();
 sg13g2_decap_8 FILLER_74_1162 ();
 sg13g2_decap_8 FILLER_74_1169 ();
 sg13g2_decap_4 FILLER_74_1176 ();
 sg13g2_fill_2 FILLER_74_1180 ();
 sg13g2_fill_2 FILLER_74_1226 ();
 sg13g2_fill_1 FILLER_74_1228 ();
 sg13g2_fill_2 FILLER_74_1270 ();
 sg13g2_fill_2 FILLER_74_1290 ();
 sg13g2_fill_1 FILLER_74_1292 ();
 sg13g2_fill_2 FILLER_74_1306 ();
 sg13g2_fill_1 FILLER_74_1378 ();
 sg13g2_decap_8 FILLER_74_1404 ();
 sg13g2_decap_4 FILLER_74_1411 ();
 sg13g2_fill_1 FILLER_74_1415 ();
 sg13g2_fill_1 FILLER_74_1445 ();
 sg13g2_fill_2 FILLER_74_1469 ();
 sg13g2_fill_2 FILLER_74_1497 ();
 sg13g2_fill_1 FILLER_74_1550 ();
 sg13g2_fill_1 FILLER_74_1569 ();
 sg13g2_decap_4 FILLER_74_1625 ();
 sg13g2_decap_4 FILLER_74_1675 ();
 sg13g2_fill_1 FILLER_74_1679 ();
 sg13g2_decap_8 FILLER_74_1735 ();
 sg13g2_fill_2 FILLER_74_1742 ();
 sg13g2_fill_1 FILLER_74_1744 ();
 sg13g2_decap_8 FILLER_74_1749 ();
 sg13g2_decap_4 FILLER_74_1756 ();
 sg13g2_fill_1 FILLER_74_1760 ();
 sg13g2_fill_1 FILLER_74_1828 ();
 sg13g2_decap_4 FILLER_74_1874 ();
 sg13g2_fill_1 FILLER_74_1878 ();
 sg13g2_decap_4 FILLER_74_1917 ();
 sg13g2_fill_2 FILLER_74_1921 ();
 sg13g2_fill_2 FILLER_74_1964 ();
 sg13g2_fill_2 FILLER_74_1986 ();
 sg13g2_fill_2 FILLER_74_2015 ();
 sg13g2_fill_2 FILLER_74_2059 ();
 sg13g2_fill_2 FILLER_74_2214 ();
 sg13g2_fill_1 FILLER_74_2216 ();
 sg13g2_decap_8 FILLER_74_2275 ();
 sg13g2_fill_1 FILLER_74_2282 ();
 sg13g2_fill_2 FILLER_74_2346 ();
 sg13g2_fill_1 FILLER_74_2348 ();
 sg13g2_fill_1 FILLER_74_2384 ();
 sg13g2_fill_2 FILLER_74_2422 ();
 sg13g2_fill_2 FILLER_74_2455 ();
 sg13g2_fill_1 FILLER_74_2457 ();
 sg13g2_fill_1 FILLER_74_2485 ();
 sg13g2_fill_1 FILLER_74_2528 ();
 sg13g2_fill_1 FILLER_74_2546 ();
 sg13g2_fill_1 FILLER_74_2589 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_68 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_192 ();
 sg13g2_fill_1 FILLER_75_194 ();
 sg13g2_fill_2 FILLER_75_311 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_1 FILLER_75_410 ();
 sg13g2_fill_2 FILLER_75_447 ();
 sg13g2_fill_2 FILLER_75_493 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_fill_2 FILLER_75_532 ();
 sg13g2_fill_1 FILLER_75_534 ();
 sg13g2_fill_2 FILLER_75_544 ();
 sg13g2_fill_2 FILLER_75_589 ();
 sg13g2_fill_2 FILLER_75_606 ();
 sg13g2_fill_1 FILLER_75_640 ();
 sg13g2_fill_1 FILLER_75_709 ();
 sg13g2_fill_1 FILLER_75_803 ();
 sg13g2_fill_2 FILLER_75_813 ();
 sg13g2_fill_1 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_decap_8 FILLER_75_855 ();
 sg13g2_decap_8 FILLER_75_862 ();
 sg13g2_decap_4 FILLER_75_869 ();
 sg13g2_fill_2 FILLER_75_873 ();
 sg13g2_fill_2 FILLER_75_888 ();
 sg13g2_fill_1 FILLER_75_890 ();
 sg13g2_decap_8 FILLER_75_897 ();
 sg13g2_decap_8 FILLER_75_904 ();
 sg13g2_decap_8 FILLER_75_911 ();
 sg13g2_decap_8 FILLER_75_918 ();
 sg13g2_fill_2 FILLER_75_925 ();
 sg13g2_fill_1 FILLER_75_927 ();
 sg13g2_decap_8 FILLER_75_940 ();
 sg13g2_decap_8 FILLER_75_947 ();
 sg13g2_fill_2 FILLER_75_954 ();
 sg13g2_decap_8 FILLER_75_960 ();
 sg13g2_fill_1 FILLER_75_967 ();
 sg13g2_decap_8 FILLER_75_979 ();
 sg13g2_decap_4 FILLER_75_986 ();
 sg13g2_fill_2 FILLER_75_990 ();
 sg13g2_decap_4 FILLER_75_997 ();
 sg13g2_fill_1 FILLER_75_1001 ();
 sg13g2_decap_8 FILLER_75_1007 ();
 sg13g2_decap_8 FILLER_75_1014 ();
 sg13g2_decap_8 FILLER_75_1021 ();
 sg13g2_fill_2 FILLER_75_1028 ();
 sg13g2_decap_8 FILLER_75_1043 ();
 sg13g2_decap_4 FILLER_75_1050 ();
 sg13g2_decap_8 FILLER_75_1060 ();
 sg13g2_decap_8 FILLER_75_1067 ();
 sg13g2_fill_2 FILLER_75_1074 ();
 sg13g2_fill_1 FILLER_75_1076 ();
 sg13g2_decap_4 FILLER_75_1101 ();
 sg13g2_decap_8 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1131 ();
 sg13g2_decap_8 FILLER_75_1138 ();
 sg13g2_fill_2 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1165 ();
 sg13g2_decap_8 FILLER_75_1172 ();
 sg13g2_fill_1 FILLER_75_1179 ();
 sg13g2_fill_2 FILLER_75_1268 ();
 sg13g2_fill_2 FILLER_75_1392 ();
 sg13g2_decap_8 FILLER_75_1404 ();
 sg13g2_fill_1 FILLER_75_1411 ();
 sg13g2_fill_2 FILLER_75_1444 ();
 sg13g2_fill_1 FILLER_75_1446 ();
 sg13g2_fill_1 FILLER_75_1482 ();
 sg13g2_fill_2 FILLER_75_1537 ();
 sg13g2_fill_1 FILLER_75_1539 ();
 sg13g2_fill_2 FILLER_75_1555 ();
 sg13g2_fill_1 FILLER_75_1557 ();
 sg13g2_fill_2 FILLER_75_1565 ();
 sg13g2_fill_1 FILLER_75_1567 ();
 sg13g2_fill_2 FILLER_75_1621 ();
 sg13g2_decap_8 FILLER_75_1647 ();
 sg13g2_decap_4 FILLER_75_1654 ();
 sg13g2_fill_2 FILLER_75_1663 ();
 sg13g2_fill_1 FILLER_75_1665 ();
 sg13g2_fill_1 FILLER_75_1675 ();
 sg13g2_fill_2 FILLER_75_1690 ();
 sg13g2_fill_2 FILLER_75_1709 ();
 sg13g2_fill_2 FILLER_75_1756 ();
 sg13g2_fill_1 FILLER_75_1758 ();
 sg13g2_fill_2 FILLER_75_1763 ();
 sg13g2_fill_1 FILLER_75_1840 ();
 sg13g2_fill_2 FILLER_75_1928 ();
 sg13g2_fill_1 FILLER_75_1930 ();
 sg13g2_fill_1 FILLER_75_1971 ();
 sg13g2_fill_2 FILLER_75_2022 ();
 sg13g2_fill_1 FILLER_75_2024 ();
 sg13g2_fill_1 FILLER_75_2045 ();
 sg13g2_fill_2 FILLER_75_2096 ();
 sg13g2_fill_1 FILLER_75_2098 ();
 sg13g2_fill_1 FILLER_75_2105 ();
 sg13g2_fill_1 FILLER_75_2115 ();
 sg13g2_fill_2 FILLER_75_2132 ();
 sg13g2_fill_2 FILLER_75_2194 ();
 sg13g2_fill_1 FILLER_75_2196 ();
 sg13g2_fill_2 FILLER_75_2225 ();
 sg13g2_fill_1 FILLER_75_2227 ();
 sg13g2_fill_1 FILLER_75_2282 ();
 sg13g2_fill_2 FILLER_75_2287 ();
 sg13g2_fill_1 FILLER_75_2289 ();
 sg13g2_fill_1 FILLER_75_2307 ();
 sg13g2_fill_2 FILLER_75_2341 ();
 sg13g2_fill_1 FILLER_75_2352 ();
 sg13g2_fill_2 FILLER_75_2385 ();
 sg13g2_fill_2 FILLER_75_2480 ();
 sg13g2_fill_2 FILLER_75_2537 ();
 sg13g2_fill_1 FILLER_75_2539 ();
 sg13g2_fill_2 FILLER_75_2639 ();
 sg13g2_fill_2 FILLER_75_2660 ();
 sg13g2_fill_2 FILLER_75_2671 ();
 sg13g2_fill_1 FILLER_75_2673 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_73 ();
 sg13g2_fill_1 FILLER_76_123 ();
 sg13g2_fill_2 FILLER_76_171 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_223 ();
 sg13g2_fill_1 FILLER_76_261 ();
 sg13g2_fill_2 FILLER_76_343 ();
 sg13g2_fill_1 FILLER_76_451 ();
 sg13g2_fill_1 FILLER_76_492 ();
 sg13g2_fill_2 FILLER_76_576 ();
 sg13g2_fill_1 FILLER_76_578 ();
 sg13g2_fill_1 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_793 ();
 sg13g2_fill_1 FILLER_76_826 ();
 sg13g2_decap_4 FILLER_76_857 ();
 sg13g2_fill_2 FILLER_76_861 ();
 sg13g2_fill_1 FILLER_76_869 ();
 sg13g2_decap_8 FILLER_76_874 ();
 sg13g2_decap_8 FILLER_76_881 ();
 sg13g2_decap_8 FILLER_76_901 ();
 sg13g2_decap_4 FILLER_76_908 ();
 sg13g2_decap_8 FILLER_76_916 ();
 sg13g2_decap_8 FILLER_76_923 ();
 sg13g2_decap_8 FILLER_76_930 ();
 sg13g2_fill_2 FILLER_76_937 ();
 sg13g2_decap_8 FILLER_76_945 ();
 sg13g2_decap_8 FILLER_76_952 ();
 sg13g2_fill_2 FILLER_76_959 ();
 sg13g2_fill_1 FILLER_76_961 ();
 sg13g2_fill_2 FILLER_76_981 ();
 sg13g2_fill_1 FILLER_76_983 ();
 sg13g2_decap_8 FILLER_76_989 ();
 sg13g2_fill_1 FILLER_76_1000 ();
 sg13g2_decap_8 FILLER_76_1011 ();
 sg13g2_decap_8 FILLER_76_1018 ();
 sg13g2_decap_4 FILLER_76_1025 ();
 sg13g2_fill_1 FILLER_76_1029 ();
 sg13g2_decap_4 FILLER_76_1043 ();
 sg13g2_fill_2 FILLER_76_1047 ();
 sg13g2_decap_8 FILLER_76_1063 ();
 sg13g2_decap_8 FILLER_76_1070 ();
 sg13g2_decap_4 FILLER_76_1077 ();
 sg13g2_fill_1 FILLER_76_1081 ();
 sg13g2_decap_8 FILLER_76_1090 ();
 sg13g2_decap_8 FILLER_76_1097 ();
 sg13g2_decap_4 FILLER_76_1104 ();
 sg13g2_decap_4 FILLER_76_1113 ();
 sg13g2_fill_1 FILLER_76_1117 ();
 sg13g2_decap_8 FILLER_76_1128 ();
 sg13g2_decap_8 FILLER_76_1135 ();
 sg13g2_decap_4 FILLER_76_1142 ();
 sg13g2_fill_2 FILLER_76_1151 ();
 sg13g2_fill_1 FILLER_76_1158 ();
 sg13g2_decap_8 FILLER_76_1165 ();
 sg13g2_decap_8 FILLER_76_1172 ();
 sg13g2_fill_2 FILLER_76_1179 ();
 sg13g2_fill_1 FILLER_76_1181 ();
 sg13g2_fill_2 FILLER_76_1282 ();
 sg13g2_decap_4 FILLER_76_1330 ();
 sg13g2_fill_1 FILLER_76_1334 ();
 sg13g2_decap_4 FILLER_76_1390 ();
 sg13g2_decap_8 FILLER_76_1399 ();
 sg13g2_fill_2 FILLER_76_1410 ();
 sg13g2_fill_1 FILLER_76_1412 ();
 sg13g2_fill_1 FILLER_76_1488 ();
 sg13g2_fill_2 FILLER_76_1516 ();
 sg13g2_decap_4 FILLER_76_1546 ();
 sg13g2_decap_4 FILLER_76_1635 ();
 sg13g2_fill_1 FILLER_76_1679 ();
 sg13g2_fill_1 FILLER_76_1704 ();
 sg13g2_fill_1 FILLER_76_1791 ();
 sg13g2_fill_2 FILLER_76_1838 ();
 sg13g2_fill_2 FILLER_76_1873 ();
 sg13g2_fill_1 FILLER_76_1897 ();
 sg13g2_fill_2 FILLER_76_1929 ();
 sg13g2_fill_2 FILLER_76_2008 ();
 sg13g2_fill_1 FILLER_76_2083 ();
 sg13g2_fill_1 FILLER_76_2089 ();
 sg13g2_fill_1 FILLER_76_2117 ();
 sg13g2_fill_2 FILLER_76_2154 ();
 sg13g2_fill_2 FILLER_76_2165 ();
 sg13g2_fill_1 FILLER_76_2167 ();
 sg13g2_fill_2 FILLER_76_2185 ();
 sg13g2_fill_1 FILLER_76_2187 ();
 sg13g2_fill_2 FILLER_76_2240 ();
 sg13g2_fill_1 FILLER_76_2264 ();
 sg13g2_fill_1 FILLER_76_2326 ();
 sg13g2_fill_2 FILLER_76_2433 ();
 sg13g2_fill_1 FILLER_76_2435 ();
 sg13g2_fill_2 FILLER_76_2449 ();
 sg13g2_fill_2 FILLER_76_2477 ();
 sg13g2_fill_1 FILLER_76_2510 ();
 sg13g2_fill_2 FILLER_76_2543 ();
 sg13g2_fill_1 FILLER_76_2545 ();
 sg13g2_fill_1 FILLER_76_2572 ();
 sg13g2_fill_2 FILLER_76_2600 ();
 sg13g2_fill_2 FILLER_76_2615 ();
 sg13g2_fill_1 FILLER_76_2617 ();
 sg13g2_fill_2 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_44 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_2 FILLER_77_410 ();
 sg13g2_fill_1 FILLER_77_564 ();
 sg13g2_fill_2 FILLER_77_602 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_fill_1 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_821 ();
 sg13g2_decap_4 FILLER_77_859 ();
 sg13g2_decap_4 FILLER_77_868 ();
 sg13g2_fill_2 FILLER_77_872 ();
 sg13g2_fill_2 FILLER_77_879 ();
 sg13g2_fill_1 FILLER_77_881 ();
 sg13g2_fill_2 FILLER_77_887 ();
 sg13g2_decap_4 FILLER_77_893 ();
 sg13g2_fill_1 FILLER_77_897 ();
 sg13g2_decap_8 FILLER_77_914 ();
 sg13g2_decap_8 FILLER_77_921 ();
 sg13g2_decap_8 FILLER_77_928 ();
 sg13g2_decap_8 FILLER_77_935 ();
 sg13g2_decap_8 FILLER_77_948 ();
 sg13g2_decap_8 FILLER_77_955 ();
 sg13g2_decap_4 FILLER_77_962 ();
 sg13g2_fill_2 FILLER_77_966 ();
 sg13g2_fill_2 FILLER_77_981 ();
 sg13g2_fill_1 FILLER_77_993 ();
 sg13g2_decap_8 FILLER_77_1014 ();
 sg13g2_decap_4 FILLER_77_1021 ();
 sg13g2_fill_2 FILLER_77_1025 ();
 sg13g2_decap_8 FILLER_77_1065 ();
 sg13g2_decap_8 FILLER_77_1072 ();
 sg13g2_decap_4 FILLER_77_1079 ();
 sg13g2_fill_2 FILLER_77_1083 ();
 sg13g2_decap_8 FILLER_77_1095 ();
 sg13g2_decap_8 FILLER_77_1102 ();
 sg13g2_fill_1 FILLER_77_1109 ();
 sg13g2_decap_8 FILLER_77_1115 ();
 sg13g2_decap_8 FILLER_77_1122 ();
 sg13g2_decap_8 FILLER_77_1129 ();
 sg13g2_decap_8 FILLER_77_1136 ();
 sg13g2_decap_8 FILLER_77_1143 ();
 sg13g2_decap_4 FILLER_77_1150 ();
 sg13g2_fill_2 FILLER_77_1154 ();
 sg13g2_decap_8 FILLER_77_1169 ();
 sg13g2_decap_8 FILLER_77_1176 ();
 sg13g2_fill_2 FILLER_77_1183 ();
 sg13g2_fill_2 FILLER_77_1229 ();
 sg13g2_decap_4 FILLER_77_1328 ();
 sg13g2_fill_1 FILLER_77_1342 ();
 sg13g2_fill_2 FILLER_77_1373 ();
 sg13g2_fill_2 FILLER_77_1398 ();
 sg13g2_fill_1 FILLER_77_1455 ();
 sg13g2_decap_8 FILLER_77_1460 ();
 sg13g2_fill_2 FILLER_77_1467 ();
 sg13g2_fill_1 FILLER_77_1469 ();
 sg13g2_decap_4 FILLER_77_1552 ();
 sg13g2_fill_1 FILLER_77_1556 ();
 sg13g2_decap_4 FILLER_77_1566 ();
 sg13g2_fill_1 FILLER_77_1570 ();
 sg13g2_fill_1 FILLER_77_1581 ();
 sg13g2_decap_4 FILLER_77_1647 ();
 sg13g2_fill_1 FILLER_77_1707 ();
 sg13g2_fill_1 FILLER_77_1804 ();
 sg13g2_fill_1 FILLER_77_1881 ();
 sg13g2_fill_2 FILLER_77_1918 ();
 sg13g2_fill_1 FILLER_77_1920 ();
 sg13g2_decap_4 FILLER_77_1930 ();
 sg13g2_fill_2 FILLER_77_1966 ();
 sg13g2_fill_1 FILLER_77_1981 ();
 sg13g2_fill_2 FILLER_77_1995 ();
 sg13g2_fill_2 FILLER_77_2010 ();
 sg13g2_fill_1 FILLER_77_2048 ();
 sg13g2_fill_2 FILLER_77_2104 ();
 sg13g2_fill_1 FILLER_77_2106 ();
 sg13g2_fill_2 FILLER_77_2139 ();
 sg13g2_fill_2 FILLER_77_2181 ();
 sg13g2_fill_1 FILLER_77_2183 ();
 sg13g2_fill_1 FILLER_77_2274 ();
 sg13g2_fill_1 FILLER_77_2326 ();
 sg13g2_fill_2 FILLER_77_2378 ();
 sg13g2_fill_2 FILLER_77_2408 ();
 sg13g2_fill_2 FILLER_77_2443 ();
 sg13g2_fill_1 FILLER_77_2445 ();
 sg13g2_fill_1 FILLER_77_2507 ();
 sg13g2_fill_2 FILLER_77_2616 ();
 sg13g2_fill_1 FILLER_77_2673 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_29 ();
 sg13g2_fill_1 FILLER_78_50 ();
 sg13g2_fill_2 FILLER_78_93 ();
 sg13g2_fill_2 FILLER_78_131 ();
 sg13g2_fill_1 FILLER_78_187 ();
 sg13g2_fill_1 FILLER_78_215 ();
 sg13g2_fill_2 FILLER_78_276 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_fill_1 FILLER_78_424 ();
 sg13g2_fill_1 FILLER_78_456 ();
 sg13g2_fill_1 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_727 ();
 sg13g2_decap_8 FILLER_78_865 ();
 sg13g2_decap_8 FILLER_78_872 ();
 sg13g2_fill_1 FILLER_78_879 ();
 sg13g2_fill_2 FILLER_78_889 ();
 sg13g2_decap_8 FILLER_78_915 ();
 sg13g2_decap_4 FILLER_78_922 ();
 sg13g2_fill_2 FILLER_78_926 ();
 sg13g2_decap_8 FILLER_78_950 ();
 sg13g2_decap_8 FILLER_78_957 ();
 sg13g2_decap_8 FILLER_78_964 ();
 sg13g2_decap_4 FILLER_78_971 ();
 sg13g2_fill_1 FILLER_78_979 ();
 sg13g2_fill_2 FILLER_78_994 ();
 sg13g2_fill_2 FILLER_78_1000 ();
 sg13g2_decap_4 FILLER_78_1025 ();
 sg13g2_fill_1 FILLER_78_1029 ();
 sg13g2_decap_4 FILLER_78_1040 ();
 sg13g2_fill_2 FILLER_78_1044 ();
 sg13g2_fill_2 FILLER_78_1051 ();
 sg13g2_decap_8 FILLER_78_1064 ();
 sg13g2_decap_4 FILLER_78_1101 ();
 sg13g2_fill_2 FILLER_78_1105 ();
 sg13g2_fill_1 FILLER_78_1111 ();
 sg13g2_decap_8 FILLER_78_1135 ();
 sg13g2_decap_8 FILLER_78_1142 ();
 sg13g2_decap_8 FILLER_78_1149 ();
 sg13g2_fill_2 FILLER_78_1156 ();
 sg13g2_fill_1 FILLER_78_1162 ();
 sg13g2_decap_8 FILLER_78_1174 ();
 sg13g2_decap_8 FILLER_78_1181 ();
 sg13g2_fill_2 FILLER_78_1315 ();
 sg13g2_decap_4 FILLER_78_1372 ();
 sg13g2_fill_2 FILLER_78_1430 ();
 sg13g2_fill_2 FILLER_78_1459 ();
 sg13g2_fill_2 FILLER_78_1561 ();
 sg13g2_fill_2 FILLER_78_1591 ();
 sg13g2_fill_1 FILLER_78_1593 ();
 sg13g2_fill_1 FILLER_78_1625 ();
 sg13g2_fill_2 FILLER_78_1666 ();
 sg13g2_fill_1 FILLER_78_1668 ();
 sg13g2_fill_2 FILLER_78_1758 ();
 sg13g2_fill_1 FILLER_78_1760 ();
 sg13g2_fill_1 FILLER_78_1794 ();
 sg13g2_fill_2 FILLER_78_1822 ();
 sg13g2_decap_8 FILLER_78_1910 ();
 sg13g2_decap_8 FILLER_78_1917 ();
 sg13g2_fill_2 FILLER_78_2050 ();
 sg13g2_fill_1 FILLER_78_2065 ();
 sg13g2_fill_2 FILLER_78_2098 ();
 sg13g2_fill_1 FILLER_78_2100 ();
 sg13g2_fill_1 FILLER_78_2110 ();
 sg13g2_fill_1 FILLER_78_2151 ();
 sg13g2_fill_1 FILLER_78_2184 ();
 sg13g2_fill_2 FILLER_78_2226 ();
 sg13g2_fill_2 FILLER_78_2261 ();
 sg13g2_fill_1 FILLER_78_2263 ();
 sg13g2_fill_1 FILLER_78_2292 ();
 sg13g2_fill_2 FILLER_78_2334 ();
 sg13g2_fill_1 FILLER_78_2336 ();
 sg13g2_fill_2 FILLER_78_2375 ();
 sg13g2_fill_2 FILLER_78_2390 ();
 sg13g2_fill_1 FILLER_78_2433 ();
 sg13g2_fill_1 FILLER_78_2511 ();
 sg13g2_fill_2 FILLER_78_2549 ();
 sg13g2_fill_2 FILLER_78_2672 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_150 ();
 sg13g2_fill_1 FILLER_79_201 ();
 sg13g2_fill_1 FILLER_79_229 ();
 sg13g2_fill_2 FILLER_79_366 ();
 sg13g2_fill_2 FILLER_79_513 ();
 sg13g2_fill_1 FILLER_79_543 ();
 sg13g2_fill_1 FILLER_79_577 ();
 sg13g2_fill_1 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_652 ();
 sg13g2_fill_2 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_8 FILLER_79_869 ();
 sg13g2_decap_8 FILLER_79_876 ();
 sg13g2_decap_4 FILLER_79_883 ();
 sg13g2_fill_1 FILLER_79_887 ();
 sg13g2_decap_8 FILLER_79_891 ();
 sg13g2_decap_8 FILLER_79_898 ();
 sg13g2_decap_8 FILLER_79_905 ();
 sg13g2_decap_8 FILLER_79_912 ();
 sg13g2_decap_8 FILLER_79_919 ();
 sg13g2_decap_8 FILLER_79_926 ();
 sg13g2_decap_8 FILLER_79_933 ();
 sg13g2_decap_8 FILLER_79_940 ();
 sg13g2_decap_8 FILLER_79_947 ();
 sg13g2_decap_8 FILLER_79_954 ();
 sg13g2_decap_8 FILLER_79_961 ();
 sg13g2_decap_8 FILLER_79_968 ();
 sg13g2_decap_8 FILLER_79_975 ();
 sg13g2_decap_8 FILLER_79_982 ();
 sg13g2_fill_2 FILLER_79_989 ();
 sg13g2_decap_8 FILLER_79_995 ();
 sg13g2_decap_8 FILLER_79_1002 ();
 sg13g2_decap_8 FILLER_79_1009 ();
 sg13g2_decap_8 FILLER_79_1016 ();
 sg13g2_decap_8 FILLER_79_1023 ();
 sg13g2_decap_4 FILLER_79_1030 ();
 sg13g2_fill_2 FILLER_79_1034 ();
 sg13g2_decap_8 FILLER_79_1041 ();
 sg13g2_decap_8 FILLER_79_1048 ();
 sg13g2_decap_8 FILLER_79_1055 ();
 sg13g2_decap_8 FILLER_79_1062 ();
 sg13g2_decap_8 FILLER_79_1069 ();
 sg13g2_decap_8 FILLER_79_1076 ();
 sg13g2_decap_8 FILLER_79_1083 ();
 sg13g2_fill_1 FILLER_79_1090 ();
 sg13g2_decap_8 FILLER_79_1095 ();
 sg13g2_decap_8 FILLER_79_1102 ();
 sg13g2_decap_8 FILLER_79_1109 ();
 sg13g2_decap_4 FILLER_79_1116 ();
 sg13g2_decap_8 FILLER_79_1129 ();
 sg13g2_decap_8 FILLER_79_1136 ();
 sg13g2_decap_8 FILLER_79_1143 ();
 sg13g2_decap_8 FILLER_79_1150 ();
 sg13g2_decap_8 FILLER_79_1157 ();
 sg13g2_decap_8 FILLER_79_1164 ();
 sg13g2_decap_8 FILLER_79_1171 ();
 sg13g2_decap_8 FILLER_79_1178 ();
 sg13g2_decap_8 FILLER_79_1185 ();
 sg13g2_decap_4 FILLER_79_1192 ();
 sg13g2_fill_1 FILLER_79_1251 ();
 sg13g2_fill_1 FILLER_79_1284 ();
 sg13g2_decap_4 FILLER_79_1341 ();
 sg13g2_decap_8 FILLER_79_1373 ();
 sg13g2_fill_1 FILLER_79_1380 ();
 sg13g2_fill_2 FILLER_79_1394 ();
 sg13g2_fill_2 FILLER_79_1452 ();
 sg13g2_fill_2 FILLER_79_1467 ();
 sg13g2_decap_8 FILLER_79_1519 ();
 sg13g2_fill_2 FILLER_79_1526 ();
 sg13g2_decap_4 FILLER_79_1566 ();
 sg13g2_fill_2 FILLER_79_1570 ();
 sg13g2_decap_4 FILLER_79_1613 ();
 sg13g2_fill_1 FILLER_79_1617 ();
 sg13g2_fill_1 FILLER_79_1717 ();
 sg13g2_fill_1 FILLER_79_1751 ();
 sg13g2_fill_2 FILLER_79_1785 ();
 sg13g2_fill_1 FILLER_79_1787 ();
 sg13g2_fill_1 FILLER_79_1864 ();
 sg13g2_fill_2 FILLER_79_1893 ();
 sg13g2_fill_2 FILLER_79_1904 ();
 sg13g2_fill_1 FILLER_79_1906 ();
 sg13g2_decap_8 FILLER_79_1916 ();
 sg13g2_decap_8 FILLER_79_1923 ();
 sg13g2_fill_1 FILLER_79_1930 ();
 sg13g2_fill_2 FILLER_79_1985 ();
 sg13g2_fill_1 FILLER_79_1987 ();
 sg13g2_decap_4 FILLER_79_1997 ();
 sg13g2_fill_1 FILLER_79_2044 ();
 sg13g2_fill_2 FILLER_79_2072 ();
 sg13g2_fill_2 FILLER_79_2082 ();
 sg13g2_fill_2 FILLER_79_2124 ();
 sg13g2_fill_1 FILLER_79_2126 ();
 sg13g2_fill_2 FILLER_79_2140 ();
 sg13g2_fill_2 FILLER_79_2288 ();
 sg13g2_fill_2 FILLER_79_2331 ();
 sg13g2_fill_2 FILLER_79_2379 ();
 sg13g2_fill_2 FILLER_79_2385 ();
 sg13g2_fill_1 FILLER_79_2387 ();
 sg13g2_fill_1 FILLER_79_2451 ();
 sg13g2_fill_2 FILLER_79_2482 ();
 sg13g2_fill_1 FILLER_79_2484 ();
 sg13g2_fill_1 FILLER_79_2513 ();
 sg13g2_fill_2 FILLER_79_2519 ();
 sg13g2_fill_1 FILLER_79_2521 ();
 sg13g2_fill_2 FILLER_79_2596 ();
 sg13g2_fill_2 FILLER_79_2672 ();
 sg13g2_fill_2 FILLER_80_127 ();
 sg13g2_fill_2 FILLER_80_143 ();
 sg13g2_fill_1 FILLER_80_145 ();
 sg13g2_fill_1 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_381 ();
 sg13g2_fill_2 FILLER_80_409 ();
 sg13g2_fill_1 FILLER_80_432 ();
 sg13g2_fill_2 FILLER_80_447 ();
 sg13g2_fill_1 FILLER_80_449 ();
 sg13g2_fill_2 FILLER_80_511 ();
 sg13g2_fill_1 FILLER_80_566 ();
 sg13g2_fill_2 FILLER_80_576 ();
 sg13g2_fill_1 FILLER_80_578 ();
 sg13g2_fill_2 FILLER_80_644 ();
 sg13g2_fill_1 FILLER_80_728 ();
 sg13g2_fill_2 FILLER_80_752 ();
 sg13g2_fill_2 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_870 ();
 sg13g2_decap_8 FILLER_80_877 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_898 ();
 sg13g2_decap_8 FILLER_80_905 ();
 sg13g2_decap_8 FILLER_80_912 ();
 sg13g2_decap_8 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_933 ();
 sg13g2_decap_8 FILLER_80_940 ();
 sg13g2_decap_8 FILLER_80_947 ();
 sg13g2_decap_8 FILLER_80_954 ();
 sg13g2_decap_8 FILLER_80_961 ();
 sg13g2_decap_8 FILLER_80_968 ();
 sg13g2_decap_8 FILLER_80_975 ();
 sg13g2_decap_8 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_decap_8 FILLER_80_1003 ();
 sg13g2_decap_8 FILLER_80_1010 ();
 sg13g2_decap_8 FILLER_80_1017 ();
 sg13g2_decap_8 FILLER_80_1024 ();
 sg13g2_decap_8 FILLER_80_1031 ();
 sg13g2_decap_8 FILLER_80_1038 ();
 sg13g2_decap_8 FILLER_80_1045 ();
 sg13g2_decap_8 FILLER_80_1052 ();
 sg13g2_decap_8 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_decap_8 FILLER_80_1073 ();
 sg13g2_decap_8 FILLER_80_1080 ();
 sg13g2_decap_8 FILLER_80_1087 ();
 sg13g2_decap_8 FILLER_80_1094 ();
 sg13g2_decap_8 FILLER_80_1101 ();
 sg13g2_decap_8 FILLER_80_1108 ();
 sg13g2_decap_8 FILLER_80_1115 ();
 sg13g2_decap_8 FILLER_80_1122 ();
 sg13g2_decap_8 FILLER_80_1129 ();
 sg13g2_decap_8 FILLER_80_1136 ();
 sg13g2_decap_8 FILLER_80_1143 ();
 sg13g2_decap_8 FILLER_80_1150 ();
 sg13g2_decap_8 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1171 ();
 sg13g2_decap_8 FILLER_80_1178 ();
 sg13g2_decap_8 FILLER_80_1185 ();
 sg13g2_decap_8 FILLER_80_1192 ();
 sg13g2_fill_2 FILLER_80_1199 ();
 sg13g2_fill_2 FILLER_80_1214 ();
 sg13g2_fill_1 FILLER_80_1216 ();
 sg13g2_fill_2 FILLER_80_1248 ();
 sg13g2_fill_2 FILLER_80_1286 ();
 sg13g2_fill_2 FILLER_80_1312 ();
 sg13g2_fill_2 FILLER_80_1326 ();
 sg13g2_fill_1 FILLER_80_1328 ();
 sg13g2_fill_1 FILLER_80_1338 ();
 sg13g2_decap_4 FILLER_80_1357 ();
 sg13g2_fill_1 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1408 ();
 sg13g2_fill_2 FILLER_80_1415 ();
 sg13g2_decap_8 FILLER_80_1430 ();
 sg13g2_decap_8 FILLER_80_1437 ();
 sg13g2_decap_8 FILLER_80_1444 ();
 sg13g2_decap_4 FILLER_80_1451 ();
 sg13g2_fill_2 FILLER_80_1455 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_fill_2 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1512 ();
 sg13g2_decap_8 FILLER_80_1519 ();
 sg13g2_fill_2 FILLER_80_1526 ();
 sg13g2_decap_4 FILLER_80_1550 ();
 sg13g2_fill_1 FILLER_80_1554 ();
 sg13g2_fill_2 FILLER_80_1591 ();
 sg13g2_fill_2 FILLER_80_1602 ();
 sg13g2_fill_1 FILLER_80_1604 ();
 sg13g2_decap_8 FILLER_80_1614 ();
 sg13g2_decap_8 FILLER_80_1621 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_4 FILLER_80_1649 ();
 sg13g2_fill_2 FILLER_80_1653 ();
 sg13g2_decap_8 FILLER_80_1668 ();
 sg13g2_decap_8 FILLER_80_1675 ();
 sg13g2_decap_8 FILLER_80_1682 ();
 sg13g2_fill_2 FILLER_80_1689 ();
 sg13g2_fill_1 FILLER_80_1700 ();
 sg13g2_fill_1 FILLER_80_1718 ();
 sg13g2_fill_1 FILLER_80_1776 ();
 sg13g2_fill_2 FILLER_80_1803 ();
 sg13g2_fill_1 FILLER_80_1805 ();
 sg13g2_fill_2 FILLER_80_1820 ();
 sg13g2_fill_1 FILLER_80_1822 ();
 sg13g2_fill_2 FILLER_80_1832 ();
 sg13g2_fill_1 FILLER_80_1839 ();
 sg13g2_fill_2 FILLER_80_1864 ();
 sg13g2_fill_1 FILLER_80_1892 ();
 sg13g2_decap_8 FILLER_80_1902 ();
 sg13g2_decap_8 FILLER_80_1909 ();
 sg13g2_decap_8 FILLER_80_1916 ();
 sg13g2_decap_8 FILLER_80_1923 ();
 sg13g2_decap_8 FILLER_80_1930 ();
 sg13g2_decap_8 FILLER_80_1937 ();
 sg13g2_fill_2 FILLER_80_1944 ();
 sg13g2_fill_2 FILLER_80_1950 ();
 sg13g2_fill_1 FILLER_80_1952 ();
 sg13g2_fill_1 FILLER_80_1962 ();
 sg13g2_fill_2 FILLER_80_1971 ();
 sg13g2_decap_8 FILLER_80_1986 ();
 sg13g2_decap_8 FILLER_80_1993 ();
 sg13g2_decap_8 FILLER_80_2000 ();
 sg13g2_decap_8 FILLER_80_2007 ();
 sg13g2_decap_4 FILLER_80_2023 ();
 sg13g2_fill_1 FILLER_80_2027 ();
 sg13g2_decap_8 FILLER_80_2037 ();
 sg13g2_fill_1 FILLER_80_2044 ();
 sg13g2_decap_8 FILLER_80_2071 ();
 sg13g2_decap_4 FILLER_80_2078 ();
 sg13g2_fill_2 FILLER_80_2082 ();
 sg13g2_fill_1 FILLER_80_2088 ();
 sg13g2_fill_2 FILLER_80_2120 ();
 sg13g2_fill_2 FILLER_80_2144 ();
 sg13g2_fill_1 FILLER_80_2146 ();
 sg13g2_fill_1 FILLER_80_2151 ();
 sg13g2_fill_2 FILLER_80_2157 ();
 sg13g2_fill_2 FILLER_80_2181 ();
 sg13g2_fill_1 FILLER_80_2213 ();
 sg13g2_fill_2 FILLER_80_2223 ();
 sg13g2_fill_1 FILLER_80_2225 ();
 sg13g2_fill_2 FILLER_80_2299 ();
 sg13g2_fill_1 FILLER_80_2354 ();
 sg13g2_decap_8 FILLER_80_2377 ();
 sg13g2_fill_2 FILLER_80_2384 ();
 sg13g2_fill_1 FILLER_80_2386 ();
 sg13g2_fill_2 FILLER_80_2450 ();
 sg13g2_fill_1 FILLER_80_2470 ();
 sg13g2_fill_1 FILLER_80_2511 ();
 sg13g2_fill_1 FILLER_80_2529 ();
 sg13g2_fill_1 FILLER_80_2539 ();
 sg13g2_fill_1 FILLER_80_2583 ();
 sg13g2_fill_2 FILLER_80_2588 ();
 sg13g2_fill_1 FILLER_80_2634 ();
 sg13g2_fill_2 FILLER_80_2643 ();
 sg13g2_fill_2 FILLER_80_2672 ();
 assign uio_oe[0] = net77;
 assign uio_oe[3] = net78;
 assign uio_oe[6] = net79;
endmodule
