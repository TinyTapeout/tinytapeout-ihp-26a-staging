module tt_um_mlyoung_wedgetail (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire net64;
 wire _024_;
 wire net65;
 wire _026_;
 wire net66;
 wire _028_;
 wire net67;
 wire _030_;
 wire net68;
 wire _032_;
 wire net69;
 wire _034_;
 wire net70;
 wire _036_;
 wire clk_regs;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire \dpll.clk8x_fout ;
 wire \dpll.clk_fout ;
 wire \dpll.id_decrement ;
 wire \dpll.id_decrement_done ;
 wire \dpll.id_increment ;
 wire \dpll.id_increment_done ;
 wire \dpll.id_out ;
 wire \dpll.k_count[0] ;
 wire \dpll.k_count[1] ;
 wire \dpll.k_count[2] ;
 wire \dpll.k_count[3] ;
 wire \dpll.k_count[4] ;
 wire \dpll.k_count[5] ;
 wire \dpll.k_count[6] ;
 wire \dpll.k_count[7] ;
 wire \dpll.k_count_borrow ;
 wire \dpll.k_count_carry ;
 wire \dpll.n_count[0] ;
 wire \dpll.n_count[1] ;
 wire \dpll.n_count[2] ;
 wire \dpll.n_count[4] ;
 wire \dpll.n_count[5] ;
 wire \mod_ro_128.fabric[0] ;
 wire \mod_ro_128.fabric[100] ;
 wire \mod_ro_128.fabric[101] ;
 wire \mod_ro_128.fabric[102] ;
 wire \mod_ro_128.fabric[103] ;
 wire \mod_ro_128.fabric[104] ;
 wire \mod_ro_128.fabric[105] ;
 wire \mod_ro_128.fabric[106] ;
 wire \mod_ro_128.fabric[107] ;
 wire \mod_ro_128.fabric[108] ;
 wire \mod_ro_128.fabric[109] ;
 wire \mod_ro_128.fabric[10] ;
 wire \mod_ro_128.fabric[110] ;
 wire \mod_ro_128.fabric[111] ;
 wire \mod_ro_128.fabric[112] ;
 wire \mod_ro_128.fabric[113] ;
 wire \mod_ro_128.fabric[114] ;
 wire \mod_ro_128.fabric[115] ;
 wire \mod_ro_128.fabric[116] ;
 wire \mod_ro_128.fabric[117] ;
 wire \mod_ro_128.fabric[118] ;
 wire \mod_ro_128.fabric[119] ;
 wire \mod_ro_128.fabric[11] ;
 wire \mod_ro_128.fabric[120] ;
 wire \mod_ro_128.fabric[121] ;
 wire \mod_ro_128.fabric[122] ;
 wire \mod_ro_128.fabric[123] ;
 wire \mod_ro_128.fabric[124] ;
 wire \mod_ro_128.fabric[125] ;
 wire \mod_ro_128.fabric[126] ;
 wire \mod_ro_128.fabric[127] ;
 wire \mod_ro_128.fabric[128] ;
 wire \mod_ro_128.fabric[12] ;
 wire \mod_ro_128.fabric[13] ;
 wire \mod_ro_128.fabric[14] ;
 wire \mod_ro_128.fabric[15] ;
 wire \mod_ro_128.fabric[16] ;
 wire \mod_ro_128.fabric[17] ;
 wire \mod_ro_128.fabric[18] ;
 wire \mod_ro_128.fabric[19] ;
 wire \mod_ro_128.fabric[1] ;
 wire \mod_ro_128.fabric[20] ;
 wire \mod_ro_128.fabric[21] ;
 wire \mod_ro_128.fabric[22] ;
 wire \mod_ro_128.fabric[23] ;
 wire \mod_ro_128.fabric[24] ;
 wire \mod_ro_128.fabric[25] ;
 wire \mod_ro_128.fabric[26] ;
 wire \mod_ro_128.fabric[27] ;
 wire \mod_ro_128.fabric[28] ;
 wire \mod_ro_128.fabric[29] ;
 wire \mod_ro_128.fabric[2] ;
 wire \mod_ro_128.fabric[30] ;
 wire \mod_ro_128.fabric[31] ;
 wire \mod_ro_128.fabric[32] ;
 wire \mod_ro_128.fabric[33] ;
 wire \mod_ro_128.fabric[34] ;
 wire \mod_ro_128.fabric[35] ;
 wire \mod_ro_128.fabric[36] ;
 wire \mod_ro_128.fabric[37] ;
 wire \mod_ro_128.fabric[38] ;
 wire \mod_ro_128.fabric[39] ;
 wire \mod_ro_128.fabric[3] ;
 wire \mod_ro_128.fabric[40] ;
 wire \mod_ro_128.fabric[41] ;
 wire \mod_ro_128.fabric[42] ;
 wire \mod_ro_128.fabric[43] ;
 wire \mod_ro_128.fabric[44] ;
 wire \mod_ro_128.fabric[45] ;
 wire \mod_ro_128.fabric[46] ;
 wire \mod_ro_128.fabric[47] ;
 wire \mod_ro_128.fabric[48] ;
 wire \mod_ro_128.fabric[49] ;
 wire \mod_ro_128.fabric[4] ;
 wire \mod_ro_128.fabric[50] ;
 wire \mod_ro_128.fabric[51] ;
 wire \mod_ro_128.fabric[52] ;
 wire \mod_ro_128.fabric[53] ;
 wire \mod_ro_128.fabric[54] ;
 wire \mod_ro_128.fabric[55] ;
 wire \mod_ro_128.fabric[56] ;
 wire \mod_ro_128.fabric[57] ;
 wire \mod_ro_128.fabric[58] ;
 wire \mod_ro_128.fabric[59] ;
 wire \mod_ro_128.fabric[5] ;
 wire \mod_ro_128.fabric[60] ;
 wire \mod_ro_128.fabric[61] ;
 wire \mod_ro_128.fabric[62] ;
 wire \mod_ro_128.fabric[63] ;
 wire \mod_ro_128.fabric[64] ;
 wire \mod_ro_128.fabric[65] ;
 wire \mod_ro_128.fabric[66] ;
 wire \mod_ro_128.fabric[67] ;
 wire \mod_ro_128.fabric[68] ;
 wire \mod_ro_128.fabric[69] ;
 wire \mod_ro_128.fabric[6] ;
 wire \mod_ro_128.fabric[70] ;
 wire \mod_ro_128.fabric[71] ;
 wire \mod_ro_128.fabric[72] ;
 wire \mod_ro_128.fabric[73] ;
 wire \mod_ro_128.fabric[74] ;
 wire \mod_ro_128.fabric[75] ;
 wire \mod_ro_128.fabric[76] ;
 wire \mod_ro_128.fabric[77] ;
 wire \mod_ro_128.fabric[78] ;
 wire \mod_ro_128.fabric[79] ;
 wire \mod_ro_128.fabric[7] ;
 wire \mod_ro_128.fabric[80] ;
 wire \mod_ro_128.fabric[81] ;
 wire \mod_ro_128.fabric[82] ;
 wire \mod_ro_128.fabric[83] ;
 wire \mod_ro_128.fabric[84] ;
 wire \mod_ro_128.fabric[85] ;
 wire \mod_ro_128.fabric[86] ;
 wire \mod_ro_128.fabric[87] ;
 wire \mod_ro_128.fabric[88] ;
 wire \mod_ro_128.fabric[89] ;
 wire \mod_ro_128.fabric[8] ;
 wire \mod_ro_128.fabric[90] ;
 wire \mod_ro_128.fabric[91] ;
 wire \mod_ro_128.fabric[92] ;
 wire \mod_ro_128.fabric[93] ;
 wire \mod_ro_128.fabric[94] ;
 wire \mod_ro_128.fabric[95] ;
 wire \mod_ro_128.fabric[96] ;
 wire \mod_ro_128.fabric[97] ;
 wire \mod_ro_128.fabric[98] ;
 wire \mod_ro_128.fabric[99] ;
 wire \mod_ro_128.fabric[9] ;
 wire \mod_ro_16.fabric[0] ;
 wire \mod_ro_16.fabric[10] ;
 wire \mod_ro_16.fabric[11] ;
 wire \mod_ro_16.fabric[12] ;
 wire \mod_ro_16.fabric[13] ;
 wire \mod_ro_16.fabric[14] ;
 wire \mod_ro_16.fabric[15] ;
 wire \mod_ro_16.fabric[16] ;
 wire \mod_ro_16.fabric[1] ;
 wire \mod_ro_16.fabric[2] ;
 wire \mod_ro_16.fabric[3] ;
 wire \mod_ro_16.fabric[4] ;
 wire \mod_ro_16.fabric[5] ;
 wire \mod_ro_16.fabric[6] ;
 wire \mod_ro_16.fabric[7] ;
 wire \mod_ro_16.fabric[8] ;
 wire \mod_ro_16.fabric[9] ;
 wire \mod_ro_256.fabric[0] ;
 wire \mod_ro_256.fabric[100] ;
 wire \mod_ro_256.fabric[101] ;
 wire \mod_ro_256.fabric[102] ;
 wire \mod_ro_256.fabric[103] ;
 wire \mod_ro_256.fabric[104] ;
 wire \mod_ro_256.fabric[105] ;
 wire \mod_ro_256.fabric[106] ;
 wire \mod_ro_256.fabric[107] ;
 wire \mod_ro_256.fabric[108] ;
 wire \mod_ro_256.fabric[109] ;
 wire \mod_ro_256.fabric[10] ;
 wire \mod_ro_256.fabric[110] ;
 wire \mod_ro_256.fabric[111] ;
 wire \mod_ro_256.fabric[112] ;
 wire \mod_ro_256.fabric[113] ;
 wire \mod_ro_256.fabric[114] ;
 wire \mod_ro_256.fabric[115] ;
 wire \mod_ro_256.fabric[116] ;
 wire \mod_ro_256.fabric[117] ;
 wire \mod_ro_256.fabric[118] ;
 wire \mod_ro_256.fabric[119] ;
 wire \mod_ro_256.fabric[11] ;
 wire \mod_ro_256.fabric[120] ;
 wire \mod_ro_256.fabric[121] ;
 wire \mod_ro_256.fabric[122] ;
 wire \mod_ro_256.fabric[123] ;
 wire \mod_ro_256.fabric[124] ;
 wire \mod_ro_256.fabric[125] ;
 wire \mod_ro_256.fabric[126] ;
 wire \mod_ro_256.fabric[127] ;
 wire \mod_ro_256.fabric[128] ;
 wire \mod_ro_256.fabric[129] ;
 wire \mod_ro_256.fabric[12] ;
 wire \mod_ro_256.fabric[130] ;
 wire \mod_ro_256.fabric[131] ;
 wire \mod_ro_256.fabric[132] ;
 wire \mod_ro_256.fabric[133] ;
 wire \mod_ro_256.fabric[134] ;
 wire \mod_ro_256.fabric[135] ;
 wire \mod_ro_256.fabric[136] ;
 wire \mod_ro_256.fabric[137] ;
 wire \mod_ro_256.fabric[138] ;
 wire \mod_ro_256.fabric[139] ;
 wire \mod_ro_256.fabric[13] ;
 wire \mod_ro_256.fabric[140] ;
 wire \mod_ro_256.fabric[141] ;
 wire \mod_ro_256.fabric[142] ;
 wire \mod_ro_256.fabric[143] ;
 wire \mod_ro_256.fabric[144] ;
 wire \mod_ro_256.fabric[145] ;
 wire \mod_ro_256.fabric[146] ;
 wire \mod_ro_256.fabric[147] ;
 wire \mod_ro_256.fabric[148] ;
 wire \mod_ro_256.fabric[149] ;
 wire \mod_ro_256.fabric[14] ;
 wire \mod_ro_256.fabric[150] ;
 wire \mod_ro_256.fabric[151] ;
 wire \mod_ro_256.fabric[152] ;
 wire \mod_ro_256.fabric[153] ;
 wire \mod_ro_256.fabric[154] ;
 wire \mod_ro_256.fabric[155] ;
 wire \mod_ro_256.fabric[156] ;
 wire \mod_ro_256.fabric[157] ;
 wire \mod_ro_256.fabric[158] ;
 wire \mod_ro_256.fabric[159] ;
 wire \mod_ro_256.fabric[15] ;
 wire \mod_ro_256.fabric[160] ;
 wire \mod_ro_256.fabric[161] ;
 wire \mod_ro_256.fabric[162] ;
 wire \mod_ro_256.fabric[163] ;
 wire \mod_ro_256.fabric[164] ;
 wire \mod_ro_256.fabric[165] ;
 wire \mod_ro_256.fabric[166] ;
 wire \mod_ro_256.fabric[167] ;
 wire \mod_ro_256.fabric[168] ;
 wire \mod_ro_256.fabric[169] ;
 wire \mod_ro_256.fabric[16] ;
 wire \mod_ro_256.fabric[170] ;
 wire \mod_ro_256.fabric[171] ;
 wire \mod_ro_256.fabric[172] ;
 wire \mod_ro_256.fabric[173] ;
 wire \mod_ro_256.fabric[174] ;
 wire \mod_ro_256.fabric[175] ;
 wire \mod_ro_256.fabric[176] ;
 wire \mod_ro_256.fabric[177] ;
 wire \mod_ro_256.fabric[178] ;
 wire \mod_ro_256.fabric[179] ;
 wire \mod_ro_256.fabric[17] ;
 wire \mod_ro_256.fabric[180] ;
 wire \mod_ro_256.fabric[181] ;
 wire \mod_ro_256.fabric[182] ;
 wire \mod_ro_256.fabric[183] ;
 wire \mod_ro_256.fabric[184] ;
 wire \mod_ro_256.fabric[185] ;
 wire \mod_ro_256.fabric[186] ;
 wire \mod_ro_256.fabric[187] ;
 wire \mod_ro_256.fabric[188] ;
 wire \mod_ro_256.fabric[189] ;
 wire \mod_ro_256.fabric[18] ;
 wire \mod_ro_256.fabric[190] ;
 wire \mod_ro_256.fabric[191] ;
 wire \mod_ro_256.fabric[192] ;
 wire \mod_ro_256.fabric[193] ;
 wire \mod_ro_256.fabric[194] ;
 wire \mod_ro_256.fabric[195] ;
 wire \mod_ro_256.fabric[196] ;
 wire \mod_ro_256.fabric[197] ;
 wire \mod_ro_256.fabric[198] ;
 wire \mod_ro_256.fabric[199] ;
 wire \mod_ro_256.fabric[19] ;
 wire \mod_ro_256.fabric[1] ;
 wire \mod_ro_256.fabric[200] ;
 wire \mod_ro_256.fabric[201] ;
 wire \mod_ro_256.fabric[202] ;
 wire \mod_ro_256.fabric[203] ;
 wire \mod_ro_256.fabric[204] ;
 wire \mod_ro_256.fabric[205] ;
 wire \mod_ro_256.fabric[206] ;
 wire \mod_ro_256.fabric[207] ;
 wire \mod_ro_256.fabric[208] ;
 wire \mod_ro_256.fabric[209] ;
 wire \mod_ro_256.fabric[20] ;
 wire \mod_ro_256.fabric[210] ;
 wire \mod_ro_256.fabric[211] ;
 wire \mod_ro_256.fabric[212] ;
 wire \mod_ro_256.fabric[213] ;
 wire \mod_ro_256.fabric[214] ;
 wire \mod_ro_256.fabric[215] ;
 wire \mod_ro_256.fabric[216] ;
 wire \mod_ro_256.fabric[217] ;
 wire \mod_ro_256.fabric[218] ;
 wire \mod_ro_256.fabric[219] ;
 wire \mod_ro_256.fabric[21] ;
 wire \mod_ro_256.fabric[220] ;
 wire \mod_ro_256.fabric[221] ;
 wire \mod_ro_256.fabric[222] ;
 wire \mod_ro_256.fabric[223] ;
 wire \mod_ro_256.fabric[224] ;
 wire \mod_ro_256.fabric[225] ;
 wire \mod_ro_256.fabric[226] ;
 wire \mod_ro_256.fabric[227] ;
 wire \mod_ro_256.fabric[228] ;
 wire \mod_ro_256.fabric[229] ;
 wire \mod_ro_256.fabric[22] ;
 wire \mod_ro_256.fabric[230] ;
 wire \mod_ro_256.fabric[231] ;
 wire \mod_ro_256.fabric[232] ;
 wire \mod_ro_256.fabric[233] ;
 wire \mod_ro_256.fabric[234] ;
 wire \mod_ro_256.fabric[235] ;
 wire \mod_ro_256.fabric[236] ;
 wire \mod_ro_256.fabric[237] ;
 wire \mod_ro_256.fabric[238] ;
 wire \mod_ro_256.fabric[239] ;
 wire \mod_ro_256.fabric[23] ;
 wire \mod_ro_256.fabric[240] ;
 wire \mod_ro_256.fabric[241] ;
 wire \mod_ro_256.fabric[242] ;
 wire \mod_ro_256.fabric[243] ;
 wire \mod_ro_256.fabric[244] ;
 wire \mod_ro_256.fabric[245] ;
 wire \mod_ro_256.fabric[246] ;
 wire \mod_ro_256.fabric[247] ;
 wire \mod_ro_256.fabric[248] ;
 wire \mod_ro_256.fabric[249] ;
 wire \mod_ro_256.fabric[24] ;
 wire \mod_ro_256.fabric[250] ;
 wire \mod_ro_256.fabric[251] ;
 wire \mod_ro_256.fabric[252] ;
 wire \mod_ro_256.fabric[253] ;
 wire \mod_ro_256.fabric[254] ;
 wire \mod_ro_256.fabric[255] ;
 wire \mod_ro_256.fabric[256] ;
 wire \mod_ro_256.fabric[25] ;
 wire \mod_ro_256.fabric[26] ;
 wire \mod_ro_256.fabric[27] ;
 wire \mod_ro_256.fabric[28] ;
 wire \mod_ro_256.fabric[29] ;
 wire \mod_ro_256.fabric[2] ;
 wire \mod_ro_256.fabric[30] ;
 wire \mod_ro_256.fabric[31] ;
 wire \mod_ro_256.fabric[32] ;
 wire \mod_ro_256.fabric[33] ;
 wire \mod_ro_256.fabric[34] ;
 wire \mod_ro_256.fabric[35] ;
 wire \mod_ro_256.fabric[36] ;
 wire \mod_ro_256.fabric[37] ;
 wire \mod_ro_256.fabric[38] ;
 wire \mod_ro_256.fabric[39] ;
 wire \mod_ro_256.fabric[3] ;
 wire \mod_ro_256.fabric[40] ;
 wire \mod_ro_256.fabric[41] ;
 wire \mod_ro_256.fabric[42] ;
 wire \mod_ro_256.fabric[43] ;
 wire \mod_ro_256.fabric[44] ;
 wire \mod_ro_256.fabric[45] ;
 wire \mod_ro_256.fabric[46] ;
 wire \mod_ro_256.fabric[47] ;
 wire \mod_ro_256.fabric[48] ;
 wire \mod_ro_256.fabric[49] ;
 wire \mod_ro_256.fabric[4] ;
 wire \mod_ro_256.fabric[50] ;
 wire \mod_ro_256.fabric[51] ;
 wire \mod_ro_256.fabric[52] ;
 wire \mod_ro_256.fabric[53] ;
 wire \mod_ro_256.fabric[54] ;
 wire \mod_ro_256.fabric[55] ;
 wire \mod_ro_256.fabric[56] ;
 wire \mod_ro_256.fabric[57] ;
 wire \mod_ro_256.fabric[58] ;
 wire \mod_ro_256.fabric[59] ;
 wire \mod_ro_256.fabric[5] ;
 wire \mod_ro_256.fabric[60] ;
 wire \mod_ro_256.fabric[61] ;
 wire \mod_ro_256.fabric[62] ;
 wire \mod_ro_256.fabric[63] ;
 wire \mod_ro_256.fabric[64] ;
 wire \mod_ro_256.fabric[65] ;
 wire \mod_ro_256.fabric[66] ;
 wire \mod_ro_256.fabric[67] ;
 wire \mod_ro_256.fabric[68] ;
 wire \mod_ro_256.fabric[69] ;
 wire \mod_ro_256.fabric[6] ;
 wire \mod_ro_256.fabric[70] ;
 wire \mod_ro_256.fabric[71] ;
 wire \mod_ro_256.fabric[72] ;
 wire \mod_ro_256.fabric[73] ;
 wire \mod_ro_256.fabric[74] ;
 wire \mod_ro_256.fabric[75] ;
 wire \mod_ro_256.fabric[76] ;
 wire \mod_ro_256.fabric[77] ;
 wire \mod_ro_256.fabric[78] ;
 wire \mod_ro_256.fabric[79] ;
 wire \mod_ro_256.fabric[7] ;
 wire \mod_ro_256.fabric[80] ;
 wire \mod_ro_256.fabric[81] ;
 wire \mod_ro_256.fabric[82] ;
 wire \mod_ro_256.fabric[83] ;
 wire \mod_ro_256.fabric[84] ;
 wire \mod_ro_256.fabric[85] ;
 wire \mod_ro_256.fabric[86] ;
 wire \mod_ro_256.fabric[87] ;
 wire \mod_ro_256.fabric[88] ;
 wire \mod_ro_256.fabric[89] ;
 wire \mod_ro_256.fabric[8] ;
 wire \mod_ro_256.fabric[90] ;
 wire \mod_ro_256.fabric[91] ;
 wire \mod_ro_256.fabric[92] ;
 wire \mod_ro_256.fabric[93] ;
 wire \mod_ro_256.fabric[94] ;
 wire \mod_ro_256.fabric[95] ;
 wire \mod_ro_256.fabric[96] ;
 wire \mod_ro_256.fabric[97] ;
 wire \mod_ro_256.fabric[98] ;
 wire \mod_ro_256.fabric[99] ;
 wire \mod_ro_256.fabric[9] ;
 wire \mod_ro_256_drive4.fabric[0] ;
 wire \mod_ro_256_drive4.fabric[100] ;
 wire \mod_ro_256_drive4.fabric[101] ;
 wire \mod_ro_256_drive4.fabric[102] ;
 wire \mod_ro_256_drive4.fabric[103] ;
 wire \mod_ro_256_drive4.fabric[104] ;
 wire \mod_ro_256_drive4.fabric[105] ;
 wire \mod_ro_256_drive4.fabric[106] ;
 wire \mod_ro_256_drive4.fabric[107] ;
 wire \mod_ro_256_drive4.fabric[108] ;
 wire \mod_ro_256_drive4.fabric[109] ;
 wire \mod_ro_256_drive4.fabric[10] ;
 wire \mod_ro_256_drive4.fabric[110] ;
 wire \mod_ro_256_drive4.fabric[111] ;
 wire \mod_ro_256_drive4.fabric[112] ;
 wire \mod_ro_256_drive4.fabric[113] ;
 wire \mod_ro_256_drive4.fabric[114] ;
 wire \mod_ro_256_drive4.fabric[115] ;
 wire \mod_ro_256_drive4.fabric[116] ;
 wire \mod_ro_256_drive4.fabric[117] ;
 wire \mod_ro_256_drive4.fabric[118] ;
 wire \mod_ro_256_drive4.fabric[119] ;
 wire \mod_ro_256_drive4.fabric[11] ;
 wire \mod_ro_256_drive4.fabric[120] ;
 wire \mod_ro_256_drive4.fabric[121] ;
 wire \mod_ro_256_drive4.fabric[122] ;
 wire \mod_ro_256_drive4.fabric[123] ;
 wire \mod_ro_256_drive4.fabric[124] ;
 wire \mod_ro_256_drive4.fabric[125] ;
 wire \mod_ro_256_drive4.fabric[126] ;
 wire \mod_ro_256_drive4.fabric[127] ;
 wire \mod_ro_256_drive4.fabric[128] ;
 wire \mod_ro_256_drive4.fabric[129] ;
 wire \mod_ro_256_drive4.fabric[12] ;
 wire \mod_ro_256_drive4.fabric[130] ;
 wire \mod_ro_256_drive4.fabric[131] ;
 wire \mod_ro_256_drive4.fabric[132] ;
 wire \mod_ro_256_drive4.fabric[133] ;
 wire \mod_ro_256_drive4.fabric[134] ;
 wire \mod_ro_256_drive4.fabric[135] ;
 wire \mod_ro_256_drive4.fabric[136] ;
 wire \mod_ro_256_drive4.fabric[137] ;
 wire \mod_ro_256_drive4.fabric[138] ;
 wire \mod_ro_256_drive4.fabric[139] ;
 wire \mod_ro_256_drive4.fabric[13] ;
 wire \mod_ro_256_drive4.fabric[140] ;
 wire \mod_ro_256_drive4.fabric[141] ;
 wire \mod_ro_256_drive4.fabric[142] ;
 wire \mod_ro_256_drive4.fabric[143] ;
 wire \mod_ro_256_drive4.fabric[144] ;
 wire \mod_ro_256_drive4.fabric[145] ;
 wire \mod_ro_256_drive4.fabric[146] ;
 wire \mod_ro_256_drive4.fabric[147] ;
 wire \mod_ro_256_drive4.fabric[148] ;
 wire \mod_ro_256_drive4.fabric[149] ;
 wire \mod_ro_256_drive4.fabric[14] ;
 wire \mod_ro_256_drive4.fabric[150] ;
 wire \mod_ro_256_drive4.fabric[151] ;
 wire \mod_ro_256_drive4.fabric[152] ;
 wire \mod_ro_256_drive4.fabric[153] ;
 wire \mod_ro_256_drive4.fabric[154] ;
 wire \mod_ro_256_drive4.fabric[155] ;
 wire \mod_ro_256_drive4.fabric[156] ;
 wire \mod_ro_256_drive4.fabric[157] ;
 wire \mod_ro_256_drive4.fabric[158] ;
 wire \mod_ro_256_drive4.fabric[159] ;
 wire \mod_ro_256_drive4.fabric[15] ;
 wire \mod_ro_256_drive4.fabric[160] ;
 wire \mod_ro_256_drive4.fabric[161] ;
 wire \mod_ro_256_drive4.fabric[162] ;
 wire \mod_ro_256_drive4.fabric[163] ;
 wire \mod_ro_256_drive4.fabric[164] ;
 wire \mod_ro_256_drive4.fabric[165] ;
 wire \mod_ro_256_drive4.fabric[166] ;
 wire \mod_ro_256_drive4.fabric[167] ;
 wire \mod_ro_256_drive4.fabric[168] ;
 wire \mod_ro_256_drive4.fabric[169] ;
 wire \mod_ro_256_drive4.fabric[16] ;
 wire \mod_ro_256_drive4.fabric[170] ;
 wire \mod_ro_256_drive4.fabric[171] ;
 wire \mod_ro_256_drive4.fabric[172] ;
 wire \mod_ro_256_drive4.fabric[173] ;
 wire \mod_ro_256_drive4.fabric[174] ;
 wire \mod_ro_256_drive4.fabric[175] ;
 wire \mod_ro_256_drive4.fabric[176] ;
 wire \mod_ro_256_drive4.fabric[177] ;
 wire \mod_ro_256_drive4.fabric[178] ;
 wire \mod_ro_256_drive4.fabric[179] ;
 wire \mod_ro_256_drive4.fabric[17] ;
 wire \mod_ro_256_drive4.fabric[180] ;
 wire \mod_ro_256_drive4.fabric[181] ;
 wire \mod_ro_256_drive4.fabric[182] ;
 wire \mod_ro_256_drive4.fabric[183] ;
 wire \mod_ro_256_drive4.fabric[184] ;
 wire \mod_ro_256_drive4.fabric[185] ;
 wire \mod_ro_256_drive4.fabric[186] ;
 wire \mod_ro_256_drive4.fabric[187] ;
 wire \mod_ro_256_drive4.fabric[188] ;
 wire \mod_ro_256_drive4.fabric[189] ;
 wire \mod_ro_256_drive4.fabric[18] ;
 wire \mod_ro_256_drive4.fabric[190] ;
 wire \mod_ro_256_drive4.fabric[191] ;
 wire \mod_ro_256_drive4.fabric[192] ;
 wire \mod_ro_256_drive4.fabric[193] ;
 wire \mod_ro_256_drive4.fabric[194] ;
 wire \mod_ro_256_drive4.fabric[195] ;
 wire \mod_ro_256_drive4.fabric[196] ;
 wire \mod_ro_256_drive4.fabric[197] ;
 wire \mod_ro_256_drive4.fabric[198] ;
 wire \mod_ro_256_drive4.fabric[199] ;
 wire \mod_ro_256_drive4.fabric[19] ;
 wire \mod_ro_256_drive4.fabric[1] ;
 wire \mod_ro_256_drive4.fabric[200] ;
 wire \mod_ro_256_drive4.fabric[201] ;
 wire \mod_ro_256_drive4.fabric[202] ;
 wire \mod_ro_256_drive4.fabric[203] ;
 wire \mod_ro_256_drive4.fabric[204] ;
 wire \mod_ro_256_drive4.fabric[205] ;
 wire \mod_ro_256_drive4.fabric[206] ;
 wire \mod_ro_256_drive4.fabric[207] ;
 wire \mod_ro_256_drive4.fabric[208] ;
 wire \mod_ro_256_drive4.fabric[209] ;
 wire \mod_ro_256_drive4.fabric[20] ;
 wire \mod_ro_256_drive4.fabric[210] ;
 wire \mod_ro_256_drive4.fabric[211] ;
 wire \mod_ro_256_drive4.fabric[212] ;
 wire \mod_ro_256_drive4.fabric[213] ;
 wire \mod_ro_256_drive4.fabric[214] ;
 wire \mod_ro_256_drive4.fabric[215] ;
 wire \mod_ro_256_drive4.fabric[216] ;
 wire \mod_ro_256_drive4.fabric[217] ;
 wire \mod_ro_256_drive4.fabric[218] ;
 wire \mod_ro_256_drive4.fabric[219] ;
 wire \mod_ro_256_drive4.fabric[21] ;
 wire \mod_ro_256_drive4.fabric[220] ;
 wire \mod_ro_256_drive4.fabric[221] ;
 wire \mod_ro_256_drive4.fabric[222] ;
 wire \mod_ro_256_drive4.fabric[223] ;
 wire \mod_ro_256_drive4.fabric[224] ;
 wire \mod_ro_256_drive4.fabric[225] ;
 wire \mod_ro_256_drive4.fabric[226] ;
 wire \mod_ro_256_drive4.fabric[227] ;
 wire \mod_ro_256_drive4.fabric[228] ;
 wire \mod_ro_256_drive4.fabric[229] ;
 wire \mod_ro_256_drive4.fabric[22] ;
 wire \mod_ro_256_drive4.fabric[230] ;
 wire \mod_ro_256_drive4.fabric[231] ;
 wire \mod_ro_256_drive4.fabric[232] ;
 wire \mod_ro_256_drive4.fabric[233] ;
 wire \mod_ro_256_drive4.fabric[234] ;
 wire \mod_ro_256_drive4.fabric[235] ;
 wire \mod_ro_256_drive4.fabric[236] ;
 wire \mod_ro_256_drive4.fabric[237] ;
 wire \mod_ro_256_drive4.fabric[238] ;
 wire \mod_ro_256_drive4.fabric[239] ;
 wire \mod_ro_256_drive4.fabric[23] ;
 wire \mod_ro_256_drive4.fabric[240] ;
 wire \mod_ro_256_drive4.fabric[241] ;
 wire \mod_ro_256_drive4.fabric[242] ;
 wire \mod_ro_256_drive4.fabric[243] ;
 wire \mod_ro_256_drive4.fabric[244] ;
 wire \mod_ro_256_drive4.fabric[245] ;
 wire \mod_ro_256_drive4.fabric[246] ;
 wire \mod_ro_256_drive4.fabric[247] ;
 wire \mod_ro_256_drive4.fabric[248] ;
 wire \mod_ro_256_drive4.fabric[249] ;
 wire \mod_ro_256_drive4.fabric[24] ;
 wire \mod_ro_256_drive4.fabric[250] ;
 wire \mod_ro_256_drive4.fabric[251] ;
 wire \mod_ro_256_drive4.fabric[252] ;
 wire \mod_ro_256_drive4.fabric[253] ;
 wire \mod_ro_256_drive4.fabric[254] ;
 wire \mod_ro_256_drive4.fabric[255] ;
 wire \mod_ro_256_drive4.fabric[256] ;
 wire \mod_ro_256_drive4.fabric[25] ;
 wire \mod_ro_256_drive4.fabric[26] ;
 wire \mod_ro_256_drive4.fabric[27] ;
 wire \mod_ro_256_drive4.fabric[28] ;
 wire \mod_ro_256_drive4.fabric[29] ;
 wire \mod_ro_256_drive4.fabric[2] ;
 wire \mod_ro_256_drive4.fabric[30] ;
 wire \mod_ro_256_drive4.fabric[31] ;
 wire \mod_ro_256_drive4.fabric[32] ;
 wire \mod_ro_256_drive4.fabric[33] ;
 wire \mod_ro_256_drive4.fabric[34] ;
 wire \mod_ro_256_drive4.fabric[35] ;
 wire \mod_ro_256_drive4.fabric[36] ;
 wire \mod_ro_256_drive4.fabric[37] ;
 wire \mod_ro_256_drive4.fabric[38] ;
 wire \mod_ro_256_drive4.fabric[39] ;
 wire \mod_ro_256_drive4.fabric[3] ;
 wire \mod_ro_256_drive4.fabric[40] ;
 wire \mod_ro_256_drive4.fabric[41] ;
 wire \mod_ro_256_drive4.fabric[42] ;
 wire \mod_ro_256_drive4.fabric[43] ;
 wire \mod_ro_256_drive4.fabric[44] ;
 wire \mod_ro_256_drive4.fabric[45] ;
 wire \mod_ro_256_drive4.fabric[46] ;
 wire \mod_ro_256_drive4.fabric[47] ;
 wire \mod_ro_256_drive4.fabric[48] ;
 wire \mod_ro_256_drive4.fabric[49] ;
 wire \mod_ro_256_drive4.fabric[4] ;
 wire \mod_ro_256_drive4.fabric[50] ;
 wire \mod_ro_256_drive4.fabric[51] ;
 wire \mod_ro_256_drive4.fabric[52] ;
 wire \mod_ro_256_drive4.fabric[53] ;
 wire \mod_ro_256_drive4.fabric[54] ;
 wire \mod_ro_256_drive4.fabric[55] ;
 wire \mod_ro_256_drive4.fabric[56] ;
 wire \mod_ro_256_drive4.fabric[57] ;
 wire \mod_ro_256_drive4.fabric[58] ;
 wire \mod_ro_256_drive4.fabric[59] ;
 wire \mod_ro_256_drive4.fabric[5] ;
 wire \mod_ro_256_drive4.fabric[60] ;
 wire \mod_ro_256_drive4.fabric[61] ;
 wire \mod_ro_256_drive4.fabric[62] ;
 wire \mod_ro_256_drive4.fabric[63] ;
 wire \mod_ro_256_drive4.fabric[64] ;
 wire \mod_ro_256_drive4.fabric[65] ;
 wire \mod_ro_256_drive4.fabric[66] ;
 wire \mod_ro_256_drive4.fabric[67] ;
 wire \mod_ro_256_drive4.fabric[68] ;
 wire \mod_ro_256_drive4.fabric[69] ;
 wire \mod_ro_256_drive4.fabric[6] ;
 wire \mod_ro_256_drive4.fabric[70] ;
 wire \mod_ro_256_drive4.fabric[71] ;
 wire \mod_ro_256_drive4.fabric[72] ;
 wire \mod_ro_256_drive4.fabric[73] ;
 wire \mod_ro_256_drive4.fabric[74] ;
 wire \mod_ro_256_drive4.fabric[75] ;
 wire \mod_ro_256_drive4.fabric[76] ;
 wire \mod_ro_256_drive4.fabric[77] ;
 wire \mod_ro_256_drive4.fabric[78] ;
 wire \mod_ro_256_drive4.fabric[79] ;
 wire \mod_ro_256_drive4.fabric[7] ;
 wire \mod_ro_256_drive4.fabric[80] ;
 wire \mod_ro_256_drive4.fabric[81] ;
 wire \mod_ro_256_drive4.fabric[82] ;
 wire \mod_ro_256_drive4.fabric[83] ;
 wire \mod_ro_256_drive4.fabric[84] ;
 wire \mod_ro_256_drive4.fabric[85] ;
 wire \mod_ro_256_drive4.fabric[86] ;
 wire \mod_ro_256_drive4.fabric[87] ;
 wire \mod_ro_256_drive4.fabric[88] ;
 wire \mod_ro_256_drive4.fabric[89] ;
 wire \mod_ro_256_drive4.fabric[8] ;
 wire \mod_ro_256_drive4.fabric[90] ;
 wire \mod_ro_256_drive4.fabric[91] ;
 wire \mod_ro_256_drive4.fabric[92] ;
 wire \mod_ro_256_drive4.fabric[93] ;
 wire \mod_ro_256_drive4.fabric[94] ;
 wire \mod_ro_256_drive4.fabric[95] ;
 wire \mod_ro_256_drive4.fabric[96] ;
 wire \mod_ro_256_drive4.fabric[97] ;
 wire \mod_ro_256_drive4.fabric[98] ;
 wire \mod_ro_256_drive4.fabric[99] ;
 wire \mod_ro_256_drive4.fabric[9] ;
 wire \mod_ro_31.fabric[0] ;
 wire \mod_ro_31.fabric[10] ;
 wire \mod_ro_31.fabric[11] ;
 wire \mod_ro_31.fabric[12] ;
 wire \mod_ro_31.fabric[13] ;
 wire \mod_ro_31.fabric[14] ;
 wire \mod_ro_31.fabric[15] ;
 wire \mod_ro_31.fabric[16] ;
 wire \mod_ro_31.fabric[17] ;
 wire \mod_ro_31.fabric[18] ;
 wire \mod_ro_31.fabric[19] ;
 wire \mod_ro_31.fabric[1] ;
 wire \mod_ro_31.fabric[20] ;
 wire \mod_ro_31.fabric[21] ;
 wire \mod_ro_31.fabric[22] ;
 wire \mod_ro_31.fabric[23] ;
 wire \mod_ro_31.fabric[24] ;
 wire \mod_ro_31.fabric[25] ;
 wire \mod_ro_31.fabric[26] ;
 wire \mod_ro_31.fabric[27] ;
 wire \mod_ro_31.fabric[28] ;
 wire \mod_ro_31.fabric[29] ;
 wire \mod_ro_31.fabric[2] ;
 wire \mod_ro_31.fabric[30] ;
 wire \mod_ro_31.fabric[31] ;
 wire \mod_ro_31.fabric[3] ;
 wire \mod_ro_31.fabric[4] ;
 wire \mod_ro_31.fabric[5] ;
 wire \mod_ro_31.fabric[6] ;
 wire \mod_ro_31.fabric[7] ;
 wire \mod_ro_31.fabric[8] ;
 wire \mod_ro_31.fabric[9] ;
 wire \mod_ro_32_1.fabric[0] ;
 wire \mod_ro_32_1.fabric[10] ;
 wire \mod_ro_32_1.fabric[11] ;
 wire \mod_ro_32_1.fabric[12] ;
 wire \mod_ro_32_1.fabric[13] ;
 wire \mod_ro_32_1.fabric[14] ;
 wire \mod_ro_32_1.fabric[15] ;
 wire \mod_ro_32_1.fabric[16] ;
 wire \mod_ro_32_1.fabric[17] ;
 wire \mod_ro_32_1.fabric[18] ;
 wire \mod_ro_32_1.fabric[19] ;
 wire \mod_ro_32_1.fabric[1] ;
 wire \mod_ro_32_1.fabric[20] ;
 wire \mod_ro_32_1.fabric[21] ;
 wire \mod_ro_32_1.fabric[22] ;
 wire \mod_ro_32_1.fabric[23] ;
 wire \mod_ro_32_1.fabric[24] ;
 wire \mod_ro_32_1.fabric[25] ;
 wire \mod_ro_32_1.fabric[26] ;
 wire \mod_ro_32_1.fabric[27] ;
 wire \mod_ro_32_1.fabric[28] ;
 wire \mod_ro_32_1.fabric[29] ;
 wire \mod_ro_32_1.fabric[2] ;
 wire \mod_ro_32_1.fabric[30] ;
 wire \mod_ro_32_1.fabric[31] ;
 wire \mod_ro_32_1.fabric[32] ;
 wire \mod_ro_32_1.fabric[3] ;
 wire \mod_ro_32_1.fabric[4] ;
 wire \mod_ro_32_1.fabric[5] ;
 wire \mod_ro_32_1.fabric[6] ;
 wire \mod_ro_32_1.fabric[7] ;
 wire \mod_ro_32_1.fabric[8] ;
 wire \mod_ro_32_1.fabric[9] ;
 wire \mod_ro_32_2.fabric[0] ;
 wire \mod_ro_32_2.fabric[10] ;
 wire \mod_ro_32_2.fabric[11] ;
 wire \mod_ro_32_2.fabric[12] ;
 wire \mod_ro_32_2.fabric[13] ;
 wire \mod_ro_32_2.fabric[14] ;
 wire \mod_ro_32_2.fabric[15] ;
 wire \mod_ro_32_2.fabric[16] ;
 wire \mod_ro_32_2.fabric[17] ;
 wire \mod_ro_32_2.fabric[18] ;
 wire \mod_ro_32_2.fabric[19] ;
 wire \mod_ro_32_2.fabric[1] ;
 wire \mod_ro_32_2.fabric[20] ;
 wire \mod_ro_32_2.fabric[21] ;
 wire \mod_ro_32_2.fabric[22] ;
 wire \mod_ro_32_2.fabric[23] ;
 wire \mod_ro_32_2.fabric[24] ;
 wire \mod_ro_32_2.fabric[25] ;
 wire \mod_ro_32_2.fabric[26] ;
 wire \mod_ro_32_2.fabric[27] ;
 wire \mod_ro_32_2.fabric[28] ;
 wire \mod_ro_32_2.fabric[29] ;
 wire \mod_ro_32_2.fabric[2] ;
 wire \mod_ro_32_2.fabric[30] ;
 wire \mod_ro_32_2.fabric[31] ;
 wire \mod_ro_32_2.fabric[32] ;
 wire \mod_ro_32_2.fabric[3] ;
 wire \mod_ro_32_2.fabric[4] ;
 wire \mod_ro_32_2.fabric[5] ;
 wire \mod_ro_32_2.fabric[6] ;
 wire \mod_ro_32_2.fabric[7] ;
 wire \mod_ro_32_2.fabric[8] ;
 wire \mod_ro_32_2.fabric[9] ;
 wire \mod_ro_32_drive4.fabric[0] ;
 wire \mod_ro_32_drive4.fabric[10] ;
 wire \mod_ro_32_drive4.fabric[11] ;
 wire \mod_ro_32_drive4.fabric[12] ;
 wire \mod_ro_32_drive4.fabric[13] ;
 wire \mod_ro_32_drive4.fabric[14] ;
 wire \mod_ro_32_drive4.fabric[15] ;
 wire \mod_ro_32_drive4.fabric[16] ;
 wire \mod_ro_32_drive4.fabric[17] ;
 wire \mod_ro_32_drive4.fabric[18] ;
 wire \mod_ro_32_drive4.fabric[19] ;
 wire \mod_ro_32_drive4.fabric[1] ;
 wire \mod_ro_32_drive4.fabric[20] ;
 wire \mod_ro_32_drive4.fabric[21] ;
 wire \mod_ro_32_drive4.fabric[22] ;
 wire \mod_ro_32_drive4.fabric[23] ;
 wire \mod_ro_32_drive4.fabric[24] ;
 wire \mod_ro_32_drive4.fabric[25] ;
 wire \mod_ro_32_drive4.fabric[26] ;
 wire \mod_ro_32_drive4.fabric[27] ;
 wire \mod_ro_32_drive4.fabric[28] ;
 wire \mod_ro_32_drive4.fabric[29] ;
 wire \mod_ro_32_drive4.fabric[2] ;
 wire \mod_ro_32_drive4.fabric[30] ;
 wire \mod_ro_32_drive4.fabric[31] ;
 wire \mod_ro_32_drive4.fabric[32] ;
 wire \mod_ro_32_drive4.fabric[3] ;
 wire \mod_ro_32_drive4.fabric[4] ;
 wire \mod_ro_32_drive4.fabric[5] ;
 wire \mod_ro_32_drive4.fabric[6] ;
 wire \mod_ro_32_drive4.fabric[7] ;
 wire \mod_ro_32_drive4.fabric[8] ;
 wire \mod_ro_32_drive4.fabric[9] ;
 wire \mod_ro_32_raw.fabric[0] ;
 wire \mod_ro_32_raw.fabric[10] ;
 wire \mod_ro_32_raw.fabric[11] ;
 wire \mod_ro_32_raw.fabric[12] ;
 wire \mod_ro_32_raw.fabric[13] ;
 wire \mod_ro_32_raw.fabric[14] ;
 wire \mod_ro_32_raw.fabric[15] ;
 wire \mod_ro_32_raw.fabric[16] ;
 wire \mod_ro_32_raw.fabric[17] ;
 wire \mod_ro_32_raw.fabric[18] ;
 wire \mod_ro_32_raw.fabric[19] ;
 wire \mod_ro_32_raw.fabric[1] ;
 wire \mod_ro_32_raw.fabric[20] ;
 wire \mod_ro_32_raw.fabric[21] ;
 wire \mod_ro_32_raw.fabric[22] ;
 wire \mod_ro_32_raw.fabric[23] ;
 wire \mod_ro_32_raw.fabric[24] ;
 wire \mod_ro_32_raw.fabric[25] ;
 wire \mod_ro_32_raw.fabric[26] ;
 wire \mod_ro_32_raw.fabric[27] ;
 wire \mod_ro_32_raw.fabric[28] ;
 wire \mod_ro_32_raw.fabric[29] ;
 wire \mod_ro_32_raw.fabric[2] ;
 wire \mod_ro_32_raw.fabric[30] ;
 wire \mod_ro_32_raw.fabric[31] ;
 wire \mod_ro_32_raw.fabric[32] ;
 wire \mod_ro_32_raw.fabric[3] ;
 wire \mod_ro_32_raw.fabric[4] ;
 wire \mod_ro_32_raw.fabric[5] ;
 wire \mod_ro_32_raw.fabric[6] ;
 wire \mod_ro_32_raw.fabric[7] ;
 wire \mod_ro_32_raw.fabric[8] ;
 wire \mod_ro_32_raw.fabric[9] ;
 wire \mod_ro_64.fabric[0] ;
 wire \mod_ro_64.fabric[10] ;
 wire \mod_ro_64.fabric[11] ;
 wire \mod_ro_64.fabric[12] ;
 wire \mod_ro_64.fabric[13] ;
 wire \mod_ro_64.fabric[14] ;
 wire \mod_ro_64.fabric[15] ;
 wire \mod_ro_64.fabric[16] ;
 wire \mod_ro_64.fabric[17] ;
 wire \mod_ro_64.fabric[18] ;
 wire \mod_ro_64.fabric[19] ;
 wire \mod_ro_64.fabric[1] ;
 wire \mod_ro_64.fabric[20] ;
 wire \mod_ro_64.fabric[21] ;
 wire \mod_ro_64.fabric[22] ;
 wire \mod_ro_64.fabric[23] ;
 wire \mod_ro_64.fabric[24] ;
 wire \mod_ro_64.fabric[25] ;
 wire \mod_ro_64.fabric[26] ;
 wire \mod_ro_64.fabric[27] ;
 wire \mod_ro_64.fabric[28] ;
 wire \mod_ro_64.fabric[29] ;
 wire \mod_ro_64.fabric[2] ;
 wire \mod_ro_64.fabric[30] ;
 wire \mod_ro_64.fabric[31] ;
 wire \mod_ro_64.fabric[32] ;
 wire \mod_ro_64.fabric[33] ;
 wire \mod_ro_64.fabric[34] ;
 wire \mod_ro_64.fabric[35] ;
 wire \mod_ro_64.fabric[36] ;
 wire \mod_ro_64.fabric[37] ;
 wire \mod_ro_64.fabric[38] ;
 wire \mod_ro_64.fabric[39] ;
 wire \mod_ro_64.fabric[3] ;
 wire \mod_ro_64.fabric[40] ;
 wire \mod_ro_64.fabric[41] ;
 wire \mod_ro_64.fabric[42] ;
 wire \mod_ro_64.fabric[43] ;
 wire \mod_ro_64.fabric[44] ;
 wire \mod_ro_64.fabric[45] ;
 wire \mod_ro_64.fabric[46] ;
 wire \mod_ro_64.fabric[47] ;
 wire \mod_ro_64.fabric[48] ;
 wire \mod_ro_64.fabric[49] ;
 wire \mod_ro_64.fabric[4] ;
 wire \mod_ro_64.fabric[50] ;
 wire \mod_ro_64.fabric[51] ;
 wire \mod_ro_64.fabric[52] ;
 wire \mod_ro_64.fabric[53] ;
 wire \mod_ro_64.fabric[54] ;
 wire \mod_ro_64.fabric[55] ;
 wire \mod_ro_64.fabric[56] ;
 wire \mod_ro_64.fabric[57] ;
 wire \mod_ro_64.fabric[58] ;
 wire \mod_ro_64.fabric[59] ;
 wire \mod_ro_64.fabric[5] ;
 wire \mod_ro_64.fabric[60] ;
 wire \mod_ro_64.fabric[61] ;
 wire \mod_ro_64.fabric[62] ;
 wire \mod_ro_64.fabric[63] ;
 wire \mod_ro_64.fabric[64] ;
 wire \mod_ro_64.fabric[6] ;
 wire \mod_ro_64.fabric[7] ;
 wire \mod_ro_64.fabric[8] ;
 wire \mod_ro_64.fabric[9] ;
 wire \mod_ro_prog.fabric[0] ;
 wire \mod_ro_prog.fabric[1] ;
 wire \mod_ro_prog.fabric[2] ;
 wire \mod_ro_prog.fabric[3] ;
 wire \mod_ro_prog.fabric[4] ;
 wire \mod_ro_prog.fabric[5] ;
 wire \mod_ro_prog.fabric[6] ;
 wire \mod_ro_prog.fabric[7] ;
 wire \mod_ro_prog.fabric[8] ;
 wire \mod_ro_prog.osc_gen[0].inv.i_en ;
 wire \mod_ro_prog.osc_gen[0].inv.inverted ;
 wire \mod_ro_prog.osc_gen[1].inv.i_en ;
 wire \mod_ro_prog.osc_gen[1].inv.inverted ;
 wire \mod_ro_prog.osc_gen[2].inv.i_en ;
 wire \mod_ro_prog.osc_gen[2].inv.inverted ;
 wire \mod_ro_prog.osc_gen[3].inv.i_en ;
 wire \mod_ro_prog.osc_gen[3].inv.inverted ;
 wire \mod_ro_prog.osc_gen[4].inv.i_en ;
 wire \mod_ro_prog.osc_gen[4].inv.inverted ;
 wire \mod_ro_prog.osc_gen[5].inv.i_en ;
 wire \mod_ro_prog.osc_gen[5].inv.inverted ;
 wire \mod_ro_prog.osc_gen[6].inv.i_en ;
 wire \mod_ro_prog.osc_gen[6].inv.inverted ;
 wire \mod_ro_prog.osc_gen[7].inv.i_en ;
 wire \mod_ro_prog.osc_gen[7].inv.inverted ;
 wire o_miso;
 wire o_rosc_mux_out;
 wire \reg_echo[2] ;
 wire \reg_echo[3] ;
 wire \reg_echo[4] ;
 wire \reg_echo[5] ;
 wire \reg_echo[6] ;
 wire \spi_decoder_mod.o_reg_wdata[1] ;
 wire \spi_decoder_mod.o_reg_wdata[2] ;
 wire \spi_decoder_mod.o_reg_wdata[3] ;
 wire \spi_decoder_mod.o_reg_wdata[4] ;
 wire \spi_decoder_mod.o_reg_wdata[5] ;
 wire \spi_decoder_mod.o_reg_wdata[6] ;
 wire \spi_decoder_mod.o_reg_wdata[7] ;
 wire \spi_decoder_mod.shift_cnt[0] ;
 wire \spi_decoder_mod.shift_cnt[1] ;
 wire \spi_decoder_mod.shift_cnt[2] ;
 wire \spi_decoder_mod.shift_out_reg[0] ;
 wire \spi_decoder_mod.shift_out_reg[1] ;
 wire \spi_decoder_mod.shift_out_reg[2] ;
 wire \spi_decoder_mod.shift_out_reg[3] ;
 wire \spi_decoder_mod.shift_out_reg[4] ;
 wire \spi_decoder_mod.shift_out_reg[5] ;
 wire \spi_decoder_mod.shift_out_reg[6] ;
 wire \spi_decoder_mod.spi_state[1] ;
 wire \spi_decoder_mod.spi_state[2] ;
 wire \spi_decoder_mod.spi_state[3] ;
 wire \spi_decoder_mod.start ;
 wire \spi_decoder_mod.write ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire [0:0] \spi_regfile_mod.SYS_CTRL_RESET_q ;
 wire [0:0] \spi_regfile_mod.addr ;

 sg13g2_inv_1 _245_ (.Y(_092_),
    .A(net163));
 sg13g2_inv_1 _246_ (.Y(_093_),
    .A(net144));
 sg13g2_inv_2 _247_ (.Y(_094_),
    .A(net39));
 sg13g2_inv_1 _248_ (.Y(_095_),
    .A(net162));
 sg13g2_inv_1 _249_ (.Y(_096_),
    .A(net104));
 sg13g2_inv_1 _250_ (.Y(_097_),
    .A(net166));
 sg13g2_inv_1 _251_ (.Y(_036_),
    .A(net46));
 sg13g2_inv_1 _252_ (.Y(_011_),
    .A(net79));
 sg13g2_inv_1 _253_ (.Y(_098_),
    .A(net5));
 sg13g2_inv_4 _254_ (.A(net47),
    .Y(_099_));
 sg13g2_inv_1 _454__2 (.Y(net64),
    .A(clknet_1_1__leaf_clk));
 sg13g2_and3_2 _256_ (.X(_100_),
    .A(net79),
    .B(net85),
    .C(net98));
 sg13g2_o21ai_1 _257_ (.B1(_100_),
    .Y(_101_),
    .A1(\spi_decoder_mod.spi_state[1] ),
    .A2(net123));
 sg13g2_nor2_1 _258_ (.A(net123),
    .B(net5),
    .Y(_102_));
 sg13g2_a21oi_1 _259_ (.A1(net166),
    .A2(net123),
    .Y(_103_),
    .B1(_102_));
 sg13g2_nor2_1 _260_ (.A(_101_),
    .B(_103_),
    .Y(_104_));
 sg13g2_a21oi_1 _261_ (.A1(_097_),
    .A2(_101_),
    .Y(_070_),
    .B1(_104_));
 sg13g2_a21o_1 _262_ (.A2(_098_),
    .A1(net93),
    .B1(net112),
    .X(_054_));
 sg13g2_nand2b_1 _263_ (.Y(_053_),
    .B(net77),
    .A_N(net84));
 sg13g2_nand2b_1 _264_ (.Y(_017_),
    .B(net84),
    .A_N(net77));
 sg13g2_nand2b_1 _265_ (.Y(_105_),
    .B(\spi_decoder_mod.spi_state[1] ),
    .A_N(_100_));
 sg13g2_nand2b_1 _266_ (.Y(_001_),
    .B(_105_),
    .A_N(net93));
 sg13g2_a21o_1 _267_ (.A2(_100_),
    .A1(\spi_decoder_mod.spi_state[1] ),
    .B1(net123),
    .X(_002_));
 sg13g2_nor2b_1 _268_ (.A(net1),
    .B_N(net2),
    .Y(_106_));
 sg13g2_nor2b_1 _269_ (.A(net2),
    .B_N(net1),
    .Y(_107_));
 sg13g2_nor2_1 _270_ (.A(net1),
    .B(net2),
    .Y(_108_));
 sg13g2_nand2_1 _271_ (.Y(_109_),
    .A(\mod_ro_32_drive4.fabric[0] ),
    .B(_108_));
 sg13g2_a22oi_1 _272_ (.Y(_110_),
    .B1(_107_),
    .B2(\mod_ro_256.fabric[0] ),
    .A2(_106_),
    .A1(\mod_ro_256_drive4.fabric[0] ));
 sg13g2_nand2b_1 _273_ (.Y(_111_),
    .B(net4),
    .A_N(net3));
 sg13g2_a21oi_1 _274_ (.A1(_109_),
    .A2(_110_),
    .Y(_112_),
    .B1(_111_));
 sg13g2_nor2_1 _275_ (.A(net3),
    .B(net4),
    .Y(_113_));
 sg13g2_nand2_1 _276_ (.Y(_114_),
    .A(\mod_ro_16.fabric[0] ),
    .B(_113_));
 sg13g2_nand2b_1 _277_ (.Y(_115_),
    .B(net3),
    .A_N(net4));
 sg13g2_nand2_1 _278_ (.Y(_116_),
    .A(\mod_ro_32_1.fabric[0] ),
    .B(\mod_ro_32_2.fabric[0] ));
 sg13g2_or2_1 _279_ (.X(_117_),
    .B(_116_),
    .A(_115_));
 sg13g2_nand2_1 _280_ (.Y(_118_),
    .A(net1),
    .B(net2));
 sg13g2_a21oi_1 _281_ (.A1(_114_),
    .A2(_117_),
    .Y(_119_),
    .B1(_118_));
 sg13g2_and2_1 _282_ (.A(\mod_ro_32_2.fabric[0] ),
    .B(_107_),
    .X(_120_));
 sg13g2_a221oi_1 _283_ (.B2(\mod_ro_32_1.fabric[0] ),
    .C1(_120_),
    .B1(_108_),
    .A1(\mod_ro_64.fabric[0] ),
    .Y(_121_),
    .A2(_106_));
 sg13g2_nor2b_1 _284_ (.A(_121_),
    .B_N(_113_),
    .Y(_122_));
 sg13g2_o21ai_1 _285_ (.B1(_108_),
    .Y(_123_),
    .A1(\mod_ro_32_1.fabric[0] ),
    .A2(\mod_ro_32_2.fabric[0] ));
 sg13g2_a22oi_1 _286_ (.Y(_124_),
    .B1(_107_),
    .B2(\mod_ro_31.fabric[0] ),
    .A2(_106_),
    .A1(\mod_ro_128.fabric[0] ));
 sg13g2_a21oi_1 _287_ (.A1(_123_),
    .A2(_124_),
    .Y(_125_),
    .B1(_115_));
 sg13g2_or4_1 _288_ (.A(_112_),
    .B(_119_),
    .C(_122_),
    .D(_125_),
    .X(o_rosc_mux_out));
 sg13g2_nor3_1 _289_ (.A(\spi_decoder_mod.write ),
    .B(\spi_decoder_mod.shift_cnt[0] ),
    .C(\spi_decoder_mod.shift_cnt[1] ),
    .Y(_126_));
 sg13g2_nand3b_1 _290_ (.B(\spi_decoder_mod.spi_state[3] ),
    .C(_126_),
    .Y(_127_),
    .A_N(\spi_decoder_mod.shift_cnt[2] ));
 sg13g2_nor2_2 _291_ (.A(\spi_regfile_mod.addr [0]),
    .B(net38),
    .Y(_128_));
 sg13g2_nor2_2 _292_ (.A(_097_),
    .B(net38),
    .Y(_129_));
 sg13g2_a22oi_1 _293_ (.Y(_130_),
    .B1(_129_),
    .B2(\mod_ro_prog.osc_gen[0].inv.i_en ),
    .A2(_128_),
    .A1(\spi_regfile_mod.SYS_CTRL_RESET_q [0]));
 sg13g2_inv_1 _294_ (.Y(_003_),
    .A(_130_));
 sg13g2_nor3_1 _295_ (.A(\spi_regfile_mod.addr [0]),
    .B(_015_),
    .C(net38),
    .Y(_131_));
 sg13g2_a221oi_1 _296_ (.B2(\mod_ro_prog.osc_gen[1].inv.i_en ),
    .C1(_131_),
    .B1(_129_),
    .A1(net149),
    .Y(_132_),
    .A2(net38));
 sg13g2_inv_1 _297_ (.Y(_004_),
    .A(_132_));
 sg13g2_nor3_1 _298_ (.A(\spi_regfile_mod.addr [0]),
    .B(_016_),
    .C(_127_),
    .Y(_133_));
 sg13g2_a221oi_1 _299_ (.B2(\mod_ro_prog.osc_gen[2].inv.i_en ),
    .C1(_133_),
    .B1(_129_),
    .A1(net150),
    .Y(_134_),
    .A2(_127_));
 sg13g2_inv_1 _300_ (.Y(_005_),
    .A(_134_));
 sg13g2_nand2_1 _301_ (.Y(_135_),
    .A(\reg_echo[2] ),
    .B(_128_));
 sg13g2_a22oi_1 _302_ (.Y(_136_),
    .B1(_129_),
    .B2(\mod_ro_prog.osc_gen[3].inv.i_en ),
    .A2(_127_),
    .A1(net148));
 sg13g2_nand2_1 _303_ (.Y(_006_),
    .A(_135_),
    .B(_136_));
 sg13g2_nand2_1 _304_ (.Y(_137_),
    .A(\mod_ro_prog.osc_gen[4].inv.i_en ),
    .B(_129_));
 sg13g2_a22oi_1 _305_ (.Y(_138_),
    .B1(_128_),
    .B2(\reg_echo[3] ),
    .A2(net38),
    .A1(net153));
 sg13g2_nand2_1 _306_ (.Y(_007_),
    .A(_137_),
    .B(_138_));
 sg13g2_nand2_1 _307_ (.Y(_139_),
    .A(\mod_ro_prog.osc_gen[5].inv.i_en ),
    .B(_129_));
 sg13g2_a22oi_1 _308_ (.Y(_140_),
    .B1(_128_),
    .B2(\reg_echo[4] ),
    .A2(net38),
    .A1(net147));
 sg13g2_nand2_1 _309_ (.Y(_008_),
    .A(_139_),
    .B(_140_));
 sg13g2_nand2_1 _310_ (.Y(_141_),
    .A(\mod_ro_prog.osc_gen[6].inv.i_en ),
    .B(_129_));
 sg13g2_a22oi_1 _311_ (.Y(_142_),
    .B1(_128_),
    .B2(\reg_echo[5] ),
    .A2(net38),
    .A1(net142));
 sg13g2_nand2_1 _312_ (.Y(_009_),
    .A(_141_),
    .B(_142_));
 sg13g2_nand2_1 _313_ (.Y(_143_),
    .A(\mod_ro_prog.osc_gen[7].inv.i_en ),
    .B(_129_));
 sg13g2_a22oi_1 _314_ (.Y(_144_),
    .B1(_128_),
    .B2(\reg_echo[6] ),
    .A2(net38),
    .A1(net152));
 sg13g2_nand2_1 _315_ (.Y(_010_),
    .A(_143_),
    .B(_144_));
 sg13g2_mux2_1 _316_ (.A0(\mod_ro_prog.fabric[0] ),
    .A1(\mod_ro_prog.osc_gen[0].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[0].inv.i_en ),
    .X(\mod_ro_prog.fabric[1] ));
 sg13g2_mux2_1 _317_ (.A0(\mod_ro_prog.fabric[1] ),
    .A1(\mod_ro_prog.osc_gen[1].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[1].inv.i_en ),
    .X(\mod_ro_prog.fabric[2] ));
 sg13g2_mux2_1 _318_ (.A0(\mod_ro_prog.fabric[2] ),
    .A1(\mod_ro_prog.osc_gen[2].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[2].inv.i_en ),
    .X(\mod_ro_prog.fabric[3] ));
 sg13g2_mux2_1 _319_ (.A0(\mod_ro_prog.fabric[3] ),
    .A1(\mod_ro_prog.osc_gen[3].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[3].inv.i_en ),
    .X(\mod_ro_prog.fabric[4] ));
 sg13g2_mux2_1 _320_ (.A0(\mod_ro_prog.fabric[4] ),
    .A1(\mod_ro_prog.osc_gen[4].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[4].inv.i_en ),
    .X(\mod_ro_prog.fabric[5] ));
 sg13g2_mux2_1 _321_ (.A0(\mod_ro_prog.fabric[5] ),
    .A1(\mod_ro_prog.osc_gen[5].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[5].inv.i_en ),
    .X(\mod_ro_prog.fabric[6] ));
 sg13g2_mux2_1 _322_ (.A0(\mod_ro_prog.fabric[6] ),
    .A1(\mod_ro_prog.osc_gen[6].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[6].inv.i_en ),
    .X(\mod_ro_prog.fabric[7] ));
 sg13g2_mux2_1 _323_ (.A0(\mod_ro_prog.fabric[7] ),
    .A1(\mod_ro_prog.osc_gen[7].inv.inverted ),
    .S(\mod_ro_prog.osc_gen[7].inv.i_en ),
    .X(\mod_ro_prog.fabric[8] ));
 sg13g2_xor2_1 _324_ (.B(net85),
    .A(net79),
    .X(_012_));
 sg13g2_a21oi_1 _325_ (.A1(net79),
    .A2(net85),
    .Y(_145_),
    .B1(net98));
 sg13g2_nor2_1 _326_ (.A(_100_),
    .B(_145_),
    .Y(_013_));
 sg13g2_nor2_1 _327_ (.A(\spi_decoder_mod.start ),
    .B(net77),
    .Y(_000_));
 sg13g2_nand3_1 _328_ (.B(net123),
    .C(_100_),
    .A(net112),
    .Y(_146_));
 sg13g2_nor2_2 _329_ (.A(\spi_regfile_mod.addr [0]),
    .B(_146_),
    .Y(_147_));
 sg13g2_nor2_1 _330_ (.A(net109),
    .B(net36),
    .Y(_148_));
 sg13g2_a21oi_1 _331_ (.A1(_098_),
    .A2(net36),
    .Y(_051_),
    .B1(net110));
 sg13g2_nand2_1 _332_ (.Y(_149_),
    .A(net113),
    .B(net42));
 sg13g2_nor2_1 _333_ (.A(net106),
    .B(net42),
    .Y(_150_));
 sg13g2_a21oi_1 _334_ (.A1(net113),
    .A2(net42),
    .Y(_151_),
    .B1(net107));
 sg13g2_nor2_1 _335_ (.A(_099_),
    .B(_151_),
    .Y(_052_));
 sg13g2_nor2_1 _336_ (.A(net90),
    .B(net36),
    .Y(_152_));
 sg13g2_a21oi_1 _337_ (.A1(net75),
    .A2(net36),
    .Y(_055_),
    .B1(net91));
 sg13g2_nor2_1 _338_ (.A(net101),
    .B(_147_),
    .Y(_153_));
 sg13g2_a21oi_1 _339_ (.A1(net76),
    .A2(_147_),
    .Y(_056_),
    .B1(net102));
 sg13g2_mux2_1 _340_ (.A0(net132),
    .A1(net71),
    .S(_147_),
    .X(_057_));
 sg13g2_mux2_1 _341_ (.A0(net134),
    .A1(net73),
    .S(net36),
    .X(_058_));
 sg13g2_mux2_1 _342_ (.A0(net136),
    .A1(net74),
    .S(net36),
    .X(_059_));
 sg13g2_mux2_1 _343_ (.A0(net121),
    .A1(net72),
    .S(net36),
    .X(_060_));
 sg13g2_mux2_1 _344_ (.A0(net130),
    .A1(\spi_decoder_mod.o_reg_wdata[7] ),
    .S(net36),
    .X(_061_));
 sg13g2_or2_1 _345_ (.X(_154_),
    .B(_146_),
    .A(_097_));
 sg13g2_nand2_1 _346_ (.Y(_155_),
    .A(net116),
    .B(net35));
 sg13g2_o21ai_1 _347_ (.B1(_155_),
    .Y(_062_),
    .A1(_098_),
    .A2(net35));
 sg13g2_mux2_1 _348_ (.A0(net75),
    .A1(net156),
    .S(net35),
    .X(_063_));
 sg13g2_mux2_1 _349_ (.A0(net76),
    .A1(net161),
    .S(net35),
    .X(_064_));
 sg13g2_mux2_1 _350_ (.A0(net71),
    .A1(net146),
    .S(_154_),
    .X(_065_));
 sg13g2_mux2_1 _351_ (.A0(net73),
    .A1(net155),
    .S(net35),
    .X(_066_));
 sg13g2_mux2_1 _352_ (.A0(net74),
    .A1(net157),
    .S(net35),
    .X(_067_));
 sg13g2_mux2_1 _353_ (.A0(net72),
    .A1(net154),
    .S(net35),
    .X(_068_));
 sg13g2_mux2_1 _354_ (.A0(net140),
    .A1(\mod_ro_prog.osc_gen[7].inv.i_en ),
    .S(net35),
    .X(_069_));
 sg13g2_o21ai_1 _355_ (.B1(net47),
    .Y(_156_),
    .A1(net42),
    .A2(net99));
 sg13g2_a21oi_1 _356_ (.A1(net42),
    .A2(net99),
    .Y(_071_),
    .B1(_156_));
 sg13g2_a21oi_1 _357_ (.A1(net42),
    .A2(\dpll.n_count[0] ),
    .Y(_157_),
    .B1(net95));
 sg13g2_nand3_1 _358_ (.B(net95),
    .C(net99),
    .A(net143),
    .Y(_158_));
 sg13g2_nand2_1 _359_ (.Y(_159_),
    .A(net47),
    .B(_158_));
 sg13g2_nor2_1 _360_ (.A(net96),
    .B(_159_),
    .Y(_072_));
 sg13g2_or2_1 _361_ (.X(_160_),
    .B(_158_),
    .A(_096_));
 sg13g2_nand2_1 _362_ (.Y(_161_),
    .A(net48),
    .B(_160_));
 sg13g2_a21oi_1 _363_ (.A1(_096_),
    .A2(_158_),
    .Y(_073_),
    .B1(_161_));
 sg13g2_and2_1 _364_ (.A(_095_),
    .B(_160_),
    .X(_162_));
 sg13g2_nor2_2 _365_ (.A(_095_),
    .B(_160_),
    .Y(_163_));
 sg13g2_nor3_1 _366_ (.A(_099_),
    .B(_162_),
    .C(_163_),
    .Y(_074_));
 sg13g2_xnor2_1 _367_ (.Y(_164_),
    .A(net158),
    .B(_163_));
 sg13g2_nor2_1 _368_ (.A(_099_),
    .B(_164_),
    .Y(_075_));
 sg13g2_a21oi_1 _369_ (.A1(net158),
    .A2(_163_),
    .Y(_165_),
    .B1(net41));
 sg13g2_nand3_1 _370_ (.B(net158),
    .C(_163_),
    .A(net41),
    .Y(_166_));
 sg13g2_nand2_1 _371_ (.Y(_167_),
    .A(net48),
    .B(_166_));
 sg13g2_nor2_1 _372_ (.A(net159),
    .B(_167_),
    .Y(_076_));
 sg13g2_o21ai_1 _373_ (.B1(net48),
    .Y(_168_),
    .A1(_093_),
    .A2(_166_));
 sg13g2_a21oi_1 _374_ (.A1(_093_),
    .A2(_166_),
    .Y(_077_),
    .B1(_168_));
 sg13g2_nand2b_1 _375_ (.Y(_169_),
    .B(net80),
    .A_N(net42));
 sg13g2_a21oi_1 _376_ (.A1(net114),
    .A2(_169_),
    .Y(_078_),
    .B1(_099_));
 sg13g2_nor2b_1 _377_ (.A(net82),
    .B_N(net42),
    .Y(_170_));
 sg13g2_nor3_1 _378_ (.A(_099_),
    .B(net107),
    .C(_170_),
    .Y(_079_));
 sg13g2_o21ai_1 _379_ (.B1(net47),
    .Y(_171_),
    .A1(\dpll.id_decrement ),
    .A2(\dpll.k_count_borrow ));
 sg13g2_a21oi_1 _380_ (.A1(\dpll.id_decrement ),
    .A2(net82),
    .Y(_080_),
    .B1(_171_));
 sg13g2_o21ai_1 _381_ (.B1(net47),
    .Y(_172_),
    .A1(\dpll.id_increment ),
    .A2(\dpll.k_count_carry ));
 sg13g2_a21oi_1 _382_ (.A1(\dpll.id_increment ),
    .A2(net80),
    .Y(_081_),
    .B1(_172_));
 sg13g2_xor2_1 _383_ (.B(net6),
    .A(net144),
    .X(_173_));
 sg13g2_nor2_2 _384_ (.A(_099_),
    .B(_173_),
    .Y(_174_));
 sg13g2_nor2_1 _385_ (.A(_092_),
    .B(_174_),
    .Y(_175_));
 sg13g2_nand2_2 _386_ (.Y(_176_),
    .A(net48),
    .B(_173_));
 sg13g2_a21oi_1 _387_ (.A1(_092_),
    .A2(_176_),
    .Y(_082_),
    .B1(_175_));
 sg13g2_nand2_1 _388_ (.Y(_177_),
    .A(net125),
    .B(_174_));
 sg13g2_nor2b_1 _389_ (.A(net40),
    .B_N(\dpll.k_count[1] ),
    .Y(_178_));
 sg13g2_xnor2_1 _390_ (.Y(_179_),
    .A(net125),
    .B(net40));
 sg13g2_xnor2_1 _391_ (.Y(_180_),
    .A(\dpll.k_count[0] ),
    .B(_179_));
 sg13g2_o21ai_1 _392_ (.B1(net126),
    .Y(_083_),
    .A1(_176_),
    .A2(_180_));
 sg13g2_nand2_1 _393_ (.Y(_181_),
    .A(net138),
    .B(net37));
 sg13g2_nor2b_1 _394_ (.A(net39),
    .B_N(net138),
    .Y(_182_));
 sg13g2_xnor2_1 _395_ (.Y(_183_),
    .A(net138),
    .B(net39));
 sg13g2_a21o_2 _396_ (.A2(_179_),
    .A1(\dpll.k_count[0] ),
    .B1(_178_),
    .X(_184_));
 sg13g2_xnor2_1 _397_ (.Y(_185_),
    .A(_183_),
    .B(_184_));
 sg13g2_o21ai_1 _398_ (.B1(_181_),
    .Y(_084_),
    .A1(_176_),
    .A2(_185_));
 sg13g2_a21oi_1 _399_ (.A1(_183_),
    .A2(_184_),
    .Y(_186_),
    .B1(_182_));
 sg13g2_nor2_1 _400_ (.A(\dpll.k_count[3] ),
    .B(_094_),
    .Y(_187_));
 sg13g2_xor2_1 _401_ (.B(net39),
    .A(net151),
    .X(_188_));
 sg13g2_xnor2_1 _402_ (.Y(_189_),
    .A(_186_),
    .B(_188_));
 sg13g2_nand2_1 _403_ (.Y(_190_),
    .A(net151),
    .B(net37));
 sg13g2_o21ai_1 _404_ (.B1(_190_),
    .Y(_085_),
    .A1(_176_),
    .A2(_189_));
 sg13g2_nand2_1 _405_ (.Y(_191_),
    .A(net128),
    .B(net37));
 sg13g2_nor2b_1 _406_ (.A(net39),
    .B_N(\dpll.k_count[4] ),
    .Y(_192_));
 sg13g2_xor2_1 _407_ (.B(net39),
    .A(net128),
    .X(_193_));
 sg13g2_a221oi_1 _408_ (.B2(_184_),
    .C1(_182_),
    .B1(_183_),
    .A1(\dpll.k_count[3] ),
    .Y(_194_),
    .A2(_094_));
 sg13g2_nor2_1 _409_ (.A(_187_),
    .B(_194_),
    .Y(_195_));
 sg13g2_nor3_1 _410_ (.A(_187_),
    .B(_193_),
    .C(_194_),
    .Y(_196_));
 sg13g2_xor2_1 _411_ (.B(_195_),
    .A(_193_),
    .X(_197_));
 sg13g2_o21ai_1 _412_ (.B1(_191_),
    .Y(_086_),
    .A1(_176_),
    .A2(_197_));
 sg13g2_xnor2_1 _413_ (.Y(_198_),
    .A(net164),
    .B(net39));
 sg13g2_nor3_1 _414_ (.A(_192_),
    .B(_196_),
    .C(_198_),
    .Y(_199_));
 sg13g2_o21ai_1 _415_ (.B1(_198_),
    .Y(_200_),
    .A1(_192_),
    .A2(_196_));
 sg13g2_nor2_1 _416_ (.A(_176_),
    .B(_199_),
    .Y(_201_));
 sg13g2_a22oi_1 _417_ (.Y(_202_),
    .B1(_200_),
    .B2(_201_),
    .A2(net37),
    .A1(net164));
 sg13g2_inv_1 _418_ (.Y(_087_),
    .A(net165));
 sg13g2_nand2_1 _419_ (.Y(_203_),
    .A(net119),
    .B(net37));
 sg13g2_nand2_1 _420_ (.Y(_204_),
    .A(\dpll.k_count[6] ),
    .B(_094_));
 sg13g2_xor2_1 _421_ (.B(net39),
    .A(net119),
    .X(_205_));
 sg13g2_nor2b_1 _422_ (.A(_193_),
    .B_N(_198_),
    .Y(_206_));
 sg13g2_a221oi_1 _423_ (.B2(_206_),
    .C1(_192_),
    .B1(_195_),
    .A1(\dpll.k_count[5] ),
    .Y(_207_),
    .A2(_094_));
 sg13g2_xnor2_1 _424_ (.Y(_208_),
    .A(_205_),
    .B(_207_));
 sg13g2_o21ai_1 _425_ (.B1(_203_),
    .Y(_088_),
    .A1(_176_),
    .A2(_208_));
 sg13g2_nand2_1 _426_ (.Y(_209_),
    .A(net117),
    .B(net37));
 sg13g2_o21ai_1 _427_ (.B1(_204_),
    .Y(_210_),
    .A1(_205_),
    .A2(_207_));
 sg13g2_xnor2_1 _428_ (.Y(_211_),
    .A(net117),
    .B(net41));
 sg13g2_xnor2_1 _429_ (.Y(_212_),
    .A(_210_),
    .B(_211_));
 sg13g2_o21ai_1 _430_ (.B1(_209_),
    .Y(_089_),
    .A1(_176_),
    .A2(_212_));
 sg13g2_nand2_1 _431_ (.Y(_213_),
    .A(_094_),
    .B(net47));
 sg13g2_nor4_1 _432_ (.A(\dpll.k_count[3] ),
    .B(\dpll.k_count[2] ),
    .C(\dpll.k_count[1] ),
    .D(\dpll.k_count[0] ),
    .Y(_214_));
 sg13g2_nor4_1 _433_ (.A(\dpll.k_count[7] ),
    .B(\dpll.k_count[6] ),
    .C(\dpll.k_count[5] ),
    .D(\dpll.k_count[4] ),
    .Y(_215_));
 sg13g2_a21oi_1 _434_ (.A1(_214_),
    .A2(_215_),
    .Y(_216_),
    .B1(_213_));
 sg13g2_a21oi_1 _435_ (.A1(_094_),
    .A2(net47),
    .Y(_217_),
    .B1(net86));
 sg13g2_nor3_1 _436_ (.A(net37),
    .B(_216_),
    .C(_217_),
    .Y(_090_));
 sg13g2_nand3_1 _437_ (.B(\dpll.k_count[2] ),
    .C(\dpll.k_count[1] ),
    .A(\dpll.k_count[3] ),
    .Y(_218_));
 sg13g2_nand4_1 _438_ (.B(\dpll.k_count[6] ),
    .C(\dpll.k_count[5] ),
    .A(\dpll.k_count[7] ),
    .Y(_219_),
    .D(\dpll.k_count[4] ));
 sg13g2_nor3_1 _439_ (.A(_092_),
    .B(_218_),
    .C(_219_),
    .Y(_220_));
 sg13g2_nor3_1 _440_ (.A(_094_),
    .B(_099_),
    .C(_220_),
    .Y(_221_));
 sg13g2_a21oi_1 _441_ (.A1(net40),
    .A2(net47),
    .Y(_222_),
    .B1(net88));
 sg13g2_nor3_1 _442_ (.A(net37),
    .B(_221_),
    .C(_222_),
    .Y(_091_));
 sg13g2_inv_1 _443_ (.Y(_034_),
    .A(net43));
 sg13g2_inv_1 _444_ (.Y(_032_),
    .A(net43));
 sg13g2_inv_1 _445_ (.Y(_030_),
    .A(net43));
 sg13g2_inv_1 _446_ (.Y(_028_),
    .A(net44));
 sg13g2_inv_1 _447_ (.Y(_026_),
    .A(net44));
 sg13g2_inv_1 _448_ (.Y(_024_),
    .A(net44));
 sg13g2_inv_1 _449_ (.Y(_022_),
    .A(net43));
 sg13g2_inv_1 _450_ (.Y(_018_),
    .A(net43));
 sg13g2_inv_1 _451_ (.Y(_019_),
    .A(net45));
 sg13g2_inv_1 _452_ (.Y(_020_),
    .A(net46));
 sg13g2_inv_1 _453_ (.Y(_021_),
    .A(net45));
 sg13g2_inv_1 _455__3 (.Y(net65),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _456__4 (.Y(net66),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _457__5 (.Y(net67),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _458__6 (.Y(net68),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _459__7 (.Y(net69),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _460__8 (.Y(net70),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_inv_1 _461_ (.Y(_038_),
    .A(net45));
 sg13g2_inv_1 _462_ (.Y(_039_),
    .A(net44));
 sg13g2_inv_1 _463_ (.Y(_040_),
    .A(net44));
 sg13g2_inv_1 _464_ (.Y(_041_),
    .A(net46));
 sg13g2_inv_1 _465_ (.Y(_042_),
    .A(net45));
 sg13g2_inv_1 _466_ (.Y(_043_),
    .A(net44));
 sg13g2_inv_1 _467_ (.Y(_044_),
    .A(net44));
 sg13g2_inv_1 _468_ (.Y(_045_),
    .A(net44));
 sg13g2_inv_1 _469_ (.Y(_046_),
    .A(net43));
 sg13g2_inv_1 _470_ (.Y(_047_),
    .A(net43));
 sg13g2_inv_1 _471_ (.Y(_048_),
    .A(net43));
 sg13g2_inv_1 _472_ (.Y(_049_),
    .A(net45));
 sg13g2_inv_1 _473_ (.Y(_050_),
    .A(net45));
 sg13g2_dfrbpq_1 _474_ (.RESET_B(net49),
    .D(net111),
    .Q(\spi_regfile_mod.SYS_CTRL_RESET_q [0]),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _475_ (.RESET_B(_018_),
    .D(_017_),
    .Q(_014_),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _476_ (.RESET_B(_019_),
    .D(net94),
    .Q(\spi_decoder_mod.spi_state[1] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _477_ (.RESET_B(_020_),
    .D(net78),
    .Q(\spi_decoder_mod.spi_state[2] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_2 _478_ (.RESET_B(_021_),
    .D(net124),
    .Q(\spi_decoder_mod.spi_state[3] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _479_ (.RESET_B(_022_),
    .D(_003_),
    .Q(\spi_decoder_mod.shift_out_reg[0] ),
    .CLK(net63));
 sg13g2_dfrbpq_1 _480_ (.RESET_B(_024_),
    .D(_004_),
    .Q(\spi_decoder_mod.shift_out_reg[1] ),
    .CLK(net64));
 sg13g2_dfrbpq_1 _481_ (.RESET_B(_026_),
    .D(_005_),
    .Q(\spi_decoder_mod.shift_out_reg[2] ),
    .CLK(net65));
 sg13g2_dfrbpq_1 _482_ (.RESET_B(_028_),
    .D(_006_),
    .Q(\spi_decoder_mod.shift_out_reg[3] ),
    .CLK(net66));
 sg13g2_dfrbpq_1 _483_ (.RESET_B(_030_),
    .D(_007_),
    .Q(\spi_decoder_mod.shift_out_reg[4] ),
    .CLK(net67));
 sg13g2_dfrbpq_1 _484_ (.RESET_B(_032_),
    .D(_008_),
    .Q(\spi_decoder_mod.shift_out_reg[5] ),
    .CLK(net68));
 sg13g2_dfrbpq_1 _485_ (.RESET_B(_034_),
    .D(_009_),
    .Q(\spi_decoder_mod.shift_out_reg[6] ),
    .CLK(net69));
 sg13g2_dfrbpq_1 _486_ (.RESET_B(_036_),
    .D(_010_),
    .Q(o_miso),
    .CLK(net70));
 sg13g2_dfrbpq_1 _487_ (.RESET_B(net31),
    .D(_052_),
    .Q(\dpll.id_out ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _488_ (.RESET_B(_038_),
    .D(_011_),
    .Q(\spi_decoder_mod.shift_cnt[0] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_2 _489_ (.RESET_B(_039_),
    .D(_012_),
    .Q(\spi_decoder_mod.shift_cnt[1] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _490_ (.RESET_B(_040_),
    .D(_013_),
    .Q(\spi_decoder_mod.shift_cnt[2] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _491_ (.RESET_B(_041_),
    .D(_053_),
    .Q(\spi_decoder_mod.start ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _492_ (.RESET_B(_042_),
    .D(net5),
    .Q(\spi_decoder_mod.o_reg_wdata[1] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _493_ (.RESET_B(_043_),
    .D(net75),
    .Q(\spi_decoder_mod.o_reg_wdata[2] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _494_ (.RESET_B(_044_),
    .D(net76),
    .Q(\spi_decoder_mod.o_reg_wdata[3] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _495_ (.RESET_B(_045_),
    .D(net71),
    .Q(\spi_decoder_mod.o_reg_wdata[4] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _496_ (.RESET_B(_046_),
    .D(net73),
    .Q(\spi_decoder_mod.o_reg_wdata[5] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _497_ (.RESET_B(_047_),
    .D(net74),
    .Q(\spi_decoder_mod.o_reg_wdata[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _498_ (.RESET_B(_048_),
    .D(net72),
    .Q(\spi_decoder_mod.o_reg_wdata[7] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _499_ (.RESET_B(_049_),
    .D(_054_),
    .Q(\spi_decoder_mod.write ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _500_ (.RESET_B(net50),
    .D(net92),
    .Q(_015_),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _501_ (.RESET_B(net50),
    .D(net103),
    .Q(_016_),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _502_ (.RESET_B(net50),
    .D(net133),
    .Q(\reg_echo[2] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _503_ (.RESET_B(net49),
    .D(net135),
    .Q(\reg_echo[3] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _504_ (.RESET_B(net49),
    .D(net137),
    .Q(\reg_echo[4] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _505_ (.RESET_B(net49),
    .D(net122),
    .Q(\reg_echo[5] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _506_ (.RESET_B(net49),
    .D(net131),
    .Q(\reg_echo[6] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _507_ (.RESET_B(net50),
    .D(_062_),
    .Q(\mod_ro_prog.osc_gen[0].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _508_ (.RESET_B(net50),
    .D(_063_),
    .Q(\mod_ro_prog.osc_gen[1].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _509_ (.RESET_B(net50),
    .D(_064_),
    .Q(\mod_ro_prog.osc_gen[2].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _510_ (.RESET_B(net50),
    .D(_065_),
    .Q(\mod_ro_prog.osc_gen[3].inv.i_en ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _511_ (.RESET_B(net49),
    .D(_066_),
    .Q(\mod_ro_prog.osc_gen[4].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _512_ (.RESET_B(net49),
    .D(_067_),
    .Q(\mod_ro_prog.osc_gen[5].inv.i_en ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _513_ (.RESET_B(net48),
    .D(_068_),
    .Q(\mod_ro_prog.osc_gen[6].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _514_ (.RESET_B(net49),
    .D(net141),
    .Q(\mod_ro_prog.osc_gen[7].inv.i_en ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_2 _515_ (.RESET_B(_050_),
    .D(net167),
    .Q(\spi_regfile_mod.addr [0]),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_2 _516_ (.RESET_B(net61),
    .D(net100),
    .Q(\dpll.n_count[0] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _517_ (.RESET_B(net59),
    .D(net97),
    .Q(\dpll.n_count[1] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _518_ (.RESET_B(net57),
    .D(net105),
    .Q(\dpll.n_count[2] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _519_ (.RESET_B(net55),
    .D(_074_),
    .Q(\dpll.clk8x_fout ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _520_ (.RESET_B(net53),
    .D(_075_),
    .Q(\dpll.n_count[4] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _521_ (.RESET_B(net51),
    .D(net160),
    .Q(\dpll.n_count[5] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _522_ (.RESET_B(net34),
    .D(net145),
    .Q(\dpll.clk_fout ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _523_ (.RESET_B(net32),
    .D(net115),
    .Q(\dpll.id_increment_done ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _524_ (.RESET_B(net29),
    .D(net108),
    .Q(\dpll.id_decrement_done ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net27),
    .D(net83),
    .Q(\dpll.id_decrement ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _526_ (.RESET_B(net25),
    .D(net81),
    .Q(\dpll.id_increment ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _527_ (.RESET_B(net60),
    .D(_082_),
    .Q(\dpll.k_count[0] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_2 _528_ (.RESET_B(net56),
    .D(net127),
    .Q(\dpll.k_count[1] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _529_ (.RESET_B(net52),
    .D(net139),
    .Q(\dpll.k_count[2] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _530_ (.RESET_B(net33),
    .D(_085_),
    .Q(\dpll.k_count[3] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _531_ (.RESET_B(net28),
    .D(net129),
    .Q(\dpll.k_count[4] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _532_ (.RESET_B(net62),
    .D(_087_),
    .Q(\dpll.k_count[5] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _533_ (.RESET_B(net54),
    .D(net120),
    .Q(\dpll.k_count[6] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _534_ (.RESET_B(net30),
    .D(net118),
    .Q(\dpll.k_count[7] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net58),
    .D(net87),
    .Q(\dpll.k_count_borrow ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net26),
    .D(net89),
    .Q(\dpll.k_count_carry ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_tiehi _536__26 (.L_HI(net26));
 sg13g2_tiehi _525__27 (.L_HI(net27));
 sg13g2_tiehi _531__28 (.L_HI(net28));
 sg13g2_tiehi _524__29 (.L_HI(net29));
 sg13g2_tiehi _534__30 (.L_HI(net30));
 sg13g2_tiehi _487__31 (.L_HI(net31));
 sg13g2_tiehi _523__32 (.L_HI(net32));
 sg13g2_tiehi _530__33 (.L_HI(net33));
 sg13g2_tiehi _522__34 (.L_HI(net34));
 sg13g2_tiehi _521__35 (.L_HI(net51));
 sg13g2_tiehi _529__36 (.L_HI(net52));
 sg13g2_tiehi _520__37 (.L_HI(net53));
 sg13g2_tiehi _533__38 (.L_HI(net54));
 sg13g2_tiehi _519__39 (.L_HI(net55));
 sg13g2_tiehi _528__40 (.L_HI(net56));
 sg13g2_tiehi _518__41 (.L_HI(net57));
 sg13g2_tiehi _535__42 (.L_HI(net58));
 sg13g2_tiehi _517__43 (.L_HI(net59));
 sg13g2_tiehi _527__44 (.L_HI(net60));
 sg13g2_tiehi _516__45 (.L_HI(net61));
 sg13g2_tiehi _532__46 (.L_HI(net62));
 sg13g2_inv_1 _255__1 (.Y(net63),
    .A(clknet_1_1__leaf_clk));
 sg13g2_tielo tt_um_mlyoung_wedgetail_8 (.L_LO(net8));
 sg13g2_tielo tt_um_mlyoung_wedgetail_9 (.L_LO(net9));
 sg13g2_tielo tt_um_mlyoung_wedgetail_10 (.L_LO(net10));
 sg13g2_tielo tt_um_mlyoung_wedgetail_11 (.L_LO(net11));
 sg13g2_tielo tt_um_mlyoung_wedgetail_12 (.L_LO(net12));
 sg13g2_tielo tt_um_mlyoung_wedgetail_13 (.L_LO(net13));
 sg13g2_tielo tt_um_mlyoung_wedgetail_14 (.L_LO(net14));
 sg13g2_tielo tt_um_mlyoung_wedgetail_15 (.L_LO(net15));
 sg13g2_tielo tt_um_mlyoung_wedgetail_16 (.L_LO(net16));
 sg13g2_tielo tt_um_mlyoung_wedgetail_17 (.L_LO(net17));
 sg13g2_tielo tt_um_mlyoung_wedgetail_18 (.L_LO(net18));
 sg13g2_tielo tt_um_mlyoung_wedgetail_19 (.L_LO(net19));
 sg13g2_tielo tt_um_mlyoung_wedgetail_20 (.L_LO(net20));
 sg13g2_tielo tt_um_mlyoung_wedgetail_21 (.L_LO(net21));
 sg13g2_tielo tt_um_mlyoung_wedgetail_22 (.L_LO(net22));
 sg13g2_tielo tt_um_mlyoung_wedgetail_23 (.L_LO(net23));
 sg13g2_tielo tt_um_mlyoung_wedgetail_24 (.L_LO(net24));
 sg13g2_tiehi _526__25 (.L_HI(net25));
 sg13g2_buf_1 _577_ (.A(o_rosc_mux_out),
    .X(uo_out[0]));
 sg13g2_buf_1 _578_ (.A(\mod_ro_32_raw.fabric[0] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _579_ (.A(\dpll.clk_fout ),
    .X(uo_out[3]));
 sg13g2_buf_1 _580_ (.A(\dpll.clk8x_fout ),
    .X(uo_out[4]));
 sg13g2_buf_1 _581_ (.A(o_miso),
    .X(uo_out[5]));
 sg13g2_buf_1 _582_ (.A(\mod_ro_prog.fabric[0] ),
    .X(uo_out[6]));
 sg13g2_inv_1 \mod_ro_128.feedback  (.Y(\mod_ro_128.fabric[0] ),
    .A(\mod_ro_128.fabric[128] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[0].inv  (.Y(\mod_ro_128.fabric[1] ),
    .A(\mod_ro_128.fabric[0] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[100].inv  (.Y(\mod_ro_128.fabric[101] ),
    .A(\mod_ro_128.fabric[100] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[101].inv  (.Y(\mod_ro_128.fabric[102] ),
    .A(\mod_ro_128.fabric[101] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[102].inv  (.Y(\mod_ro_128.fabric[103] ),
    .A(\mod_ro_128.fabric[102] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[103].inv  (.Y(\mod_ro_128.fabric[104] ),
    .A(\mod_ro_128.fabric[103] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[104].inv  (.Y(\mod_ro_128.fabric[105] ),
    .A(\mod_ro_128.fabric[104] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[105].inv  (.Y(\mod_ro_128.fabric[106] ),
    .A(\mod_ro_128.fabric[105] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[106].inv  (.Y(\mod_ro_128.fabric[107] ),
    .A(\mod_ro_128.fabric[106] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[107].inv  (.Y(\mod_ro_128.fabric[108] ),
    .A(\mod_ro_128.fabric[107] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[108].inv  (.Y(\mod_ro_128.fabric[109] ),
    .A(\mod_ro_128.fabric[108] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[109].inv  (.Y(\mod_ro_128.fabric[110] ),
    .A(\mod_ro_128.fabric[109] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[10].inv  (.Y(\mod_ro_128.fabric[11] ),
    .A(\mod_ro_128.fabric[10] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[110].inv  (.Y(\mod_ro_128.fabric[111] ),
    .A(\mod_ro_128.fabric[110] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[111].inv  (.Y(\mod_ro_128.fabric[112] ),
    .A(\mod_ro_128.fabric[111] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[112].inv  (.Y(\mod_ro_128.fabric[113] ),
    .A(\mod_ro_128.fabric[112] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[113].inv  (.Y(\mod_ro_128.fabric[114] ),
    .A(\mod_ro_128.fabric[113] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[114].inv  (.Y(\mod_ro_128.fabric[115] ),
    .A(\mod_ro_128.fabric[114] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[115].inv  (.Y(\mod_ro_128.fabric[116] ),
    .A(\mod_ro_128.fabric[115] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[116].inv  (.Y(\mod_ro_128.fabric[117] ),
    .A(\mod_ro_128.fabric[116] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[117].inv  (.Y(\mod_ro_128.fabric[118] ),
    .A(\mod_ro_128.fabric[117] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[118].inv  (.Y(\mod_ro_128.fabric[119] ),
    .A(\mod_ro_128.fabric[118] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[119].inv  (.Y(\mod_ro_128.fabric[120] ),
    .A(\mod_ro_128.fabric[119] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[11].inv  (.Y(\mod_ro_128.fabric[12] ),
    .A(\mod_ro_128.fabric[11] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[120].inv  (.Y(\mod_ro_128.fabric[121] ),
    .A(\mod_ro_128.fabric[120] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[121].inv  (.Y(\mod_ro_128.fabric[122] ),
    .A(\mod_ro_128.fabric[121] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[122].inv  (.Y(\mod_ro_128.fabric[123] ),
    .A(\mod_ro_128.fabric[122] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[123].inv  (.Y(\mod_ro_128.fabric[124] ),
    .A(\mod_ro_128.fabric[123] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[124].inv  (.Y(\mod_ro_128.fabric[125] ),
    .A(\mod_ro_128.fabric[124] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[125].inv  (.Y(\mod_ro_128.fabric[126] ),
    .A(\mod_ro_128.fabric[125] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[126].inv  (.Y(\mod_ro_128.fabric[127] ),
    .A(\mod_ro_128.fabric[126] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[127].inv  (.Y(\mod_ro_128.fabric[128] ),
    .A(\mod_ro_128.fabric[127] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[12].inv  (.Y(\mod_ro_128.fabric[13] ),
    .A(\mod_ro_128.fabric[12] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[13].inv  (.Y(\mod_ro_128.fabric[14] ),
    .A(\mod_ro_128.fabric[13] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[14].inv  (.Y(\mod_ro_128.fabric[15] ),
    .A(\mod_ro_128.fabric[14] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[15].inv  (.Y(\mod_ro_128.fabric[16] ),
    .A(\mod_ro_128.fabric[15] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[16].inv  (.Y(\mod_ro_128.fabric[17] ),
    .A(\mod_ro_128.fabric[16] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[17].inv  (.Y(\mod_ro_128.fabric[18] ),
    .A(\mod_ro_128.fabric[17] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[18].inv  (.Y(\mod_ro_128.fabric[19] ),
    .A(\mod_ro_128.fabric[18] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[19].inv  (.Y(\mod_ro_128.fabric[20] ),
    .A(\mod_ro_128.fabric[19] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[1].inv  (.Y(\mod_ro_128.fabric[2] ),
    .A(\mod_ro_128.fabric[1] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[20].inv  (.Y(\mod_ro_128.fabric[21] ),
    .A(\mod_ro_128.fabric[20] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[21].inv  (.Y(\mod_ro_128.fabric[22] ),
    .A(\mod_ro_128.fabric[21] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[22].inv  (.Y(\mod_ro_128.fabric[23] ),
    .A(\mod_ro_128.fabric[22] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[23].inv  (.Y(\mod_ro_128.fabric[24] ),
    .A(\mod_ro_128.fabric[23] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[24].inv  (.Y(\mod_ro_128.fabric[25] ),
    .A(\mod_ro_128.fabric[24] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[25].inv  (.Y(\mod_ro_128.fabric[26] ),
    .A(\mod_ro_128.fabric[25] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[26].inv  (.Y(\mod_ro_128.fabric[27] ),
    .A(\mod_ro_128.fabric[26] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[27].inv  (.Y(\mod_ro_128.fabric[28] ),
    .A(\mod_ro_128.fabric[27] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[28].inv  (.Y(\mod_ro_128.fabric[29] ),
    .A(\mod_ro_128.fabric[28] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[29].inv  (.Y(\mod_ro_128.fabric[30] ),
    .A(\mod_ro_128.fabric[29] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[2].inv  (.Y(\mod_ro_128.fabric[3] ),
    .A(\mod_ro_128.fabric[2] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[30].inv  (.Y(\mod_ro_128.fabric[31] ),
    .A(\mod_ro_128.fabric[30] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[31].inv  (.Y(\mod_ro_128.fabric[32] ),
    .A(\mod_ro_128.fabric[31] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[32].inv  (.Y(\mod_ro_128.fabric[33] ),
    .A(\mod_ro_128.fabric[32] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[33].inv  (.Y(\mod_ro_128.fabric[34] ),
    .A(\mod_ro_128.fabric[33] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[34].inv  (.Y(\mod_ro_128.fabric[35] ),
    .A(\mod_ro_128.fabric[34] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[35].inv  (.Y(\mod_ro_128.fabric[36] ),
    .A(\mod_ro_128.fabric[35] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[36].inv  (.Y(\mod_ro_128.fabric[37] ),
    .A(\mod_ro_128.fabric[36] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[37].inv  (.Y(\mod_ro_128.fabric[38] ),
    .A(\mod_ro_128.fabric[37] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[38].inv  (.Y(\mod_ro_128.fabric[39] ),
    .A(\mod_ro_128.fabric[38] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[39].inv  (.Y(\mod_ro_128.fabric[40] ),
    .A(\mod_ro_128.fabric[39] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[3].inv  (.Y(\mod_ro_128.fabric[4] ),
    .A(\mod_ro_128.fabric[3] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[40].inv  (.Y(\mod_ro_128.fabric[41] ),
    .A(\mod_ro_128.fabric[40] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[41].inv  (.Y(\mod_ro_128.fabric[42] ),
    .A(\mod_ro_128.fabric[41] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[42].inv  (.Y(\mod_ro_128.fabric[43] ),
    .A(\mod_ro_128.fabric[42] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[43].inv  (.Y(\mod_ro_128.fabric[44] ),
    .A(\mod_ro_128.fabric[43] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[44].inv  (.Y(\mod_ro_128.fabric[45] ),
    .A(\mod_ro_128.fabric[44] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[45].inv  (.Y(\mod_ro_128.fabric[46] ),
    .A(\mod_ro_128.fabric[45] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[46].inv  (.Y(\mod_ro_128.fabric[47] ),
    .A(\mod_ro_128.fabric[46] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[47].inv  (.Y(\mod_ro_128.fabric[48] ),
    .A(\mod_ro_128.fabric[47] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[48].inv  (.Y(\mod_ro_128.fabric[49] ),
    .A(\mod_ro_128.fabric[48] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[49].inv  (.Y(\mod_ro_128.fabric[50] ),
    .A(\mod_ro_128.fabric[49] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[4].inv  (.Y(\mod_ro_128.fabric[5] ),
    .A(\mod_ro_128.fabric[4] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[50].inv  (.Y(\mod_ro_128.fabric[51] ),
    .A(\mod_ro_128.fabric[50] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[51].inv  (.Y(\mod_ro_128.fabric[52] ),
    .A(\mod_ro_128.fabric[51] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[52].inv  (.Y(\mod_ro_128.fabric[53] ),
    .A(\mod_ro_128.fabric[52] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[53].inv  (.Y(\mod_ro_128.fabric[54] ),
    .A(\mod_ro_128.fabric[53] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[54].inv  (.Y(\mod_ro_128.fabric[55] ),
    .A(\mod_ro_128.fabric[54] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[55].inv  (.Y(\mod_ro_128.fabric[56] ),
    .A(\mod_ro_128.fabric[55] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[56].inv  (.Y(\mod_ro_128.fabric[57] ),
    .A(\mod_ro_128.fabric[56] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[57].inv  (.Y(\mod_ro_128.fabric[58] ),
    .A(\mod_ro_128.fabric[57] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[58].inv  (.Y(\mod_ro_128.fabric[59] ),
    .A(\mod_ro_128.fabric[58] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[59].inv  (.Y(\mod_ro_128.fabric[60] ),
    .A(\mod_ro_128.fabric[59] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[5].inv  (.Y(\mod_ro_128.fabric[6] ),
    .A(\mod_ro_128.fabric[5] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[60].inv  (.Y(\mod_ro_128.fabric[61] ),
    .A(\mod_ro_128.fabric[60] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[61].inv  (.Y(\mod_ro_128.fabric[62] ),
    .A(\mod_ro_128.fabric[61] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[62].inv  (.Y(\mod_ro_128.fabric[63] ),
    .A(\mod_ro_128.fabric[62] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[63].inv  (.Y(\mod_ro_128.fabric[64] ),
    .A(\mod_ro_128.fabric[63] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[64].inv  (.Y(\mod_ro_128.fabric[65] ),
    .A(\mod_ro_128.fabric[64] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[65].inv  (.Y(\mod_ro_128.fabric[66] ),
    .A(\mod_ro_128.fabric[65] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[66].inv  (.Y(\mod_ro_128.fabric[67] ),
    .A(\mod_ro_128.fabric[66] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[67].inv  (.Y(\mod_ro_128.fabric[68] ),
    .A(\mod_ro_128.fabric[67] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[68].inv  (.Y(\mod_ro_128.fabric[69] ),
    .A(\mod_ro_128.fabric[68] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[69].inv  (.Y(\mod_ro_128.fabric[70] ),
    .A(\mod_ro_128.fabric[69] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[6].inv  (.Y(\mod_ro_128.fabric[7] ),
    .A(\mod_ro_128.fabric[6] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[70].inv  (.Y(\mod_ro_128.fabric[71] ),
    .A(\mod_ro_128.fabric[70] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[71].inv  (.Y(\mod_ro_128.fabric[72] ),
    .A(\mod_ro_128.fabric[71] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[72].inv  (.Y(\mod_ro_128.fabric[73] ),
    .A(\mod_ro_128.fabric[72] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[73].inv  (.Y(\mod_ro_128.fabric[74] ),
    .A(\mod_ro_128.fabric[73] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[74].inv  (.Y(\mod_ro_128.fabric[75] ),
    .A(\mod_ro_128.fabric[74] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[75].inv  (.Y(\mod_ro_128.fabric[76] ),
    .A(\mod_ro_128.fabric[75] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[76].inv  (.Y(\mod_ro_128.fabric[77] ),
    .A(\mod_ro_128.fabric[76] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[77].inv  (.Y(\mod_ro_128.fabric[78] ),
    .A(\mod_ro_128.fabric[77] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[78].inv  (.Y(\mod_ro_128.fabric[79] ),
    .A(\mod_ro_128.fabric[78] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[79].inv  (.Y(\mod_ro_128.fabric[80] ),
    .A(\mod_ro_128.fabric[79] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[7].inv  (.Y(\mod_ro_128.fabric[8] ),
    .A(\mod_ro_128.fabric[7] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[80].inv  (.Y(\mod_ro_128.fabric[81] ),
    .A(\mod_ro_128.fabric[80] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[81].inv  (.Y(\mod_ro_128.fabric[82] ),
    .A(\mod_ro_128.fabric[81] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[82].inv  (.Y(\mod_ro_128.fabric[83] ),
    .A(\mod_ro_128.fabric[82] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[83].inv  (.Y(\mod_ro_128.fabric[84] ),
    .A(\mod_ro_128.fabric[83] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[84].inv  (.Y(\mod_ro_128.fabric[85] ),
    .A(\mod_ro_128.fabric[84] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[85].inv  (.Y(\mod_ro_128.fabric[86] ),
    .A(\mod_ro_128.fabric[85] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[86].inv  (.Y(\mod_ro_128.fabric[87] ),
    .A(\mod_ro_128.fabric[86] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[87].inv  (.Y(\mod_ro_128.fabric[88] ),
    .A(\mod_ro_128.fabric[87] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[88].inv  (.Y(\mod_ro_128.fabric[89] ),
    .A(\mod_ro_128.fabric[88] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[89].inv  (.Y(\mod_ro_128.fabric[90] ),
    .A(\mod_ro_128.fabric[89] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[8].inv  (.Y(\mod_ro_128.fabric[9] ),
    .A(\mod_ro_128.fabric[8] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[90].inv  (.Y(\mod_ro_128.fabric[91] ),
    .A(\mod_ro_128.fabric[90] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[91].inv  (.Y(\mod_ro_128.fabric[92] ),
    .A(\mod_ro_128.fabric[91] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[92].inv  (.Y(\mod_ro_128.fabric[93] ),
    .A(\mod_ro_128.fabric[92] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[93].inv  (.Y(\mod_ro_128.fabric[94] ),
    .A(\mod_ro_128.fabric[93] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[94].inv  (.Y(\mod_ro_128.fabric[95] ),
    .A(\mod_ro_128.fabric[94] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[95].inv  (.Y(\mod_ro_128.fabric[96] ),
    .A(\mod_ro_128.fabric[95] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[96].inv  (.Y(\mod_ro_128.fabric[97] ),
    .A(\mod_ro_128.fabric[96] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[97].inv  (.Y(\mod_ro_128.fabric[98] ),
    .A(\mod_ro_128.fabric[97] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[98].inv  (.Y(\mod_ro_128.fabric[99] ),
    .A(\mod_ro_128.fabric[98] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[99].inv  (.Y(\mod_ro_128.fabric[100] ),
    .A(\mod_ro_128.fabric[99] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[9].inv  (.Y(\mod_ro_128.fabric[10] ),
    .A(\mod_ro_128.fabric[9] ));
 sg13g2_inv_1 \mod_ro_16.feedback  (.Y(\mod_ro_16.fabric[0] ),
    .A(\mod_ro_16.fabric[16] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[0].inv  (.Y(\mod_ro_16.fabric[1] ),
    .A(\mod_ro_16.fabric[0] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[10].inv  (.Y(\mod_ro_16.fabric[11] ),
    .A(\mod_ro_16.fabric[10] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[11].inv  (.Y(\mod_ro_16.fabric[12] ),
    .A(\mod_ro_16.fabric[11] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[12].inv  (.Y(\mod_ro_16.fabric[13] ),
    .A(\mod_ro_16.fabric[12] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[13].inv  (.Y(\mod_ro_16.fabric[14] ),
    .A(\mod_ro_16.fabric[13] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[14].inv  (.Y(\mod_ro_16.fabric[15] ),
    .A(\mod_ro_16.fabric[14] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[15].inv  (.Y(\mod_ro_16.fabric[16] ),
    .A(\mod_ro_16.fabric[15] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[1].inv  (.Y(\mod_ro_16.fabric[2] ),
    .A(\mod_ro_16.fabric[1] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[2].inv  (.Y(\mod_ro_16.fabric[3] ),
    .A(\mod_ro_16.fabric[2] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[3].inv  (.Y(\mod_ro_16.fabric[4] ),
    .A(\mod_ro_16.fabric[3] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[4].inv  (.Y(\mod_ro_16.fabric[5] ),
    .A(\mod_ro_16.fabric[4] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[5].inv  (.Y(\mod_ro_16.fabric[6] ),
    .A(\mod_ro_16.fabric[5] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[6].inv  (.Y(\mod_ro_16.fabric[7] ),
    .A(\mod_ro_16.fabric[6] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[7].inv  (.Y(\mod_ro_16.fabric[8] ),
    .A(\mod_ro_16.fabric[7] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[8].inv  (.Y(\mod_ro_16.fabric[9] ),
    .A(\mod_ro_16.fabric[8] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[9].inv  (.Y(\mod_ro_16.fabric[10] ),
    .A(\mod_ro_16.fabric[9] ));
 sg13g2_inv_1 \mod_ro_256.feedback  (.Y(\mod_ro_256.fabric[0] ),
    .A(\mod_ro_256.fabric[256] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[0].inv  (.Y(\mod_ro_256.fabric[1] ),
    .A(\mod_ro_256.fabric[0] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[100].inv  (.Y(\mod_ro_256.fabric[101] ),
    .A(\mod_ro_256.fabric[100] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[101].inv  (.Y(\mod_ro_256.fabric[102] ),
    .A(\mod_ro_256.fabric[101] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[102].inv  (.Y(\mod_ro_256.fabric[103] ),
    .A(\mod_ro_256.fabric[102] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[103].inv  (.Y(\mod_ro_256.fabric[104] ),
    .A(\mod_ro_256.fabric[103] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[104].inv  (.Y(\mod_ro_256.fabric[105] ),
    .A(\mod_ro_256.fabric[104] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[105].inv  (.Y(\mod_ro_256.fabric[106] ),
    .A(\mod_ro_256.fabric[105] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[106].inv  (.Y(\mod_ro_256.fabric[107] ),
    .A(\mod_ro_256.fabric[106] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[107].inv  (.Y(\mod_ro_256.fabric[108] ),
    .A(\mod_ro_256.fabric[107] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[108].inv  (.Y(\mod_ro_256.fabric[109] ),
    .A(\mod_ro_256.fabric[108] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[109].inv  (.Y(\mod_ro_256.fabric[110] ),
    .A(\mod_ro_256.fabric[109] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[10].inv  (.Y(\mod_ro_256.fabric[11] ),
    .A(\mod_ro_256.fabric[10] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[110].inv  (.Y(\mod_ro_256.fabric[111] ),
    .A(\mod_ro_256.fabric[110] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[111].inv  (.Y(\mod_ro_256.fabric[112] ),
    .A(\mod_ro_256.fabric[111] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[112].inv  (.Y(\mod_ro_256.fabric[113] ),
    .A(\mod_ro_256.fabric[112] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[113].inv  (.Y(\mod_ro_256.fabric[114] ),
    .A(\mod_ro_256.fabric[113] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[114].inv  (.Y(\mod_ro_256.fabric[115] ),
    .A(\mod_ro_256.fabric[114] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[115].inv  (.Y(\mod_ro_256.fabric[116] ),
    .A(\mod_ro_256.fabric[115] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[116].inv  (.Y(\mod_ro_256.fabric[117] ),
    .A(\mod_ro_256.fabric[116] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[117].inv  (.Y(\mod_ro_256.fabric[118] ),
    .A(\mod_ro_256.fabric[117] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[118].inv  (.Y(\mod_ro_256.fabric[119] ),
    .A(\mod_ro_256.fabric[118] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[119].inv  (.Y(\mod_ro_256.fabric[120] ),
    .A(\mod_ro_256.fabric[119] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[11].inv  (.Y(\mod_ro_256.fabric[12] ),
    .A(\mod_ro_256.fabric[11] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[120].inv  (.Y(\mod_ro_256.fabric[121] ),
    .A(\mod_ro_256.fabric[120] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[121].inv  (.Y(\mod_ro_256.fabric[122] ),
    .A(\mod_ro_256.fabric[121] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[122].inv  (.Y(\mod_ro_256.fabric[123] ),
    .A(\mod_ro_256.fabric[122] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[123].inv  (.Y(\mod_ro_256.fabric[124] ),
    .A(\mod_ro_256.fabric[123] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[124].inv  (.Y(\mod_ro_256.fabric[125] ),
    .A(\mod_ro_256.fabric[124] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[125].inv  (.Y(\mod_ro_256.fabric[126] ),
    .A(\mod_ro_256.fabric[125] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[126].inv  (.Y(\mod_ro_256.fabric[127] ),
    .A(\mod_ro_256.fabric[126] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[127].inv  (.Y(\mod_ro_256.fabric[128] ),
    .A(\mod_ro_256.fabric[127] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[128].inv  (.Y(\mod_ro_256.fabric[129] ),
    .A(\mod_ro_256.fabric[128] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[129].inv  (.Y(\mod_ro_256.fabric[130] ),
    .A(\mod_ro_256.fabric[129] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[12].inv  (.Y(\mod_ro_256.fabric[13] ),
    .A(\mod_ro_256.fabric[12] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[130].inv  (.Y(\mod_ro_256.fabric[131] ),
    .A(\mod_ro_256.fabric[130] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[131].inv  (.Y(\mod_ro_256.fabric[132] ),
    .A(\mod_ro_256.fabric[131] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[132].inv  (.Y(\mod_ro_256.fabric[133] ),
    .A(\mod_ro_256.fabric[132] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[133].inv  (.Y(\mod_ro_256.fabric[134] ),
    .A(\mod_ro_256.fabric[133] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[134].inv  (.Y(\mod_ro_256.fabric[135] ),
    .A(\mod_ro_256.fabric[134] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[135].inv  (.Y(\mod_ro_256.fabric[136] ),
    .A(\mod_ro_256.fabric[135] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[136].inv  (.Y(\mod_ro_256.fabric[137] ),
    .A(\mod_ro_256.fabric[136] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[137].inv  (.Y(\mod_ro_256.fabric[138] ),
    .A(\mod_ro_256.fabric[137] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[138].inv  (.Y(\mod_ro_256.fabric[139] ),
    .A(\mod_ro_256.fabric[138] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[139].inv  (.Y(\mod_ro_256.fabric[140] ),
    .A(\mod_ro_256.fabric[139] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[13].inv  (.Y(\mod_ro_256.fabric[14] ),
    .A(\mod_ro_256.fabric[13] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[140].inv  (.Y(\mod_ro_256.fabric[141] ),
    .A(\mod_ro_256.fabric[140] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[141].inv  (.Y(\mod_ro_256.fabric[142] ),
    .A(\mod_ro_256.fabric[141] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[142].inv  (.Y(\mod_ro_256.fabric[143] ),
    .A(\mod_ro_256.fabric[142] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[143].inv  (.Y(\mod_ro_256.fabric[144] ),
    .A(\mod_ro_256.fabric[143] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[144].inv  (.Y(\mod_ro_256.fabric[145] ),
    .A(\mod_ro_256.fabric[144] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[145].inv  (.Y(\mod_ro_256.fabric[146] ),
    .A(\mod_ro_256.fabric[145] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[146].inv  (.Y(\mod_ro_256.fabric[147] ),
    .A(\mod_ro_256.fabric[146] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[147].inv  (.Y(\mod_ro_256.fabric[148] ),
    .A(\mod_ro_256.fabric[147] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[148].inv  (.Y(\mod_ro_256.fabric[149] ),
    .A(\mod_ro_256.fabric[148] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[149].inv  (.Y(\mod_ro_256.fabric[150] ),
    .A(\mod_ro_256.fabric[149] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[14].inv  (.Y(\mod_ro_256.fabric[15] ),
    .A(\mod_ro_256.fabric[14] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[150].inv  (.Y(\mod_ro_256.fabric[151] ),
    .A(\mod_ro_256.fabric[150] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[151].inv  (.Y(\mod_ro_256.fabric[152] ),
    .A(\mod_ro_256.fabric[151] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[152].inv  (.Y(\mod_ro_256.fabric[153] ),
    .A(\mod_ro_256.fabric[152] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[153].inv  (.Y(\mod_ro_256.fabric[154] ),
    .A(\mod_ro_256.fabric[153] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[154].inv  (.Y(\mod_ro_256.fabric[155] ),
    .A(\mod_ro_256.fabric[154] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[155].inv  (.Y(\mod_ro_256.fabric[156] ),
    .A(\mod_ro_256.fabric[155] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[156].inv  (.Y(\mod_ro_256.fabric[157] ),
    .A(\mod_ro_256.fabric[156] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[157].inv  (.Y(\mod_ro_256.fabric[158] ),
    .A(\mod_ro_256.fabric[157] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[158].inv  (.Y(\mod_ro_256.fabric[159] ),
    .A(\mod_ro_256.fabric[158] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[159].inv  (.Y(\mod_ro_256.fabric[160] ),
    .A(\mod_ro_256.fabric[159] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[15].inv  (.Y(\mod_ro_256.fabric[16] ),
    .A(\mod_ro_256.fabric[15] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[160].inv  (.Y(\mod_ro_256.fabric[161] ),
    .A(\mod_ro_256.fabric[160] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[161].inv  (.Y(\mod_ro_256.fabric[162] ),
    .A(\mod_ro_256.fabric[161] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[162].inv  (.Y(\mod_ro_256.fabric[163] ),
    .A(\mod_ro_256.fabric[162] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[163].inv  (.Y(\mod_ro_256.fabric[164] ),
    .A(\mod_ro_256.fabric[163] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[164].inv  (.Y(\mod_ro_256.fabric[165] ),
    .A(\mod_ro_256.fabric[164] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[165].inv  (.Y(\mod_ro_256.fabric[166] ),
    .A(\mod_ro_256.fabric[165] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[166].inv  (.Y(\mod_ro_256.fabric[167] ),
    .A(\mod_ro_256.fabric[166] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[167].inv  (.Y(\mod_ro_256.fabric[168] ),
    .A(\mod_ro_256.fabric[167] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[168].inv  (.Y(\mod_ro_256.fabric[169] ),
    .A(\mod_ro_256.fabric[168] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[169].inv  (.Y(\mod_ro_256.fabric[170] ),
    .A(\mod_ro_256.fabric[169] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[16].inv  (.Y(\mod_ro_256.fabric[17] ),
    .A(\mod_ro_256.fabric[16] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[170].inv  (.Y(\mod_ro_256.fabric[171] ),
    .A(\mod_ro_256.fabric[170] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[171].inv  (.Y(\mod_ro_256.fabric[172] ),
    .A(\mod_ro_256.fabric[171] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[172].inv  (.Y(\mod_ro_256.fabric[173] ),
    .A(\mod_ro_256.fabric[172] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[173].inv  (.Y(\mod_ro_256.fabric[174] ),
    .A(\mod_ro_256.fabric[173] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[174].inv  (.Y(\mod_ro_256.fabric[175] ),
    .A(\mod_ro_256.fabric[174] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[175].inv  (.Y(\mod_ro_256.fabric[176] ),
    .A(\mod_ro_256.fabric[175] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[176].inv  (.Y(\mod_ro_256.fabric[177] ),
    .A(\mod_ro_256.fabric[176] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[177].inv  (.Y(\mod_ro_256.fabric[178] ),
    .A(\mod_ro_256.fabric[177] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[178].inv  (.Y(\mod_ro_256.fabric[179] ),
    .A(\mod_ro_256.fabric[178] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[179].inv  (.Y(\mod_ro_256.fabric[180] ),
    .A(\mod_ro_256.fabric[179] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[17].inv  (.Y(\mod_ro_256.fabric[18] ),
    .A(\mod_ro_256.fabric[17] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[180].inv  (.Y(\mod_ro_256.fabric[181] ),
    .A(\mod_ro_256.fabric[180] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[181].inv  (.Y(\mod_ro_256.fabric[182] ),
    .A(\mod_ro_256.fabric[181] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[182].inv  (.Y(\mod_ro_256.fabric[183] ),
    .A(\mod_ro_256.fabric[182] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[183].inv  (.Y(\mod_ro_256.fabric[184] ),
    .A(\mod_ro_256.fabric[183] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[184].inv  (.Y(\mod_ro_256.fabric[185] ),
    .A(\mod_ro_256.fabric[184] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[185].inv  (.Y(\mod_ro_256.fabric[186] ),
    .A(\mod_ro_256.fabric[185] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[186].inv  (.Y(\mod_ro_256.fabric[187] ),
    .A(\mod_ro_256.fabric[186] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[187].inv  (.Y(\mod_ro_256.fabric[188] ),
    .A(\mod_ro_256.fabric[187] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[188].inv  (.Y(\mod_ro_256.fabric[189] ),
    .A(\mod_ro_256.fabric[188] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[189].inv  (.Y(\mod_ro_256.fabric[190] ),
    .A(\mod_ro_256.fabric[189] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[18].inv  (.Y(\mod_ro_256.fabric[19] ),
    .A(\mod_ro_256.fabric[18] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[190].inv  (.Y(\mod_ro_256.fabric[191] ),
    .A(\mod_ro_256.fabric[190] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[191].inv  (.Y(\mod_ro_256.fabric[192] ),
    .A(\mod_ro_256.fabric[191] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[192].inv  (.Y(\mod_ro_256.fabric[193] ),
    .A(\mod_ro_256.fabric[192] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[193].inv  (.Y(\mod_ro_256.fabric[194] ),
    .A(\mod_ro_256.fabric[193] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[194].inv  (.Y(\mod_ro_256.fabric[195] ),
    .A(\mod_ro_256.fabric[194] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[195].inv  (.Y(\mod_ro_256.fabric[196] ),
    .A(\mod_ro_256.fabric[195] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[196].inv  (.Y(\mod_ro_256.fabric[197] ),
    .A(\mod_ro_256.fabric[196] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[197].inv  (.Y(\mod_ro_256.fabric[198] ),
    .A(\mod_ro_256.fabric[197] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[198].inv  (.Y(\mod_ro_256.fabric[199] ),
    .A(\mod_ro_256.fabric[198] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[199].inv  (.Y(\mod_ro_256.fabric[200] ),
    .A(\mod_ro_256.fabric[199] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[19].inv  (.Y(\mod_ro_256.fabric[20] ),
    .A(\mod_ro_256.fabric[19] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[1].inv  (.Y(\mod_ro_256.fabric[2] ),
    .A(\mod_ro_256.fabric[1] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[200].inv  (.Y(\mod_ro_256.fabric[201] ),
    .A(\mod_ro_256.fabric[200] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[201].inv  (.Y(\mod_ro_256.fabric[202] ),
    .A(\mod_ro_256.fabric[201] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[202].inv  (.Y(\mod_ro_256.fabric[203] ),
    .A(\mod_ro_256.fabric[202] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[203].inv  (.Y(\mod_ro_256.fabric[204] ),
    .A(\mod_ro_256.fabric[203] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[204].inv  (.Y(\mod_ro_256.fabric[205] ),
    .A(\mod_ro_256.fabric[204] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[205].inv  (.Y(\mod_ro_256.fabric[206] ),
    .A(\mod_ro_256.fabric[205] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[206].inv  (.Y(\mod_ro_256.fabric[207] ),
    .A(\mod_ro_256.fabric[206] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[207].inv  (.Y(\mod_ro_256.fabric[208] ),
    .A(\mod_ro_256.fabric[207] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[208].inv  (.Y(\mod_ro_256.fabric[209] ),
    .A(\mod_ro_256.fabric[208] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[209].inv  (.Y(\mod_ro_256.fabric[210] ),
    .A(\mod_ro_256.fabric[209] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[20].inv  (.Y(\mod_ro_256.fabric[21] ),
    .A(\mod_ro_256.fabric[20] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[210].inv  (.Y(\mod_ro_256.fabric[211] ),
    .A(\mod_ro_256.fabric[210] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[211].inv  (.Y(\mod_ro_256.fabric[212] ),
    .A(\mod_ro_256.fabric[211] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[212].inv  (.Y(\mod_ro_256.fabric[213] ),
    .A(\mod_ro_256.fabric[212] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[213].inv  (.Y(\mod_ro_256.fabric[214] ),
    .A(\mod_ro_256.fabric[213] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[214].inv  (.Y(\mod_ro_256.fabric[215] ),
    .A(\mod_ro_256.fabric[214] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[215].inv  (.Y(\mod_ro_256.fabric[216] ),
    .A(\mod_ro_256.fabric[215] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[216].inv  (.Y(\mod_ro_256.fabric[217] ),
    .A(\mod_ro_256.fabric[216] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[217].inv  (.Y(\mod_ro_256.fabric[218] ),
    .A(\mod_ro_256.fabric[217] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[218].inv  (.Y(\mod_ro_256.fabric[219] ),
    .A(\mod_ro_256.fabric[218] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[219].inv  (.Y(\mod_ro_256.fabric[220] ),
    .A(\mod_ro_256.fabric[219] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[21].inv  (.Y(\mod_ro_256.fabric[22] ),
    .A(\mod_ro_256.fabric[21] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[220].inv  (.Y(\mod_ro_256.fabric[221] ),
    .A(\mod_ro_256.fabric[220] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[221].inv  (.Y(\mod_ro_256.fabric[222] ),
    .A(\mod_ro_256.fabric[221] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[222].inv  (.Y(\mod_ro_256.fabric[223] ),
    .A(\mod_ro_256.fabric[222] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[223].inv  (.Y(\mod_ro_256.fabric[224] ),
    .A(\mod_ro_256.fabric[223] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[224].inv  (.Y(\mod_ro_256.fabric[225] ),
    .A(\mod_ro_256.fabric[224] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[225].inv  (.Y(\mod_ro_256.fabric[226] ),
    .A(\mod_ro_256.fabric[225] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[226].inv  (.Y(\mod_ro_256.fabric[227] ),
    .A(\mod_ro_256.fabric[226] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[227].inv  (.Y(\mod_ro_256.fabric[228] ),
    .A(\mod_ro_256.fabric[227] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[228].inv  (.Y(\mod_ro_256.fabric[229] ),
    .A(\mod_ro_256.fabric[228] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[229].inv  (.Y(\mod_ro_256.fabric[230] ),
    .A(\mod_ro_256.fabric[229] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[22].inv  (.Y(\mod_ro_256.fabric[23] ),
    .A(\mod_ro_256.fabric[22] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[230].inv  (.Y(\mod_ro_256.fabric[231] ),
    .A(\mod_ro_256.fabric[230] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[231].inv  (.Y(\mod_ro_256.fabric[232] ),
    .A(\mod_ro_256.fabric[231] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[232].inv  (.Y(\mod_ro_256.fabric[233] ),
    .A(\mod_ro_256.fabric[232] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[233].inv  (.Y(\mod_ro_256.fabric[234] ),
    .A(\mod_ro_256.fabric[233] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[234].inv  (.Y(\mod_ro_256.fabric[235] ),
    .A(\mod_ro_256.fabric[234] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[235].inv  (.Y(\mod_ro_256.fabric[236] ),
    .A(\mod_ro_256.fabric[235] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[236].inv  (.Y(\mod_ro_256.fabric[237] ),
    .A(\mod_ro_256.fabric[236] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[237].inv  (.Y(\mod_ro_256.fabric[238] ),
    .A(\mod_ro_256.fabric[237] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[238].inv  (.Y(\mod_ro_256.fabric[239] ),
    .A(\mod_ro_256.fabric[238] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[239].inv  (.Y(\mod_ro_256.fabric[240] ),
    .A(\mod_ro_256.fabric[239] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[23].inv  (.Y(\mod_ro_256.fabric[24] ),
    .A(\mod_ro_256.fabric[23] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[240].inv  (.Y(\mod_ro_256.fabric[241] ),
    .A(\mod_ro_256.fabric[240] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[241].inv  (.Y(\mod_ro_256.fabric[242] ),
    .A(\mod_ro_256.fabric[241] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[242].inv  (.Y(\mod_ro_256.fabric[243] ),
    .A(\mod_ro_256.fabric[242] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[243].inv  (.Y(\mod_ro_256.fabric[244] ),
    .A(\mod_ro_256.fabric[243] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[244].inv  (.Y(\mod_ro_256.fabric[245] ),
    .A(\mod_ro_256.fabric[244] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[245].inv  (.Y(\mod_ro_256.fabric[246] ),
    .A(\mod_ro_256.fabric[245] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[246].inv  (.Y(\mod_ro_256.fabric[247] ),
    .A(\mod_ro_256.fabric[246] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[247].inv  (.Y(\mod_ro_256.fabric[248] ),
    .A(\mod_ro_256.fabric[247] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[248].inv  (.Y(\mod_ro_256.fabric[249] ),
    .A(\mod_ro_256.fabric[248] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[249].inv  (.Y(\mod_ro_256.fabric[250] ),
    .A(\mod_ro_256.fabric[249] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[24].inv  (.Y(\mod_ro_256.fabric[25] ),
    .A(\mod_ro_256.fabric[24] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[250].inv  (.Y(\mod_ro_256.fabric[251] ),
    .A(\mod_ro_256.fabric[250] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[251].inv  (.Y(\mod_ro_256.fabric[252] ),
    .A(\mod_ro_256.fabric[251] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[252].inv  (.Y(\mod_ro_256.fabric[253] ),
    .A(\mod_ro_256.fabric[252] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[253].inv  (.Y(\mod_ro_256.fabric[254] ),
    .A(\mod_ro_256.fabric[253] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[254].inv  (.Y(\mod_ro_256.fabric[255] ),
    .A(\mod_ro_256.fabric[254] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[255].inv  (.Y(\mod_ro_256.fabric[256] ),
    .A(\mod_ro_256.fabric[255] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[25].inv  (.Y(\mod_ro_256.fabric[26] ),
    .A(\mod_ro_256.fabric[25] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[26].inv  (.Y(\mod_ro_256.fabric[27] ),
    .A(\mod_ro_256.fabric[26] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[27].inv  (.Y(\mod_ro_256.fabric[28] ),
    .A(\mod_ro_256.fabric[27] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[28].inv  (.Y(\mod_ro_256.fabric[29] ),
    .A(\mod_ro_256.fabric[28] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[29].inv  (.Y(\mod_ro_256.fabric[30] ),
    .A(\mod_ro_256.fabric[29] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[2].inv  (.Y(\mod_ro_256.fabric[3] ),
    .A(\mod_ro_256.fabric[2] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[30].inv  (.Y(\mod_ro_256.fabric[31] ),
    .A(\mod_ro_256.fabric[30] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[31].inv  (.Y(\mod_ro_256.fabric[32] ),
    .A(\mod_ro_256.fabric[31] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[32].inv  (.Y(\mod_ro_256.fabric[33] ),
    .A(\mod_ro_256.fabric[32] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[33].inv  (.Y(\mod_ro_256.fabric[34] ),
    .A(\mod_ro_256.fabric[33] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[34].inv  (.Y(\mod_ro_256.fabric[35] ),
    .A(\mod_ro_256.fabric[34] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[35].inv  (.Y(\mod_ro_256.fabric[36] ),
    .A(\mod_ro_256.fabric[35] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[36].inv  (.Y(\mod_ro_256.fabric[37] ),
    .A(\mod_ro_256.fabric[36] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[37].inv  (.Y(\mod_ro_256.fabric[38] ),
    .A(\mod_ro_256.fabric[37] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[38].inv  (.Y(\mod_ro_256.fabric[39] ),
    .A(\mod_ro_256.fabric[38] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[39].inv  (.Y(\mod_ro_256.fabric[40] ),
    .A(\mod_ro_256.fabric[39] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[3].inv  (.Y(\mod_ro_256.fabric[4] ),
    .A(\mod_ro_256.fabric[3] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[40].inv  (.Y(\mod_ro_256.fabric[41] ),
    .A(\mod_ro_256.fabric[40] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[41].inv  (.Y(\mod_ro_256.fabric[42] ),
    .A(\mod_ro_256.fabric[41] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[42].inv  (.Y(\mod_ro_256.fabric[43] ),
    .A(\mod_ro_256.fabric[42] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[43].inv  (.Y(\mod_ro_256.fabric[44] ),
    .A(\mod_ro_256.fabric[43] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[44].inv  (.Y(\mod_ro_256.fabric[45] ),
    .A(\mod_ro_256.fabric[44] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[45].inv  (.Y(\mod_ro_256.fabric[46] ),
    .A(\mod_ro_256.fabric[45] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[46].inv  (.Y(\mod_ro_256.fabric[47] ),
    .A(\mod_ro_256.fabric[46] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[47].inv  (.Y(\mod_ro_256.fabric[48] ),
    .A(\mod_ro_256.fabric[47] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[48].inv  (.Y(\mod_ro_256.fabric[49] ),
    .A(\mod_ro_256.fabric[48] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[49].inv  (.Y(\mod_ro_256.fabric[50] ),
    .A(\mod_ro_256.fabric[49] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[4].inv  (.Y(\mod_ro_256.fabric[5] ),
    .A(\mod_ro_256.fabric[4] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[50].inv  (.Y(\mod_ro_256.fabric[51] ),
    .A(\mod_ro_256.fabric[50] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[51].inv  (.Y(\mod_ro_256.fabric[52] ),
    .A(\mod_ro_256.fabric[51] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[52].inv  (.Y(\mod_ro_256.fabric[53] ),
    .A(\mod_ro_256.fabric[52] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[53].inv  (.Y(\mod_ro_256.fabric[54] ),
    .A(\mod_ro_256.fabric[53] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[54].inv  (.Y(\mod_ro_256.fabric[55] ),
    .A(\mod_ro_256.fabric[54] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[55].inv  (.Y(\mod_ro_256.fabric[56] ),
    .A(\mod_ro_256.fabric[55] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[56].inv  (.Y(\mod_ro_256.fabric[57] ),
    .A(\mod_ro_256.fabric[56] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[57].inv  (.Y(\mod_ro_256.fabric[58] ),
    .A(\mod_ro_256.fabric[57] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[58].inv  (.Y(\mod_ro_256.fabric[59] ),
    .A(\mod_ro_256.fabric[58] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[59].inv  (.Y(\mod_ro_256.fabric[60] ),
    .A(\mod_ro_256.fabric[59] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[5].inv  (.Y(\mod_ro_256.fabric[6] ),
    .A(\mod_ro_256.fabric[5] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[60].inv  (.Y(\mod_ro_256.fabric[61] ),
    .A(\mod_ro_256.fabric[60] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[61].inv  (.Y(\mod_ro_256.fabric[62] ),
    .A(\mod_ro_256.fabric[61] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[62].inv  (.Y(\mod_ro_256.fabric[63] ),
    .A(\mod_ro_256.fabric[62] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[63].inv  (.Y(\mod_ro_256.fabric[64] ),
    .A(\mod_ro_256.fabric[63] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[64].inv  (.Y(\mod_ro_256.fabric[65] ),
    .A(\mod_ro_256.fabric[64] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[65].inv  (.Y(\mod_ro_256.fabric[66] ),
    .A(\mod_ro_256.fabric[65] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[66].inv  (.Y(\mod_ro_256.fabric[67] ),
    .A(\mod_ro_256.fabric[66] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[67].inv  (.Y(\mod_ro_256.fabric[68] ),
    .A(\mod_ro_256.fabric[67] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[68].inv  (.Y(\mod_ro_256.fabric[69] ),
    .A(\mod_ro_256.fabric[68] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[69].inv  (.Y(\mod_ro_256.fabric[70] ),
    .A(\mod_ro_256.fabric[69] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[6].inv  (.Y(\mod_ro_256.fabric[7] ),
    .A(\mod_ro_256.fabric[6] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[70].inv  (.Y(\mod_ro_256.fabric[71] ),
    .A(\mod_ro_256.fabric[70] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[71].inv  (.Y(\mod_ro_256.fabric[72] ),
    .A(\mod_ro_256.fabric[71] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[72].inv  (.Y(\mod_ro_256.fabric[73] ),
    .A(\mod_ro_256.fabric[72] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[73].inv  (.Y(\mod_ro_256.fabric[74] ),
    .A(\mod_ro_256.fabric[73] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[74].inv  (.Y(\mod_ro_256.fabric[75] ),
    .A(\mod_ro_256.fabric[74] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[75].inv  (.Y(\mod_ro_256.fabric[76] ),
    .A(\mod_ro_256.fabric[75] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[76].inv  (.Y(\mod_ro_256.fabric[77] ),
    .A(\mod_ro_256.fabric[76] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[77].inv  (.Y(\mod_ro_256.fabric[78] ),
    .A(\mod_ro_256.fabric[77] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[78].inv  (.Y(\mod_ro_256.fabric[79] ),
    .A(\mod_ro_256.fabric[78] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[79].inv  (.Y(\mod_ro_256.fabric[80] ),
    .A(\mod_ro_256.fabric[79] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[7].inv  (.Y(\mod_ro_256.fabric[8] ),
    .A(\mod_ro_256.fabric[7] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[80].inv  (.Y(\mod_ro_256.fabric[81] ),
    .A(\mod_ro_256.fabric[80] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[81].inv  (.Y(\mod_ro_256.fabric[82] ),
    .A(\mod_ro_256.fabric[81] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[82].inv  (.Y(\mod_ro_256.fabric[83] ),
    .A(\mod_ro_256.fabric[82] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[83].inv  (.Y(\mod_ro_256.fabric[84] ),
    .A(\mod_ro_256.fabric[83] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[84].inv  (.Y(\mod_ro_256.fabric[85] ),
    .A(\mod_ro_256.fabric[84] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[85].inv  (.Y(\mod_ro_256.fabric[86] ),
    .A(\mod_ro_256.fabric[85] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[86].inv  (.Y(\mod_ro_256.fabric[87] ),
    .A(\mod_ro_256.fabric[86] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[87].inv  (.Y(\mod_ro_256.fabric[88] ),
    .A(\mod_ro_256.fabric[87] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[88].inv  (.Y(\mod_ro_256.fabric[89] ),
    .A(\mod_ro_256.fabric[88] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[89].inv  (.Y(\mod_ro_256.fabric[90] ),
    .A(\mod_ro_256.fabric[89] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[8].inv  (.Y(\mod_ro_256.fabric[9] ),
    .A(\mod_ro_256.fabric[8] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[90].inv  (.Y(\mod_ro_256.fabric[91] ),
    .A(\mod_ro_256.fabric[90] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[91].inv  (.Y(\mod_ro_256.fabric[92] ),
    .A(\mod_ro_256.fabric[91] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[92].inv  (.Y(\mod_ro_256.fabric[93] ),
    .A(\mod_ro_256.fabric[92] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[93].inv  (.Y(\mod_ro_256.fabric[94] ),
    .A(\mod_ro_256.fabric[93] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[94].inv  (.Y(\mod_ro_256.fabric[95] ),
    .A(\mod_ro_256.fabric[94] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[95].inv  (.Y(\mod_ro_256.fabric[96] ),
    .A(\mod_ro_256.fabric[95] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[96].inv  (.Y(\mod_ro_256.fabric[97] ),
    .A(\mod_ro_256.fabric[96] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[97].inv  (.Y(\mod_ro_256.fabric[98] ),
    .A(\mod_ro_256.fabric[97] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[98].inv  (.Y(\mod_ro_256.fabric[99] ),
    .A(\mod_ro_256.fabric[98] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[99].inv  (.Y(\mod_ro_256.fabric[100] ),
    .A(\mod_ro_256.fabric[99] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[9].inv  (.Y(\mod_ro_256.fabric[10] ),
    .A(\mod_ro_256.fabric[9] ));
 sg13g2_inv_1 \mod_ro_256_drive4.feedback  (.Y(\mod_ro_256_drive4.fabric[0] ),
    .A(\mod_ro_256_drive4.fabric[256] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[0].inv  (.Y(\mod_ro_256_drive4.fabric[1] ),
    .A(\mod_ro_256_drive4.fabric[0] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[100].inv  (.Y(\mod_ro_256_drive4.fabric[101] ),
    .A(\mod_ro_256_drive4.fabric[100] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[101].inv  (.Y(\mod_ro_256_drive4.fabric[102] ),
    .A(\mod_ro_256_drive4.fabric[101] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[102].inv  (.Y(\mod_ro_256_drive4.fabric[103] ),
    .A(\mod_ro_256_drive4.fabric[102] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[103].inv  (.Y(\mod_ro_256_drive4.fabric[104] ),
    .A(\mod_ro_256_drive4.fabric[103] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[104].inv  (.Y(\mod_ro_256_drive4.fabric[105] ),
    .A(\mod_ro_256_drive4.fabric[104] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[105].inv  (.Y(\mod_ro_256_drive4.fabric[106] ),
    .A(\mod_ro_256_drive4.fabric[105] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[106].inv  (.Y(\mod_ro_256_drive4.fabric[107] ),
    .A(\mod_ro_256_drive4.fabric[106] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[107].inv  (.Y(\mod_ro_256_drive4.fabric[108] ),
    .A(\mod_ro_256_drive4.fabric[107] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[108].inv  (.Y(\mod_ro_256_drive4.fabric[109] ),
    .A(\mod_ro_256_drive4.fabric[108] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[109].inv  (.Y(\mod_ro_256_drive4.fabric[110] ),
    .A(\mod_ro_256_drive4.fabric[109] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[10].inv  (.Y(\mod_ro_256_drive4.fabric[11] ),
    .A(\mod_ro_256_drive4.fabric[10] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[110].inv  (.Y(\mod_ro_256_drive4.fabric[111] ),
    .A(\mod_ro_256_drive4.fabric[110] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[111].inv  (.Y(\mod_ro_256_drive4.fabric[112] ),
    .A(\mod_ro_256_drive4.fabric[111] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[112].inv  (.Y(\mod_ro_256_drive4.fabric[113] ),
    .A(\mod_ro_256_drive4.fabric[112] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[113].inv  (.Y(\mod_ro_256_drive4.fabric[114] ),
    .A(\mod_ro_256_drive4.fabric[113] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[114].inv  (.Y(\mod_ro_256_drive4.fabric[115] ),
    .A(\mod_ro_256_drive4.fabric[114] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[115].inv  (.Y(\mod_ro_256_drive4.fabric[116] ),
    .A(\mod_ro_256_drive4.fabric[115] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[116].inv  (.Y(\mod_ro_256_drive4.fabric[117] ),
    .A(\mod_ro_256_drive4.fabric[116] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[117].inv  (.Y(\mod_ro_256_drive4.fabric[118] ),
    .A(\mod_ro_256_drive4.fabric[117] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[118].inv  (.Y(\mod_ro_256_drive4.fabric[119] ),
    .A(\mod_ro_256_drive4.fabric[118] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[119].inv  (.Y(\mod_ro_256_drive4.fabric[120] ),
    .A(\mod_ro_256_drive4.fabric[119] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[11].inv  (.Y(\mod_ro_256_drive4.fabric[12] ),
    .A(\mod_ro_256_drive4.fabric[11] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[120].inv  (.Y(\mod_ro_256_drive4.fabric[121] ),
    .A(\mod_ro_256_drive4.fabric[120] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[121].inv  (.Y(\mod_ro_256_drive4.fabric[122] ),
    .A(\mod_ro_256_drive4.fabric[121] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[122].inv  (.Y(\mod_ro_256_drive4.fabric[123] ),
    .A(\mod_ro_256_drive4.fabric[122] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[123].inv  (.Y(\mod_ro_256_drive4.fabric[124] ),
    .A(\mod_ro_256_drive4.fabric[123] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[124].inv  (.Y(\mod_ro_256_drive4.fabric[125] ),
    .A(\mod_ro_256_drive4.fabric[124] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[125].inv  (.Y(\mod_ro_256_drive4.fabric[126] ),
    .A(\mod_ro_256_drive4.fabric[125] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[126].inv  (.Y(\mod_ro_256_drive4.fabric[127] ),
    .A(\mod_ro_256_drive4.fabric[126] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[127].inv  (.Y(\mod_ro_256_drive4.fabric[128] ),
    .A(\mod_ro_256_drive4.fabric[127] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[128].inv  (.Y(\mod_ro_256_drive4.fabric[129] ),
    .A(\mod_ro_256_drive4.fabric[128] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[129].inv  (.Y(\mod_ro_256_drive4.fabric[130] ),
    .A(\mod_ro_256_drive4.fabric[129] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[12].inv  (.Y(\mod_ro_256_drive4.fabric[13] ),
    .A(\mod_ro_256_drive4.fabric[12] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[130].inv  (.Y(\mod_ro_256_drive4.fabric[131] ),
    .A(\mod_ro_256_drive4.fabric[130] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[131].inv  (.Y(\mod_ro_256_drive4.fabric[132] ),
    .A(\mod_ro_256_drive4.fabric[131] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[132].inv  (.Y(\mod_ro_256_drive4.fabric[133] ),
    .A(\mod_ro_256_drive4.fabric[132] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[133].inv  (.Y(\mod_ro_256_drive4.fabric[134] ),
    .A(\mod_ro_256_drive4.fabric[133] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[134].inv  (.Y(\mod_ro_256_drive4.fabric[135] ),
    .A(\mod_ro_256_drive4.fabric[134] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[135].inv  (.Y(\mod_ro_256_drive4.fabric[136] ),
    .A(\mod_ro_256_drive4.fabric[135] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[136].inv  (.Y(\mod_ro_256_drive4.fabric[137] ),
    .A(\mod_ro_256_drive4.fabric[136] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[137].inv  (.Y(\mod_ro_256_drive4.fabric[138] ),
    .A(\mod_ro_256_drive4.fabric[137] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[138].inv  (.Y(\mod_ro_256_drive4.fabric[139] ),
    .A(\mod_ro_256_drive4.fabric[138] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[139].inv  (.Y(\mod_ro_256_drive4.fabric[140] ),
    .A(\mod_ro_256_drive4.fabric[139] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[13].inv  (.Y(\mod_ro_256_drive4.fabric[14] ),
    .A(\mod_ro_256_drive4.fabric[13] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[140].inv  (.Y(\mod_ro_256_drive4.fabric[141] ),
    .A(\mod_ro_256_drive4.fabric[140] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[141].inv  (.Y(\mod_ro_256_drive4.fabric[142] ),
    .A(\mod_ro_256_drive4.fabric[141] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[142].inv  (.Y(\mod_ro_256_drive4.fabric[143] ),
    .A(\mod_ro_256_drive4.fabric[142] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[143].inv  (.Y(\mod_ro_256_drive4.fabric[144] ),
    .A(\mod_ro_256_drive4.fabric[143] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[144].inv  (.Y(\mod_ro_256_drive4.fabric[145] ),
    .A(\mod_ro_256_drive4.fabric[144] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[145].inv  (.Y(\mod_ro_256_drive4.fabric[146] ),
    .A(\mod_ro_256_drive4.fabric[145] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[146].inv  (.Y(\mod_ro_256_drive4.fabric[147] ),
    .A(\mod_ro_256_drive4.fabric[146] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[147].inv  (.Y(\mod_ro_256_drive4.fabric[148] ),
    .A(\mod_ro_256_drive4.fabric[147] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[148].inv  (.Y(\mod_ro_256_drive4.fabric[149] ),
    .A(\mod_ro_256_drive4.fabric[148] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[149].inv  (.Y(\mod_ro_256_drive4.fabric[150] ),
    .A(\mod_ro_256_drive4.fabric[149] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[14].inv  (.Y(\mod_ro_256_drive4.fabric[15] ),
    .A(\mod_ro_256_drive4.fabric[14] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[150].inv  (.Y(\mod_ro_256_drive4.fabric[151] ),
    .A(\mod_ro_256_drive4.fabric[150] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[151].inv  (.Y(\mod_ro_256_drive4.fabric[152] ),
    .A(\mod_ro_256_drive4.fabric[151] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[152].inv  (.Y(\mod_ro_256_drive4.fabric[153] ),
    .A(\mod_ro_256_drive4.fabric[152] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[153].inv  (.Y(\mod_ro_256_drive4.fabric[154] ),
    .A(\mod_ro_256_drive4.fabric[153] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[154].inv  (.Y(\mod_ro_256_drive4.fabric[155] ),
    .A(\mod_ro_256_drive4.fabric[154] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[155].inv  (.Y(\mod_ro_256_drive4.fabric[156] ),
    .A(\mod_ro_256_drive4.fabric[155] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[156].inv  (.Y(\mod_ro_256_drive4.fabric[157] ),
    .A(\mod_ro_256_drive4.fabric[156] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[157].inv  (.Y(\mod_ro_256_drive4.fabric[158] ),
    .A(\mod_ro_256_drive4.fabric[157] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[158].inv  (.Y(\mod_ro_256_drive4.fabric[159] ),
    .A(\mod_ro_256_drive4.fabric[158] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[159].inv  (.Y(\mod_ro_256_drive4.fabric[160] ),
    .A(\mod_ro_256_drive4.fabric[159] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[15].inv  (.Y(\mod_ro_256_drive4.fabric[16] ),
    .A(\mod_ro_256_drive4.fabric[15] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[160].inv  (.Y(\mod_ro_256_drive4.fabric[161] ),
    .A(\mod_ro_256_drive4.fabric[160] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[161].inv  (.Y(\mod_ro_256_drive4.fabric[162] ),
    .A(\mod_ro_256_drive4.fabric[161] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[162].inv  (.Y(\mod_ro_256_drive4.fabric[163] ),
    .A(\mod_ro_256_drive4.fabric[162] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[163].inv  (.Y(\mod_ro_256_drive4.fabric[164] ),
    .A(\mod_ro_256_drive4.fabric[163] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[164].inv  (.Y(\mod_ro_256_drive4.fabric[165] ),
    .A(\mod_ro_256_drive4.fabric[164] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[165].inv  (.Y(\mod_ro_256_drive4.fabric[166] ),
    .A(\mod_ro_256_drive4.fabric[165] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[166].inv  (.Y(\mod_ro_256_drive4.fabric[167] ),
    .A(\mod_ro_256_drive4.fabric[166] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[167].inv  (.Y(\mod_ro_256_drive4.fabric[168] ),
    .A(\mod_ro_256_drive4.fabric[167] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[168].inv  (.Y(\mod_ro_256_drive4.fabric[169] ),
    .A(\mod_ro_256_drive4.fabric[168] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[169].inv  (.Y(\mod_ro_256_drive4.fabric[170] ),
    .A(\mod_ro_256_drive4.fabric[169] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[16].inv  (.Y(\mod_ro_256_drive4.fabric[17] ),
    .A(\mod_ro_256_drive4.fabric[16] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[170].inv  (.Y(\mod_ro_256_drive4.fabric[171] ),
    .A(\mod_ro_256_drive4.fabric[170] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[171].inv  (.Y(\mod_ro_256_drive4.fabric[172] ),
    .A(\mod_ro_256_drive4.fabric[171] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[172].inv  (.Y(\mod_ro_256_drive4.fabric[173] ),
    .A(\mod_ro_256_drive4.fabric[172] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[173].inv  (.Y(\mod_ro_256_drive4.fabric[174] ),
    .A(\mod_ro_256_drive4.fabric[173] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[174].inv  (.Y(\mod_ro_256_drive4.fabric[175] ),
    .A(\mod_ro_256_drive4.fabric[174] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[175].inv  (.Y(\mod_ro_256_drive4.fabric[176] ),
    .A(\mod_ro_256_drive4.fabric[175] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[176].inv  (.Y(\mod_ro_256_drive4.fabric[177] ),
    .A(\mod_ro_256_drive4.fabric[176] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[177].inv  (.Y(\mod_ro_256_drive4.fabric[178] ),
    .A(\mod_ro_256_drive4.fabric[177] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[178].inv  (.Y(\mod_ro_256_drive4.fabric[179] ),
    .A(\mod_ro_256_drive4.fabric[178] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[179].inv  (.Y(\mod_ro_256_drive4.fabric[180] ),
    .A(\mod_ro_256_drive4.fabric[179] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[17].inv  (.Y(\mod_ro_256_drive4.fabric[18] ),
    .A(\mod_ro_256_drive4.fabric[17] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[180].inv  (.Y(\mod_ro_256_drive4.fabric[181] ),
    .A(\mod_ro_256_drive4.fabric[180] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[181].inv  (.Y(\mod_ro_256_drive4.fabric[182] ),
    .A(\mod_ro_256_drive4.fabric[181] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[182].inv  (.Y(\mod_ro_256_drive4.fabric[183] ),
    .A(\mod_ro_256_drive4.fabric[182] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[183].inv  (.Y(\mod_ro_256_drive4.fabric[184] ),
    .A(\mod_ro_256_drive4.fabric[183] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[184].inv  (.Y(\mod_ro_256_drive4.fabric[185] ),
    .A(\mod_ro_256_drive4.fabric[184] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[185].inv  (.Y(\mod_ro_256_drive4.fabric[186] ),
    .A(\mod_ro_256_drive4.fabric[185] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[186].inv  (.Y(\mod_ro_256_drive4.fabric[187] ),
    .A(\mod_ro_256_drive4.fabric[186] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[187].inv  (.Y(\mod_ro_256_drive4.fabric[188] ),
    .A(\mod_ro_256_drive4.fabric[187] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[188].inv  (.Y(\mod_ro_256_drive4.fabric[189] ),
    .A(\mod_ro_256_drive4.fabric[188] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[189].inv  (.Y(\mod_ro_256_drive4.fabric[190] ),
    .A(\mod_ro_256_drive4.fabric[189] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[18].inv  (.Y(\mod_ro_256_drive4.fabric[19] ),
    .A(\mod_ro_256_drive4.fabric[18] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[190].inv  (.Y(\mod_ro_256_drive4.fabric[191] ),
    .A(\mod_ro_256_drive4.fabric[190] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[191].inv  (.Y(\mod_ro_256_drive4.fabric[192] ),
    .A(\mod_ro_256_drive4.fabric[191] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[192].inv  (.Y(\mod_ro_256_drive4.fabric[193] ),
    .A(\mod_ro_256_drive4.fabric[192] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[193].inv  (.Y(\mod_ro_256_drive4.fabric[194] ),
    .A(\mod_ro_256_drive4.fabric[193] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[194].inv  (.Y(\mod_ro_256_drive4.fabric[195] ),
    .A(\mod_ro_256_drive4.fabric[194] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[195].inv  (.Y(\mod_ro_256_drive4.fabric[196] ),
    .A(\mod_ro_256_drive4.fabric[195] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[196].inv  (.Y(\mod_ro_256_drive4.fabric[197] ),
    .A(\mod_ro_256_drive4.fabric[196] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[197].inv  (.Y(\mod_ro_256_drive4.fabric[198] ),
    .A(\mod_ro_256_drive4.fabric[197] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[198].inv  (.Y(\mod_ro_256_drive4.fabric[199] ),
    .A(\mod_ro_256_drive4.fabric[198] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[199].inv  (.Y(\mod_ro_256_drive4.fabric[200] ),
    .A(\mod_ro_256_drive4.fabric[199] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[19].inv  (.Y(\mod_ro_256_drive4.fabric[20] ),
    .A(\mod_ro_256_drive4.fabric[19] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[1].inv  (.Y(\mod_ro_256_drive4.fabric[2] ),
    .A(\mod_ro_256_drive4.fabric[1] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[200].inv  (.Y(\mod_ro_256_drive4.fabric[201] ),
    .A(\mod_ro_256_drive4.fabric[200] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[201].inv  (.Y(\mod_ro_256_drive4.fabric[202] ),
    .A(\mod_ro_256_drive4.fabric[201] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[202].inv  (.Y(\mod_ro_256_drive4.fabric[203] ),
    .A(\mod_ro_256_drive4.fabric[202] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[203].inv  (.Y(\mod_ro_256_drive4.fabric[204] ),
    .A(\mod_ro_256_drive4.fabric[203] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[204].inv  (.Y(\mod_ro_256_drive4.fabric[205] ),
    .A(\mod_ro_256_drive4.fabric[204] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[205].inv  (.Y(\mod_ro_256_drive4.fabric[206] ),
    .A(\mod_ro_256_drive4.fabric[205] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[206].inv  (.Y(\mod_ro_256_drive4.fabric[207] ),
    .A(\mod_ro_256_drive4.fabric[206] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[207].inv  (.Y(\mod_ro_256_drive4.fabric[208] ),
    .A(\mod_ro_256_drive4.fabric[207] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[208].inv  (.Y(\mod_ro_256_drive4.fabric[209] ),
    .A(\mod_ro_256_drive4.fabric[208] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[209].inv  (.Y(\mod_ro_256_drive4.fabric[210] ),
    .A(\mod_ro_256_drive4.fabric[209] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[20].inv  (.Y(\mod_ro_256_drive4.fabric[21] ),
    .A(\mod_ro_256_drive4.fabric[20] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[210].inv  (.Y(\mod_ro_256_drive4.fabric[211] ),
    .A(\mod_ro_256_drive4.fabric[210] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[211].inv  (.Y(\mod_ro_256_drive4.fabric[212] ),
    .A(\mod_ro_256_drive4.fabric[211] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[212].inv  (.Y(\mod_ro_256_drive4.fabric[213] ),
    .A(\mod_ro_256_drive4.fabric[212] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[213].inv  (.Y(\mod_ro_256_drive4.fabric[214] ),
    .A(\mod_ro_256_drive4.fabric[213] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[214].inv  (.Y(\mod_ro_256_drive4.fabric[215] ),
    .A(\mod_ro_256_drive4.fabric[214] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[215].inv  (.Y(\mod_ro_256_drive4.fabric[216] ),
    .A(\mod_ro_256_drive4.fabric[215] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[216].inv  (.Y(\mod_ro_256_drive4.fabric[217] ),
    .A(\mod_ro_256_drive4.fabric[216] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[217].inv  (.Y(\mod_ro_256_drive4.fabric[218] ),
    .A(\mod_ro_256_drive4.fabric[217] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[218].inv  (.Y(\mod_ro_256_drive4.fabric[219] ),
    .A(\mod_ro_256_drive4.fabric[218] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[219].inv  (.Y(\mod_ro_256_drive4.fabric[220] ),
    .A(\mod_ro_256_drive4.fabric[219] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[21].inv  (.Y(\mod_ro_256_drive4.fabric[22] ),
    .A(\mod_ro_256_drive4.fabric[21] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[220].inv  (.Y(\mod_ro_256_drive4.fabric[221] ),
    .A(\mod_ro_256_drive4.fabric[220] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[221].inv  (.Y(\mod_ro_256_drive4.fabric[222] ),
    .A(\mod_ro_256_drive4.fabric[221] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[222].inv  (.Y(\mod_ro_256_drive4.fabric[223] ),
    .A(\mod_ro_256_drive4.fabric[222] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[223].inv  (.Y(\mod_ro_256_drive4.fabric[224] ),
    .A(\mod_ro_256_drive4.fabric[223] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[224].inv  (.Y(\mod_ro_256_drive4.fabric[225] ),
    .A(\mod_ro_256_drive4.fabric[224] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[225].inv  (.Y(\mod_ro_256_drive4.fabric[226] ),
    .A(\mod_ro_256_drive4.fabric[225] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[226].inv  (.Y(\mod_ro_256_drive4.fabric[227] ),
    .A(\mod_ro_256_drive4.fabric[226] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[227].inv  (.Y(\mod_ro_256_drive4.fabric[228] ),
    .A(\mod_ro_256_drive4.fabric[227] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[228].inv  (.Y(\mod_ro_256_drive4.fabric[229] ),
    .A(\mod_ro_256_drive4.fabric[228] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[229].inv  (.Y(\mod_ro_256_drive4.fabric[230] ),
    .A(\mod_ro_256_drive4.fabric[229] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[22].inv  (.Y(\mod_ro_256_drive4.fabric[23] ),
    .A(\mod_ro_256_drive4.fabric[22] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[230].inv  (.Y(\mod_ro_256_drive4.fabric[231] ),
    .A(\mod_ro_256_drive4.fabric[230] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[231].inv  (.Y(\mod_ro_256_drive4.fabric[232] ),
    .A(\mod_ro_256_drive4.fabric[231] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[232].inv  (.Y(\mod_ro_256_drive4.fabric[233] ),
    .A(\mod_ro_256_drive4.fabric[232] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[233].inv  (.Y(\mod_ro_256_drive4.fabric[234] ),
    .A(\mod_ro_256_drive4.fabric[233] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[234].inv  (.Y(\mod_ro_256_drive4.fabric[235] ),
    .A(\mod_ro_256_drive4.fabric[234] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[235].inv  (.Y(\mod_ro_256_drive4.fabric[236] ),
    .A(\mod_ro_256_drive4.fabric[235] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[236].inv  (.Y(\mod_ro_256_drive4.fabric[237] ),
    .A(\mod_ro_256_drive4.fabric[236] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[237].inv  (.Y(\mod_ro_256_drive4.fabric[238] ),
    .A(\mod_ro_256_drive4.fabric[237] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[238].inv  (.Y(\mod_ro_256_drive4.fabric[239] ),
    .A(\mod_ro_256_drive4.fabric[238] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[239].inv  (.Y(\mod_ro_256_drive4.fabric[240] ),
    .A(\mod_ro_256_drive4.fabric[239] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[23].inv  (.Y(\mod_ro_256_drive4.fabric[24] ),
    .A(\mod_ro_256_drive4.fabric[23] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[240].inv  (.Y(\mod_ro_256_drive4.fabric[241] ),
    .A(\mod_ro_256_drive4.fabric[240] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[241].inv  (.Y(\mod_ro_256_drive4.fabric[242] ),
    .A(\mod_ro_256_drive4.fabric[241] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[242].inv  (.Y(\mod_ro_256_drive4.fabric[243] ),
    .A(\mod_ro_256_drive4.fabric[242] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[243].inv  (.Y(\mod_ro_256_drive4.fabric[244] ),
    .A(\mod_ro_256_drive4.fabric[243] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[244].inv  (.Y(\mod_ro_256_drive4.fabric[245] ),
    .A(\mod_ro_256_drive4.fabric[244] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[245].inv  (.Y(\mod_ro_256_drive4.fabric[246] ),
    .A(\mod_ro_256_drive4.fabric[245] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[246].inv  (.Y(\mod_ro_256_drive4.fabric[247] ),
    .A(\mod_ro_256_drive4.fabric[246] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[247].inv  (.Y(\mod_ro_256_drive4.fabric[248] ),
    .A(\mod_ro_256_drive4.fabric[247] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[248].inv  (.Y(\mod_ro_256_drive4.fabric[249] ),
    .A(\mod_ro_256_drive4.fabric[248] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[249].inv  (.Y(\mod_ro_256_drive4.fabric[250] ),
    .A(\mod_ro_256_drive4.fabric[249] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[24].inv  (.Y(\mod_ro_256_drive4.fabric[25] ),
    .A(\mod_ro_256_drive4.fabric[24] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[250].inv  (.Y(\mod_ro_256_drive4.fabric[251] ),
    .A(\mod_ro_256_drive4.fabric[250] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[251].inv  (.Y(\mod_ro_256_drive4.fabric[252] ),
    .A(\mod_ro_256_drive4.fabric[251] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[252].inv  (.Y(\mod_ro_256_drive4.fabric[253] ),
    .A(\mod_ro_256_drive4.fabric[252] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[253].inv  (.Y(\mod_ro_256_drive4.fabric[254] ),
    .A(\mod_ro_256_drive4.fabric[253] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[254].inv  (.Y(\mod_ro_256_drive4.fabric[255] ),
    .A(\mod_ro_256_drive4.fabric[254] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[255].inv  (.Y(\mod_ro_256_drive4.fabric[256] ),
    .A(\mod_ro_256_drive4.fabric[255] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[25].inv  (.Y(\mod_ro_256_drive4.fabric[26] ),
    .A(\mod_ro_256_drive4.fabric[25] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[26].inv  (.Y(\mod_ro_256_drive4.fabric[27] ),
    .A(\mod_ro_256_drive4.fabric[26] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[27].inv  (.Y(\mod_ro_256_drive4.fabric[28] ),
    .A(\mod_ro_256_drive4.fabric[27] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[28].inv  (.Y(\mod_ro_256_drive4.fabric[29] ),
    .A(\mod_ro_256_drive4.fabric[28] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[29].inv  (.Y(\mod_ro_256_drive4.fabric[30] ),
    .A(\mod_ro_256_drive4.fabric[29] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[2].inv  (.Y(\mod_ro_256_drive4.fabric[3] ),
    .A(\mod_ro_256_drive4.fabric[2] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[30].inv  (.Y(\mod_ro_256_drive4.fabric[31] ),
    .A(\mod_ro_256_drive4.fabric[30] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[31].inv  (.Y(\mod_ro_256_drive4.fabric[32] ),
    .A(\mod_ro_256_drive4.fabric[31] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[32].inv  (.Y(\mod_ro_256_drive4.fabric[33] ),
    .A(\mod_ro_256_drive4.fabric[32] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[33].inv  (.Y(\mod_ro_256_drive4.fabric[34] ),
    .A(\mod_ro_256_drive4.fabric[33] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[34].inv  (.Y(\mod_ro_256_drive4.fabric[35] ),
    .A(\mod_ro_256_drive4.fabric[34] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[35].inv  (.Y(\mod_ro_256_drive4.fabric[36] ),
    .A(\mod_ro_256_drive4.fabric[35] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[36].inv  (.Y(\mod_ro_256_drive4.fabric[37] ),
    .A(\mod_ro_256_drive4.fabric[36] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[37].inv  (.Y(\mod_ro_256_drive4.fabric[38] ),
    .A(\mod_ro_256_drive4.fabric[37] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[38].inv  (.Y(\mod_ro_256_drive4.fabric[39] ),
    .A(\mod_ro_256_drive4.fabric[38] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[39].inv  (.Y(\mod_ro_256_drive4.fabric[40] ),
    .A(\mod_ro_256_drive4.fabric[39] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[3].inv  (.Y(\mod_ro_256_drive4.fabric[4] ),
    .A(\mod_ro_256_drive4.fabric[3] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[40].inv  (.Y(\mod_ro_256_drive4.fabric[41] ),
    .A(\mod_ro_256_drive4.fabric[40] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[41].inv  (.Y(\mod_ro_256_drive4.fabric[42] ),
    .A(\mod_ro_256_drive4.fabric[41] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[42].inv  (.Y(\mod_ro_256_drive4.fabric[43] ),
    .A(\mod_ro_256_drive4.fabric[42] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[43].inv  (.Y(\mod_ro_256_drive4.fabric[44] ),
    .A(\mod_ro_256_drive4.fabric[43] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[44].inv  (.Y(\mod_ro_256_drive4.fabric[45] ),
    .A(\mod_ro_256_drive4.fabric[44] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[45].inv  (.Y(\mod_ro_256_drive4.fabric[46] ),
    .A(\mod_ro_256_drive4.fabric[45] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[46].inv  (.Y(\mod_ro_256_drive4.fabric[47] ),
    .A(\mod_ro_256_drive4.fabric[46] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[47].inv  (.Y(\mod_ro_256_drive4.fabric[48] ),
    .A(\mod_ro_256_drive4.fabric[47] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[48].inv  (.Y(\mod_ro_256_drive4.fabric[49] ),
    .A(\mod_ro_256_drive4.fabric[48] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[49].inv  (.Y(\mod_ro_256_drive4.fabric[50] ),
    .A(\mod_ro_256_drive4.fabric[49] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[4].inv  (.Y(\mod_ro_256_drive4.fabric[5] ),
    .A(\mod_ro_256_drive4.fabric[4] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[50].inv  (.Y(\mod_ro_256_drive4.fabric[51] ),
    .A(\mod_ro_256_drive4.fabric[50] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[51].inv  (.Y(\mod_ro_256_drive4.fabric[52] ),
    .A(\mod_ro_256_drive4.fabric[51] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[52].inv  (.Y(\mod_ro_256_drive4.fabric[53] ),
    .A(\mod_ro_256_drive4.fabric[52] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[53].inv  (.Y(\mod_ro_256_drive4.fabric[54] ),
    .A(\mod_ro_256_drive4.fabric[53] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[54].inv  (.Y(\mod_ro_256_drive4.fabric[55] ),
    .A(\mod_ro_256_drive4.fabric[54] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[55].inv  (.Y(\mod_ro_256_drive4.fabric[56] ),
    .A(\mod_ro_256_drive4.fabric[55] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[56].inv  (.Y(\mod_ro_256_drive4.fabric[57] ),
    .A(\mod_ro_256_drive4.fabric[56] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[57].inv  (.Y(\mod_ro_256_drive4.fabric[58] ),
    .A(\mod_ro_256_drive4.fabric[57] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[58].inv  (.Y(\mod_ro_256_drive4.fabric[59] ),
    .A(\mod_ro_256_drive4.fabric[58] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[59].inv  (.Y(\mod_ro_256_drive4.fabric[60] ),
    .A(\mod_ro_256_drive4.fabric[59] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[5].inv  (.Y(\mod_ro_256_drive4.fabric[6] ),
    .A(\mod_ro_256_drive4.fabric[5] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[60].inv  (.Y(\mod_ro_256_drive4.fabric[61] ),
    .A(\mod_ro_256_drive4.fabric[60] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[61].inv  (.Y(\mod_ro_256_drive4.fabric[62] ),
    .A(\mod_ro_256_drive4.fabric[61] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[62].inv  (.Y(\mod_ro_256_drive4.fabric[63] ),
    .A(\mod_ro_256_drive4.fabric[62] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[63].inv  (.Y(\mod_ro_256_drive4.fabric[64] ),
    .A(\mod_ro_256_drive4.fabric[63] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[64].inv  (.Y(\mod_ro_256_drive4.fabric[65] ),
    .A(\mod_ro_256_drive4.fabric[64] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[65].inv  (.Y(\mod_ro_256_drive4.fabric[66] ),
    .A(\mod_ro_256_drive4.fabric[65] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[66].inv  (.Y(\mod_ro_256_drive4.fabric[67] ),
    .A(\mod_ro_256_drive4.fabric[66] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[67].inv  (.Y(\mod_ro_256_drive4.fabric[68] ),
    .A(\mod_ro_256_drive4.fabric[67] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[68].inv  (.Y(\mod_ro_256_drive4.fabric[69] ),
    .A(\mod_ro_256_drive4.fabric[68] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[69].inv  (.Y(\mod_ro_256_drive4.fabric[70] ),
    .A(\mod_ro_256_drive4.fabric[69] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[6].inv  (.Y(\mod_ro_256_drive4.fabric[7] ),
    .A(\mod_ro_256_drive4.fabric[6] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[70].inv  (.Y(\mod_ro_256_drive4.fabric[71] ),
    .A(\mod_ro_256_drive4.fabric[70] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[71].inv  (.Y(\mod_ro_256_drive4.fabric[72] ),
    .A(\mod_ro_256_drive4.fabric[71] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[72].inv  (.Y(\mod_ro_256_drive4.fabric[73] ),
    .A(\mod_ro_256_drive4.fabric[72] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[73].inv  (.Y(\mod_ro_256_drive4.fabric[74] ),
    .A(\mod_ro_256_drive4.fabric[73] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[74].inv  (.Y(\mod_ro_256_drive4.fabric[75] ),
    .A(\mod_ro_256_drive4.fabric[74] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[75].inv  (.Y(\mod_ro_256_drive4.fabric[76] ),
    .A(\mod_ro_256_drive4.fabric[75] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[76].inv  (.Y(\mod_ro_256_drive4.fabric[77] ),
    .A(\mod_ro_256_drive4.fabric[76] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[77].inv  (.Y(\mod_ro_256_drive4.fabric[78] ),
    .A(\mod_ro_256_drive4.fabric[77] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[78].inv  (.Y(\mod_ro_256_drive4.fabric[79] ),
    .A(\mod_ro_256_drive4.fabric[78] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[79].inv  (.Y(\mod_ro_256_drive4.fabric[80] ),
    .A(\mod_ro_256_drive4.fabric[79] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[7].inv  (.Y(\mod_ro_256_drive4.fabric[8] ),
    .A(\mod_ro_256_drive4.fabric[7] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[80].inv  (.Y(\mod_ro_256_drive4.fabric[81] ),
    .A(\mod_ro_256_drive4.fabric[80] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[81].inv  (.Y(\mod_ro_256_drive4.fabric[82] ),
    .A(\mod_ro_256_drive4.fabric[81] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[82].inv  (.Y(\mod_ro_256_drive4.fabric[83] ),
    .A(\mod_ro_256_drive4.fabric[82] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[83].inv  (.Y(\mod_ro_256_drive4.fabric[84] ),
    .A(\mod_ro_256_drive4.fabric[83] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[84].inv  (.Y(\mod_ro_256_drive4.fabric[85] ),
    .A(\mod_ro_256_drive4.fabric[84] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[85].inv  (.Y(\mod_ro_256_drive4.fabric[86] ),
    .A(\mod_ro_256_drive4.fabric[85] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[86].inv  (.Y(\mod_ro_256_drive4.fabric[87] ),
    .A(\mod_ro_256_drive4.fabric[86] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[87].inv  (.Y(\mod_ro_256_drive4.fabric[88] ),
    .A(\mod_ro_256_drive4.fabric[87] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[88].inv  (.Y(\mod_ro_256_drive4.fabric[89] ),
    .A(\mod_ro_256_drive4.fabric[88] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[89].inv  (.Y(\mod_ro_256_drive4.fabric[90] ),
    .A(\mod_ro_256_drive4.fabric[89] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[8].inv  (.Y(\mod_ro_256_drive4.fabric[9] ),
    .A(\mod_ro_256_drive4.fabric[8] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[90].inv  (.Y(\mod_ro_256_drive4.fabric[91] ),
    .A(\mod_ro_256_drive4.fabric[90] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[91].inv  (.Y(\mod_ro_256_drive4.fabric[92] ),
    .A(\mod_ro_256_drive4.fabric[91] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[92].inv  (.Y(\mod_ro_256_drive4.fabric[93] ),
    .A(\mod_ro_256_drive4.fabric[92] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[93].inv  (.Y(\mod_ro_256_drive4.fabric[94] ),
    .A(\mod_ro_256_drive4.fabric[93] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[94].inv  (.Y(\mod_ro_256_drive4.fabric[95] ),
    .A(\mod_ro_256_drive4.fabric[94] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[95].inv  (.Y(\mod_ro_256_drive4.fabric[96] ),
    .A(\mod_ro_256_drive4.fabric[95] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[96].inv  (.Y(\mod_ro_256_drive4.fabric[97] ),
    .A(\mod_ro_256_drive4.fabric[96] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[97].inv  (.Y(\mod_ro_256_drive4.fabric[98] ),
    .A(\mod_ro_256_drive4.fabric[97] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[98].inv  (.Y(\mod_ro_256_drive4.fabric[99] ),
    .A(\mod_ro_256_drive4.fabric[98] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[99].inv  (.Y(\mod_ro_256_drive4.fabric[100] ),
    .A(\mod_ro_256_drive4.fabric[99] ));
 sg13g2_inv_1 \mod_ro_256_drive4.osc_gen[9].inv  (.Y(\mod_ro_256_drive4.fabric[10] ),
    .A(\mod_ro_256_drive4.fabric[9] ));
 sg13g2_inv_1 \mod_ro_31.feedback  (.Y(\mod_ro_31.fabric[0] ),
    .A(\mod_ro_31.fabric[31] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[0].inv  (.Y(\mod_ro_31.fabric[1] ),
    .A(\mod_ro_31.fabric[0] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[10].inv  (.Y(\mod_ro_31.fabric[11] ),
    .A(\mod_ro_31.fabric[10] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[11].inv  (.Y(\mod_ro_31.fabric[12] ),
    .A(\mod_ro_31.fabric[11] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[12].inv  (.Y(\mod_ro_31.fabric[13] ),
    .A(\mod_ro_31.fabric[12] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[13].inv  (.Y(\mod_ro_31.fabric[14] ),
    .A(\mod_ro_31.fabric[13] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[14].inv  (.Y(\mod_ro_31.fabric[15] ),
    .A(\mod_ro_31.fabric[14] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[15].inv  (.Y(\mod_ro_31.fabric[16] ),
    .A(\mod_ro_31.fabric[15] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[16].inv  (.Y(\mod_ro_31.fabric[17] ),
    .A(\mod_ro_31.fabric[16] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[17].inv  (.Y(\mod_ro_31.fabric[18] ),
    .A(\mod_ro_31.fabric[17] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[18].inv  (.Y(\mod_ro_31.fabric[19] ),
    .A(\mod_ro_31.fabric[18] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[19].inv  (.Y(\mod_ro_31.fabric[20] ),
    .A(\mod_ro_31.fabric[19] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[1].inv  (.Y(\mod_ro_31.fabric[2] ),
    .A(\mod_ro_31.fabric[1] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[20].inv  (.Y(\mod_ro_31.fabric[21] ),
    .A(\mod_ro_31.fabric[20] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[21].inv  (.Y(\mod_ro_31.fabric[22] ),
    .A(\mod_ro_31.fabric[21] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[22].inv  (.Y(\mod_ro_31.fabric[23] ),
    .A(\mod_ro_31.fabric[22] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[23].inv  (.Y(\mod_ro_31.fabric[24] ),
    .A(\mod_ro_31.fabric[23] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[24].inv  (.Y(\mod_ro_31.fabric[25] ),
    .A(\mod_ro_31.fabric[24] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[25].inv  (.Y(\mod_ro_31.fabric[26] ),
    .A(\mod_ro_31.fabric[25] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[26].inv  (.Y(\mod_ro_31.fabric[27] ),
    .A(\mod_ro_31.fabric[26] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[27].inv  (.Y(\mod_ro_31.fabric[28] ),
    .A(\mod_ro_31.fabric[27] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[28].inv  (.Y(\mod_ro_31.fabric[29] ),
    .A(\mod_ro_31.fabric[28] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[29].inv  (.Y(\mod_ro_31.fabric[30] ),
    .A(\mod_ro_31.fabric[29] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[2].inv  (.Y(\mod_ro_31.fabric[3] ),
    .A(\mod_ro_31.fabric[2] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[30].inv  (.Y(\mod_ro_31.fabric[31] ),
    .A(\mod_ro_31.fabric[30] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[3].inv  (.Y(\mod_ro_31.fabric[4] ),
    .A(\mod_ro_31.fabric[3] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[4].inv  (.Y(\mod_ro_31.fabric[5] ),
    .A(\mod_ro_31.fabric[4] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[5].inv  (.Y(\mod_ro_31.fabric[6] ),
    .A(\mod_ro_31.fabric[5] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[6].inv  (.Y(\mod_ro_31.fabric[7] ),
    .A(\mod_ro_31.fabric[6] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[7].inv  (.Y(\mod_ro_31.fabric[8] ),
    .A(\mod_ro_31.fabric[7] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[8].inv  (.Y(\mod_ro_31.fabric[9] ),
    .A(\mod_ro_31.fabric[8] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[9].inv  (.Y(\mod_ro_31.fabric[10] ),
    .A(\mod_ro_31.fabric[9] ));
 sg13g2_inv_2 \mod_ro_32_1.feedback  (.Y(\mod_ro_32_1.fabric[0] ),
    .A(\mod_ro_32_1.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[0].inv  (.Y(\mod_ro_32_1.fabric[1] ),
    .A(\mod_ro_32_1.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[10].inv  (.Y(\mod_ro_32_1.fabric[11] ),
    .A(\mod_ro_32_1.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[11].inv  (.Y(\mod_ro_32_1.fabric[12] ),
    .A(\mod_ro_32_1.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[12].inv  (.Y(\mod_ro_32_1.fabric[13] ),
    .A(\mod_ro_32_1.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[13].inv  (.Y(\mod_ro_32_1.fabric[14] ),
    .A(\mod_ro_32_1.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[14].inv  (.Y(\mod_ro_32_1.fabric[15] ),
    .A(\mod_ro_32_1.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[15].inv  (.Y(\mod_ro_32_1.fabric[16] ),
    .A(\mod_ro_32_1.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[16].inv  (.Y(\mod_ro_32_1.fabric[17] ),
    .A(\mod_ro_32_1.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[17].inv  (.Y(\mod_ro_32_1.fabric[18] ),
    .A(\mod_ro_32_1.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[18].inv  (.Y(\mod_ro_32_1.fabric[19] ),
    .A(\mod_ro_32_1.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[19].inv  (.Y(\mod_ro_32_1.fabric[20] ),
    .A(\mod_ro_32_1.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[1].inv  (.Y(\mod_ro_32_1.fabric[2] ),
    .A(\mod_ro_32_1.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[20].inv  (.Y(\mod_ro_32_1.fabric[21] ),
    .A(\mod_ro_32_1.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[21].inv  (.Y(\mod_ro_32_1.fabric[22] ),
    .A(\mod_ro_32_1.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[22].inv  (.Y(\mod_ro_32_1.fabric[23] ),
    .A(\mod_ro_32_1.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[23].inv  (.Y(\mod_ro_32_1.fabric[24] ),
    .A(\mod_ro_32_1.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[24].inv  (.Y(\mod_ro_32_1.fabric[25] ),
    .A(\mod_ro_32_1.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[25].inv  (.Y(\mod_ro_32_1.fabric[26] ),
    .A(\mod_ro_32_1.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[26].inv  (.Y(\mod_ro_32_1.fabric[27] ),
    .A(\mod_ro_32_1.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[27].inv  (.Y(\mod_ro_32_1.fabric[28] ),
    .A(\mod_ro_32_1.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[28].inv  (.Y(\mod_ro_32_1.fabric[29] ),
    .A(\mod_ro_32_1.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[29].inv  (.Y(\mod_ro_32_1.fabric[30] ),
    .A(\mod_ro_32_1.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[2].inv  (.Y(\mod_ro_32_1.fabric[3] ),
    .A(\mod_ro_32_1.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[30].inv  (.Y(\mod_ro_32_1.fabric[31] ),
    .A(\mod_ro_32_1.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[31].inv  (.Y(\mod_ro_32_1.fabric[32] ),
    .A(\mod_ro_32_1.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[3].inv  (.Y(\mod_ro_32_1.fabric[4] ),
    .A(\mod_ro_32_1.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[4].inv  (.Y(\mod_ro_32_1.fabric[5] ),
    .A(\mod_ro_32_1.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[5].inv  (.Y(\mod_ro_32_1.fabric[6] ),
    .A(\mod_ro_32_1.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[6].inv  (.Y(\mod_ro_32_1.fabric[7] ),
    .A(\mod_ro_32_1.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[7].inv  (.Y(\mod_ro_32_1.fabric[8] ),
    .A(\mod_ro_32_1.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[8].inv  (.Y(\mod_ro_32_1.fabric[9] ),
    .A(\mod_ro_32_1.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[9].inv  (.Y(\mod_ro_32_1.fabric[10] ),
    .A(\mod_ro_32_1.fabric[9] ));
 sg13g2_inv_2 \mod_ro_32_2.feedback  (.Y(\mod_ro_32_2.fabric[0] ),
    .A(\mod_ro_32_2.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[0].inv  (.Y(\mod_ro_32_2.fabric[1] ),
    .A(\mod_ro_32_2.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[10].inv  (.Y(\mod_ro_32_2.fabric[11] ),
    .A(\mod_ro_32_2.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[11].inv  (.Y(\mod_ro_32_2.fabric[12] ),
    .A(\mod_ro_32_2.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[12].inv  (.Y(\mod_ro_32_2.fabric[13] ),
    .A(\mod_ro_32_2.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[13].inv  (.Y(\mod_ro_32_2.fabric[14] ),
    .A(\mod_ro_32_2.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[14].inv  (.Y(\mod_ro_32_2.fabric[15] ),
    .A(\mod_ro_32_2.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[15].inv  (.Y(\mod_ro_32_2.fabric[16] ),
    .A(\mod_ro_32_2.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[16].inv  (.Y(\mod_ro_32_2.fabric[17] ),
    .A(\mod_ro_32_2.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[17].inv  (.Y(\mod_ro_32_2.fabric[18] ),
    .A(\mod_ro_32_2.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[18].inv  (.Y(\mod_ro_32_2.fabric[19] ),
    .A(\mod_ro_32_2.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[19].inv  (.Y(\mod_ro_32_2.fabric[20] ),
    .A(\mod_ro_32_2.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[1].inv  (.Y(\mod_ro_32_2.fabric[2] ),
    .A(\mod_ro_32_2.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[20].inv  (.Y(\mod_ro_32_2.fabric[21] ),
    .A(\mod_ro_32_2.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[21].inv  (.Y(\mod_ro_32_2.fabric[22] ),
    .A(\mod_ro_32_2.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[22].inv  (.Y(\mod_ro_32_2.fabric[23] ),
    .A(\mod_ro_32_2.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[23].inv  (.Y(\mod_ro_32_2.fabric[24] ),
    .A(\mod_ro_32_2.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[24].inv  (.Y(\mod_ro_32_2.fabric[25] ),
    .A(\mod_ro_32_2.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[25].inv  (.Y(\mod_ro_32_2.fabric[26] ),
    .A(\mod_ro_32_2.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[26].inv  (.Y(\mod_ro_32_2.fabric[27] ),
    .A(\mod_ro_32_2.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[27].inv  (.Y(\mod_ro_32_2.fabric[28] ),
    .A(\mod_ro_32_2.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[28].inv  (.Y(\mod_ro_32_2.fabric[29] ),
    .A(\mod_ro_32_2.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[29].inv  (.Y(\mod_ro_32_2.fabric[30] ),
    .A(\mod_ro_32_2.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[2].inv  (.Y(\mod_ro_32_2.fabric[3] ),
    .A(\mod_ro_32_2.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[30].inv  (.Y(\mod_ro_32_2.fabric[31] ),
    .A(\mod_ro_32_2.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[31].inv  (.Y(\mod_ro_32_2.fabric[32] ),
    .A(\mod_ro_32_2.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[3].inv  (.Y(\mod_ro_32_2.fabric[4] ),
    .A(\mod_ro_32_2.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[4].inv  (.Y(\mod_ro_32_2.fabric[5] ),
    .A(\mod_ro_32_2.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[5].inv  (.Y(\mod_ro_32_2.fabric[6] ),
    .A(\mod_ro_32_2.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[6].inv  (.Y(\mod_ro_32_2.fabric[7] ),
    .A(\mod_ro_32_2.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[7].inv  (.Y(\mod_ro_32_2.fabric[8] ),
    .A(\mod_ro_32_2.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[8].inv  (.Y(\mod_ro_32_2.fabric[9] ),
    .A(\mod_ro_32_2.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[9].inv  (.Y(\mod_ro_32_2.fabric[10] ),
    .A(\mod_ro_32_2.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_drive4.feedback  (.Y(\mod_ro_32_drive4.fabric[0] ),
    .A(\mod_ro_32_drive4.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[0].inv  (.Y(\mod_ro_32_drive4.fabric[1] ),
    .A(\mod_ro_32_drive4.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[10].inv  (.Y(\mod_ro_32_drive4.fabric[11] ),
    .A(\mod_ro_32_drive4.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[11].inv  (.Y(\mod_ro_32_drive4.fabric[12] ),
    .A(\mod_ro_32_drive4.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[12].inv  (.Y(\mod_ro_32_drive4.fabric[13] ),
    .A(\mod_ro_32_drive4.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[13].inv  (.Y(\mod_ro_32_drive4.fabric[14] ),
    .A(\mod_ro_32_drive4.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[14].inv  (.Y(\mod_ro_32_drive4.fabric[15] ),
    .A(\mod_ro_32_drive4.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[15].inv  (.Y(\mod_ro_32_drive4.fabric[16] ),
    .A(\mod_ro_32_drive4.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[16].inv  (.Y(\mod_ro_32_drive4.fabric[17] ),
    .A(\mod_ro_32_drive4.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[17].inv  (.Y(\mod_ro_32_drive4.fabric[18] ),
    .A(\mod_ro_32_drive4.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[18].inv  (.Y(\mod_ro_32_drive4.fabric[19] ),
    .A(\mod_ro_32_drive4.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[19].inv  (.Y(\mod_ro_32_drive4.fabric[20] ),
    .A(\mod_ro_32_drive4.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[1].inv  (.Y(\mod_ro_32_drive4.fabric[2] ),
    .A(\mod_ro_32_drive4.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[20].inv  (.Y(\mod_ro_32_drive4.fabric[21] ),
    .A(\mod_ro_32_drive4.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[21].inv  (.Y(\mod_ro_32_drive4.fabric[22] ),
    .A(\mod_ro_32_drive4.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[22].inv  (.Y(\mod_ro_32_drive4.fabric[23] ),
    .A(\mod_ro_32_drive4.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[23].inv  (.Y(\mod_ro_32_drive4.fabric[24] ),
    .A(\mod_ro_32_drive4.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[24].inv  (.Y(\mod_ro_32_drive4.fabric[25] ),
    .A(\mod_ro_32_drive4.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[25].inv  (.Y(\mod_ro_32_drive4.fabric[26] ),
    .A(\mod_ro_32_drive4.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[26].inv  (.Y(\mod_ro_32_drive4.fabric[27] ),
    .A(\mod_ro_32_drive4.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[27].inv  (.Y(\mod_ro_32_drive4.fabric[28] ),
    .A(\mod_ro_32_drive4.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[28].inv  (.Y(\mod_ro_32_drive4.fabric[29] ),
    .A(\mod_ro_32_drive4.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[29].inv  (.Y(\mod_ro_32_drive4.fabric[30] ),
    .A(\mod_ro_32_drive4.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[2].inv  (.Y(\mod_ro_32_drive4.fabric[3] ),
    .A(\mod_ro_32_drive4.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[30].inv  (.Y(\mod_ro_32_drive4.fabric[31] ),
    .A(\mod_ro_32_drive4.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[31].inv  (.Y(\mod_ro_32_drive4.fabric[32] ),
    .A(\mod_ro_32_drive4.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[3].inv  (.Y(\mod_ro_32_drive4.fabric[4] ),
    .A(\mod_ro_32_drive4.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[4].inv  (.Y(\mod_ro_32_drive4.fabric[5] ),
    .A(\mod_ro_32_drive4.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[5].inv  (.Y(\mod_ro_32_drive4.fabric[6] ),
    .A(\mod_ro_32_drive4.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[6].inv  (.Y(\mod_ro_32_drive4.fabric[7] ),
    .A(\mod_ro_32_drive4.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[7].inv  (.Y(\mod_ro_32_drive4.fabric[8] ),
    .A(\mod_ro_32_drive4.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[8].inv  (.Y(\mod_ro_32_drive4.fabric[9] ),
    .A(\mod_ro_32_drive4.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_drive4.osc_gen[9].inv  (.Y(\mod_ro_32_drive4.fabric[10] ),
    .A(\mod_ro_32_drive4.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_raw.feedback  (.Y(\mod_ro_32_raw.fabric[0] ),
    .A(\mod_ro_32_raw.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[0].inv  (.Y(\mod_ro_32_raw.fabric[1] ),
    .A(\mod_ro_32_raw.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[10].inv  (.Y(\mod_ro_32_raw.fabric[11] ),
    .A(\mod_ro_32_raw.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[11].inv  (.Y(\mod_ro_32_raw.fabric[12] ),
    .A(\mod_ro_32_raw.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[12].inv  (.Y(\mod_ro_32_raw.fabric[13] ),
    .A(\mod_ro_32_raw.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[13].inv  (.Y(\mod_ro_32_raw.fabric[14] ),
    .A(\mod_ro_32_raw.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[14].inv  (.Y(\mod_ro_32_raw.fabric[15] ),
    .A(\mod_ro_32_raw.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[15].inv  (.Y(\mod_ro_32_raw.fabric[16] ),
    .A(\mod_ro_32_raw.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[16].inv  (.Y(\mod_ro_32_raw.fabric[17] ),
    .A(\mod_ro_32_raw.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[17].inv  (.Y(\mod_ro_32_raw.fabric[18] ),
    .A(\mod_ro_32_raw.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[18].inv  (.Y(\mod_ro_32_raw.fabric[19] ),
    .A(\mod_ro_32_raw.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[19].inv  (.Y(\mod_ro_32_raw.fabric[20] ),
    .A(\mod_ro_32_raw.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[1].inv  (.Y(\mod_ro_32_raw.fabric[2] ),
    .A(\mod_ro_32_raw.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[20].inv  (.Y(\mod_ro_32_raw.fabric[21] ),
    .A(\mod_ro_32_raw.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[21].inv  (.Y(\mod_ro_32_raw.fabric[22] ),
    .A(\mod_ro_32_raw.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[22].inv  (.Y(\mod_ro_32_raw.fabric[23] ),
    .A(\mod_ro_32_raw.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[23].inv  (.Y(\mod_ro_32_raw.fabric[24] ),
    .A(\mod_ro_32_raw.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[24].inv  (.Y(\mod_ro_32_raw.fabric[25] ),
    .A(\mod_ro_32_raw.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[25].inv  (.Y(\mod_ro_32_raw.fabric[26] ),
    .A(\mod_ro_32_raw.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[26].inv  (.Y(\mod_ro_32_raw.fabric[27] ),
    .A(\mod_ro_32_raw.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[27].inv  (.Y(\mod_ro_32_raw.fabric[28] ),
    .A(\mod_ro_32_raw.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[28].inv  (.Y(\mod_ro_32_raw.fabric[29] ),
    .A(\mod_ro_32_raw.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[29].inv  (.Y(\mod_ro_32_raw.fabric[30] ),
    .A(\mod_ro_32_raw.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[2].inv  (.Y(\mod_ro_32_raw.fabric[3] ),
    .A(\mod_ro_32_raw.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[30].inv  (.Y(\mod_ro_32_raw.fabric[31] ),
    .A(\mod_ro_32_raw.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[31].inv  (.Y(\mod_ro_32_raw.fabric[32] ),
    .A(\mod_ro_32_raw.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[3].inv  (.Y(\mod_ro_32_raw.fabric[4] ),
    .A(\mod_ro_32_raw.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[4].inv  (.Y(\mod_ro_32_raw.fabric[5] ),
    .A(\mod_ro_32_raw.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[5].inv  (.Y(\mod_ro_32_raw.fabric[6] ),
    .A(\mod_ro_32_raw.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[6].inv  (.Y(\mod_ro_32_raw.fabric[7] ),
    .A(\mod_ro_32_raw.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[7].inv  (.Y(\mod_ro_32_raw.fabric[8] ),
    .A(\mod_ro_32_raw.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[8].inv  (.Y(\mod_ro_32_raw.fabric[9] ),
    .A(\mod_ro_32_raw.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[9].inv  (.Y(\mod_ro_32_raw.fabric[10] ),
    .A(\mod_ro_32_raw.fabric[9] ));
 sg13g2_inv_1 \mod_ro_64.feedback  (.Y(\mod_ro_64.fabric[0] ),
    .A(\mod_ro_64.fabric[64] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[0].inv  (.Y(\mod_ro_64.fabric[1] ),
    .A(\mod_ro_64.fabric[0] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[10].inv  (.Y(\mod_ro_64.fabric[11] ),
    .A(\mod_ro_64.fabric[10] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[11].inv  (.Y(\mod_ro_64.fabric[12] ),
    .A(\mod_ro_64.fabric[11] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[12].inv  (.Y(\mod_ro_64.fabric[13] ),
    .A(\mod_ro_64.fabric[12] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[13].inv  (.Y(\mod_ro_64.fabric[14] ),
    .A(\mod_ro_64.fabric[13] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[14].inv  (.Y(\mod_ro_64.fabric[15] ),
    .A(\mod_ro_64.fabric[14] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[15].inv  (.Y(\mod_ro_64.fabric[16] ),
    .A(\mod_ro_64.fabric[15] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[16].inv  (.Y(\mod_ro_64.fabric[17] ),
    .A(\mod_ro_64.fabric[16] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[17].inv  (.Y(\mod_ro_64.fabric[18] ),
    .A(\mod_ro_64.fabric[17] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[18].inv  (.Y(\mod_ro_64.fabric[19] ),
    .A(\mod_ro_64.fabric[18] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[19].inv  (.Y(\mod_ro_64.fabric[20] ),
    .A(\mod_ro_64.fabric[19] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[1].inv  (.Y(\mod_ro_64.fabric[2] ),
    .A(\mod_ro_64.fabric[1] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[20].inv  (.Y(\mod_ro_64.fabric[21] ),
    .A(\mod_ro_64.fabric[20] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[21].inv  (.Y(\mod_ro_64.fabric[22] ),
    .A(\mod_ro_64.fabric[21] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[22].inv  (.Y(\mod_ro_64.fabric[23] ),
    .A(\mod_ro_64.fabric[22] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[23].inv  (.Y(\mod_ro_64.fabric[24] ),
    .A(\mod_ro_64.fabric[23] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[24].inv  (.Y(\mod_ro_64.fabric[25] ),
    .A(\mod_ro_64.fabric[24] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[25].inv  (.Y(\mod_ro_64.fabric[26] ),
    .A(\mod_ro_64.fabric[25] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[26].inv  (.Y(\mod_ro_64.fabric[27] ),
    .A(\mod_ro_64.fabric[26] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[27].inv  (.Y(\mod_ro_64.fabric[28] ),
    .A(\mod_ro_64.fabric[27] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[28].inv  (.Y(\mod_ro_64.fabric[29] ),
    .A(\mod_ro_64.fabric[28] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[29].inv  (.Y(\mod_ro_64.fabric[30] ),
    .A(\mod_ro_64.fabric[29] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[2].inv  (.Y(\mod_ro_64.fabric[3] ),
    .A(\mod_ro_64.fabric[2] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[30].inv  (.Y(\mod_ro_64.fabric[31] ),
    .A(\mod_ro_64.fabric[30] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[31].inv  (.Y(\mod_ro_64.fabric[32] ),
    .A(\mod_ro_64.fabric[31] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[32].inv  (.Y(\mod_ro_64.fabric[33] ),
    .A(\mod_ro_64.fabric[32] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[33].inv  (.Y(\mod_ro_64.fabric[34] ),
    .A(\mod_ro_64.fabric[33] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[34].inv  (.Y(\mod_ro_64.fabric[35] ),
    .A(\mod_ro_64.fabric[34] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[35].inv  (.Y(\mod_ro_64.fabric[36] ),
    .A(\mod_ro_64.fabric[35] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[36].inv  (.Y(\mod_ro_64.fabric[37] ),
    .A(\mod_ro_64.fabric[36] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[37].inv  (.Y(\mod_ro_64.fabric[38] ),
    .A(\mod_ro_64.fabric[37] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[38].inv  (.Y(\mod_ro_64.fabric[39] ),
    .A(\mod_ro_64.fabric[38] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[39].inv  (.Y(\mod_ro_64.fabric[40] ),
    .A(\mod_ro_64.fabric[39] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[3].inv  (.Y(\mod_ro_64.fabric[4] ),
    .A(\mod_ro_64.fabric[3] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[40].inv  (.Y(\mod_ro_64.fabric[41] ),
    .A(\mod_ro_64.fabric[40] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[41].inv  (.Y(\mod_ro_64.fabric[42] ),
    .A(\mod_ro_64.fabric[41] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[42].inv  (.Y(\mod_ro_64.fabric[43] ),
    .A(\mod_ro_64.fabric[42] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[43].inv  (.Y(\mod_ro_64.fabric[44] ),
    .A(\mod_ro_64.fabric[43] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[44].inv  (.Y(\mod_ro_64.fabric[45] ),
    .A(\mod_ro_64.fabric[44] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[45].inv  (.Y(\mod_ro_64.fabric[46] ),
    .A(\mod_ro_64.fabric[45] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[46].inv  (.Y(\mod_ro_64.fabric[47] ),
    .A(\mod_ro_64.fabric[46] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[47].inv  (.Y(\mod_ro_64.fabric[48] ),
    .A(\mod_ro_64.fabric[47] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[48].inv  (.Y(\mod_ro_64.fabric[49] ),
    .A(\mod_ro_64.fabric[48] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[49].inv  (.Y(\mod_ro_64.fabric[50] ),
    .A(\mod_ro_64.fabric[49] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[4].inv  (.Y(\mod_ro_64.fabric[5] ),
    .A(\mod_ro_64.fabric[4] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[50].inv  (.Y(\mod_ro_64.fabric[51] ),
    .A(\mod_ro_64.fabric[50] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[51].inv  (.Y(\mod_ro_64.fabric[52] ),
    .A(\mod_ro_64.fabric[51] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[52].inv  (.Y(\mod_ro_64.fabric[53] ),
    .A(\mod_ro_64.fabric[52] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[53].inv  (.Y(\mod_ro_64.fabric[54] ),
    .A(\mod_ro_64.fabric[53] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[54].inv  (.Y(\mod_ro_64.fabric[55] ),
    .A(\mod_ro_64.fabric[54] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[55].inv  (.Y(\mod_ro_64.fabric[56] ),
    .A(\mod_ro_64.fabric[55] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[56].inv  (.Y(\mod_ro_64.fabric[57] ),
    .A(\mod_ro_64.fabric[56] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[57].inv  (.Y(\mod_ro_64.fabric[58] ),
    .A(\mod_ro_64.fabric[57] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[58].inv  (.Y(\mod_ro_64.fabric[59] ),
    .A(\mod_ro_64.fabric[58] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[59].inv  (.Y(\mod_ro_64.fabric[60] ),
    .A(\mod_ro_64.fabric[59] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[5].inv  (.Y(\mod_ro_64.fabric[6] ),
    .A(\mod_ro_64.fabric[5] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[60].inv  (.Y(\mod_ro_64.fabric[61] ),
    .A(\mod_ro_64.fabric[60] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[61].inv  (.Y(\mod_ro_64.fabric[62] ),
    .A(\mod_ro_64.fabric[61] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[62].inv  (.Y(\mod_ro_64.fabric[63] ),
    .A(\mod_ro_64.fabric[62] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[63].inv  (.Y(\mod_ro_64.fabric[64] ),
    .A(\mod_ro_64.fabric[63] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[6].inv  (.Y(\mod_ro_64.fabric[7] ),
    .A(\mod_ro_64.fabric[6] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[7].inv  (.Y(\mod_ro_64.fabric[8] ),
    .A(\mod_ro_64.fabric[7] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[8].inv  (.Y(\mod_ro_64.fabric[9] ),
    .A(\mod_ro_64.fabric[8] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[9].inv  (.Y(\mod_ro_64.fabric[10] ),
    .A(\mod_ro_64.fabric[9] ));
 sg13g2_inv_1 \mod_ro_prog.feedback  (.Y(\mod_ro_prog.fabric[0] ),
    .A(\mod_ro_prog.fabric[8] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[0].inv.inv  (.Y(\mod_ro_prog.osc_gen[0].inv.inverted ),
    .A(\mod_ro_prog.fabric[0] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[1].inv.inv  (.Y(\mod_ro_prog.osc_gen[1].inv.inverted ),
    .A(\mod_ro_prog.fabric[1] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[2].inv.inv  (.Y(\mod_ro_prog.osc_gen[2].inv.inverted ),
    .A(\mod_ro_prog.fabric[2] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[3].inv.inv  (.Y(\mod_ro_prog.osc_gen[3].inv.inverted ),
    .A(\mod_ro_prog.fabric[3] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[4].inv.inv  (.Y(\mod_ro_prog.osc_gen[4].inv.inverted ),
    .A(\mod_ro_prog.fabric[4] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[5].inv.inv  (.Y(\mod_ro_prog.osc_gen[5].inv.inverted ),
    .A(\mod_ro_prog.fabric[5] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[6].inv.inv  (.Y(\mod_ro_prog.osc_gen[6].inv.inverted ),
    .A(\mod_ro_prog.fabric[6] ));
 sg13g2_inv_1 \mod_ro_prog.osc_gen[7].inv.inv  (.Y(\mod_ro_prog.osc_gen[7].inv.inverted ),
    .A(\mod_ro_prog.fabric[7] ));
 sg13g2_buf_8 fanout35 (.A(_154_),
    .X(net35));
 sg13g2_buf_8 fanout36 (.A(_147_),
    .X(net36));
 sg13g2_buf_8 fanout37 (.A(_174_),
    .X(net37));
 sg13g2_buf_8 fanout38 (.A(_127_),
    .X(net38));
 sg13g2_buf_8 fanout39 (.A(net40),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(\dpll.n_count[5] ),
    .X(net41));
 sg13g2_buf_8 fanout42 (.A(net143),
    .X(net42));
 sg13g2_buf_8 fanout43 (.A(net46),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(net46),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45));
 sg13g2_buf_8 fanout46 (.A(ui_in[6]),
    .X(net46));
 sg13g2_buf_8 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_8 fanout48 (.A(rst_n),
    .X(net48));
 sg13g2_buf_8 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_8 fanout50 (.A(rst_n),
    .X(net50));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_tielo tt_um_mlyoung_wedgetail_7 (.L_LO(net7));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_decoder_mod.o_reg_wdata[3] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold2 (.A(\spi_decoder_mod.o_reg_wdata[6] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spi_decoder_mod.o_reg_wdata[4] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold4 (.A(\spi_decoder_mod.o_reg_wdata[5] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold5 (.A(\spi_decoder_mod.o_reg_wdata[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold6 (.A(\spi_decoder_mod.o_reg_wdata[2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold7 (.A(_014_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold8 (.A(_000_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold9 (.A(\spi_decoder_mod.shift_cnt[0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold10 (.A(\dpll.id_increment_done ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold11 (.A(_081_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold12 (.A(\dpll.id_decrement_done ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold13 (.A(_080_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold14 (.A(\spi_decoder_mod.start ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold15 (.A(\spi_decoder_mod.shift_cnt[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dpll.k_count_borrow ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold17 (.A(_090_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold18 (.A(\dpll.k_count_carry ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold19 (.A(_091_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold20 (.A(_015_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold21 (.A(_152_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold22 (.A(_055_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold23 (.A(\spi_decoder_mod.spi_state[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold24 (.A(_001_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold25 (.A(\dpll.n_count[1] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold26 (.A(_157_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold27 (.A(_072_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold28 (.A(\spi_decoder_mod.shift_cnt[2] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold29 (.A(\dpll.n_count[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold30 (.A(_071_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold31 (.A(_016_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold32 (.A(_153_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold33 (.A(_056_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dpll.n_count[2] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold35 (.A(_073_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dpll.id_decrement ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold37 (.A(_150_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold38 (.A(_079_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold39 (.A(\spi_regfile_mod.SYS_CTRL_RESET_q [0]),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold40 (.A(_148_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold41 (.A(_051_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold42 (.A(\spi_decoder_mod.write ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold43 (.A(\dpll.id_increment ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold44 (.A(_149_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold45 (.A(_078_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mod_ro_prog.osc_gen[0].inv.i_en ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold47 (.A(\dpll.k_count[7] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold48 (.A(_089_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold49 (.A(\dpll.k_count[6] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold50 (.A(_088_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold51 (.A(\reg_echo[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold52 (.A(_060_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold53 (.A(\spi_decoder_mod.spi_state[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold54 (.A(_002_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold55 (.A(\dpll.k_count[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold56 (.A(_177_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold57 (.A(_083_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold58 (.A(\dpll.k_count[4] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold59 (.A(_086_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold60 (.A(\reg_echo[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold61 (.A(_061_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold62 (.A(\reg_echo[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold63 (.A(_057_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold64 (.A(\reg_echo[3] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold65 (.A(_058_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold66 (.A(\reg_echo[4] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold67 (.A(_059_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold68 (.A(\dpll.k_count[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold69 (.A(_084_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold70 (.A(\spi_decoder_mod.o_reg_wdata[7] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold71 (.A(_069_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold72 (.A(\spi_decoder_mod.shift_out_reg[5] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold73 (.A(\dpll.id_out ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold74 (.A(\dpll.clk_fout ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold75 (.A(_077_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mod_ro_prog.osc_gen[3].inv.i_en ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold77 (.A(\spi_decoder_mod.shift_out_reg[4] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold78 (.A(\spi_decoder_mod.shift_out_reg[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold79 (.A(\spi_decoder_mod.shift_out_reg[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold80 (.A(\spi_decoder_mod.shift_out_reg[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold81 (.A(\dpll.k_count[3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold82 (.A(\spi_decoder_mod.shift_out_reg[6] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold83 (.A(\spi_decoder_mod.shift_out_reg[3] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mod_ro_prog.osc_gen[6].inv.i_en ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mod_ro_prog.osc_gen[4].inv.i_en ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mod_ro_prog.osc_gen[1].inv.i_en ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mod_ro_prog.osc_gen[5].inv.i_en ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold88 (.A(\dpll.n_count[4] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold89 (.A(_165_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold90 (.A(_076_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mod_ro_prog.osc_gen[2].inv.i_en ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold92 (.A(\dpll.clk8x_fout ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold93 (.A(\dpll.k_count[0] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold94 (.A(\dpll.k_count[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold95 (.A(_202_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold96 (.A(\spi_regfile_mod.addr [0]),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold97 (.A(_070_),
    .X(net167));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_4 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_240 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_fill_2 FILLER_0_359 ();
 sg13g2_fill_1 FILLER_0_361 ();
 sg13g2_fill_1 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_4 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_193 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_fill_2 FILLER_1_230 ();
 sg13g2_decap_4 FILLER_1_244 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_decap_8 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_276 ();
 sg13g2_fill_2 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_285 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_318 ();
 sg13g2_fill_2 FILLER_1_325 ();
 sg13g2_fill_1 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_4 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_140 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_4 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_4 FILLER_2_207 ();
 sg13g2_fill_1 FILLER_2_211 ();
 sg13g2_decap_8 FILLER_2_218 ();
 sg13g2_decap_4 FILLER_2_225 ();
 sg13g2_decap_8 FILLER_2_241 ();
 sg13g2_decap_4 FILLER_2_248 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_fill_2 FILLER_2_280 ();
 sg13g2_fill_1 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_4 FILLER_2_296 ();
 sg13g2_fill_2 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_2_319 ();
 sg13g2_fill_2 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_fill_2 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_4 FILLER_2_354 ();
 sg13g2_fill_2 FILLER_2_358 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_decap_4 FILLER_2_373 ();
 sg13g2_fill_1 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_150 ();
 sg13g2_decap_8 FILLER_3_157 ();
 sg13g2_decap_8 FILLER_3_164 ();
 sg13g2_fill_2 FILLER_3_171 ();
 sg13g2_decap_4 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_4 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_4 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_fill_2 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_decap_4 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_decap_4 FILLER_4_241 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_314 ();
 sg13g2_decap_4 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_4 FILLER_4_352 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_4 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_169 ();
 sg13g2_fill_1 FILLER_5_176 ();
 sg13g2_decap_4 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_4 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_4 FILLER_5_371 ();
 sg13g2_fill_2 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_4 FILLER_6_147 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_4 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_192 ();
 sg13g2_decap_8 FILLER_6_199 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_4 FILLER_6_234 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_fill_1 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_4 FILLER_6_287 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_2 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_4 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_164 ();
 sg13g2_decap_8 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_fill_1 FILLER_7_190 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_253 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_262 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_fill_2 FILLER_7_295 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_decap_4 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_fill_2 FILLER_7_357 ();
 sg13g2_fill_1 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_fill_2 FILLER_7_392 ();
 sg13g2_fill_1 FILLER_7_394 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_4 FILLER_8_140 ();
 sg13g2_fill_2 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_232 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_4 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_297 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_4 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_332 ();
 sg13g2_decap_4 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_4 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_fill_2 FILLER_8_393 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_195 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_377 ();
 sg13g2_decap_4 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_394 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_decap_8 FILLER_10_148 ();
 sg13g2_decap_4 FILLER_10_155 ();
 sg13g2_fill_2 FILLER_10_159 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_4 FILLER_10_228 ();
 sg13g2_fill_1 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_4 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_fill_2 FILLER_10_360 ();
 sg13g2_fill_1 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_4 FILLER_10_385 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_8 FILLER_11_157 ();
 sg13g2_decap_8 FILLER_11_164 ();
 sg13g2_decap_8 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_216 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_237 ();
 sg13g2_fill_2 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_fill_1 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_fill_1 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_4 FILLER_12_342 ();
 sg13g2_fill_2 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_177 ();
 sg13g2_decap_8 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_4 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_4 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_fill_2 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_4 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_4 FILLER_14_347 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_fill_1 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_fill_2 FILLER_15_339 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_4 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_4 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_306 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_4 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_4 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_4 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_fill_2 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_4 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_fill_2 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_fill_2 FILLER_19_386 ();
 sg13g2_fill_1 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_4 FILLER_20_39 ();
 sg13g2_fill_2 FILLER_20_43 ();
 sg13g2_fill_2 FILLER_20_50 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_106 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_decap_8 FILLER_20_118 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_decap_8 FILLER_20_202 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_4 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_4 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_13 ();
 sg13g2_decap_4 FILLER_21_20 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_167 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_37 ();
 sg13g2_decap_8 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_decap_4 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_decap_4 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_66 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_decap_8 FILLER_23_136 ();
 sg13g2_decap_4 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_4 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_decap_4 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_392 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_30 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_decap_4 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_4 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_64 ();
 sg13g2_decap_8 FILLER_25_71 ();
 sg13g2_decap_4 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_163 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_4 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_fill_1 FILLER_26_45 ();
 sg13g2_decap_4 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_decap_4 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_4 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_391 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_68 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_141 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_decap_8 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_4 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_decap_4 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_4 FILLER_28_388 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_40 ();
 sg13g2_decap_4 FILLER_29_66 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_decap_4 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_decap_4 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_decap_4 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_4 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_decap_4 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_104 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_125 ();
 sg13g2_decap_4 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_decap_4 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_decap_4 FILLER_30_388 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_decap_4 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_4 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_4 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_4 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_4 FILLER_32_183 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_227 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_decap_4 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_decap_4 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_4 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_37 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_1 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_fill_2 FILLER_33_196 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_286 ();
 sg13g2_decap_4 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_4 FILLER_33_387 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_decap_4 FILLER_34_276 ();
 sg13g2_fill_2 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_4 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_25 ();
 sg13g2_decap_8 FILLER_35_68 ();
 sg13g2_decap_4 FILLER_35_75 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_158 ();
 sg13g2_fill_2 FILLER_35_162 ();
 sg13g2_decap_8 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_decap_4 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_385 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_113 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_122 ();
 sg13g2_decap_4 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_148 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_103 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_393 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_decap_4 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_392 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
 assign uo_out[1] = net23;
 assign uo_out[7] = net24;
endmodule
