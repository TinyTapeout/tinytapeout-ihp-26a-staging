module tt_um_herald (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire clknet_leaf_0_clk;
 wire \byte_counter[0] ;
 wire \byte_counter[1] ;
 wire \cmd_reg[0] ;
 wire \cmd_reg[1] ;
 wire \cmd_reg[2] ;
 wire \cmd_reg[3] ;
 wire \cmd_reg[4] ;
 wire \cmd_reg[5] ;
 wire \cmd_reg[6] ;
 wire \cmd_reg[7] ;
 wire \cordic_atan2_result[0] ;
 wire \cordic_atan2_result[10] ;
 wire \cordic_atan2_result[11] ;
 wire \cordic_atan2_result[12] ;
 wire \cordic_atan2_result[13] ;
 wire \cordic_atan2_result[14] ;
 wire \cordic_atan2_result[15] ;
 wire \cordic_atan2_result[1] ;
 wire \cordic_atan2_result[2] ;
 wire \cordic_atan2_result[3] ;
 wire \cordic_atan2_result[4] ;
 wire \cordic_atan2_result[5] ;
 wire \cordic_atan2_result[6] ;
 wire \cordic_atan2_result[7] ;
 wire \cordic_atan2_result[8] ;
 wire \cordic_atan2_result[9] ;
 wire cordic_busy;
 wire cordic_en_atan2;
 wire cordic_en_get_atan2;
 wire cordic_en_get_sin_cos;
 wire cordic_en_get_sqrt;
 wire cordic_en_sin_cos;
 wire cordic_en_sqrt;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[1] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[2] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[3] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[4] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[5] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[6] ;
 wire \cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[7] ;
 wire \cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[23] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[24] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[25] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[26] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[27] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[28] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[29] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[30] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[31] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ;
 wire \cordic_inst.cordic_state[0] ;
 wire \cordic_inst.cordic_state[23] ;
 wire \cordic_inst.cordic_state[24] ;
 wire \cordic_inst.cordic_state[25] ;
 wire \cordic_inst.cordic_state[26] ;
 wire \cordic_inst.cordic_state[27] ;
 wire \cordic_inst.cordic_state[28] ;
 wire \cordic_inst.cordic_state[29] ;
 wire \cordic_inst.cordic_state[30] ;
 wire \cordic_inst.cordic_state[31] ;
 wire \cordic_inst.cordic_state[32] ;
 wire \cordic_inst.cordic_state[33] ;
 wire \cordic_inst.cordic_state[34] ;
 wire \cordic_inst.cordic_state[35] ;
 wire \cordic_inst.cordic_state[36] ;
 wire \cordic_inst.cordic_state[37] ;
 wire \cordic_inst.cordic_state[38] ;
 wire \cordic_inst.cordic_state[39] ;
 wire \cordic_inst.cordic_state[3] ;
 wire \cordic_inst.cordic_state[40] ;
 wire \cordic_inst.cordic_state[41] ;
 wire \cordic_inst.cordic_state[42] ;
 wire \cordic_inst.cordic_state[43] ;
 wire \cordic_inst.cordic_state[44] ;
 wire \cordic_inst.cordic_state[45] ;
 wire \cordic_inst.cordic_state[46] ;
 wire \cordic_inst.cordic_state[47] ;
 wire \cordic_inst.cordic_state[48] ;
 wire \cordic_inst.cordic_state[49] ;
 wire \cordic_inst.cordic_state[4] ;
 wire \cordic_inst.cordic_state[50] ;
 wire \cordic_inst.cordic_state[51] ;
 wire \cordic_inst.cordic_state[52] ;
 wire \cordic_inst.cordic_state[53] ;
 wire \cordic_inst.cordic_state[54] ;
 wire \cordic_inst.cordic_state[5] ;
 wire \cordic_inst.cordic_state[6] ;
 wire \cordic_inst.current_op[0] ;
 wire \cordic_inst.current_op[1] ;
 wire \cordic_inst.current_op[2] ;
 wire \cordic_inst.operation_pending ;
 wire \cordic_inst.result_ready ;
 wire \exec_phase[1] ;
 wire \exec_phase[2] ;
 wire mac_en_clear;
 wire mac_en_get_mac;
 wire mac_en_get_multiply;
 wire mac_en_mac;
 wire mac_en_multiply;
 wire \mac_inst.RDY_get_mac ;
 wire \mac_inst.RDY_get_multiply ;
 wire \mac_inst.accumulator[0] ;
 wire \mac_inst.accumulator[10] ;
 wire \mac_inst.accumulator[11] ;
 wire \mac_inst.accumulator[12] ;
 wire \mac_inst.accumulator[13] ;
 wire \mac_inst.accumulator[14] ;
 wire \mac_inst.accumulator[15] ;
 wire \mac_inst.accumulator[1] ;
 wire \mac_inst.accumulator[2] ;
 wire \mac_inst.accumulator[3] ;
 wire \mac_inst.accumulator[4] ;
 wire \mac_inst.accumulator[5] ;
 wire \mac_inst.accumulator[6] ;
 wire \mac_inst.accumulator[7] ;
 wire \mac_inst.accumulator[8] ;
 wire \mac_inst.accumulator[9] ;
 wire \mac_inst.get_multiply[0] ;
 wire \mac_inst.get_multiply[10] ;
 wire \mac_inst.get_multiply[11] ;
 wire \mac_inst.get_multiply[12] ;
 wire \mac_inst.get_multiply[13] ;
 wire \mac_inst.get_multiply[14] ;
 wire \mac_inst.get_multiply[15] ;
 wire \mac_inst.get_multiply[1] ;
 wire \mac_inst.get_multiply[2] ;
 wire \mac_inst.get_multiply[3] ;
 wire \mac_inst.get_multiply[4] ;
 wire \mac_inst.get_multiply[5] ;
 wire \mac_inst.get_multiply[6] ;
 wire \mac_inst.get_multiply[7] ;
 wire \mac_inst.get_multiply[8] ;
 wire \mac_inst.get_multiply[9] ;
 wire rd_prev;
 wire \result_reg[0] ;
 wire \result_reg[10] ;
 wire \result_reg[11] ;
 wire \result_reg[12] ;
 wire \result_reg[13] ;
 wire \result_reg[14] ;
 wire \result_reg[15] ;
 wire \result_reg[16] ;
 wire \result_reg[17] ;
 wire \result_reg[18] ;
 wire \result_reg[19] ;
 wire \result_reg[1] ;
 wire \result_reg[20] ;
 wire \result_reg[21] ;
 wire \result_reg[22] ;
 wire \result_reg[23] ;
 wire \result_reg[24] ;
 wire \result_reg[25] ;
 wire \result_reg[26] ;
 wire \result_reg[27] ;
 wire \result_reg[28] ;
 wire \result_reg[29] ;
 wire \result_reg[2] ;
 wire \result_reg[30] ;
 wire \result_reg[31] ;
 wire \result_reg[3] ;
 wire \result_reg[4] ;
 wire \result_reg[5] ;
 wire \result_reg[6] ;
 wire \result_reg[7] ;
 wire \result_reg[8] ;
 wire \result_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire wr_prev;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;

 sg13g2_inv_2 _2708_ (.Y(_2189_),
    .A(\mac_inst.RDY_get_mac ));
 sg13g2_inv_2 _2709_ (.Y(_2190_),
    .A(\mac_inst.RDY_get_multiply ));
 sg13g2_inv_1 _2710_ (.Y(_2191_),
    .A(\mac_inst.accumulator[13] ));
 sg13g2_inv_1 _2711_ (.Y(_2192_),
    .A(\mac_inst.accumulator[12] ));
 sg13g2_inv_1 _2712_ (.Y(_2193_),
    .A(net205));
 sg13g2_inv_1 _2713_ (.Y(_2194_),
    .A(net202));
 sg13g2_inv_2 _2714_ (.Y(_2195_),
    .A(net673));
 sg13g2_inv_1 _2715_ (.Y(_2196_),
    .A(net150));
 sg13g2_inv_1 _2716_ (.Y(_2197_),
    .A(net145));
 sg13g2_inv_1 _2717_ (.Y(_2198_),
    .A(net146));
 sg13g2_inv_1 _2718_ (.Y(_2199_),
    .A(net151));
 sg13g2_inv_1 _2719_ (.Y(_2200_),
    .A(net154));
 sg13g2_inv_1 _2720_ (.Y(_2201_),
    .A(net141));
 sg13g2_inv_1 _2721_ (.Y(_2202_),
    .A(net142));
 sg13g2_inv_1 _2722_ (.Y(_2203_),
    .A(\cordic_inst.result_ready ));
 sg13g2_inv_1 _2723_ (.Y(_2204_),
    .A(\cordic_inst.cordic_state[51] ));
 sg13g2_inv_1 _2724_ (.Y(_2205_),
    .A(net341));
 sg13g2_inv_1 _2725_ (.Y(_2206_),
    .A(net314));
 sg13g2_inv_2 _2726_ (.Y(_2207_),
    .A(net405));
 sg13g2_inv_2 _2727_ (.Y(_2208_),
    .A(net406));
 sg13g2_inv_1 _2728_ (.Y(_2209_),
    .A(\cordic_atan2_result[6] ));
 sg13g2_inv_1 _2729_ (.Y(_2210_),
    .A(net654));
 sg13g2_inv_2 _2730_ (.Y(_2211_),
    .A(net659));
 sg13g2_inv_2 _2731_ (.Y(_2212_),
    .A(net382));
 sg13g2_inv_1 _2732_ (.Y(_2213_),
    .A(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ));
 sg13g2_inv_1 _2733_ (.Y(_2214_),
    .A(net250));
 sg13g2_inv_4 _2734_ (.A(net788),
    .Y(_2215_));
 sg13g2_inv_2 _2735_ (.Y(_2216_),
    .A(net677));
 sg13g2_inv_4 _2736_ (.A(net670),
    .Y(_2217_));
 sg13g2_inv_2 _2737_ (.Y(_2218_),
    .A(net738));
 sg13g2_inv_2 _2738_ (.Y(_2219_),
    .A(net734));
 sg13g2_inv_4 _2739_ (.A(net725),
    .Y(_2220_));
 sg13g2_inv_2 _2740_ (.Y(_2221_),
    .A(net719));
 sg13g2_inv_1 _2741_ (.Y(_2222_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[5] ));
 sg13g2_inv_1 _2742_ (.Y(_2223_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[7] ));
 sg13g2_inv_1 _2743_ (.Y(_2224_),
    .A(net711));
 sg13g2_inv_4 _2744_ (.A(net746),
    .Y(_2225_));
 sg13g2_inv_2 _2745_ (.Y(_2226_),
    .A(net744));
 sg13g2_inv_2 _2746_ (.Y(_2227_),
    .A(net640));
 sg13g2_inv_1 _2747_ (.Y(_2228_),
    .A(net634));
 sg13g2_inv_2 _2748_ (.Y(_2229_),
    .A(net624));
 sg13g2_inv_4 _2749_ (.A(net620),
    .Y(_2230_));
 sg13g2_inv_1 _2750_ (.Y(_2231_),
    .A(net618));
 sg13g2_inv_1 _2751_ (.Y(_2232_),
    .A(net708));
 sg13g2_inv_4 _2752_ (.A(net687),
    .Y(_2233_));
 sg13g2_inv_1 _2753_ (.Y(_2234_),
    .A(net642));
 sg13g2_nor2_1 _2754_ (.A(net332),
    .B(net344),
    .Y(_2235_));
 sg13g2_and2_1 _2755_ (.A(net741),
    .B(_2235_),
    .X(_2236_));
 sg13g2_nand2_2 _2756_ (.Y(_2237_),
    .A(net741),
    .B(_2235_));
 sg13g2_nor2_1 _2757_ (.A(net217),
    .B(net176),
    .Y(_2238_));
 sg13g2_nand3b_1 _2758_ (.B(net271),
    .C(_2238_),
    .Y(_2239_),
    .A_N(net258));
 sg13g2_nor2_1 _2759_ (.A(net138),
    .B(net320),
    .Y(_2240_));
 sg13g2_nor4_2 _2760_ (.A(\cmd_reg[1] ),
    .B(net138),
    .C(\cmd_reg[2] ),
    .Y(_2241_),
    .D(_2239_));
 sg13g2_nand3b_1 _2761_ (.B(_2240_),
    .C(net317),
    .Y(_2242_),
    .A_N(net740));
 sg13g2_nand3b_1 _2762_ (.B(_2238_),
    .C(net258),
    .Y(_2243_),
    .A_N(net271));
 sg13g2_nor2_1 _2763_ (.A(_2242_),
    .B(_2243_),
    .Y(_2244_));
 sg13g2_or2_1 _2764_ (.X(_2245_),
    .B(_2243_),
    .A(_2242_));
 sg13g2_nor4_2 _2765_ (.A(net317),
    .B(net138),
    .C(net320),
    .Y(_2246_),
    .D(_2243_));
 sg13g2_nor2_1 _2766_ (.A(_2244_),
    .B(_2246_),
    .Y(_2247_));
 sg13g2_and2_1 _2767_ (.A(net740),
    .B(_2246_),
    .X(_2248_));
 sg13g2_nand2_1 _2768_ (.Y(_2249_),
    .A(net740),
    .B(_2246_));
 sg13g2_nor2_1 _2769_ (.A(_2241_),
    .B(net572),
    .Y(_2250_));
 sg13g2_nor3_1 _2770_ (.A(_2241_),
    .B(_2244_),
    .C(net572),
    .Y(_2251_));
 sg13g2_nand2_2 _2771_ (.Y(_2252_),
    .A(_2245_),
    .B(net555));
 sg13g2_nor2b_2 _2772_ (.A(net740),
    .B_N(_2246_),
    .Y(_2253_));
 sg13g2_nand2b_2 _2773_ (.Y(_2254_),
    .B(_2246_),
    .A_N(net740));
 sg13g2_o21ai_1 _2774_ (.B1(_2236_),
    .Y(_2255_),
    .A1(_2252_),
    .A2(_2253_));
 sg13g2_nor2b_2 _2775_ (.A(net379),
    .B_N(\state[0] ),
    .Y(_2256_));
 sg13g2_nor2b_2 _2776_ (.A(net741),
    .B_N(_2256_),
    .Y(_2257_));
 sg13g2_nand2b_1 _2777_ (.Y(_2258_),
    .B(_2256_),
    .A_N(net741));
 sg13g2_or2_1 _2778_ (.X(_2259_),
    .B(_2242_),
    .A(_2239_));
 sg13g2_and2_1 _2779_ (.A(_2257_),
    .B(_2259_),
    .X(_2260_));
 sg13g2_nor3_2 _2780_ (.A(net741),
    .B(net332),
    .C(\state[1] ),
    .Y(_2261_));
 sg13g2_nor2_1 _2781_ (.A(net741),
    .B(_2235_),
    .Y(_2262_));
 sg13g2_nor2b_2 _2782_ (.A(net315),
    .B_N(net9),
    .Y(_2263_));
 sg13g2_nand2b_2 _2783_ (.Y(_2264_),
    .B(net9),
    .A_N(wr_prev));
 sg13g2_nor2b_1 _2784_ (.A(net763),
    .B_N(net765),
    .Y(_2265_));
 sg13g2_nand2_1 _2785_ (.Y(_2266_),
    .A(_2263_),
    .B(_2265_));
 sg13g2_nor2b_2 _2786_ (.A(net741),
    .B_N(net344),
    .Y(_2267_));
 sg13g2_nand2_1 _2787_ (.Y(_2268_),
    .A(_2266_),
    .B(_2267_));
 sg13g2_nor2b_1 _2788_ (.A(_2260_),
    .B_N(_2268_),
    .Y(_2269_));
 sg13g2_o21ai_1 _2789_ (.B1(_2269_),
    .Y(_2270_),
    .A1(_2236_),
    .A2(_2262_));
 sg13g2_nor2b_2 _2790_ (.A(net332),
    .B_N(_2267_),
    .Y(_2271_));
 sg13g2_inv_1 _2791_ (.Y(_2272_),
    .A(_2271_));
 sg13g2_nor2_1 _2792_ (.A(_2266_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_a21o_1 _2793_ (.A2(net569),
    .A1(_2252_),
    .B1(_2270_),
    .X(_2274_));
 sg13g2_nor2_1 _2794_ (.A(_2236_),
    .B(_2274_),
    .Y(_2275_));
 sg13g2_a21oi_1 _2795_ (.A1(_2234_),
    .A2(_2255_),
    .Y(_0018_),
    .B1(_2275_));
 sg13g2_and2_1 _2796_ (.A(net740),
    .B(_2241_),
    .X(_2276_));
 sg13g2_nand2_1 _2797_ (.Y(_2277_),
    .A(net740),
    .B(net139));
 sg13g2_nor3_1 _2798_ (.A(net133),
    .B(_2237_),
    .C(_2277_),
    .Y(_0010_));
 sg13g2_nor2b_1 _2799_ (.A(\cmd_reg[0] ),
    .B_N(_2241_),
    .Y(_2278_));
 sg13g2_nand2b_2 _2800_ (.Y(_2279_),
    .B(net139),
    .A_N(net135));
 sg13g2_nor3_1 _2801_ (.A(net133),
    .B(_2237_),
    .C(_2279_),
    .Y(_0011_));
 sg13g2_nor3_1 _2802_ (.A(net642),
    .B(net592),
    .C(_2245_),
    .Y(_0006_));
 sg13g2_nor3_1 _2803_ (.A(net133),
    .B(_2237_),
    .C(net136),
    .Y(_0001_));
 sg13g2_nor2b_1 _2804_ (.A(net679),
    .B_N(cordic_en_atan2),
    .Y(_2280_));
 sg13g2_nor2_2 _2805_ (.A(net682),
    .B(net676),
    .Y(_2281_));
 sg13g2_nor2_2 _2806_ (.A(net685),
    .B(net683),
    .Y(_2282_));
 sg13g2_nor3_2 _2807_ (.A(net685),
    .B(net683),
    .C(net681),
    .Y(_2283_));
 sg13g2_nand2_2 _2808_ (.Y(_2284_),
    .A(_2216_),
    .B(_2282_));
 sg13g2_nand2_2 _2809_ (.Y(_2285_),
    .A(net784),
    .B(net600));
 sg13g2_a21oi_1 _2810_ (.A1(net152),
    .A2(net600),
    .Y(_2286_),
    .B1(net603));
 sg13g2_nor2_1 _2811_ (.A(net769),
    .B(net153),
    .Y(_0014_));
 sg13g2_nor2_2 _2812_ (.A(\cordic_inst.cordic_state[0] ),
    .B(_2212_),
    .Y(_2287_));
 sg13g2_nand2b_2 _2813_ (.Y(_2288_),
    .B(cordic_busy),
    .A_N(\cordic_inst.cordic_state[0] ));
 sg13g2_nor2_2 _2814_ (.A(net684),
    .B(_2288_),
    .Y(_2289_));
 sg13g2_or2_1 _2815_ (.X(_2290_),
    .B(_2288_),
    .A(net684));
 sg13g2_nand2_2 _2816_ (.Y(_2291_),
    .A(_2282_),
    .B(_2287_));
 sg13g2_nor2_2 _2817_ (.A(net675),
    .B(net584),
    .Y(_2292_));
 sg13g2_nand2_2 _2818_ (.Y(_2293_),
    .A(_2281_),
    .B(net590));
 sg13g2_a21o_2 _2819_ (.A2(net665),
    .A1(net660),
    .B1(net658),
    .X(_2294_));
 sg13g2_nand2_2 _2820_ (.Y(_2295_),
    .A(net669),
    .B(_2287_));
 sg13g2_nand2_2 _2821_ (.Y(_2296_),
    .A(net658),
    .B(net660));
 sg13g2_nor2_1 _2822_ (.A(_2295_),
    .B(_2296_),
    .Y(_2297_));
 sg13g2_nor2_1 _2823_ (.A(_2293_),
    .B(_2297_),
    .Y(_2298_));
 sg13g2_nor2_2 _2824_ (.A(_2284_),
    .B(_2287_),
    .Y(_2299_));
 sg13g2_nand2_2 _2825_ (.Y(_2300_),
    .A(_2283_),
    .B(_2288_));
 sg13g2_a21o_1 _2826_ (.A2(net578),
    .A1(net658),
    .B1(net770),
    .X(_2301_));
 sg13g2_a21oi_2 _2827_ (.B1(_2301_),
    .Y(_2302_),
    .A2(_2298_),
    .A1(_2294_));
 sg13g2_inv_1 _2828_ (.Y(_0111_),
    .A(_2302_));
 sg13g2_xnor2_1 _2829_ (.Y(_2303_),
    .A(net660),
    .B(_2295_));
 sg13g2_and2_1 _2830_ (.A(net600),
    .B(_2303_),
    .X(_2304_));
 sg13g2_nand2b_1 _2831_ (.Y(_2305_),
    .B(_2302_),
    .A_N(_2304_));
 sg13g2_nor2_1 _2832_ (.A(net654),
    .B(_2297_),
    .Y(_2306_));
 sg13g2_nor3_2 _2833_ (.A(_2210_),
    .B(_2295_),
    .C(_2296_),
    .Y(_2307_));
 sg13g2_nor3_2 _2834_ (.A(_2285_),
    .B(_2306_),
    .C(_2307_),
    .Y(_0112_));
 sg13g2_nand2b_2 _2835_ (.Y(_2308_),
    .B(_2302_),
    .A_N(_0112_));
 sg13g2_xor2_1 _2836_ (.B(_2288_),
    .A(net665),
    .X(_2309_));
 sg13g2_o21ai_1 _2837_ (.B1(net776),
    .Y(_0109_),
    .A1(_2284_),
    .A2(_2309_));
 sg13g2_nor2_1 _2838_ (.A(_2308_),
    .B(_0109_),
    .Y(_2310_));
 sg13g2_o21ai_1 _2839_ (.B1(_2305_),
    .Y(_0000_),
    .A1(_2308_),
    .A2(_0109_));
 sg13g2_nand2b_2 _2840_ (.Y(_2311_),
    .B(net642),
    .A_N(\exec_phase[2] ));
 sg13g2_or2_1 _2841_ (.X(_2312_),
    .B(_2311_),
    .A(_2214_));
 sg13g2_or2_1 _2842_ (.X(_2313_),
    .B(_2312_),
    .A(net592));
 sg13g2_nor2_1 _2843_ (.A(_2277_),
    .B(_2313_),
    .Y(_0008_));
 sg13g2_nor2_1 _2844_ (.A(_2279_),
    .B(_2313_),
    .Y(_0009_));
 sg13g2_nor2_1 _2845_ (.A(_2245_),
    .B(_2313_),
    .Y(_0004_));
 sg13g2_nor2_1 _2846_ (.A(net136),
    .B(_2313_),
    .Y(_0002_));
 sg13g2_nor2_1 _2847_ (.A(_2254_),
    .B(_2313_),
    .Y(_0003_));
 sg13g2_nor2_1 _2848_ (.A(net592),
    .B(_2259_),
    .Y(_2314_));
 sg13g2_nor3_1 _2849_ (.A(net642),
    .B(net592),
    .C(_2259_),
    .Y(_0007_));
 sg13g2_a21oi_1 _2850_ (.A1(net155),
    .A2(_2282_),
    .Y(_2315_),
    .B1(net681));
 sg13g2_nor2_1 _2851_ (.A(net770),
    .B(net156),
    .Y(_0013_));
 sg13g2_nand3_1 _2852_ (.B(_2190_),
    .C(_2241_),
    .A(_2189_),
    .Y(_2316_));
 sg13g2_o21ai_1 _2853_ (.B1(_2316_),
    .Y(_2317_),
    .A1(cordic_busy),
    .A2(_2247_));
 sg13g2_nand3_1 _2854_ (.B(_2236_),
    .C(_2317_),
    .A(\exec_phase[2] ),
    .Y(_2318_));
 sg13g2_a21oi_1 _2855_ (.A1(_2214_),
    .A2(_2318_),
    .Y(_0015_),
    .B1(_2275_));
 sg13g2_o21ai_1 _2856_ (.B1(_2281_),
    .Y(_2319_),
    .A1(net684),
    .A2(net310));
 sg13g2_nand2_1 _2857_ (.Y(_0012_),
    .A(net783),
    .B(net311));
 sg13g2_nor2_1 _2858_ (.A(net592),
    .B(_2317_),
    .Y(_2320_));
 sg13g2_o21ai_1 _2859_ (.B1(net254),
    .Y(_2321_),
    .A1(_2274_),
    .A2(_2320_));
 sg13g2_o21ai_1 _2860_ (.B1(net255),
    .Y(_0016_),
    .A1(net642),
    .A2(_2255_));
 sg13g2_nor3_1 _2861_ (.A(net642),
    .B(net592),
    .C(_2254_),
    .Y(_0005_));
 sg13g2_nor2_1 _2862_ (.A(\exec_phase[1] ),
    .B(_2311_),
    .Y(_2322_));
 sg13g2_o21ai_1 _2863_ (.B1(net642),
    .Y(_2323_),
    .A1(\exec_phase[1] ),
    .A2(\exec_phase[2] ));
 sg13g2_o21ai_1 _2864_ (.B1(_2323_),
    .Y(_2324_),
    .A1(net572),
    .A2(net563));
 sg13g2_a22oi_1 _2865_ (.Y(_2325_),
    .B1(_2253_),
    .B2(_2311_),
    .A2(net572),
    .A1(\exec_phase[2] ));
 sg13g2_a21oi_1 _2866_ (.A1(_2324_),
    .A2(_2325_),
    .Y(_2326_),
    .B1(net592));
 sg13g2_a21oi_1 _2867_ (.A1(_2253_),
    .A2(_2322_),
    .Y(_2327_),
    .B1(net567));
 sg13g2_o21ai_1 _2868_ (.B1(_2236_),
    .Y(_2328_),
    .A1(_2189_),
    .A2(_2312_));
 sg13g2_nand3_1 _2869_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[0] ),
    .A(\cordic_inst.result_ready ),
    .Y(_2329_));
 sg13g2_nand2_1 _2870_ (.Y(_2330_),
    .A(_0003_),
    .B(_2329_));
 sg13g2_o21ai_1 _2871_ (.B1(_2330_),
    .Y(_2331_),
    .A1(_2327_),
    .A2(_2328_));
 sg13g2_nand3_1 _2872_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[1] ),
    .A(\cordic_inst.result_ready ),
    .Y(_2332_));
 sg13g2_nor2_1 _2873_ (.A(_2312_),
    .B(_2332_),
    .Y(_2333_));
 sg13g2_nor3_1 _2874_ (.A(net592),
    .B(_2245_),
    .C(_2333_),
    .Y(_2334_));
 sg13g2_and2_1 _2875_ (.A(_2260_),
    .B(_2264_),
    .X(_2335_));
 sg13g2_nor4_1 _2876_ (.A(_2326_),
    .B(_2331_),
    .C(_2334_),
    .D(_2335_),
    .Y(_2336_));
 sg13g2_nand2_2 _2877_ (.Y(_2337_),
    .A(net741),
    .B(_2256_));
 sg13g2_xnor2_1 _2878_ (.Y(_2338_),
    .A(net763),
    .B(_2253_));
 sg13g2_nand2_1 _2879_ (.Y(_2339_),
    .A(net765),
    .B(_2338_));
 sg13g2_nand3_1 _2880_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[2] ),
    .A(\cordic_inst.result_ready ),
    .Y(_2340_));
 sg13g2_a22oi_1 _2881_ (.Y(_2341_),
    .B1(_2340_),
    .B2(net572),
    .A2(net563),
    .A1(_2190_));
 sg13g2_nor2_1 _2882_ (.A(_2313_),
    .B(_2341_),
    .Y(_2342_));
 sg13g2_nand4_1 _2883_ (.B(net642),
    .C(_2236_),
    .A(\exec_phase[2] ),
    .Y(_2343_),
    .D(net565));
 sg13g2_nor2b_1 _2884_ (.A(_2342_),
    .B_N(_2343_),
    .Y(_2344_));
 sg13g2_nand3_1 _2885_ (.B(_2251_),
    .C(_2254_),
    .A(_2236_),
    .Y(_2345_));
 sg13g2_o21ai_1 _2886_ (.B1(net344),
    .Y(_2346_),
    .A1(\state[2] ),
    .A2(_2264_));
 sg13g2_nor2b_2 _2887_ (.A(rd_prev),
    .B_N(net10),
    .Y(_2347_));
 sg13g2_nand3_1 _2888_ (.B(_2345_),
    .C(_2346_),
    .A(_2344_),
    .Y(_2348_));
 sg13g2_and2_1 _2889_ (.A(_2339_),
    .B(_2347_),
    .X(_2349_));
 sg13g2_o21ai_1 _2890_ (.B1(_2336_),
    .Y(_2350_),
    .A1(_2337_),
    .A2(_2349_));
 sg13g2_nor3_1 _2891_ (.A(_2275_),
    .B(_2348_),
    .C(_2350_),
    .Y(_2351_));
 sg13g2_nor2_1 _2892_ (.A(_2256_),
    .B(_2267_),
    .Y(_2352_));
 sg13g2_o21ai_1 _2893_ (.B1(_2258_),
    .Y(_2353_),
    .A1(net765),
    .A2(_2352_));
 sg13g2_mux2_1 _2894_ (.A0(net765),
    .A1(_2353_),
    .S(_2351_),
    .X(_0019_));
 sg13g2_nor2b_1 _2895_ (.A(net765),
    .B_N(net763),
    .Y(_2354_));
 sg13g2_a21oi_1 _2896_ (.A1(_2265_),
    .A2(_2272_),
    .Y(_2355_),
    .B1(_2354_));
 sg13g2_nor3_1 _2897_ (.A(_2257_),
    .B(_2352_),
    .C(_2355_),
    .Y(_2356_));
 sg13g2_mux2_1 _2898_ (.A0(net763),
    .A1(_2356_),
    .S(_2351_),
    .X(_0020_));
 sg13g2_mux2_1 _2899_ (.A0(net762),
    .A1(net1),
    .S(net568),
    .X(_0021_));
 sg13g2_mux2_1 _2900_ (.A0(net759),
    .A1(net2),
    .S(net568),
    .X(_0022_));
 sg13g2_mux2_1 _2901_ (.A0(net756),
    .A1(net3),
    .S(net568),
    .X(_0023_));
 sg13g2_mux2_1 _2902_ (.A0(net753),
    .A1(net4),
    .S(net568),
    .X(_0024_));
 sg13g2_mux2_1 _2903_ (.A0(net750),
    .A1(net5),
    .S(net569),
    .X(_0025_));
 sg13g2_mux2_1 _2904_ (.A0(net748),
    .A1(net6),
    .S(net569),
    .X(_0026_));
 sg13g2_nand2_1 _2905_ (.Y(_2357_),
    .A(net7),
    .B(net568));
 sg13g2_o21ai_1 _2906_ (.B1(_2357_),
    .Y(_0027_),
    .A1(_2225_),
    .A2(net568));
 sg13g2_nand2_1 _2907_ (.Y(_2358_),
    .A(net8),
    .B(net568));
 sg13g2_o21ai_1 _2908_ (.B1(_2358_),
    .Y(_0028_),
    .A1(_2226_),
    .A2(net568));
 sg13g2_nor2_2 _2909_ (.A(net659),
    .B(net664),
    .Y(_2359_));
 sg13g2_nand2_1 _2910_ (.Y(_2360_),
    .A(net652),
    .B(net656));
 sg13g2_nor2_1 _2911_ (.A(_2359_),
    .B(_2360_),
    .Y(_2361_));
 sg13g2_nand2_1 _2912_ (.Y(_2362_),
    .A(net776),
    .B(_2304_));
 sg13g2_inv_1 _2913_ (.Y(_0110_),
    .A(_2362_));
 sg13g2_nand2_1 _2914_ (.Y(_2363_),
    .A(_2309_),
    .B(_0110_));
 sg13g2_nor2_1 _2915_ (.A(_2308_),
    .B(_2363_),
    .Y(_0029_));
 sg13g2_nand2_1 _2916_ (.Y(_2364_),
    .A(_0109_),
    .B(_2362_));
 sg13g2_nor2_1 _2917_ (.A(_2308_),
    .B(_2364_),
    .Y(_0030_));
 sg13g2_inv_1 _2918_ (.Y(_2365_),
    .A(_0030_));
 sg13g2_nor2_1 _2919_ (.A(_2304_),
    .B(_2308_),
    .Y(_0164_));
 sg13g2_or2_1 _2920_ (.X(_2366_),
    .B(_0109_),
    .A(_2304_));
 sg13g2_nand2_1 _2921_ (.Y(_2367_),
    .A(\cordic_inst.cordic_state[39] ),
    .B(net553));
 sg13g2_nand2_1 _2922_ (.Y(_2368_),
    .A(\cordic_atan2_result[0] ),
    .B(net571));
 sg13g2_a22oi_1 _2923_ (.Y(_2369_),
    .B1(net563),
    .B2(net142),
    .A2(net567),
    .A1(\mac_inst.accumulator[0] ));
 sg13g2_nand3_1 _2924_ (.B(_2368_),
    .C(_2369_),
    .A(_2367_),
    .Y(_2370_));
 sg13g2_a22oi_1 _2925_ (.Y(_2371_),
    .B1(_2332_),
    .B2(_2244_),
    .A2(_2329_),
    .A1(_2253_));
 sg13g2_a21oi_1 _2926_ (.A1(_2341_),
    .A2(_2371_),
    .Y(_2372_),
    .B1(_2312_));
 sg13g2_nand2_1 _2927_ (.Y(_2373_),
    .A(_2247_),
    .B(_2279_));
 sg13g2_a221oi_1 _2928_ (.B2(_2311_),
    .C1(_2255_),
    .B1(_2373_),
    .A1(_2252_),
    .Y(_2374_),
    .A2(_2322_));
 sg13g2_nor2_1 _2929_ (.A(_2331_),
    .B(_2372_),
    .Y(_2375_));
 sg13g2_nand2_1 _2930_ (.Y(_2376_),
    .A(_2374_),
    .B(_2375_));
 sg13g2_mux2_1 _2931_ (.A0(_2370_),
    .A1(net232),
    .S(net546),
    .X(_0031_));
 sg13g2_a22oi_1 _2932_ (.Y(_2377_),
    .B1(net567),
    .B2(\mac_inst.accumulator[1] ),
    .A2(net573),
    .A1(\cordic_atan2_result[1] ));
 sg13g2_a22oi_1 _2933_ (.Y(_2378_),
    .B1(net563),
    .B2(\mac_inst.get_multiply[1] ),
    .A2(net555),
    .A1(\cordic_inst.cordic_state[40] ));
 sg13g2_a21oi_1 _2934_ (.A1(_2377_),
    .A2(_2378_),
    .Y(_2379_),
    .B1(net547));
 sg13g2_a21o_1 _2935_ (.A2(net546),
    .A1(net159),
    .B1(_2379_),
    .X(_0032_));
 sg13g2_a22oi_1 _2936_ (.Y(_2380_),
    .B1(net565),
    .B2(\mac_inst.get_multiply[2] ),
    .A2(net566),
    .A1(\mac_inst.accumulator[2] ));
 sg13g2_a22oi_1 _2937_ (.Y(_2381_),
    .B1(net555),
    .B2(\cordic_inst.cordic_state[41] ),
    .A2(net572),
    .A1(\cordic_atan2_result[2] ));
 sg13g2_nand2_2 _2938_ (.Y(_2382_),
    .A(_2380_),
    .B(_2381_));
 sg13g2_mux2_1 _2939_ (.A0(_2382_),
    .A1(net194),
    .S(net545),
    .X(_0033_));
 sg13g2_a22oi_1 _2940_ (.Y(_2383_),
    .B1(net564),
    .B2(net141),
    .A2(net566),
    .A1(\mac_inst.accumulator[3] ));
 sg13g2_a22oi_1 _2941_ (.Y(_2384_),
    .B1(net555),
    .B2(\cordic_inst.cordic_state[42] ),
    .A2(net572),
    .A1(\cordic_atan2_result[3] ));
 sg13g2_nand2_2 _2942_ (.Y(_2385_),
    .A(_2383_),
    .B(_2384_));
 sg13g2_mux2_1 _2943_ (.A0(_2385_),
    .A1(net209),
    .S(net545),
    .X(_0034_));
 sg13g2_nand2_1 _2944_ (.Y(_2386_),
    .A(\cordic_inst.cordic_state[43] ),
    .B(net553));
 sg13g2_nand2_1 _2945_ (.Y(_2387_),
    .A(\mac_inst.accumulator[4] ),
    .B(net566));
 sg13g2_a22oi_1 _2946_ (.Y(_2388_),
    .B1(net563),
    .B2(\mac_inst.get_multiply[4] ),
    .A2(net570),
    .A1(\cordic_atan2_result[4] ));
 sg13g2_nand3_1 _2947_ (.B(_2387_),
    .C(_2388_),
    .A(_2386_),
    .Y(_2389_));
 sg13g2_mux2_1 _2948_ (.A0(_2389_),
    .A1(net180),
    .S(net547),
    .X(_0035_));
 sg13g2_nand2_1 _2949_ (.Y(_2390_),
    .A(\cordic_inst.cordic_state[44] ),
    .B(net553));
 sg13g2_a22oi_1 _2950_ (.Y(_2391_),
    .B1(net567),
    .B2(\mac_inst.accumulator[5] ),
    .A2(net570),
    .A1(\cordic_atan2_result[5] ));
 sg13g2_nand2_1 _2951_ (.Y(_2392_),
    .A(net154),
    .B(net563));
 sg13g2_nand3_1 _2952_ (.B(_2391_),
    .C(_2392_),
    .A(_2390_),
    .Y(_2393_));
 sg13g2_mux2_1 _2953_ (.A0(_2393_),
    .A1(net228),
    .S(net546),
    .X(_0036_));
 sg13g2_a22oi_1 _2954_ (.Y(_2394_),
    .B1(net564),
    .B2(net151),
    .A2(net566),
    .A1(\mac_inst.accumulator[6] ));
 sg13g2_a22oi_1 _2955_ (.Y(_2395_),
    .B1(net554),
    .B2(\cordic_inst.cordic_state[45] ),
    .A2(net570),
    .A1(\cordic_atan2_result[6] ));
 sg13g2_nand2_2 _2956_ (.Y(_2396_),
    .A(_2394_),
    .B(_2395_));
 sg13g2_mux2_1 _2957_ (.A0(_2396_),
    .A1(net198),
    .S(net545),
    .X(_0037_));
 sg13g2_nand2_1 _2958_ (.Y(_2397_),
    .A(\cordic_inst.cordic_state[46] ),
    .B(net554));
 sg13g2_nand2_1 _2959_ (.Y(_2398_),
    .A(\cordic_atan2_result[7] ),
    .B(net570));
 sg13g2_a22oi_1 _2960_ (.Y(_2399_),
    .B1(net564),
    .B2(\mac_inst.get_multiply[7] ),
    .A2(_2276_),
    .A1(\mac_inst.accumulator[7] ));
 sg13g2_nand3_1 _2961_ (.B(_2398_),
    .C(_2399_),
    .A(_2397_),
    .Y(_2400_));
 sg13g2_mux2_1 _2962_ (.A0(_2400_),
    .A1(net174),
    .S(net547),
    .X(_0038_));
 sg13g2_a22oi_1 _2963_ (.Y(_2401_),
    .B1(net564),
    .B2(\mac_inst.get_multiply[8] ),
    .A2(_2276_),
    .A1(\mac_inst.accumulator[8] ));
 sg13g2_a22oi_1 _2964_ (.Y(_2402_),
    .B1(net554),
    .B2(\cordic_inst.cordic_state[47] ),
    .A2(net570),
    .A1(\cordic_atan2_result[8] ));
 sg13g2_nand2_1 _2965_ (.Y(_2403_),
    .A(_2401_),
    .B(_2402_));
 sg13g2_mux2_1 _2966_ (.A0(_2403_),
    .A1(net215),
    .S(net545),
    .X(_0039_));
 sg13g2_a22oi_1 _2967_ (.Y(_2404_),
    .B1(net564),
    .B2(net145),
    .A2(net567),
    .A1(\mac_inst.accumulator[9] ));
 sg13g2_a22oi_1 _2968_ (.Y(_2405_),
    .B1(net554),
    .B2(\cordic_inst.cordic_state[48] ),
    .A2(net570),
    .A1(\cordic_atan2_result[9] ));
 sg13g2_nand2_1 _2969_ (.Y(_2406_),
    .A(_2404_),
    .B(_2405_));
 sg13g2_mux2_1 _2970_ (.A0(_2406_),
    .A1(net196),
    .S(net546),
    .X(_0040_));
 sg13g2_nand2_1 _2971_ (.Y(_2407_),
    .A(\cordic_inst.cordic_state[49] ),
    .B(net553));
 sg13g2_nand2_1 _2972_ (.Y(_2408_),
    .A(\mac_inst.get_multiply[10] ),
    .B(net564));
 sg13g2_a22oi_1 _2973_ (.Y(_2409_),
    .B1(net567),
    .B2(\mac_inst.accumulator[10] ),
    .A2(net570),
    .A1(\cordic_atan2_result[10] ));
 sg13g2_nand3_1 _2974_ (.B(_2408_),
    .C(_2409_),
    .A(_2407_),
    .Y(_2410_));
 sg13g2_mux2_1 _2975_ (.A0(_2410_),
    .A1(net204),
    .S(net545),
    .X(_0041_));
 sg13g2_a22oi_1 _2976_ (.Y(_2411_),
    .B1(net567),
    .B2(\mac_inst.accumulator[11] ),
    .A2(net571),
    .A1(\cordic_atan2_result[11] ));
 sg13g2_a22oi_1 _2977_ (.Y(_2412_),
    .B1(net563),
    .B2(\mac_inst.get_multiply[11] ),
    .A2(net554),
    .A1(\cordic_inst.cordic_state[50] ));
 sg13g2_a21oi_2 _2978_ (.B1(net547),
    .Y(_2413_),
    .A2(_2412_),
    .A1(_2411_));
 sg13g2_a21o_1 _2979_ (.A2(net545),
    .A1(net157),
    .B1(_2413_),
    .X(_0042_));
 sg13g2_a22oi_1 _2980_ (.Y(_2414_),
    .B1(net564),
    .B2(\mac_inst.get_multiply[12] ),
    .A2(net566),
    .A1(\mac_inst.accumulator[12] ));
 sg13g2_a22oi_1 _2981_ (.Y(_2415_),
    .B1(net553),
    .B2(\cordic_inst.cordic_state[51] ),
    .A2(net571),
    .A1(\cordic_atan2_result[12] ));
 sg13g2_nand2_2 _2982_ (.Y(_2416_),
    .A(_2414_),
    .B(_2415_));
 sg13g2_mux2_1 _2983_ (.A0(_2416_),
    .A1(net186),
    .S(net547),
    .X(_0043_));
 sg13g2_nand2_1 _2984_ (.Y(_2417_),
    .A(\cordic_inst.cordic_state[52] ),
    .B(net553));
 sg13g2_a22oi_1 _2985_ (.Y(_2418_),
    .B1(net563),
    .B2(\mac_inst.get_multiply[13] ),
    .A2(net572),
    .A1(\cordic_atan2_result[13] ));
 sg13g2_nand2_1 _2986_ (.Y(_2419_),
    .A(\mac_inst.accumulator[13] ),
    .B(net566));
 sg13g2_nand3_1 _2987_ (.B(_2418_),
    .C(_2419_),
    .A(_2417_),
    .Y(_2420_));
 sg13g2_mux2_1 _2988_ (.A0(_2420_),
    .A1(net184),
    .S(net545),
    .X(_0044_));
 sg13g2_a22oi_1 _2989_ (.Y(_2421_),
    .B1(net564),
    .B2(\mac_inst.get_multiply[14] ),
    .A2(net566),
    .A1(\mac_inst.accumulator[14] ));
 sg13g2_a22oi_1 _2990_ (.Y(_2422_),
    .B1(net553),
    .B2(\cordic_inst.cordic_state[53] ),
    .A2(net570),
    .A1(\cordic_atan2_result[14] ));
 sg13g2_nand2_2 _2991_ (.Y(_2423_),
    .A(_2421_),
    .B(_2422_));
 sg13g2_mux2_1 _2992_ (.A0(_2423_),
    .A1(net178),
    .S(net545),
    .X(_0045_));
 sg13g2_a22oi_1 _2993_ (.Y(_2424_),
    .B1(net565),
    .B2(\mac_inst.get_multiply[15] ),
    .A2(net566),
    .A1(net164));
 sg13g2_a22oi_1 _2994_ (.Y(_2425_),
    .B1(net553),
    .B2(net645),
    .A2(net571),
    .A1(\cordic_atan2_result[15] ));
 sg13g2_nand2_1 _2995_ (.Y(_2426_),
    .A(_2424_),
    .B(_2425_));
 sg13g2_mux2_1 _2996_ (.A0(_2426_),
    .A1(net238),
    .S(net547),
    .X(_0046_));
 sg13g2_or2_1 _2997_ (.X(_2427_),
    .B(_0112_),
    .A(_2302_));
 sg13g2_nor3_1 _2998_ (.A(_2309_),
    .B(_2362_),
    .C(_2427_),
    .Y(_0048_));
 sg13g2_nor2_1 _2999_ (.A(_2364_),
    .B(_2427_),
    .Y(_0049_));
 sg13g2_nor2_1 _3000_ (.A(_2366_),
    .B(_2427_),
    .Y(_0050_));
 sg13g2_nor2_1 _3001_ (.A(_0029_),
    .B(_0030_),
    .Y(_2428_));
 sg13g2_nand2b_1 _3002_ (.Y(_0051_),
    .B(_2428_),
    .A_N(_0048_));
 sg13g2_o21ai_1 _3003_ (.B1(_2365_),
    .Y(_0052_),
    .A1(_0112_),
    .A2(_2363_));
 sg13g2_or2_1 _3004_ (.X(_0053_),
    .B(_0049_),
    .A(_2310_));
 sg13g2_nand2b_1 _3005_ (.Y(_0054_),
    .B(_2428_),
    .A_N(_0050_));
 sg13g2_nor2_2 _3006_ (.A(_2256_),
    .B(_2261_),
    .Y(_2429_));
 sg13g2_or2_1 _3007_ (.X(_2430_),
    .B(net763),
    .A(net765));
 sg13g2_and2_1 _3008_ (.A(net766),
    .B(net764),
    .X(_2431_));
 sg13g2_nor2b_2 _3009_ (.A(_2337_),
    .B_N(_2347_),
    .Y(_2432_));
 sg13g2_mux4_1 _3010_ (.S0(net765),
    .A0(net232),
    .A1(net215),
    .A2(net256),
    .A3(net147),
    .S1(net763),
    .X(_2433_));
 sg13g2_a22oi_1 _3011_ (.Y(_2434_),
    .B1(_2432_),
    .B2(_2433_),
    .A2(_2429_),
    .A1(net269));
 sg13g2_inv_1 _3012_ (.Y(_0055_),
    .A(net270));
 sg13g2_mux4_1 _3013_ (.S0(net766),
    .A0(net159),
    .A1(net196),
    .A2(net236),
    .A3(net190),
    .S1(net764),
    .X(_2435_));
 sg13g2_a22oi_1 _3014_ (.Y(_2436_),
    .B1(_2432_),
    .B2(_2435_),
    .A2(_2429_),
    .A1(net282));
 sg13g2_inv_1 _3015_ (.Y(_0056_),
    .A(net283));
 sg13g2_mux4_1 _3016_ (.S0(net766),
    .A0(net194),
    .A1(net204),
    .A2(net221),
    .A3(net192),
    .S1(net764),
    .X(_2437_));
 sg13g2_a22oi_1 _3017_ (.Y(_2438_),
    .B1(_2432_),
    .B2(_2437_),
    .A2(_2429_),
    .A1(net280));
 sg13g2_inv_1 _3018_ (.Y(_0057_),
    .A(net281));
 sg13g2_mux4_1 _3019_ (.S0(net766),
    .A0(net209),
    .A1(net157),
    .A2(net182),
    .A3(net226),
    .S1(net764),
    .X(_2439_));
 sg13g2_a22oi_1 _3020_ (.Y(_2440_),
    .B1(_2432_),
    .B2(_2439_),
    .A2(_2429_),
    .A1(net267));
 sg13g2_inv_1 _3021_ (.Y(_0058_),
    .A(net268));
 sg13g2_mux4_1 _3022_ (.S0(net765),
    .A0(net180),
    .A1(net186),
    .A2(net213),
    .A3(net161),
    .S1(net763),
    .X(_2441_));
 sg13g2_a22oi_1 _3023_ (.Y(_2442_),
    .B1(_2432_),
    .B2(_2441_),
    .A2(_2429_),
    .A1(net275));
 sg13g2_inv_1 _3024_ (.Y(_0059_),
    .A(net276));
 sg13g2_mux4_1 _3025_ (.S0(net766),
    .A0(net228),
    .A1(net184),
    .A2(net172),
    .A3(net207),
    .S1(net764),
    .X(_2443_));
 sg13g2_a22oi_1 _3026_ (.Y(_2444_),
    .B1(_2432_),
    .B2(_2443_),
    .A2(_2429_),
    .A1(net284));
 sg13g2_inv_1 _3027_ (.Y(_0060_),
    .A(net285));
 sg13g2_mux4_1 _3028_ (.S0(net766),
    .A0(net198),
    .A1(net178),
    .A2(net240),
    .A3(net200),
    .S1(net764),
    .X(_2445_));
 sg13g2_a22oi_1 _3029_ (.Y(_2446_),
    .B1(_2432_),
    .B2(_2445_),
    .A2(_2429_),
    .A1(net312));
 sg13g2_inv_1 _3030_ (.Y(_0061_),
    .A(net313));
 sg13g2_nand2b_1 _3031_ (.Y(_2447_),
    .B(net238),
    .A_N(net763));
 sg13g2_a22oi_1 _3032_ (.Y(_2448_),
    .B1(_2431_),
    .B2(net170),
    .A2(_2354_),
    .A1(net188));
 sg13g2_nand3_1 _3033_ (.B(_2447_),
    .C(_2448_),
    .A(_2430_),
    .Y(_2449_));
 sg13g2_or2_1 _3034_ (.X(_2450_),
    .B(_2430_),
    .A(net174));
 sg13g2_nand4_1 _3035_ (.B(_2347_),
    .C(_2449_),
    .A(_2256_),
    .Y(_2451_),
    .D(_2450_));
 sg13g2_a21oi_1 _3036_ (.A1(net299),
    .A2(_2429_),
    .Y(_2452_),
    .B1(_2257_));
 sg13g2_nand2_1 _3037_ (.Y(_0062_),
    .A(_2451_),
    .B(net300));
 sg13g2_nand2_1 _3038_ (.Y(_2453_),
    .A(_2339_),
    .B(_2432_));
 sg13g2_o21ai_1 _3039_ (.B1(_2268_),
    .Y(_2454_),
    .A1(_2337_),
    .A2(_2347_));
 sg13g2_nand3_1 _3040_ (.B(_2190_),
    .C(_2234_),
    .A(_2189_),
    .Y(_2455_));
 sg13g2_a221oi_1 _3041_ (.B2(_2455_),
    .C1(_2454_),
    .B1(_2314_),
    .A1(_2261_),
    .Y(_2456_),
    .A2(_2264_));
 sg13g2_nand4_1 _3042_ (.B(_2344_),
    .C(_2453_),
    .A(_2336_),
    .Y(_2457_),
    .D(_2456_));
 sg13g2_a21oi_1 _3043_ (.A1(_2252_),
    .A2(_2271_),
    .Y(_2458_),
    .B1(_2261_));
 sg13g2_a21oi_1 _3044_ (.A1(_2255_),
    .A2(_2458_),
    .Y(_2459_),
    .B1(_2457_));
 sg13g2_a21o_1 _3045_ (.A2(_2457_),
    .A1(net332),
    .B1(_2459_),
    .X(_0063_));
 sg13g2_a21oi_1 _3046_ (.A1(_2252_),
    .A2(_2271_),
    .Y(_2460_),
    .B1(_2260_));
 sg13g2_o21ai_1 _3047_ (.B1(_2268_),
    .Y(_0064_),
    .A1(_2457_),
    .A2(_2460_));
 sg13g2_nand2_2 _3048_ (.Y(_2461_),
    .A(net332),
    .B(_2267_));
 sg13g2_o21ai_1 _3049_ (.B1(_2461_),
    .Y(_2462_),
    .A1(_2258_),
    .A2(_2259_));
 sg13g2_a21oi_1 _3050_ (.A1(_2251_),
    .A2(_2271_),
    .Y(_2463_),
    .B1(_2462_));
 sg13g2_nand2_1 _3051_ (.Y(_2464_),
    .A(_2255_),
    .B(_2463_));
 sg13g2_mux2_1 _3052_ (.A0(_2464_),
    .A1(net298),
    .S(_2457_),
    .X(_0065_));
 sg13g2_nand2_2 _3053_ (.Y(_2465_),
    .A(net380),
    .B(_2263_));
 sg13g2_mux2_1 _3054_ (.A0(net1),
    .A1(net740),
    .S(_2465_),
    .X(_0066_));
 sg13g2_mux2_1 _3055_ (.A0(net2),
    .A1(net317),
    .S(_2465_),
    .X(_0067_));
 sg13g2_mux2_1 _3056_ (.A0(net3),
    .A1(net320),
    .S(_2465_),
    .X(_0068_));
 sg13g2_mux2_1 _3057_ (.A0(net4),
    .A1(net138),
    .S(_2465_),
    .X(_0069_));
 sg13g2_mux2_1 _3058_ (.A0(net5),
    .A1(net258),
    .S(_2465_),
    .X(_0070_));
 sg13g2_mux2_1 _3059_ (.A0(net6),
    .A1(net271),
    .S(_2465_),
    .X(_0071_));
 sg13g2_mux2_1 _3060_ (.A0(net7),
    .A1(net176),
    .S(_2465_),
    .X(_0072_));
 sg13g2_mux2_1 _3061_ (.A0(net8),
    .A1(net217),
    .S(_2465_),
    .X(_0073_));
 sg13g2_nand2_2 _3062_ (.Y(_2466_),
    .A(_2260_),
    .B(_2263_));
 sg13g2_nor2_1 _3063_ (.A(net1),
    .B(net551),
    .Y(_2467_));
 sg13g2_a21oi_1 _3064_ (.A1(_2218_),
    .A2(net551),
    .Y(_0074_),
    .B1(_2467_));
 sg13g2_nor2_1 _3065_ (.A(net2),
    .B(net552),
    .Y(_2468_));
 sg13g2_a21oi_1 _3066_ (.A1(_2219_),
    .A2(net551),
    .Y(_0075_),
    .B1(_2468_));
 sg13g2_mux2_1 _3067_ (.A0(net3),
    .A1(net728),
    .S(net552),
    .X(_0076_));
 sg13g2_nor2_1 _3068_ (.A(net4),
    .B(net551),
    .Y(_2469_));
 sg13g2_a21oi_1 _3069_ (.A1(_2220_),
    .A2(net551),
    .Y(_0077_),
    .B1(_2469_));
 sg13g2_nor2_1 _3070_ (.A(net5),
    .B(net552),
    .Y(_2470_));
 sg13g2_a21oi_1 _3071_ (.A1(_2221_),
    .A2(net551),
    .Y(_0078_),
    .B1(_2470_));
 sg13g2_mux2_1 _3072_ (.A0(net6),
    .A1(net718),
    .S(net552),
    .X(_0079_));
 sg13g2_mux2_1 _3073_ (.A0(net7),
    .A1(net712),
    .S(net552),
    .X(_0080_));
 sg13g2_nor2_1 _3074_ (.A(net8),
    .B(net551),
    .Y(_2471_));
 sg13g2_a21oi_1 _3075_ (.A1(_2224_),
    .A2(net551),
    .Y(_0081_),
    .B1(_2471_));
 sg13g2_nor2_2 _3076_ (.A(_2266_),
    .B(_2461_),
    .Y(_2472_));
 sg13g2_nand2_1 _3077_ (.Y(_2473_),
    .A(net1),
    .B(net577));
 sg13g2_o21ai_1 _3078_ (.B1(_2473_),
    .Y(_0082_),
    .A1(_2232_),
    .A2(net577));
 sg13g2_mux2_1 _3079_ (.A0(net703),
    .A1(net2),
    .S(_2472_),
    .X(_0083_));
 sg13g2_mux2_1 _3080_ (.A0(net700),
    .A1(net3),
    .S(net577),
    .X(_0084_));
 sg13g2_mux2_1 _3081_ (.A0(net697),
    .A1(net4),
    .S(net577),
    .X(_0085_));
 sg13g2_mux2_1 _3082_ (.A0(net693),
    .A1(net5),
    .S(_2472_),
    .X(_0086_));
 sg13g2_mux2_1 _3083_ (.A0(net690),
    .A1(net6),
    .S(net577),
    .X(_0087_));
 sg13g2_mux2_1 _3084_ (.A0(net688),
    .A1(net7),
    .S(net577),
    .X(_0088_));
 sg13g2_nand2_1 _3085_ (.Y(_2474_),
    .A(net8),
    .B(net577));
 sg13g2_o21ai_1 _3086_ (.B1(_2474_),
    .Y(_0089_),
    .A1(_2233_),
    .A2(net577));
 sg13g2_nor3_1 _3087_ (.A(_2254_),
    .B(_2313_),
    .C(_2329_),
    .Y(_2475_));
 sg13g2_mux2_1 _3088_ (.A0(net256),
    .A1(\cordic_inst.cordic_state[23] ),
    .S(net548),
    .X(_0090_));
 sg13g2_mux2_1 _3089_ (.A0(net236),
    .A1(\cordic_inst.cordic_state[24] ),
    .S(net548),
    .X(_0091_));
 sg13g2_mux2_1 _3090_ (.A0(net221),
    .A1(\cordic_inst.cordic_state[25] ),
    .S(net549),
    .X(_0092_));
 sg13g2_mux2_1 _3091_ (.A0(net182),
    .A1(\cordic_inst.cordic_state[26] ),
    .S(net548),
    .X(_0093_));
 sg13g2_mux2_1 _3092_ (.A0(net213),
    .A1(\cordic_inst.cordic_state[27] ),
    .S(net550),
    .X(_0094_));
 sg13g2_mux2_1 _3093_ (.A0(net172),
    .A1(\cordic_inst.cordic_state[28] ),
    .S(net549),
    .X(_0095_));
 sg13g2_mux2_1 _3094_ (.A0(net240),
    .A1(\cordic_inst.cordic_state[29] ),
    .S(net548),
    .X(_0096_));
 sg13g2_mux2_1 _3095_ (.A0(net188),
    .A1(\cordic_inst.cordic_state[30] ),
    .S(net550),
    .X(_0097_));
 sg13g2_nor2_1 _3096_ (.A(net147),
    .B(net550),
    .Y(_2476_));
 sg13g2_a21oi_1 _3097_ (.A1(_2208_),
    .A2(net550),
    .Y(_0098_),
    .B1(net148));
 sg13g2_mux2_1 _3098_ (.A0(net190),
    .A1(\cordic_inst.cordic_state[32] ),
    .S(net549),
    .X(_0099_));
 sg13g2_mux2_1 _3099_ (.A0(net192),
    .A1(\cordic_inst.cordic_state[33] ),
    .S(net548),
    .X(_0100_));
 sg13g2_mux2_1 _3100_ (.A0(net226),
    .A1(\cordic_inst.cordic_state[34] ),
    .S(net548),
    .X(_0101_));
 sg13g2_nor2_1 _3101_ (.A(net161),
    .B(net550),
    .Y(_2477_));
 sg13g2_a21oi_1 _3102_ (.A1(_2207_),
    .A2(net550),
    .Y(_0102_),
    .B1(net162));
 sg13g2_mux2_1 _3103_ (.A0(net207),
    .A1(\cordic_inst.cordic_state[36] ),
    .S(net548),
    .X(_0103_));
 sg13g2_mux2_1 _3104_ (.A0(net200),
    .A1(\cordic_inst.cordic_state[37] ),
    .S(net548),
    .X(_0104_));
 sg13g2_mux2_1 _3105_ (.A0(net170),
    .A1(\cordic_inst.cordic_state[38] ),
    .S(net550),
    .X(_0105_));
 sg13g2_nand2b_1 _3106_ (.Y(_2478_),
    .B(net304),
    .A_N(net684));
 sg13g2_nand3_1 _3107_ (.B(_2281_),
    .C(_2478_),
    .A(net775),
    .Y(_0106_));
 sg13g2_o21ai_1 _3108_ (.B1(net600),
    .Y(_2479_),
    .A1(_2212_),
    .A2(_2307_));
 sg13g2_and2_1 _3109_ (.A(net783),
    .B(_2479_),
    .X(_0107_));
 sg13g2_nor2_1 _3110_ (.A(net296),
    .B(_2307_),
    .Y(_2480_));
 sg13g2_nor2_1 _3111_ (.A(_2285_),
    .B(net297),
    .Y(_0108_));
 sg13g2_and2_1 _3112_ (.A(_2281_),
    .B(net589),
    .X(_2481_));
 sg13g2_nand2_1 _3113_ (.Y(_2482_),
    .A(\cordic_atan2_result[0] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ));
 sg13g2_xnor2_1 _3114_ (.Y(_2483_),
    .A(net328),
    .B(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ));
 sg13g2_a22oi_1 _3115_ (.Y(_2484_),
    .B1(net591),
    .B2(_2483_),
    .A2(_2218_),
    .A1(net685));
 sg13g2_a22oi_1 _3116_ (.Y(_2485_),
    .B1(net576),
    .B2(_2484_),
    .A2(net583),
    .A1(net328));
 sg13g2_nand2_1 _3117_ (.Y(_0113_),
    .A(net792),
    .B(net329));
 sg13g2_nand2_1 _3118_ (.Y(_2486_),
    .A(\cordic_atan2_result[15] ),
    .B(_2213_));
 sg13g2_nor4_1 _3119_ (.A(net650),
    .B(net651),
    .C(\cordic_inst.cordic_state[31] ),
    .D(\cordic_inst.cordic_state[30] ),
    .Y(_2487_));
 sg13g2_nor4_1 _3120_ (.A(\cordic_inst.cordic_state[37] ),
    .B(\cordic_inst.cordic_state[36] ),
    .C(\cordic_inst.cordic_state[35] ),
    .D(net649),
    .Y(_2488_));
 sg13g2_nor4_1 _3121_ (.A(\cordic_inst.cordic_state[29] ),
    .B(\cordic_inst.cordic_state[28] ),
    .C(\cordic_inst.cordic_state[27] ),
    .D(\cordic_inst.cordic_state[26] ),
    .Y(_2489_));
 sg13g2_nor3_1 _3122_ (.A(\cordic_inst.cordic_state[25] ),
    .B(\cordic_inst.cordic_state[24] ),
    .C(\cordic_inst.cordic_state[23] ),
    .Y(_2490_));
 sg13g2_and3_2 _3123_ (.X(_2491_),
    .A(_2487_),
    .B(_2488_),
    .C(_2490_));
 sg13g2_nand2b_1 _3124_ (.Y(_2492_),
    .B(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .A_N(net648));
 sg13g2_a21oi_1 _3125_ (.A1(_2489_),
    .A2(_2491_),
    .Y(_2493_),
    .B1(_2492_));
 sg13g2_a21o_1 _3126_ (.A2(_2491_),
    .A1(_2489_),
    .B1(_2492_),
    .X(_2494_));
 sg13g2_and2_1 _3127_ (.A(_2486_),
    .B(_2494_),
    .X(_2495_));
 sg13g2_nand2_1 _3128_ (.Y(_2496_),
    .A(_2486_),
    .B(_2494_));
 sg13g2_nand3_1 _3129_ (.B(_2486_),
    .C(_2494_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ),
    .Y(_2497_));
 sg13g2_xnor2_1 _3130_ (.Y(_2498_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[1] ),
    .B(_2497_));
 sg13g2_nand2_1 _3131_ (.Y(_2499_),
    .A(\cordic_atan2_result[1] ),
    .B(_2498_));
 sg13g2_xnor2_1 _3132_ (.Y(_2500_),
    .A(\cordic_atan2_result[1] ),
    .B(_2498_));
 sg13g2_or2_1 _3133_ (.X(_2501_),
    .B(_2500_),
    .A(_2482_));
 sg13g2_a21oi_1 _3134_ (.A1(_2482_),
    .A2(_2500_),
    .Y(_2502_),
    .B1(_2290_));
 sg13g2_a22oi_1 _3135_ (.Y(_2503_),
    .B1(_2501_),
    .B2(_2502_),
    .A2(net734),
    .A1(net685));
 sg13g2_inv_1 _3136_ (.Y(_2504_),
    .A(_2503_));
 sg13g2_a22oi_1 _3137_ (.Y(_2505_),
    .B1(net576),
    .B2(_2504_),
    .A2(net583),
    .A1(net302));
 sg13g2_nor2_1 _3138_ (.A(net769),
    .B(net303),
    .Y(_0114_));
 sg13g2_or2_1 _3139_ (.X(_2506_),
    .B(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[1] ),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ));
 sg13g2_a21o_2 _3140_ (.A2(_2506_),
    .A1(net562),
    .B1(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[2] ),
    .X(_2507_));
 sg13g2_nand3_1 _3141_ (.B(net562),
    .C(_2506_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[2] ),
    .Y(_2508_));
 sg13g2_and2_1 _3142_ (.A(_2507_),
    .B(_2508_),
    .X(_2509_));
 sg13g2_xnor2_1 _3143_ (.Y(_2510_),
    .A(\cordic_atan2_result[2] ),
    .B(_2509_));
 sg13g2_a21oi_1 _3144_ (.A1(_2499_),
    .A2(_2501_),
    .Y(_2511_),
    .B1(_2510_));
 sg13g2_nand3_1 _3145_ (.B(_2501_),
    .C(_2510_),
    .A(_2499_),
    .Y(_2512_));
 sg13g2_nand2b_1 _3146_ (.Y(_2513_),
    .B(_2512_),
    .A_N(_2511_));
 sg13g2_and2_1 _3147_ (.A(net684),
    .B(_2281_),
    .X(_2514_));
 sg13g2_nand2_1 _3148_ (.Y(_2515_),
    .A(net728),
    .B(_2514_));
 sg13g2_a22oi_1 _3149_ (.Y(_2516_),
    .B1(_2515_),
    .B2(_2293_),
    .A2(_2513_),
    .A1(net590));
 sg13g2_a21oi_1 _3150_ (.A1(net330),
    .A2(net582),
    .Y(_2517_),
    .B1(_2516_));
 sg13g2_nand2_1 _3151_ (.Y(_0115_),
    .A(net783),
    .B(_2517_));
 sg13g2_a21o_1 _3152_ (.A2(_2509_),
    .A1(\cordic_atan2_result[2] ),
    .B1(_2511_),
    .X(_2518_));
 sg13g2_nand2_1 _3153_ (.Y(_2519_),
    .A(net562),
    .B(_2507_));
 sg13g2_xor2_1 _3154_ (.B(_2519_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[3] ),
    .X(_2520_));
 sg13g2_nor2b_1 _3155_ (.A(_2520_),
    .B_N(\cordic_atan2_result[3] ),
    .Y(_2521_));
 sg13g2_xnor2_1 _3156_ (.Y(_2522_),
    .A(\cordic_atan2_result[3] ),
    .B(_2520_));
 sg13g2_o21ai_1 _3157_ (.B1(net590),
    .Y(_2523_),
    .A1(_2518_),
    .A2(_2522_));
 sg13g2_a21oi_1 _3158_ (.A1(_2518_),
    .A2(_2522_),
    .Y(_2524_),
    .B1(_2523_));
 sg13g2_a21o_1 _3159_ (.A2(net723),
    .A1(net684),
    .B1(_2524_),
    .X(_2525_));
 sg13g2_a22oi_1 _3160_ (.Y(_2526_),
    .B1(net576),
    .B2(_2525_),
    .A2(net578),
    .A1(net309));
 sg13g2_nor2_1 _3161_ (.A(net770),
    .B(_2526_),
    .Y(_0116_));
 sg13g2_a21oi_1 _3162_ (.A1(_2518_),
    .A2(_2522_),
    .Y(_2527_),
    .B1(_2521_));
 sg13g2_o21ai_1 _3163_ (.B1(net562),
    .Y(_2528_),
    .A1(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[3] ),
    .A2(_2507_));
 sg13g2_xnor2_1 _3164_ (.Y(_2529_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[4] ),
    .B(_2528_));
 sg13g2_xor2_1 _3165_ (.B(_2529_),
    .A(net334),
    .X(_2530_));
 sg13g2_nor2b_1 _3166_ (.A(_2527_),
    .B_N(_2530_),
    .Y(_2531_));
 sg13g2_xnor2_1 _3167_ (.Y(_2532_),
    .A(_2527_),
    .B(_2530_));
 sg13g2_nor2_1 _3168_ (.A(_2290_),
    .B(_2532_),
    .Y(_2533_));
 sg13g2_a21oi_1 _3169_ (.A1(net719),
    .A2(_2514_),
    .Y(_2534_),
    .B1(_2292_));
 sg13g2_a21oi_1 _3170_ (.A1(net334),
    .A2(net582),
    .Y(_2535_),
    .B1(net769));
 sg13g2_o21ai_1 _3171_ (.B1(_2535_),
    .Y(_0117_),
    .A1(_2533_),
    .A2(_2534_));
 sg13g2_a21oi_1 _3172_ (.A1(\cordic_atan2_result[4] ),
    .A2(_2529_),
    .Y(_2536_),
    .B1(_2531_));
 sg13g2_nor3_1 _3173_ (.A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[3] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[4] ),
    .C(_2507_),
    .Y(_2537_));
 sg13g2_nor2_1 _3174_ (.A(net558),
    .B(_2537_),
    .Y(_2538_));
 sg13g2_xnor2_1 _3175_ (.Y(_2539_),
    .A(_2222_),
    .B(_2538_));
 sg13g2_nand2_1 _3176_ (.Y(_2540_),
    .A(\cordic_atan2_result[5] ),
    .B(_2539_));
 sg13g2_xnor2_1 _3177_ (.Y(_2541_),
    .A(\cordic_atan2_result[5] ),
    .B(_2539_));
 sg13g2_o21ai_1 _3178_ (.B1(net590),
    .Y(_2542_),
    .A1(_2536_),
    .A2(_2541_));
 sg13g2_a21oi_1 _3179_ (.A1(_2536_),
    .A2(_2541_),
    .Y(_2543_),
    .B1(_2542_));
 sg13g2_a21o_1 _3180_ (.A2(net718),
    .A1(net684),
    .B1(_2543_),
    .X(_2544_));
 sg13g2_a22oi_1 _3181_ (.Y(_2545_),
    .B1(net576),
    .B2(_2544_),
    .A2(net578),
    .A1(net326));
 sg13g2_nor2_1 _3182_ (.A(net770),
    .B(_2545_),
    .Y(_0118_));
 sg13g2_o21ai_1 _3183_ (.B1(_2540_),
    .Y(_2546_),
    .A1(_2536_),
    .A2(_2541_));
 sg13g2_a21oi_1 _3184_ (.A1(_2222_),
    .A2(_2537_),
    .Y(_2547_),
    .B1(net558));
 sg13g2_xnor2_1 _3185_ (.Y(_2548_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[6] ),
    .B(_2547_));
 sg13g2_or2_1 _3186_ (.X(_2549_),
    .B(_2548_),
    .A(_2209_));
 sg13g2_xnor2_1 _3187_ (.Y(_2550_),
    .A(_2209_),
    .B(_2548_));
 sg13g2_nand2b_1 _3188_ (.Y(_2551_),
    .B(_2546_),
    .A_N(_2550_));
 sg13g2_xor2_1 _3189_ (.B(_2550_),
    .A(_2546_),
    .X(_2552_));
 sg13g2_nand2_1 _3190_ (.Y(_2553_),
    .A(net712),
    .B(_2514_));
 sg13g2_a22oi_1 _3191_ (.Y(_2554_),
    .B1(_2553_),
    .B2(_2293_),
    .A2(_2552_),
    .A1(net590));
 sg13g2_a21oi_1 _3192_ (.A1(net327),
    .A2(net578),
    .Y(_2555_),
    .B1(_2554_));
 sg13g2_nand2_1 _3193_ (.Y(_0119_),
    .A(net783),
    .B(_2555_));
 sg13g2_a21oi_1 _3194_ (.A1(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[6] ),
    .A2(net562),
    .Y(_2556_),
    .B1(_2547_));
 sg13g2_xnor2_1 _3195_ (.Y(_2557_),
    .A(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[7] ),
    .B(_2556_));
 sg13g2_nand2_1 _3196_ (.Y(_2558_),
    .A(\cordic_atan2_result[7] ),
    .B(_2557_));
 sg13g2_xnor2_1 _3197_ (.Y(_2559_),
    .A(\cordic_atan2_result[7] ),
    .B(_2557_));
 sg13g2_nand3_1 _3198_ (.B(_2551_),
    .C(_2559_),
    .A(_2549_),
    .Y(_2560_));
 sg13g2_a21o_1 _3199_ (.A2(_2551_),
    .A1(_2549_),
    .B1(_2559_),
    .X(_2561_));
 sg13g2_and2_1 _3200_ (.A(net590),
    .B(_2560_),
    .X(_2562_));
 sg13g2_a22oi_1 _3201_ (.Y(_2563_),
    .B1(_2561_),
    .B2(_2562_),
    .A2(net711),
    .A1(net684));
 sg13g2_inv_1 _3202_ (.Y(_2564_),
    .A(_2563_));
 sg13g2_a22oi_1 _3203_ (.Y(_2565_),
    .B1(net576),
    .B2(_2564_),
    .A2(net578),
    .A1(net308));
 sg13g2_nor2_1 _3204_ (.A(net770),
    .B(_2565_),
    .Y(_0120_));
 sg13g2_a21oi_1 _3205_ (.A1(_2223_),
    .A2(_2556_),
    .Y(_2566_),
    .B1(net558));
 sg13g2_nand2_1 _3206_ (.Y(_2567_),
    .A(\cordic_atan2_result[8] ),
    .B(net544));
 sg13g2_xnor2_1 _3207_ (.Y(_2568_),
    .A(\cordic_atan2_result[8] ),
    .B(net544));
 sg13g2_a21o_2 _3208_ (.A2(_2561_),
    .A1(_2558_),
    .B1(_2568_),
    .X(_2569_));
 sg13g2_nand3_1 _3209_ (.B(_2561_),
    .C(_2568_),
    .A(_2558_),
    .Y(_2570_));
 sg13g2_nand2_1 _3210_ (.Y(_2571_),
    .A(_2569_),
    .B(_2570_));
 sg13g2_nand2_1 _3211_ (.Y(_2572_),
    .A(net762),
    .B(_2514_));
 sg13g2_a22oi_1 _3212_ (.Y(_2573_),
    .B1(_2572_),
    .B2(_2293_),
    .A2(_2571_),
    .A1(net590));
 sg13g2_a21oi_1 _3213_ (.A1(net337),
    .A2(net582),
    .Y(_2574_),
    .B1(_2573_));
 sg13g2_nand2_1 _3214_ (.Y(_0121_),
    .A(net775),
    .B(net338));
 sg13g2_nand2_1 _3215_ (.Y(_2575_),
    .A(net685),
    .B(net759));
 sg13g2_xnor2_1 _3216_ (.Y(_2576_),
    .A(\cordic_atan2_result[9] ),
    .B(net544));
 sg13g2_a21oi_1 _3217_ (.A1(_2567_),
    .A2(_2569_),
    .Y(_2577_),
    .B1(_2576_));
 sg13g2_nand3_1 _3218_ (.B(_2569_),
    .C(_2576_),
    .A(_2567_),
    .Y(_2578_));
 sg13g2_nand2_1 _3219_ (.Y(_2579_),
    .A(net590),
    .B(_2578_));
 sg13g2_o21ai_1 _3220_ (.B1(_2575_),
    .Y(_2580_),
    .A1(_2577_),
    .A2(_2579_));
 sg13g2_a22oi_1 _3221_ (.Y(_2581_),
    .B1(net576),
    .B2(_2580_),
    .A2(net582),
    .A1(net292));
 sg13g2_nor2_1 _3222_ (.A(net769),
    .B(net293),
    .Y(_0122_));
 sg13g2_o21ai_1 _3223_ (.B1(net544),
    .Y(_2582_),
    .A1(\cordic_atan2_result[9] ),
    .A2(\cordic_atan2_result[8] ));
 sg13g2_o21ai_1 _3224_ (.B1(_2582_),
    .Y(_2583_),
    .A1(_2569_),
    .A2(_2576_));
 sg13g2_xnor2_1 _3225_ (.Y(_2584_),
    .A(\cordic_atan2_result[10] ),
    .B(net542));
 sg13g2_nor2b_1 _3226_ (.A(_2584_),
    .B_N(_2583_),
    .Y(_2585_));
 sg13g2_xnor2_1 _3227_ (.Y(_2586_),
    .A(_2583_),
    .B(_2584_));
 sg13g2_nor2_1 _3228_ (.A(_2290_),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_a21oi_1 _3229_ (.A1(net756),
    .A2(_2514_),
    .Y(_2588_),
    .B1(_2292_));
 sg13g2_a21oi_1 _3230_ (.A1(net339),
    .A2(net581),
    .Y(_2589_),
    .B1(net769));
 sg13g2_o21ai_1 _3231_ (.B1(_2589_),
    .Y(_0123_),
    .A1(_2587_),
    .A2(_2588_));
 sg13g2_a21oi_1 _3232_ (.A1(\cordic_atan2_result[10] ),
    .A2(net542),
    .Y(_2590_),
    .B1(_2585_));
 sg13g2_xnor2_1 _3233_ (.Y(_2591_),
    .A(\cordic_atan2_result[11] ),
    .B(net542));
 sg13g2_o21ai_1 _3234_ (.B1(net591),
    .Y(_2592_),
    .A1(_2590_),
    .A2(_2591_));
 sg13g2_a21oi_1 _3235_ (.A1(_2590_),
    .A2(_2591_),
    .Y(_2593_),
    .B1(_2592_));
 sg13g2_a21o_1 _3236_ (.A2(net753),
    .A1(net685),
    .B1(_2593_),
    .X(_2594_));
 sg13g2_a22oi_1 _3237_ (.Y(_2595_),
    .B1(net576),
    .B2(_2594_),
    .A2(net581),
    .A1(net306));
 sg13g2_nor2_1 _3238_ (.A(net769),
    .B(net307),
    .Y(_0124_));
 sg13g2_or4_1 _3239_ (.A(_2569_),
    .B(_2576_),
    .C(_2584_),
    .D(_2591_),
    .X(_2596_));
 sg13g2_o21ai_1 _3240_ (.B1(net542),
    .Y(_2597_),
    .A1(\cordic_atan2_result[11] ),
    .A2(\cordic_atan2_result[10] ));
 sg13g2_nand3_1 _3241_ (.B(_2596_),
    .C(_2597_),
    .A(_2582_),
    .Y(_2598_));
 sg13g2_xnor2_1 _3242_ (.Y(_2599_),
    .A(\cordic_atan2_result[12] ),
    .B(net543));
 sg13g2_nor2b_1 _3243_ (.A(_2599_),
    .B_N(_2598_),
    .Y(_2600_));
 sg13g2_xor2_1 _3244_ (.B(_2599_),
    .A(_2598_),
    .X(_2601_));
 sg13g2_nand2_1 _3245_ (.Y(_2602_),
    .A(net750),
    .B(_2514_));
 sg13g2_a22oi_1 _3246_ (.Y(_2603_),
    .B1(_2602_),
    .B2(_2293_),
    .A2(_2601_),
    .A1(net591));
 sg13g2_a21oi_1 _3247_ (.A1(net318),
    .A2(net581),
    .Y(_2604_),
    .B1(_2603_));
 sg13g2_nand2_1 _3248_ (.Y(_0125_),
    .A(net787),
    .B(net319));
 sg13g2_a21oi_1 _3249_ (.A1(\cordic_atan2_result[12] ),
    .A2(net543),
    .Y(_2605_),
    .B1(_2600_));
 sg13g2_nand2_1 _3250_ (.Y(_0207_),
    .A(\cordic_atan2_result[13] ),
    .B(net542));
 sg13g2_nor2_1 _3251_ (.A(\cordic_atan2_result[13] ),
    .B(net543),
    .Y(_0208_));
 sg13g2_xnor2_1 _3252_ (.Y(_0209_),
    .A(\cordic_atan2_result[13] ),
    .B(net543));
 sg13g2_o21ai_1 _3253_ (.B1(net591),
    .Y(_0210_),
    .A1(_2605_),
    .A2(_0209_));
 sg13g2_a21oi_1 _3254_ (.A1(_2605_),
    .A2(_0209_),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_a21o_1 _3255_ (.A2(net748),
    .A1(net685),
    .B1(_0211_),
    .X(_0212_));
 sg13g2_a22oi_1 _3256_ (.Y(_0213_),
    .B1(net576),
    .B2(_0212_),
    .A2(net581),
    .A1(net323));
 sg13g2_nor2_1 _3257_ (.A(net772),
    .B(net324),
    .Y(_0126_));
 sg13g2_xnor2_1 _3258_ (.Y(_0214_),
    .A(\cordic_atan2_result[14] ),
    .B(net542));
 sg13g2_and2_1 _3259_ (.A(_2605_),
    .B(_0207_),
    .X(_0215_));
 sg13g2_or2_1 _3260_ (.X(_0216_),
    .B(_0215_),
    .A(_0208_));
 sg13g2_nor2_1 _3261_ (.A(_0214_),
    .B(_0216_),
    .Y(_0217_));
 sg13g2_xnor2_1 _3262_ (.Y(_0218_),
    .A(_0214_),
    .B(_0216_));
 sg13g2_nand2_1 _3263_ (.Y(_0219_),
    .A(net746),
    .B(_2514_));
 sg13g2_a22oi_1 _3264_ (.Y(_0220_),
    .B1(_0219_),
    .B2(_2293_),
    .A2(_0218_),
    .A1(net591));
 sg13g2_a21oi_1 _3265_ (.A1(net321),
    .A2(net581),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_nand2_1 _3266_ (.Y(_0127_),
    .A(net787),
    .B(net322));
 sg13g2_nand2_1 _3267_ (.Y(_0222_),
    .A(cordic_en_sin_cos),
    .B(net744));
 sg13g2_a21oi_1 _3268_ (.A1(\cordic_atan2_result[14] ),
    .A2(net542),
    .Y(_0223_),
    .B1(_0217_));
 sg13g2_xnor2_1 _3269_ (.Y(_0224_),
    .A(\cordic_atan2_result[15] ),
    .B(net542));
 sg13g2_and2_1 _3270_ (.A(_0223_),
    .B(_0224_),
    .X(_0225_));
 sg13g2_o21ai_1 _3271_ (.B1(net591),
    .Y(_0226_),
    .A1(_0223_),
    .A2(_0224_));
 sg13g2_o21ai_1 _3272_ (.B1(_0222_),
    .Y(_0227_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_a22oi_1 _3273_ (.Y(_0228_),
    .B1(_2481_),
    .B2(_0227_),
    .A2(net581),
    .A1(net342));
 sg13g2_nor2_1 _3274_ (.A(net769),
    .B(net343),
    .Y(_0128_));
 sg13g2_nor2_1 _3275_ (.A(\cordic_inst.cordic_state[53] ),
    .B(net666),
    .Y(_0229_));
 sg13g2_nor2b_1 _3276_ (.A(net645),
    .B_N(net667),
    .Y(_0230_));
 sg13g2_mux4_1 _3277_ (.S0(net666),
    .A0(\cordic_inst.cordic_state[51] ),
    .A1(\cordic_inst.cordic_state[52] ),
    .A2(\cordic_inst.cordic_state[53] ),
    .A3(net645),
    .S1(net661),
    .X(_0231_));
 sg13g2_mux4_1 _3278_ (.S0(net668),
    .A0(\cordic_inst.cordic_state[47] ),
    .A1(\cordic_inst.cordic_state[48] ),
    .A2(\cordic_inst.cordic_state[49] ),
    .A3(\cordic_inst.cordic_state[50] ),
    .S1(net661),
    .X(_0232_));
 sg13g2_mux2_1 _3279_ (.A0(_0232_),
    .A1(_0231_),
    .S(net656),
    .X(_0233_));
 sg13g2_nand2_1 _3280_ (.Y(_0234_),
    .A(net653),
    .B(_0233_));
 sg13g2_nor2_1 _3281_ (.A(net652),
    .B(net657),
    .Y(_0235_));
 sg13g2_or2_1 _3282_ (.X(_0236_),
    .B(net655),
    .A(net652));
 sg13g2_nor2_2 _3283_ (.A(net606),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_mux2_1 _3284_ (.A0(\cordic_inst.cordic_state[41] ),
    .A1(\cordic_inst.cordic_state[42] ),
    .S(net668),
    .X(_0238_));
 sg13g2_nor3_2 _3285_ (.A(net654),
    .B(net657),
    .C(net660),
    .Y(_0239_));
 sg13g2_nand2_1 _3286_ (.Y(_0240_),
    .A(net605),
    .B(net597));
 sg13g2_mux2_1 _3287_ (.A0(\cordic_inst.cordic_state[39] ),
    .A1(\cordic_inst.cordic_state[40] ),
    .S(net668),
    .X(_0241_));
 sg13g2_and2_1 _3288_ (.A(_0239_),
    .B(_0241_),
    .X(_0242_));
 sg13g2_nor2b_2 _3289_ (.A(net652),
    .B_N(net657),
    .Y(_0243_));
 sg13g2_mux2_1 _3290_ (.A0(\cordic_inst.cordic_state[45] ),
    .A1(\cordic_inst.cordic_state[46] ),
    .S(net668),
    .X(_0244_));
 sg13g2_mux2_1 _3291_ (.A0(\cordic_inst.cordic_state[43] ),
    .A1(\cordic_inst.cordic_state[44] ),
    .S(net668),
    .X(_0245_));
 sg13g2_mux2_1 _3292_ (.A0(_0244_),
    .A1(_0245_),
    .S(net606),
    .X(_0246_));
 sg13g2_a221oi_1 _3293_ (.B2(_0246_),
    .C1(_0242_),
    .B1(net596),
    .A1(_0237_),
    .Y(_0247_),
    .A2(_0238_));
 sg13g2_and2_1 _3294_ (.A(_0234_),
    .B(_0247_),
    .X(_0248_));
 sg13g2_nor2_1 _3295_ (.A(net355),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_a21oi_1 _3296_ (.A1(\cordic_inst.cordic_state[23] ),
    .A2(_0248_),
    .Y(_0250_),
    .B1(_2288_));
 sg13g2_nor2b_1 _3297_ (.A(_0249_),
    .B_N(_0250_),
    .Y(_0251_));
 sg13g2_a22oi_1 _3298_ (.Y(_0252_),
    .B1(net602),
    .B2(net738),
    .A2(net640),
    .A1(net680));
 sg13g2_o21ai_1 _3299_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_2284_),
    .A2(_0251_));
 sg13g2_o21ai_1 _3300_ (.B1(_0253_),
    .Y(_0254_),
    .A1(net355),
    .A2(net585));
 sg13g2_nand2_1 _3301_ (.Y(_0129_),
    .A(net774),
    .B(_0254_));
 sg13g2_mux2_1 _3302_ (.A0(\cordic_inst.cordic_state[50] ),
    .A1(\cordic_inst.cordic_state[51] ),
    .S(net666),
    .X(_0255_));
 sg13g2_mux2_1 _3303_ (.A0(\cordic_inst.cordic_state[48] ),
    .A1(\cordic_inst.cordic_state[49] ),
    .S(net666),
    .X(_0256_));
 sg13g2_mux4_1 _3304_ (.S0(net666),
    .A0(\cordic_inst.cordic_state[48] ),
    .A1(\cordic_inst.cordic_state[49] ),
    .A2(\cordic_inst.cordic_state[50] ),
    .A3(\cordic_inst.cordic_state[51] ),
    .S1(net661),
    .X(_0257_));
 sg13g2_mux2_1 _3305_ (.A0(\cordic_inst.cordic_state[52] ),
    .A1(\cordic_inst.cordic_state[53] ),
    .S(net666),
    .X(_0258_));
 sg13g2_nor2b_1 _3306_ (.A(net664),
    .B_N(net659),
    .Y(_0259_));
 sg13g2_a22oi_1 _3307_ (.Y(_0260_),
    .B1(_0259_),
    .B2(net643),
    .A2(_0258_),
    .A1(net605));
 sg13g2_nor2_1 _3308_ (.A(net656),
    .B(_0257_),
    .Y(_0261_));
 sg13g2_a21oi_1 _3309_ (.A1(net656),
    .A2(_0260_),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_mux2_1 _3310_ (.A0(\cordic_inst.cordic_state[46] ),
    .A1(\cordic_inst.cordic_state[47] ),
    .S(net667),
    .X(_0263_));
 sg13g2_nor2_1 _3311_ (.A(\cordic_inst.cordic_state[44] ),
    .B(net666),
    .Y(_0264_));
 sg13g2_a21oi_1 _3312_ (.A1(_2205_),
    .A2(net667),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_mux2_1 _3313_ (.A0(_0263_),
    .A1(_0265_),
    .S(net606),
    .X(_0266_));
 sg13g2_mux2_1 _3314_ (.A0(\cordic_inst.cordic_state[40] ),
    .A1(\cordic_inst.cordic_state[41] ),
    .S(net668),
    .X(_0267_));
 sg13g2_nand2_1 _3315_ (.Y(_0268_),
    .A(_0239_),
    .B(_0267_));
 sg13g2_and2_1 _3316_ (.A(net644),
    .B(net653),
    .X(_0269_));
 sg13g2_nand2b_1 _3317_ (.Y(_0270_),
    .B(_0269_),
    .A_N(_2296_));
 sg13g2_mux2_1 _3318_ (.A0(\cordic_inst.cordic_state[42] ),
    .A1(\cordic_inst.cordic_state[43] ),
    .S(net668),
    .X(_0271_));
 sg13g2_nand3_1 _3319_ (.B(net598),
    .C(_0271_),
    .A(net661),
    .Y(_0272_));
 sg13g2_nand3_1 _3320_ (.B(_0270_),
    .C(_0272_),
    .A(_0268_),
    .Y(_0273_));
 sg13g2_a221oi_1 _3321_ (.B2(net596),
    .C1(_0273_),
    .B1(_0266_),
    .A1(net652),
    .Y(_0274_),
    .A2(_0262_));
 sg13g2_a221oi_1 _3322_ (.B2(_0247_),
    .C1(_2493_),
    .B1(_0234_),
    .A1(\cordic_atan2_result[15] ),
    .Y(_0275_),
    .A2(_2213_));
 sg13g2_xor2_1 _3323_ (.B(_0275_),
    .A(_0274_),
    .X(_0276_));
 sg13g2_nand2_1 _3324_ (.Y(_0277_),
    .A(\cordic_inst.cordic_state[24] ),
    .B(_0276_));
 sg13g2_xor2_1 _3325_ (.B(_0276_),
    .A(net364),
    .X(_0278_));
 sg13g2_nand2b_1 _3326_ (.Y(_0279_),
    .B(_0249_),
    .A_N(_0278_));
 sg13g2_nand2b_1 _3327_ (.Y(_0280_),
    .B(_0278_),
    .A_N(_0249_));
 sg13g2_nand3_1 _3328_ (.B(_0279_),
    .C(_0280_),
    .A(_2292_),
    .Y(_0281_));
 sg13g2_a221oi_1 _3329_ (.B2(net734),
    .C1(net582),
    .B1(net602),
    .A1(net681),
    .Y(_0282_),
    .A2(net636));
 sg13g2_o21ai_1 _3330_ (.B1(net774),
    .Y(_0283_),
    .A1(net364),
    .A2(net586));
 sg13g2_a21oi_1 _3331_ (.A1(_0281_),
    .A2(_0282_),
    .Y(_0130_),
    .B1(_0283_));
 sg13g2_mux4_1 _3332_ (.S0(net666),
    .A0(\cordic_inst.cordic_state[49] ),
    .A1(\cordic_inst.cordic_state[50] ),
    .A2(\cordic_inst.cordic_state[51] ),
    .A3(\cordic_inst.cordic_state[52] ),
    .S1(net661),
    .X(_0284_));
 sg13g2_nor3_1 _3333_ (.A(net661),
    .B(_0229_),
    .C(_0230_),
    .Y(_0285_));
 sg13g2_mux2_1 _3334_ (.A0(_0284_),
    .A1(_0285_),
    .S(net656),
    .X(_0286_));
 sg13g2_mux4_1 _3335_ (.S0(net669),
    .A0(\cordic_inst.cordic_state[45] ),
    .A1(\cordic_inst.cordic_state[46] ),
    .A2(\cordic_inst.cordic_state[47] ),
    .A3(\cordic_inst.cordic_state[48] ),
    .S1(net661),
    .X(_0287_));
 sg13g2_nand3_1 _3336_ (.B(net598),
    .C(_0245_),
    .A(net661),
    .Y(_0288_));
 sg13g2_a22oi_1 _3337_ (.Y(_0289_),
    .B1(net596),
    .B2(_0287_),
    .A2(_0239_),
    .A1(_0238_));
 sg13g2_nand3_1 _3338_ (.B(_0288_),
    .C(_0289_),
    .A(_0270_),
    .Y(_0290_));
 sg13g2_a21oi_2 _3339_ (.B1(_0290_),
    .Y(_0291_),
    .A2(_0286_),
    .A1(net653));
 sg13g2_a21oi_1 _3340_ (.A1(_0248_),
    .A2(_0274_),
    .Y(_0292_),
    .B1(net558));
 sg13g2_xor2_1 _3341_ (.B(_0292_),
    .A(_0291_),
    .X(_0293_));
 sg13g2_nand2_1 _3342_ (.Y(_0294_),
    .A(\cordic_inst.cordic_state[25] ),
    .B(_0293_));
 sg13g2_xnor2_1 _3343_ (.Y(_0295_),
    .A(\cordic_inst.cordic_state[25] ),
    .B(_0293_));
 sg13g2_and3_1 _3344_ (.X(_0296_),
    .A(_0277_),
    .B(_0280_),
    .C(_0295_));
 sg13g2_a21o_1 _3345_ (.A2(_0280_),
    .A1(_0277_),
    .B1(_0295_),
    .X(_0297_));
 sg13g2_nand2_1 _3346_ (.Y(_0298_),
    .A(net600),
    .B(_0297_));
 sg13g2_a221oi_1 _3347_ (.B2(net728),
    .C1(net582),
    .B1(net603),
    .A1(net681),
    .Y(_0299_),
    .A2(net633));
 sg13g2_o21ai_1 _3348_ (.B1(_0299_),
    .Y(_0300_),
    .A1(_0296_),
    .A2(_0298_));
 sg13g2_o21ai_1 _3349_ (.B1(_0300_),
    .Y(_0301_),
    .A1(net392),
    .A2(net586));
 sg13g2_nand2_1 _3350_ (.Y(_0131_),
    .A(net776),
    .B(_0301_));
 sg13g2_nor2_1 _3351_ (.A(_2216_),
    .B(net629),
    .Y(_0302_));
 sg13g2_mux2_1 _3352_ (.A0(_0255_),
    .A1(_0258_),
    .S(\cordic_inst.cordic_state[4] ),
    .X(_0303_));
 sg13g2_inv_1 _3353_ (.Y(_0304_),
    .A(_0303_));
 sg13g2_nand3_1 _3354_ (.B(net656),
    .C(_2359_),
    .A(net644),
    .Y(_0305_));
 sg13g2_o21ai_1 _3355_ (.B1(_0305_),
    .Y(_0306_),
    .A1(net657),
    .A2(_0304_));
 sg13g2_mux2_1 _3356_ (.A0(_0256_),
    .A1(_0263_),
    .S(net606),
    .X(_0307_));
 sg13g2_a22oi_1 _3357_ (.Y(_0308_),
    .B1(_0271_),
    .B2(_0239_),
    .A2(_0265_),
    .A1(_0237_));
 sg13g2_a22oi_1 _3358_ (.Y(_0309_),
    .B1(net596),
    .B2(_0307_),
    .A2(_2361_),
    .A1(net644));
 sg13g2_nand2_1 _3359_ (.Y(_0310_),
    .A(_0308_),
    .B(_0309_));
 sg13g2_a21oi_1 _3360_ (.A1(net653),
    .A2(_0306_),
    .Y(_0311_),
    .B1(_0310_));
 sg13g2_nand3_1 _3361_ (.B(_0274_),
    .C(_0291_),
    .A(_0248_),
    .Y(_0312_));
 sg13g2_nand2_1 _3362_ (.Y(_0313_),
    .A(net562),
    .B(_0312_));
 sg13g2_xor2_1 _3363_ (.B(_0313_),
    .A(_0311_),
    .X(_0314_));
 sg13g2_inv_1 _3364_ (.Y(_0315_),
    .A(_0314_));
 sg13g2_nand2_1 _3365_ (.Y(_0316_),
    .A(\cordic_inst.cordic_state[26] ),
    .B(_0315_));
 sg13g2_xor2_1 _3366_ (.B(_0314_),
    .A(\cordic_inst.cordic_state[26] ),
    .X(_0317_));
 sg13g2_nand3_1 _3367_ (.B(_0297_),
    .C(_0317_),
    .A(_0294_),
    .Y(_0318_));
 sg13g2_a21o_1 _3368_ (.A2(_0297_),
    .A1(_0294_),
    .B1(_0317_),
    .X(_0319_));
 sg13g2_nor2b_1 _3369_ (.A(net584),
    .B_N(_0318_),
    .Y(_0320_));
 sg13g2_a221oi_1 _3370_ (.B2(_0320_),
    .C1(net676),
    .B1(_0319_),
    .A1(net682),
    .Y(_0321_),
    .A2(net723));
 sg13g2_o21ai_1 _3371_ (.B1(net585),
    .Y(_0322_),
    .A1(_0302_),
    .A2(_0321_));
 sg13g2_o21ai_1 _3372_ (.B1(_0322_),
    .Y(_0323_),
    .A1(net363),
    .A2(net586));
 sg13g2_nor2_1 _3373_ (.A(net770),
    .B(_0323_),
    .Y(_0132_));
 sg13g2_nand2_1 _3374_ (.Y(_0324_),
    .A(_2294_),
    .B(_0269_));
 sg13g2_nor2_2 _3375_ (.A(net608),
    .B(net656),
    .Y(_0325_));
 sg13g2_inv_2 _3376_ (.Y(_0326_),
    .A(_0325_));
 sg13g2_nand2_1 _3377_ (.Y(_0327_),
    .A(_0231_),
    .B(_0325_));
 sg13g2_a22oi_1 _3378_ (.Y(_0328_),
    .B1(_0246_),
    .B2(net598),
    .A2(net596),
    .A1(_0232_));
 sg13g2_nand3_1 _3379_ (.B(_0327_),
    .C(_0328_),
    .A(_0324_),
    .Y(_0329_));
 sg13g2_nand4_1 _3380_ (.B(_0274_),
    .C(_0291_),
    .A(_0248_),
    .Y(_0330_),
    .D(_0311_));
 sg13g2_nand2_1 _3381_ (.Y(_0331_),
    .A(net562),
    .B(_0330_));
 sg13g2_xor2_1 _3382_ (.B(_0331_),
    .A(_0329_),
    .X(_0332_));
 sg13g2_and2_1 _3383_ (.A(\cordic_inst.cordic_state[27] ),
    .B(_0332_),
    .X(_0333_));
 sg13g2_xnor2_1 _3384_ (.Y(_0334_),
    .A(\cordic_inst.cordic_state[27] ),
    .B(_0332_));
 sg13g2_nand3_1 _3385_ (.B(_0319_),
    .C(_0334_),
    .A(_0316_),
    .Y(_0335_));
 sg13g2_a21oi_1 _3386_ (.A1(_0316_),
    .A2(_0319_),
    .Y(_0336_),
    .B1(_0334_));
 sg13g2_nand2_1 _3387_ (.Y(_0337_),
    .A(_2283_),
    .B(_0335_));
 sg13g2_a221oi_1 _3388_ (.B2(net719),
    .C1(net581),
    .B1(net603),
    .A1(net681),
    .Y(_0338_),
    .A2(net625));
 sg13g2_o21ai_1 _3389_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0336_),
    .A2(_0337_));
 sg13g2_o21ai_1 _3390_ (.B1(_0339_),
    .Y(_0340_),
    .A1(net391),
    .A2(net586));
 sg13g2_nand2_1 _3391_ (.Y(_0133_),
    .A(net774),
    .B(_0340_));
 sg13g2_nor2_1 _3392_ (.A(_0260_),
    .B(_0326_),
    .Y(_0341_));
 sg13g2_a221oi_1 _3393_ (.B2(net598),
    .C1(_0341_),
    .B1(_0266_),
    .A1(net596),
    .Y(_0342_),
    .A2(_0257_));
 sg13g2_nand2_1 _3394_ (.Y(_0343_),
    .A(_0324_),
    .B(_0342_));
 sg13g2_nor2_1 _3395_ (.A(_0329_),
    .B(_0330_),
    .Y(_0344_));
 sg13g2_nor2_1 _3396_ (.A(net558),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_xor2_1 _3397_ (.B(_0345_),
    .A(_0343_),
    .X(_0346_));
 sg13g2_nand2b_1 _3398_ (.Y(_0347_),
    .B(\cordic_inst.cordic_state[28] ),
    .A_N(_0346_));
 sg13g2_xnor2_1 _3399_ (.Y(_0348_),
    .A(\cordic_inst.cordic_state[28] ),
    .B(_0346_));
 sg13g2_o21ai_1 _3400_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0333_),
    .A2(_0336_));
 sg13g2_nor3_1 _3401_ (.A(_0333_),
    .B(_0336_),
    .C(_0348_),
    .Y(_0350_));
 sg13g2_nor2_1 _3402_ (.A(net584),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_a221oi_1 _3403_ (.B2(_0351_),
    .C1(net676),
    .B1(_0349_),
    .A1(net683),
    .Y(_0352_),
    .A2(net718));
 sg13g2_a21oi_1 _3404_ (.A1(net676),
    .A2(_2230_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_nor2_1 _3405_ (.A(_2299_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_o21ai_1 _3406_ (.B1(net774),
    .Y(_0355_),
    .A1(net359),
    .A2(net586));
 sg13g2_nor2_1 _3407_ (.A(_0354_),
    .B(_0355_),
    .Y(_0134_));
 sg13g2_and2_1 _3408_ (.A(_0347_),
    .B(_0349_),
    .X(_0356_));
 sg13g2_o21ai_1 _3409_ (.B1(_2360_),
    .Y(_0357_),
    .A1(net608),
    .A2(_2359_));
 sg13g2_a22oi_1 _3410_ (.Y(_0358_),
    .B1(_0357_),
    .B2(net644),
    .A2(_0325_),
    .A1(_0285_));
 sg13g2_a22oi_1 _3411_ (.Y(_0359_),
    .B1(_0287_),
    .B2(net598),
    .A2(_0284_),
    .A1(net596));
 sg13g2_nand2_1 _3412_ (.Y(_0360_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_nand2_1 _3413_ (.Y(_0361_),
    .A(_0342_),
    .B(_0344_));
 sg13g2_nand2_1 _3414_ (.Y(_0362_),
    .A(net559),
    .B(_0361_));
 sg13g2_xor2_1 _3415_ (.B(_0362_),
    .A(_0360_),
    .X(_0363_));
 sg13g2_nand2_1 _3416_ (.Y(_0364_),
    .A(\cordic_inst.cordic_state[29] ),
    .B(_0363_));
 sg13g2_xnor2_1 _3417_ (.Y(_0365_),
    .A(\cordic_inst.cordic_state[29] ),
    .B(_0363_));
 sg13g2_xnor2_1 _3418_ (.Y(_0366_),
    .A(_0356_),
    .B(_0365_));
 sg13g2_nand2_1 _3419_ (.Y(_0367_),
    .A(_2287_),
    .B(_0366_));
 sg13g2_a221oi_1 _3420_ (.B2(_0367_),
    .C1(net675),
    .B1(_2282_),
    .A1(net682),
    .Y(_0368_),
    .A2(net712));
 sg13g2_o21ai_1 _3421_ (.B1(net588),
    .Y(_0369_),
    .A1(net604),
    .A2(net618));
 sg13g2_a21oi_1 _3422_ (.A1(net372),
    .A2(net580),
    .Y(_0370_),
    .B1(net767));
 sg13g2_o21ai_1 _3423_ (.B1(_0370_),
    .Y(_0135_),
    .A1(_0368_),
    .A2(_0369_));
 sg13g2_o21ai_1 _3424_ (.B1(_0364_),
    .Y(_0371_),
    .A1(_0356_),
    .A2(_0365_));
 sg13g2_a22oi_1 _3425_ (.Y(_0372_),
    .B1(_0307_),
    .B2(net598),
    .A2(_0303_),
    .A1(net596));
 sg13g2_nand2b_1 _3426_ (.Y(_0373_),
    .B(_0372_),
    .A_N(_0269_));
 sg13g2_or2_1 _3427_ (.X(_0374_),
    .B(_0361_),
    .A(_0360_));
 sg13g2_nand2_1 _3428_ (.Y(_0375_),
    .A(net559),
    .B(_0374_));
 sg13g2_xnor2_1 _3429_ (.Y(_0376_),
    .A(_0373_),
    .B(_0375_));
 sg13g2_nand2b_1 _3430_ (.Y(_0377_),
    .B(\cordic_inst.cordic_state[30] ),
    .A_N(_0376_));
 sg13g2_xnor2_1 _3431_ (.Y(_0378_),
    .A(\cordic_inst.cordic_state[30] ),
    .B(_0376_));
 sg13g2_nand2_1 _3432_ (.Y(_0379_),
    .A(_0371_),
    .B(_0378_));
 sg13g2_nor2_1 _3433_ (.A(_0371_),
    .B(_0378_),
    .Y(_0380_));
 sg13g2_nor2_1 _3434_ (.A(net584),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_nand2_1 _3435_ (.Y(_0382_),
    .A(_0379_),
    .B(_0381_));
 sg13g2_a21oi_1 _3436_ (.A1(net682),
    .A2(net711),
    .Y(_0383_),
    .B1(net675));
 sg13g2_nand2_1 _3437_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_o21ai_1 _3438_ (.B1(_0384_),
    .Y(_0385_),
    .A1(net604),
    .A2(net615));
 sg13g2_o21ai_1 _3439_ (.B1(net775),
    .Y(_0386_),
    .A1(net383),
    .A2(net587));
 sg13g2_a21oi_1 _3440_ (.A1(net587),
    .A2(_0385_),
    .Y(_0136_),
    .B1(_0386_));
 sg13g2_or2_1 _3441_ (.X(_0387_),
    .B(_0374_),
    .A(_0373_));
 sg13g2_nand2_1 _3442_ (.Y(_0388_),
    .A(net559),
    .B(_0387_));
 sg13g2_a21oi_1 _3443_ (.A1(net607),
    .A2(_0233_),
    .Y(_0389_),
    .B1(_0269_));
 sg13g2_xnor2_1 _3444_ (.Y(_0390_),
    .A(_0388_),
    .B(_0389_));
 sg13g2_nand2_1 _3445_ (.Y(_0391_),
    .A(\cordic_inst.cordic_state[31] ),
    .B(_0390_));
 sg13g2_xnor2_1 _3446_ (.Y(_0392_),
    .A(\cordic_inst.cordic_state[31] ),
    .B(_0390_));
 sg13g2_nand3_1 _3447_ (.B(_0379_),
    .C(_0392_),
    .A(_0377_),
    .Y(_0393_));
 sg13g2_a21o_1 _3448_ (.A2(_0379_),
    .A1(_0377_),
    .B1(_0392_),
    .X(_0394_));
 sg13g2_nand3_1 _3449_ (.B(_0393_),
    .C(_0394_),
    .A(net599),
    .Y(_0395_));
 sg13g2_a221oi_1 _3450_ (.B2(net762),
    .C1(net580),
    .B1(net601),
    .A1(net677),
    .Y(_0396_),
    .A2(net708));
 sg13g2_a22oi_1 _3451_ (.Y(_0397_),
    .B1(_0395_),
    .B2(_0396_),
    .A2(net578),
    .A1(_2208_));
 sg13g2_nand2b_1 _3452_ (.Y(_0137_),
    .B(net774),
    .A_N(_0397_));
 sg13g2_nor2_1 _3453_ (.A(net604),
    .B(net703),
    .Y(_0398_));
 sg13g2_nand2_1 _3454_ (.Y(_0399_),
    .A(net607),
    .B(_2296_));
 sg13g2_a22oi_1 _3455_ (.Y(_0400_),
    .B1(_0399_),
    .B2(net643),
    .A2(_0262_),
    .A1(net607));
 sg13g2_o21ai_1 _3456_ (.B1(net559),
    .Y(_0401_),
    .A1(_0233_),
    .A2(_0387_));
 sg13g2_xnor2_1 _3457_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_nand2_1 _3458_ (.Y(_0403_),
    .A(net651),
    .B(_0402_));
 sg13g2_xnor2_1 _3459_ (.Y(_0404_),
    .A(net651),
    .B(_0402_));
 sg13g2_nand3_1 _3460_ (.B(_0394_),
    .C(_0404_),
    .A(_0391_),
    .Y(_0405_));
 sg13g2_a21o_1 _3461_ (.A2(_0394_),
    .A1(_0391_),
    .B1(_0404_),
    .X(_0406_));
 sg13g2_nor2b_1 _3462_ (.A(net584),
    .B_N(_0405_),
    .Y(_0407_));
 sg13g2_a221oi_1 _3463_ (.B2(_0407_),
    .C1(net675),
    .B1(_0406_),
    .A1(net682),
    .Y(_0408_),
    .A2(net759));
 sg13g2_o21ai_1 _3464_ (.B1(net585),
    .Y(_0409_),
    .A1(_0398_),
    .A2(_0408_));
 sg13g2_o21ai_1 _3465_ (.B1(_0409_),
    .Y(_0410_),
    .A1(net651),
    .A2(net585));
 sg13g2_nor2_1 _3466_ (.A(net768),
    .B(_0410_),
    .Y(_0138_));
 sg13g2_a22oi_1 _3467_ (.Y(_0411_),
    .B1(_0399_),
    .B2(net643),
    .A2(_0286_),
    .A1(net607));
 sg13g2_nand2_1 _3468_ (.Y(_0412_),
    .A(_0389_),
    .B(_0400_));
 sg13g2_o21ai_1 _3469_ (.B1(net559),
    .Y(_0413_),
    .A1(_0387_),
    .A2(_0412_));
 sg13g2_xnor2_1 _3470_ (.Y(_0414_),
    .A(_0411_),
    .B(_0413_));
 sg13g2_xnor2_1 _3471_ (.Y(_0415_),
    .A(net650),
    .B(_0414_));
 sg13g2_a21oi_1 _3472_ (.A1(_0403_),
    .A2(_0406_),
    .Y(_0416_),
    .B1(_0415_));
 sg13g2_and3_1 _3473_ (.X(_0417_),
    .A(_0403_),
    .B(_0406_),
    .C(_0415_));
 sg13g2_o21ai_1 _3474_ (.B1(_2287_),
    .Y(_0418_),
    .A1(_0416_),
    .A2(_0417_));
 sg13g2_a221oi_1 _3475_ (.B2(_0418_),
    .C1(net675),
    .B1(_2282_),
    .A1(net682),
    .Y(_0419_),
    .A2(net756));
 sg13g2_o21ai_1 _3476_ (.B1(net587),
    .Y(_0420_),
    .A1(net604),
    .A2(net700));
 sg13g2_a21oi_1 _3477_ (.A1(net650),
    .A2(net578),
    .Y(_0421_),
    .B1(net768));
 sg13g2_o21ai_1 _3478_ (.B1(_0421_),
    .Y(_0139_),
    .A1(_0419_),
    .A2(_0420_));
 sg13g2_nor2_1 _3479_ (.A(net604),
    .B(net697),
    .Y(_0422_));
 sg13g2_a21o_1 _3480_ (.A2(_0414_),
    .A1(net650),
    .B1(_0416_),
    .X(_0423_));
 sg13g2_a22oi_1 _3481_ (.Y(_0424_),
    .B1(_0306_),
    .B2(net607),
    .A2(_0236_),
    .A1(net643));
 sg13g2_o21ai_1 _3482_ (.B1(_0413_),
    .Y(_0425_),
    .A1(net557),
    .A2(_0411_));
 sg13g2_xor2_1 _3483_ (.B(_0425_),
    .A(_0424_),
    .X(_0426_));
 sg13g2_nand2_1 _3484_ (.Y(_0427_),
    .A(net649),
    .B(_0426_));
 sg13g2_xor2_1 _3485_ (.B(_0426_),
    .A(net649),
    .X(_0428_));
 sg13g2_nor2_1 _3486_ (.A(_0423_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_nand2_2 _3487_ (.Y(_0430_),
    .A(_0423_),
    .B(_0428_));
 sg13g2_nor2_1 _3488_ (.A(net584),
    .B(_0429_),
    .Y(_0431_));
 sg13g2_a221oi_1 _3489_ (.B2(_0431_),
    .C1(net675),
    .B1(_0430_),
    .A1(net682),
    .Y(_0432_),
    .A2(net753));
 sg13g2_o21ai_1 _3490_ (.B1(net585),
    .Y(_0433_),
    .A1(_0422_),
    .A2(_0432_));
 sg13g2_o21ai_1 _3491_ (.B1(_0433_),
    .Y(_0434_),
    .A1(net649),
    .A2(net585));
 sg13g2_nor2_1 _3492_ (.A(net768),
    .B(_0434_),
    .Y(_0140_));
 sg13g2_mux2_1 _3493_ (.A0(net643),
    .A1(_0231_),
    .S(net597),
    .X(_0435_));
 sg13g2_nor2_1 _3494_ (.A(net557),
    .B(_0424_),
    .Y(_0436_));
 sg13g2_nor2_1 _3495_ (.A(_0425_),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_nand2b_1 _3496_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0435_));
 sg13g2_xor2_1 _3497_ (.B(_0437_),
    .A(_0435_),
    .X(_0439_));
 sg13g2_and2_1 _3498_ (.A(\cordic_inst.cordic_state[35] ),
    .B(_0439_),
    .X(_0440_));
 sg13g2_xnor2_1 _3499_ (.Y(_0441_),
    .A(\cordic_inst.cordic_state[35] ),
    .B(_0439_));
 sg13g2_nand3_1 _3500_ (.B(_0430_),
    .C(_0441_),
    .A(_0427_),
    .Y(_0442_));
 sg13g2_a21o_1 _3501_ (.A2(_0430_),
    .A1(_0427_),
    .B1(_0441_),
    .X(_0443_));
 sg13g2_nand3_1 _3502_ (.B(_0442_),
    .C(_0443_),
    .A(net599),
    .Y(_0444_));
 sg13g2_a221oi_1 _3503_ (.B2(net750),
    .C1(net580),
    .B1(net601),
    .A1(net677),
    .Y(_0445_),
    .A2(net693));
 sg13g2_a22oi_1 _3504_ (.Y(_0446_),
    .B1(_0444_),
    .B2(_0445_),
    .A2(net578),
    .A1(_2207_));
 sg13g2_nand2b_1 _3505_ (.Y(_0141_),
    .B(net774),
    .A_N(_0446_));
 sg13g2_nand2_1 _3506_ (.Y(_0447_),
    .A(net643),
    .B(_0240_));
 sg13g2_o21ai_1 _3507_ (.B1(_0447_),
    .Y(_0448_),
    .A1(_0236_),
    .A2(_0260_));
 sg13g2_nand2_1 _3508_ (.Y(_0449_),
    .A(net559),
    .B(_0438_));
 sg13g2_xor2_1 _3509_ (.B(_0449_),
    .A(_0448_),
    .X(_0450_));
 sg13g2_nand2_1 _3510_ (.Y(_0451_),
    .A(\cordic_inst.cordic_state[36] ),
    .B(_0450_));
 sg13g2_xor2_1 _3511_ (.B(_0450_),
    .A(\cordic_inst.cordic_state[36] ),
    .X(_0452_));
 sg13g2_nand2b_1 _3512_ (.Y(_0453_),
    .B(_0452_),
    .A_N(_0443_));
 sg13g2_nor2_1 _3513_ (.A(_0440_),
    .B(_0452_),
    .Y(_0454_));
 sg13g2_nand2_1 _3514_ (.Y(_0455_),
    .A(_0443_),
    .B(_0454_));
 sg13g2_nand2_1 _3515_ (.Y(_0456_),
    .A(_0440_),
    .B(_0452_));
 sg13g2_nand4_1 _3516_ (.B(_0453_),
    .C(_0455_),
    .A(_2292_),
    .Y(_0457_),
    .D(_0456_));
 sg13g2_a221oi_1 _3517_ (.B2(net748),
    .C1(net579),
    .B1(net601),
    .A1(net679),
    .Y(_0458_),
    .A2(net690));
 sg13g2_o21ai_1 _3518_ (.B1(net774),
    .Y(_0459_),
    .A1(net371),
    .A2(net585));
 sg13g2_a21oi_1 _3519_ (.A1(_0457_),
    .A2(_0458_),
    .Y(_0142_),
    .B1(_0459_));
 sg13g2_and2_1 _3520_ (.A(_0451_),
    .B(_0456_),
    .X(_0460_));
 sg13g2_a22oi_1 _3521_ (.Y(_0461_),
    .B1(_0285_),
    .B2(net597),
    .A2(_0240_),
    .A1(net643));
 sg13g2_o21ai_1 _3522_ (.B1(net559),
    .Y(_0462_),
    .A1(_0438_),
    .A2(_0448_));
 sg13g2_xnor2_1 _3523_ (.Y(_0463_),
    .A(_0461_),
    .B(_0462_));
 sg13g2_xnor2_1 _3524_ (.Y(_0464_),
    .A(\cordic_inst.cordic_state[37] ),
    .B(_0463_));
 sg13g2_nand3_1 _3525_ (.B(_0460_),
    .C(_0464_),
    .A(_0453_),
    .Y(_0465_));
 sg13g2_a21oi_1 _3526_ (.A1(_0453_),
    .A2(_0460_),
    .Y(_0466_),
    .B1(_0464_));
 sg13g2_nand2_1 _3527_ (.Y(_0467_),
    .A(net599),
    .B(_0465_));
 sg13g2_a221oi_1 _3528_ (.B2(net746),
    .C1(net579),
    .B1(net601),
    .A1(net679),
    .Y(_0468_),
    .A2(net688));
 sg13g2_o21ai_1 _3529_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0466_),
    .A2(_0467_));
 sg13g2_o21ai_1 _3530_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net389),
    .A2(net585));
 sg13g2_nand2_1 _3531_ (.Y(_0143_),
    .A(net774),
    .B(_0470_));
 sg13g2_a21oi_1 _3532_ (.A1(\cordic_inst.cordic_state[37] ),
    .A2(_0463_),
    .Y(_0471_),
    .B1(_0466_));
 sg13g2_a21oi_1 _3533_ (.A1(_0461_),
    .A2(_0462_),
    .Y(_0472_),
    .B1(net557));
 sg13g2_xnor2_1 _3534_ (.Y(_0473_),
    .A(net643),
    .B(net646));
 sg13g2_xnor2_1 _3535_ (.Y(_0474_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_a21oi_1 _3536_ (.A1(_0471_),
    .A2(_0474_),
    .Y(_0475_),
    .B1(net584));
 sg13g2_o21ai_1 _3537_ (.B1(_0475_),
    .Y(_0476_),
    .A1(_0471_),
    .A2(_0474_));
 sg13g2_a21oi_1 _3538_ (.A1(net683),
    .A2(net744),
    .Y(_0477_),
    .B1(net678));
 sg13g2_a22oi_1 _3539_ (.Y(_0478_),
    .B1(_0476_),
    .B2(_0477_),
    .A2(_2233_),
    .A1(net678));
 sg13g2_nor2_1 _3540_ (.A(net583),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_o21ai_1 _3541_ (.B1(net786),
    .Y(_0480_),
    .A1(net345),
    .A2(net589));
 sg13g2_nor2_1 _3542_ (.A(_0479_),
    .B(_0480_),
    .Y(_0144_));
 sg13g2_mux2_1 _3543_ (.A0(\cordic_inst.cordic_state[37] ),
    .A1(net646),
    .S(net662),
    .X(_0481_));
 sg13g2_mux4_1 _3544_ (.S0(net662),
    .A0(\cordic_inst.cordic_state[35] ),
    .A1(\cordic_inst.cordic_state[36] ),
    .A2(\cordic_inst.cordic_state[37] ),
    .A3(net646),
    .S1(net659),
    .X(_0482_));
 sg13g2_mux4_1 _3545_ (.S0(net662),
    .A0(\cordic_inst.cordic_state[31] ),
    .A1(net651),
    .A2(net650),
    .A3(net649),
    .S1(net659),
    .X(_0483_));
 sg13g2_mux2_1 _3546_ (.A0(_0483_),
    .A1(_0482_),
    .S(net655),
    .X(_0484_));
 sg13g2_nand2_1 _3547_ (.Y(_0485_),
    .A(net653),
    .B(_0484_));
 sg13g2_mux2_1 _3548_ (.A0(\cordic_inst.cordic_state[25] ),
    .A1(\cordic_inst.cordic_state[26] ),
    .S(net665),
    .X(_0486_));
 sg13g2_mux2_1 _3549_ (.A0(\cordic_inst.cordic_state[23] ),
    .A1(\cordic_inst.cordic_state[24] ),
    .S(net665),
    .X(_0487_));
 sg13g2_and2_1 _3550_ (.A(_0239_),
    .B(_0487_),
    .X(_0488_));
 sg13g2_mux2_1 _3551_ (.A0(\cordic_inst.cordic_state[29] ),
    .A1(\cordic_inst.cordic_state[30] ),
    .S(net663),
    .X(_0489_));
 sg13g2_mux2_1 _3552_ (.A0(\cordic_inst.cordic_state[27] ),
    .A1(\cordic_inst.cordic_state[28] ),
    .S(net664),
    .X(_0490_));
 sg13g2_mux2_1 _3553_ (.A0(_0489_),
    .A1(_0490_),
    .S(net605),
    .X(_0491_));
 sg13g2_a221oi_1 _3554_ (.B2(net595),
    .C1(_0488_),
    .B1(_0491_),
    .A1(_0237_),
    .Y(_0492_),
    .A2(_0486_));
 sg13g2_and2_1 _3555_ (.A(_0485_),
    .B(_0492_),
    .X(_0493_));
 sg13g2_nor2b_1 _3556_ (.A(_0493_),
    .B_N(\cordic_inst.cordic_state[39] ),
    .Y(_0494_));
 sg13g2_xor2_1 _3557_ (.B(_0493_),
    .A(net348),
    .X(_0495_));
 sg13g2_nand2_1 _3558_ (.Y(_0496_),
    .A(_2292_),
    .B(_0495_));
 sg13g2_a221oi_1 _3559_ (.B2(net602),
    .C1(net579),
    .B1(_2227_),
    .A1(net678),
    .Y(_0497_),
    .A2(_2218_));
 sg13g2_a22oi_1 _3560_ (.Y(_0498_),
    .B1(_0496_),
    .B2(_0497_),
    .A2(net580),
    .A1(net348));
 sg13g2_nand2_1 _3561_ (.Y(_0145_),
    .A(net775),
    .B(_0498_));
 sg13g2_mux2_1 _3562_ (.A0(\cordic_inst.cordic_state[36] ),
    .A1(\cordic_inst.cordic_state[37] ),
    .S(net662),
    .X(_0499_));
 sg13g2_a22oi_1 _3563_ (.Y(_0500_),
    .B1(_0499_),
    .B2(net605),
    .A2(_0259_),
    .A1(net646));
 sg13g2_mux2_1 _3564_ (.A0(net649),
    .A1(\cordic_inst.cordic_state[35] ),
    .S(net662),
    .X(_0501_));
 sg13g2_mux2_1 _3565_ (.A0(net651),
    .A1(net650),
    .S(net662),
    .X(_0502_));
 sg13g2_mux4_1 _3566_ (.S0(net662),
    .A0(net651),
    .A1(net650),
    .A2(net649),
    .A3(\cordic_inst.cordic_state[35] ),
    .S1(net659),
    .X(_0503_));
 sg13g2_nor2_1 _3567_ (.A(net655),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_a21oi_1 _3568_ (.A1(net655),
    .A2(_0500_),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_mux2_1 _3569_ (.A0(\cordic_inst.cordic_state[24] ),
    .A1(\cordic_inst.cordic_state[25] ),
    .S(net665),
    .X(_0506_));
 sg13g2_nand2_1 _3570_ (.Y(_0507_),
    .A(_0239_),
    .B(_0506_));
 sg13g2_mux2_1 _3571_ (.A0(\cordic_inst.cordic_state[26] ),
    .A1(\cordic_inst.cordic_state[27] ),
    .S(net665),
    .X(_0508_));
 sg13g2_nand3_1 _3572_ (.B(net597),
    .C(_0508_),
    .A(net660),
    .Y(_0509_));
 sg13g2_and2_1 _3573_ (.A(net646),
    .B(net652),
    .X(_0510_));
 sg13g2_nand2b_1 _3574_ (.Y(_0511_),
    .B(_0510_),
    .A_N(_2296_));
 sg13g2_nand3_1 _3575_ (.B(_0509_),
    .C(_0511_),
    .A(_0507_),
    .Y(_0512_));
 sg13g2_mux2_1 _3576_ (.A0(\cordic_inst.cordic_state[30] ),
    .A1(\cordic_inst.cordic_state[31] ),
    .S(net663),
    .X(_0513_));
 sg13g2_mux2_1 _3577_ (.A0(\cordic_inst.cordic_state[28] ),
    .A1(\cordic_inst.cordic_state[29] ),
    .S(net663),
    .X(_0514_));
 sg13g2_mux2_1 _3578_ (.A0(_0513_),
    .A1(_0514_),
    .S(net605),
    .X(_0515_));
 sg13g2_a221oi_1 _3579_ (.B2(net595),
    .C1(_0512_),
    .B1(_0515_),
    .A1(net652),
    .Y(_0516_),
    .A2(_0505_));
 sg13g2_a221oi_1 _3580_ (.B2(_0492_),
    .C1(_2493_),
    .B1(_0485_),
    .A1(\cordic_atan2_result[15] ),
    .Y(_0517_),
    .A2(_2213_));
 sg13g2_xnor2_1 _3581_ (.Y(_0518_),
    .A(_0516_),
    .B(_0517_));
 sg13g2_and2_1 _3582_ (.A(\cordic_inst.cordic_state[40] ),
    .B(_0518_),
    .X(_0519_));
 sg13g2_xor2_1 _3583_ (.B(_0518_),
    .A(\cordic_inst.cordic_state[40] ),
    .X(_0520_));
 sg13g2_a21oi_1 _3584_ (.A1(_0494_),
    .A2(_0520_),
    .Y(_0521_),
    .B1(_2288_));
 sg13g2_o21ai_1 _3585_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0494_),
    .A2(_0520_));
 sg13g2_nor2b_1 _3586_ (.A(net636),
    .B_N(net602),
    .Y(_0523_));
 sg13g2_a221oi_1 _3587_ (.B2(_0522_),
    .C1(_0523_),
    .B1(net599),
    .A1(net677),
    .Y(_0524_),
    .A2(_2219_));
 sg13g2_a21oi_1 _3588_ (.A1(net325),
    .A2(net581),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nor2_1 _3589_ (.A(net767),
    .B(_0525_),
    .Y(_0146_));
 sg13g2_a21oi_1 _3590_ (.A1(_0494_),
    .A2(_0520_),
    .Y(_0526_),
    .B1(_0519_));
 sg13g2_mux4_1 _3591_ (.S0(net662),
    .A0(net650),
    .A1(net649),
    .A2(\cordic_inst.cordic_state[35] ),
    .A3(\cordic_inst.cordic_state[36] ),
    .S1(net659),
    .X(_0527_));
 sg13g2_nand2_2 _3592_ (.Y(_0528_),
    .A(net605),
    .B(_0481_));
 sg13g2_nor2_1 _3593_ (.A(net655),
    .B(_0527_),
    .Y(_0529_));
 sg13g2_a21oi_1 _3594_ (.A1(net655),
    .A2(_0528_),
    .Y(_0530_),
    .B1(_0529_));
 sg13g2_mux4_1 _3595_ (.S0(net663),
    .A0(\cordic_inst.cordic_state[29] ),
    .A1(\cordic_inst.cordic_state[30] ),
    .A2(\cordic_inst.cordic_state[31] ),
    .A3(net651),
    .S1(net659),
    .X(_0531_));
 sg13g2_nand2_1 _3596_ (.Y(_0532_),
    .A(net595),
    .B(_0531_));
 sg13g2_nand2_1 _3597_ (.Y(_0533_),
    .A(_0239_),
    .B(_0486_));
 sg13g2_nand3_1 _3598_ (.B(_0532_),
    .C(_0533_),
    .A(_0511_),
    .Y(_0534_));
 sg13g2_a221oi_1 _3599_ (.B2(net652),
    .C1(_0534_),
    .B1(_0530_),
    .A1(_0237_),
    .Y(_0535_),
    .A2(_0490_));
 sg13g2_a21oi_1 _3600_ (.A1(_0493_),
    .A2(_0516_),
    .Y(_0536_),
    .B1(net557));
 sg13g2_xnor2_1 _3601_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_nand2_1 _3602_ (.Y(_0538_),
    .A(\cordic_inst.cordic_state[41] ),
    .B(_0537_));
 sg13g2_xnor2_1 _3603_ (.Y(_0539_),
    .A(\cordic_inst.cordic_state[41] ),
    .B(_0537_));
 sg13g2_xnor2_1 _3604_ (.Y(_0540_),
    .A(_0526_),
    .B(_0539_));
 sg13g2_a22oi_1 _3605_ (.Y(_0541_),
    .B1(net633),
    .B2(net603),
    .A2(net728),
    .A1(net681));
 sg13g2_o21ai_1 _3606_ (.B1(_0541_),
    .Y(_0542_),
    .A1(_2284_),
    .A2(_0540_));
 sg13g2_a21oi_1 _3607_ (.A1(net589),
    .A2(_0542_),
    .Y(_0543_),
    .B1(net769));
 sg13g2_o21ai_1 _3608_ (.B1(_0543_),
    .Y(_0147_),
    .A1(_2206_),
    .A2(net589));
 sg13g2_o21ai_1 _3609_ (.B1(_0538_),
    .Y(_0544_),
    .A1(_0526_),
    .A2(_0539_));
 sg13g2_mux2_1 _3610_ (.A0(_0499_),
    .A1(_0501_),
    .S(net605),
    .X(_0545_));
 sg13g2_nand2b_1 _3611_ (.Y(_0546_),
    .B(_0545_),
    .A_N(net655));
 sg13g2_nand3_1 _3612_ (.B(net655),
    .C(_2359_),
    .A(net646),
    .Y(_0547_));
 sg13g2_nand2_1 _3613_ (.Y(_0548_),
    .A(_0546_),
    .B(_0547_));
 sg13g2_mux2_1 _3614_ (.A0(_0502_),
    .A1(_0513_),
    .S(net605),
    .X(_0549_));
 sg13g2_a22oi_1 _3615_ (.Y(_0550_),
    .B1(_0514_),
    .B2(_0237_),
    .A2(_0508_),
    .A1(_0239_));
 sg13g2_a22oi_1 _3616_ (.Y(_0551_),
    .B1(net595),
    .B2(_0549_),
    .A2(_2361_),
    .A1(net646));
 sg13g2_nand2_1 _3617_ (.Y(_0552_),
    .A(_0550_),
    .B(_0551_));
 sg13g2_a21oi_1 _3618_ (.A1(net653),
    .A2(_0548_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_nand3_1 _3619_ (.B(_0516_),
    .C(_0535_),
    .A(_0493_),
    .Y(_0554_));
 sg13g2_nand2_1 _3620_ (.Y(_0555_),
    .A(net561),
    .B(_0554_));
 sg13g2_xor2_1 _3621_ (.B(_0555_),
    .A(_0553_),
    .X(_0556_));
 sg13g2_and2_1 _3622_ (.A(\cordic_inst.cordic_state[42] ),
    .B(_0556_),
    .X(_0557_));
 sg13g2_xor2_1 _3623_ (.B(_0556_),
    .A(\cordic_inst.cordic_state[42] ),
    .X(_0558_));
 sg13g2_a21oi_1 _3624_ (.A1(_0544_),
    .A2(_0558_),
    .Y(_0559_),
    .B1(_2288_));
 sg13g2_o21ai_1 _3625_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0544_),
    .A2(_0558_));
 sg13g2_nand2b_1 _3626_ (.Y(_0561_),
    .B(net602),
    .A_N(net629));
 sg13g2_a22oi_1 _3627_ (.Y(_0562_),
    .B1(net599),
    .B2(_0560_),
    .A2(_2220_),
    .A1(net680));
 sg13g2_a22oi_1 _3628_ (.Y(_0563_),
    .B1(_0561_),
    .B2(_0562_),
    .A2(net582),
    .A1(net336));
 sg13g2_nor2_1 _3629_ (.A(net767),
    .B(_0563_),
    .Y(_0148_));
 sg13g2_a21oi_1 _3630_ (.A1(_0544_),
    .A2(_0558_),
    .Y(_0564_),
    .B1(_0557_));
 sg13g2_a22oi_1 _3631_ (.Y(_0565_),
    .B1(_0510_),
    .B2(_2294_),
    .A2(_0483_),
    .A1(net595));
 sg13g2_a22oi_1 _3632_ (.Y(_0566_),
    .B1(_0491_),
    .B2(net597),
    .A2(_0482_),
    .A1(_0325_));
 sg13g2_nand2_2 _3633_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_nand4_1 _3634_ (.B(_0516_),
    .C(_0535_),
    .A(_0493_),
    .Y(_0568_),
    .D(_0553_));
 sg13g2_nand2_1 _3635_ (.Y(_0569_),
    .A(net561),
    .B(_0568_));
 sg13g2_xnor2_1 _3636_ (.Y(_0570_),
    .A(_0567_),
    .B(_0569_));
 sg13g2_nand2_1 _3637_ (.Y(_0571_),
    .A(\cordic_inst.cordic_state[43] ),
    .B(_0570_));
 sg13g2_xnor2_1 _3638_ (.Y(_0572_),
    .A(\cordic_inst.cordic_state[43] ),
    .B(_0570_));
 sg13g2_xor2_1 _3639_ (.B(_0572_),
    .A(_0564_),
    .X(_0573_));
 sg13g2_a221oi_1 _3640_ (.B2(net602),
    .C1(net579),
    .B1(_2229_),
    .A1(net678),
    .Y(_0574_),
    .A2(_2221_));
 sg13g2_o21ai_1 _3641_ (.B1(_0574_),
    .Y(_0575_),
    .A1(_2293_),
    .A2(_0573_));
 sg13g2_a21oi_1 _3642_ (.A1(net347),
    .A2(net583),
    .Y(_0576_),
    .B1(net767));
 sg13g2_nand2_1 _3643_ (.Y(_0149_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_nor2_1 _3644_ (.A(_2216_),
    .B(net718),
    .Y(_0577_));
 sg13g2_o21ai_1 _3645_ (.B1(_0571_),
    .Y(_0578_),
    .A1(_0564_),
    .A2(_0572_));
 sg13g2_inv_1 _3646_ (.Y(_0579_),
    .A(_0578_));
 sg13g2_nand2_1 _3647_ (.Y(_0580_),
    .A(net595),
    .B(_0503_));
 sg13g2_o21ai_1 _3648_ (.B1(_0580_),
    .Y(_0581_),
    .A1(_0326_),
    .A2(_0500_));
 sg13g2_a221oi_1 _3649_ (.B2(net598),
    .C1(_0581_),
    .B1(_0515_),
    .A1(_2294_),
    .Y(_0582_),
    .A2(_0510_));
 sg13g2_o21ai_1 _3650_ (.B1(net561),
    .Y(_0583_),
    .A1(_0567_),
    .A2(_0568_));
 sg13g2_xnor2_1 _3651_ (.Y(_0584_),
    .A(_0582_),
    .B(_0583_));
 sg13g2_inv_1 _3652_ (.Y(_0585_),
    .A(_0584_));
 sg13g2_nand2_1 _3653_ (.Y(_0586_),
    .A(\cordic_inst.cordic_state[44] ),
    .B(_0585_));
 sg13g2_xor2_1 _3654_ (.B(_0584_),
    .A(\cordic_inst.cordic_state[44] ),
    .X(_0587_));
 sg13g2_nand2b_1 _3655_ (.Y(_0588_),
    .B(_0578_),
    .A_N(_0587_));
 sg13g2_a21oi_1 _3656_ (.A1(_0579_),
    .A2(_0587_),
    .Y(_0589_),
    .B1(net584));
 sg13g2_a221oi_1 _3657_ (.B2(_0589_),
    .C1(net680),
    .B1(_0588_),
    .A1(net683),
    .Y(_0590_),
    .A2(net619));
 sg13g2_o21ai_1 _3658_ (.B1(net588),
    .Y(_0591_),
    .A1(_0577_),
    .A2(_0590_));
 sg13g2_o21ai_1 _3659_ (.B1(_0591_),
    .Y(_0592_),
    .A1(net358),
    .A2(net588));
 sg13g2_nor2_1 _3660_ (.A(net768),
    .B(_0592_),
    .Y(_0150_));
 sg13g2_nand2_1 _3661_ (.Y(_0593_),
    .A(net595),
    .B(_0527_));
 sg13g2_o21ai_1 _3662_ (.B1(_0593_),
    .Y(_0594_),
    .A1(_0326_),
    .A2(_0528_));
 sg13g2_a22oi_1 _3663_ (.Y(_0595_),
    .B1(_0531_),
    .B2(net597),
    .A2(_0357_),
    .A1(net647));
 sg13g2_nand2b_2 _3664_ (.Y(_0596_),
    .B(_0595_),
    .A_N(_0594_));
 sg13g2_a21o_1 _3665_ (.A2(_0583_),
    .A1(_0582_),
    .B1(net557),
    .X(_0597_));
 sg13g2_xnor2_1 _3666_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_nand2_1 _3667_ (.Y(_0599_),
    .A(\cordic_inst.cordic_state[45] ),
    .B(_0598_));
 sg13g2_xnor2_1 _3668_ (.Y(_0600_),
    .A(\cordic_inst.cordic_state[45] ),
    .B(_0598_));
 sg13g2_nand3_1 _3669_ (.B(_0588_),
    .C(_0600_),
    .A(_0586_),
    .Y(_0601_));
 sg13g2_a21o_1 _3670_ (.A2(_0588_),
    .A1(_0586_),
    .B1(_0600_),
    .X(_0602_));
 sg13g2_nand3_1 _3671_ (.B(_0601_),
    .C(_0602_),
    .A(net600),
    .Y(_0603_));
 sg13g2_a22oi_1 _3672_ (.Y(_0604_),
    .B1(net618),
    .B2(net601),
    .A2(net712),
    .A1(net677));
 sg13g2_nand2_1 _3673_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_a21oi_1 _3674_ (.A1(net587),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net767));
 sg13g2_o21ai_1 _3675_ (.B1(_0606_),
    .Y(_0151_),
    .A1(_2205_),
    .A2(net588));
 sg13g2_a22oi_1 _3676_ (.Y(_0607_),
    .B1(_0549_),
    .B2(net597),
    .A2(_0545_),
    .A1(net595));
 sg13g2_nand2b_2 _3677_ (.Y(_0608_),
    .B(_0607_),
    .A_N(_0510_));
 sg13g2_nand2_1 _3678_ (.Y(_0609_),
    .A(net560),
    .B(_0596_));
 sg13g2_nand2_1 _3679_ (.Y(_0610_),
    .A(_0597_),
    .B(_0609_));
 sg13g2_xor2_1 _3680_ (.B(_0610_),
    .A(_0608_),
    .X(_0611_));
 sg13g2_nand2_1 _3681_ (.Y(_0612_),
    .A(\cordic_inst.cordic_state[46] ),
    .B(_0611_));
 sg13g2_xnor2_1 _3682_ (.Y(_0613_),
    .A(\cordic_inst.cordic_state[46] ),
    .B(_0611_));
 sg13g2_a21o_1 _3683_ (.A2(_0602_),
    .A1(_0599_),
    .B1(_0613_),
    .X(_0614_));
 sg13g2_nand3_1 _3684_ (.B(_0602_),
    .C(_0613_),
    .A(_0599_),
    .Y(_0615_));
 sg13g2_nand3_1 _3685_ (.B(_0614_),
    .C(_0615_),
    .A(_2287_),
    .Y(_0616_));
 sg13g2_nand2b_1 _3686_ (.Y(_0617_),
    .B(net601),
    .A_N(net615));
 sg13g2_a22oi_1 _3687_ (.Y(_0618_),
    .B1(net599),
    .B2(_0616_),
    .A2(_2224_),
    .A1(net675));
 sg13g2_a22oi_1 _3688_ (.Y(_0619_),
    .B1(_0617_),
    .B2(_0618_),
    .A2(net580),
    .A1(net351));
 sg13g2_nor2_1 _3689_ (.A(net767),
    .B(net352),
    .Y(_0152_));
 sg13g2_a21oi_2 _3690_ (.B1(_0510_),
    .Y(_0620_),
    .A2(_0484_),
    .A1(net608));
 sg13g2_a21oi_1 _3691_ (.A1(net560),
    .A2(_0608_),
    .Y(_0621_),
    .B1(_0610_));
 sg13g2_xor2_1 _3692_ (.B(_0621_),
    .A(_0620_),
    .X(_0622_));
 sg13g2_and2_1 _3693_ (.A(\cordic_inst.cordic_state[47] ),
    .B(_0622_),
    .X(_0623_));
 sg13g2_xnor2_1 _3694_ (.Y(_0624_),
    .A(\cordic_inst.cordic_state[47] ),
    .B(_0622_));
 sg13g2_nand3_1 _3695_ (.B(_0614_),
    .C(_0624_),
    .A(_0612_),
    .Y(_0625_));
 sg13g2_a21oi_1 _3696_ (.A1(_0612_),
    .A2(_0614_),
    .Y(_0626_),
    .B1(_0624_));
 sg13g2_nand2_1 _3697_ (.Y(_0627_),
    .A(net599),
    .B(_0625_));
 sg13g2_a221oi_1 _3698_ (.B2(net601),
    .C1(net580),
    .B1(net708),
    .A1(net677),
    .Y(_0628_),
    .A2(net762));
 sg13g2_o21ai_1 _3699_ (.B1(_0628_),
    .Y(_0629_),
    .A1(_0626_),
    .A2(_0627_));
 sg13g2_o21ai_1 _3700_ (.B1(_0629_),
    .Y(_0630_),
    .A1(net374),
    .A2(net587));
 sg13g2_nand2_1 _3701_ (.Y(_0153_),
    .A(net775),
    .B(_0630_));
 sg13g2_nor2_1 _3702_ (.A(net604),
    .B(net759),
    .Y(_0631_));
 sg13g2_a22oi_1 _3703_ (.Y(_0632_),
    .B1(_0505_),
    .B2(net607),
    .A2(_0399_),
    .A1(net647));
 sg13g2_inv_1 _3704_ (.Y(_0633_),
    .A(_0632_));
 sg13g2_o21ai_1 _3705_ (.B1(_0621_),
    .Y(_0634_),
    .A1(net557),
    .A2(_0620_));
 sg13g2_xnor2_1 _3706_ (.Y(_0635_),
    .A(_0632_),
    .B(_0634_));
 sg13g2_nand2_1 _3707_ (.Y(_0636_),
    .A(\cordic_inst.cordic_state[48] ),
    .B(_0635_));
 sg13g2_xor2_1 _3708_ (.B(_0635_),
    .A(\cordic_inst.cordic_state[48] ),
    .X(_0637_));
 sg13g2_o21ai_1 _3709_ (.B1(_0637_),
    .Y(_0638_),
    .A1(_0623_),
    .A2(_0626_));
 sg13g2_nor3_1 _3710_ (.A(_0623_),
    .B(_0626_),
    .C(_0637_),
    .Y(_0639_));
 sg13g2_nor2_1 _3711_ (.A(_2291_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_a221oi_1 _3712_ (.B2(_0640_),
    .C1(net676),
    .B1(_0638_),
    .A1(net682),
    .Y(_0641_),
    .A2(net703));
 sg13g2_o21ai_1 _3713_ (.B1(net587),
    .Y(_0642_),
    .A1(_0631_),
    .A2(_0641_));
 sg13g2_o21ai_1 _3714_ (.B1(_0642_),
    .Y(_0643_),
    .A1(net361),
    .A2(net587));
 sg13g2_nor2_1 _3715_ (.A(net768),
    .B(net362),
    .Y(_0154_));
 sg13g2_a22oi_1 _3716_ (.Y(_0644_),
    .B1(_0530_),
    .B2(net607),
    .A2(_0399_),
    .A1(net647));
 sg13g2_a21oi_1 _3717_ (.A1(net560),
    .A2(_0633_),
    .Y(_0645_),
    .B1(_0634_));
 sg13g2_xor2_1 _3718_ (.B(_0645_),
    .A(_0644_),
    .X(_0646_));
 sg13g2_xnor2_1 _3719_ (.Y(_0647_),
    .A(\cordic_inst.cordic_state[49] ),
    .B(_0646_));
 sg13g2_nand3_1 _3720_ (.B(_0638_),
    .C(_0647_),
    .A(_0636_),
    .Y(_0648_));
 sg13g2_a21oi_1 _3721_ (.A1(_0636_),
    .A2(_0638_),
    .Y(_0649_),
    .B1(_0647_));
 sg13g2_nand2_1 _3722_ (.Y(_0650_),
    .A(net599),
    .B(_0648_));
 sg13g2_a221oi_1 _3723_ (.B2(net601),
    .C1(net580),
    .B1(net700),
    .A1(net675),
    .Y(_0651_),
    .A2(net756));
 sg13g2_o21ai_1 _3724_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_0649_),
    .A2(_0650_));
 sg13g2_o21ai_1 _3725_ (.B1(_0652_),
    .Y(_0653_),
    .A1(net390),
    .A2(net587));
 sg13g2_nand2_1 _3726_ (.Y(_0155_),
    .A(net775),
    .B(_0653_));
 sg13g2_nor2_1 _3727_ (.A(net604),
    .B(net753),
    .Y(_0654_));
 sg13g2_a21oi_1 _3728_ (.A1(\cordic_inst.cordic_state[49] ),
    .A2(_0646_),
    .Y(_0655_),
    .B1(_0649_));
 sg13g2_a21o_1 _3729_ (.A2(_0645_),
    .A1(_0644_),
    .B1(net557),
    .X(_0656_));
 sg13g2_a22oi_1 _3730_ (.Y(_0657_),
    .B1(_0548_),
    .B2(net607),
    .A2(_0236_),
    .A1(net647));
 sg13g2_xnor2_1 _3731_ (.Y(_0658_),
    .A(_0656_),
    .B(_0657_));
 sg13g2_nand2b_1 _3732_ (.Y(_0659_),
    .B(\cordic_inst.cordic_state[50] ),
    .A_N(_0658_));
 sg13g2_xor2_1 _3733_ (.B(_0658_),
    .A(\cordic_inst.cordic_state[50] ),
    .X(_0660_));
 sg13g2_or2_1 _3734_ (.X(_0661_),
    .B(_0660_),
    .A(_0655_));
 sg13g2_a21oi_1 _3735_ (.A1(_0655_),
    .A2(_0660_),
    .Y(_0662_),
    .B1(_2291_));
 sg13g2_a221oi_1 _3736_ (.B2(_0662_),
    .C1(net677),
    .B1(_0661_),
    .A1(cordic_en_atan2),
    .Y(_0663_),
    .A2(net697));
 sg13g2_o21ai_1 _3737_ (.B1(net588),
    .Y(_0664_),
    .A1(_0654_),
    .A2(_0663_));
 sg13g2_o21ai_1 _3738_ (.B1(_0664_),
    .Y(_0665_),
    .A1(net367),
    .A2(net588));
 sg13g2_nor2_1 _3739_ (.A(net767),
    .B(net368),
    .Y(_0156_));
 sg13g2_and2_1 _3740_ (.A(net597),
    .B(_0482_),
    .X(_0666_));
 sg13g2_a21oi_1 _3741_ (.A1(net648),
    .A2(_0236_),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_o21ai_1 _3742_ (.B1(_0656_),
    .Y(_0668_),
    .A1(net557),
    .A2(_0657_));
 sg13g2_xor2_1 _3743_ (.B(_0668_),
    .A(_0667_),
    .X(_0669_));
 sg13g2_nor2_1 _3744_ (.A(_2204_),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_xnor2_1 _3745_ (.Y(_0671_),
    .A(_2204_),
    .B(_0669_));
 sg13g2_a21oi_1 _3746_ (.A1(_0659_),
    .A2(_0661_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_and3_1 _3747_ (.X(_0673_),
    .A(_0659_),
    .B(_0661_),
    .C(_0671_));
 sg13g2_o21ai_1 _3748_ (.B1(_2287_),
    .Y(_0674_),
    .A1(_0672_),
    .A2(_0673_));
 sg13g2_a221oi_1 _3749_ (.B2(_0674_),
    .C1(net677),
    .B1(_2282_),
    .A1(cordic_en_atan2),
    .Y(_0675_),
    .A2(net693));
 sg13g2_o21ai_1 _3750_ (.B1(net588),
    .Y(_0676_),
    .A1(net604),
    .A2(net750));
 sg13g2_a21oi_1 _3751_ (.A1(net349),
    .A2(net579),
    .Y(_0677_),
    .B1(net767));
 sg13g2_o21ai_1 _3752_ (.B1(_0677_),
    .Y(_0157_),
    .A1(_0675_),
    .A2(_0676_));
 sg13g2_nand2_1 _3753_ (.Y(_0678_),
    .A(net646),
    .B(_0240_));
 sg13g2_o21ai_1 _3754_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0236_),
    .A2(_0500_));
 sg13g2_a21oi_1 _3755_ (.A1(net560),
    .A2(_0666_),
    .Y(_0680_),
    .B1(_0668_));
 sg13g2_nand2b_1 _3756_ (.Y(_0681_),
    .B(_0680_),
    .A_N(_0679_));
 sg13g2_xnor2_1 _3757_ (.Y(_0682_),
    .A(_0679_),
    .B(_0680_));
 sg13g2_xor2_1 _3758_ (.B(_0682_),
    .A(\cordic_inst.cordic_state[52] ),
    .X(_0683_));
 sg13g2_and2_1 _3759_ (.A(_0672_),
    .B(_0683_),
    .X(_0684_));
 sg13g2_nor3_1 _3760_ (.A(_0670_),
    .B(_0672_),
    .C(_0683_),
    .Y(_0685_));
 sg13g2_and2_1 _3761_ (.A(_0670_),
    .B(_0683_),
    .X(_0686_));
 sg13g2_or4_1 _3762_ (.A(_2293_),
    .B(_0684_),
    .C(_0685_),
    .D(_0686_),
    .X(_0687_));
 sg13g2_a221oi_1 _3763_ (.B2(net602),
    .C1(net579),
    .B1(net690),
    .A1(net678),
    .Y(_0688_),
    .A2(net748));
 sg13g2_o21ai_1 _3764_ (.B1(net786),
    .Y(_0689_),
    .A1(net356),
    .A2(net589));
 sg13g2_a21oi_1 _3765_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0158_),
    .B1(_0689_));
 sg13g2_a21oi_1 _3766_ (.A1(\cordic_inst.cordic_state[52] ),
    .A2(_0682_),
    .Y(_0690_),
    .B1(_0686_));
 sg13g2_nor2b_1 _3767_ (.A(_0684_),
    .B_N(_0690_),
    .Y(_0691_));
 sg13g2_nor2_1 _3768_ (.A(_0236_),
    .B(_0528_),
    .Y(_0692_));
 sg13g2_o21ai_1 _3769_ (.B1(_0678_),
    .Y(_0693_),
    .A1(_0236_),
    .A2(_0528_));
 sg13g2_nand2_1 _3770_ (.Y(_0694_),
    .A(net560),
    .B(_0681_));
 sg13g2_xnor2_1 _3771_ (.Y(_0695_),
    .A(_0693_),
    .B(_0694_));
 sg13g2_xor2_1 _3772_ (.B(_0695_),
    .A(\cordic_inst.cordic_state[53] ),
    .X(_0696_));
 sg13g2_nor2b_1 _3773_ (.A(_0691_),
    .B_N(_0696_),
    .Y(_0697_));
 sg13g2_xnor2_1 _3774_ (.Y(_0698_),
    .A(_0691_),
    .B(_0696_));
 sg13g2_o21ai_1 _3775_ (.B1(_2282_),
    .Y(_0699_),
    .A1(_2288_),
    .A2(_0698_));
 sg13g2_a21oi_1 _3776_ (.A1(net683),
    .A2(net688),
    .Y(_0700_),
    .B1(net678));
 sg13g2_a221oi_1 _3777_ (.B2(_0700_),
    .C1(net579),
    .B1(_0699_),
    .A1(net679),
    .Y(_0701_),
    .A2(_2225_));
 sg13g2_a21oi_1 _3778_ (.A1(net353),
    .A2(net583),
    .Y(_0702_),
    .B1(net773));
 sg13g2_nand2b_1 _3779_ (.Y(_0159_),
    .B(_0702_),
    .A_N(_0701_));
 sg13g2_a21o_1 _3780_ (.A2(_0695_),
    .A1(\cordic_inst.cordic_state[53] ),
    .B1(_0697_),
    .X(_0703_));
 sg13g2_o21ai_1 _3781_ (.B1(net559),
    .Y(_0704_),
    .A1(_0681_),
    .A2(_0692_));
 sg13g2_xor2_1 _3782_ (.B(_0704_),
    .A(_0473_),
    .X(_0705_));
 sg13g2_a21oi_1 _3783_ (.A1(_0703_),
    .A2(_0705_),
    .Y(_0706_),
    .B1(_2291_));
 sg13g2_o21ai_1 _3784_ (.B1(_0706_),
    .Y(_0707_),
    .A1(_0703_),
    .A2(_0705_));
 sg13g2_a21oi_1 _3785_ (.A1(net683),
    .A2(net687),
    .Y(_0708_),
    .B1(net678));
 sg13g2_a22oi_1 _3786_ (.Y(_0709_),
    .B1(_0707_),
    .B2(_0708_),
    .A2(_2226_),
    .A1(net678));
 sg13g2_nor2_1 _3787_ (.A(net579),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_o21ai_1 _3788_ (.B1(net786),
    .Y(_0711_),
    .A1(net645),
    .A2(net589));
 sg13g2_nor2_1 _3789_ (.A(_0710_),
    .B(_0711_),
    .Y(_0160_));
 sg13g2_nand3_1 _3790_ (.B(net143),
    .C(_2212_),
    .A(_2203_),
    .Y(_0712_));
 sg13g2_nand2_1 _3791_ (.Y(_0713_),
    .A(net143),
    .B(_0712_));
 sg13g2_a21oi_1 _3792_ (.A1(net600),
    .A2(net144),
    .Y(_0161_),
    .B1(net770));
 sg13g2_or4_1 _3793_ (.A(_2203_),
    .B(cordic_en_get_atan2),
    .C(cordic_en_get_sqrt),
    .D(net167),
    .X(_0714_));
 sg13g2_a21oi_1 _3794_ (.A1(_0712_),
    .A2(net168),
    .Y(_0162_),
    .B1(_2285_));
 sg13g2_nor2b_1 _3795_ (.A(_2308_),
    .B_N(_2366_),
    .Y(_0163_));
 sg13g2_nor3_2 _3796_ (.A(_2264_),
    .B(_2430_),
    .C(_2461_),
    .Y(_0715_));
 sg13g2_nand2_1 _3797_ (.Y(_0716_),
    .A(net1),
    .B(net574));
 sg13g2_o21ai_1 _3798_ (.B1(_0716_),
    .Y(_0165_),
    .A1(_2227_),
    .A2(net574));
 sg13g2_mux2_1 _3799_ (.A0(net637),
    .A1(net2),
    .S(net575),
    .X(_0166_));
 sg13g2_nand2_1 _3800_ (.Y(_0717_),
    .A(net3),
    .B(net574));
 sg13g2_o21ai_1 _3801_ (.B1(_0717_),
    .Y(_0167_),
    .A1(_2228_),
    .A2(net574));
 sg13g2_mux2_1 _3802_ (.A0(net629),
    .A1(net4),
    .S(net574),
    .X(_0168_));
 sg13g2_nand2_1 _3803_ (.Y(_0718_),
    .A(net5),
    .B(net574));
 sg13g2_o21ai_1 _3804_ (.B1(_0718_),
    .Y(_0169_),
    .A1(_2229_),
    .A2(net574));
 sg13g2_nand2_1 _3805_ (.Y(_0719_),
    .A(net6),
    .B(net575));
 sg13g2_o21ai_1 _3806_ (.B1(_0719_),
    .Y(_0170_),
    .A1(_2230_),
    .A2(net575));
 sg13g2_nand2_1 _3807_ (.Y(_0720_),
    .A(net7),
    .B(net575));
 sg13g2_o21ai_1 _3808_ (.B1(_0720_),
    .Y(_0171_),
    .A1(_2231_),
    .A2(net575));
 sg13g2_mux2_1 _3809_ (.A0(net615),
    .A1(net8),
    .S(net574),
    .X(_0172_));
 sg13g2_nor4_1 _3810_ (.A(_2218_),
    .B(_2219_),
    .C(_2229_),
    .D(_2230_),
    .Y(_0721_));
 sg13g2_nand4_1 _3811_ (.B(net732),
    .C(net624),
    .A(net737),
    .Y(_0722_),
    .D(net619));
 sg13g2_nand2_1 _3812_ (.Y(_0723_),
    .A(net727),
    .B(net629));
 sg13g2_a22oi_1 _3813_ (.Y(_0724_),
    .B1(net619),
    .B2(net737),
    .A2(net624),
    .A1(net732));
 sg13g2_nor3_1 _3814_ (.A(_0721_),
    .B(_0723_),
    .C(_0724_),
    .Y(_0725_));
 sg13g2_o21ai_1 _3815_ (.B1(_0722_),
    .Y(_0726_),
    .A1(_0723_),
    .A2(_0724_));
 sg13g2_nand2_1 _3816_ (.Y(_0727_),
    .A(net723),
    .B(net629));
 sg13g2_and4_1 _3817_ (.A(net732),
    .B(net727),
    .C(net624),
    .D(net619),
    .X(_0728_));
 sg13g2_nand4_1 _3818_ (.B(net727),
    .C(net624),
    .A(net732),
    .Y(_0729_),
    .D(net623));
 sg13g2_a22oi_1 _3819_ (.Y(_0730_),
    .B1(net619),
    .B2(net733),
    .A2(net624),
    .A1(net727));
 sg13g2_or3_1 _3820_ (.A(_0727_),
    .B(_0728_),
    .C(_0730_),
    .X(_0731_));
 sg13g2_o21ai_1 _3821_ (.B1(_0727_),
    .Y(_0732_),
    .A1(_0728_),
    .A2(_0730_));
 sg13g2_and3_1 _3822_ (.X(_0733_),
    .A(_0726_),
    .B(_0731_),
    .C(_0732_));
 sg13g2_nand2_1 _3823_ (.Y(_0734_),
    .A(net712),
    .B(net640));
 sg13g2_nand2_1 _3824_ (.Y(_0735_),
    .A(net718),
    .B(net633));
 sg13g2_nand2_1 _3825_ (.Y(_0736_),
    .A(net719),
    .B(net636));
 sg13g2_nand2_1 _3826_ (.Y(_0737_),
    .A(net719),
    .B(net633));
 sg13g2_nand2_1 _3827_ (.Y(_0738_),
    .A(net718),
    .B(net636));
 sg13g2_xor2_1 _3828_ (.B(_0738_),
    .A(_0737_),
    .X(_0739_));
 sg13g2_nand2b_1 _3829_ (.Y(_0740_),
    .B(_0739_),
    .A_N(_0734_));
 sg13g2_xnor2_1 _3830_ (.Y(_0741_),
    .A(_0734_),
    .B(_0739_));
 sg13g2_inv_1 _3831_ (.Y(_0742_),
    .A(_0741_));
 sg13g2_a21oi_1 _3832_ (.A1(_0731_),
    .A2(_0732_),
    .Y(_0743_),
    .B1(_0726_));
 sg13g2_or2_1 _3833_ (.X(_0744_),
    .B(_0743_),
    .A(_0733_));
 sg13g2_nor2_1 _3834_ (.A(_0742_),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_o21ai_1 _3835_ (.B1(_0740_),
    .Y(_0746_),
    .A1(_0737_),
    .A2(_0738_));
 sg13g2_o21ai_1 _3836_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0733_),
    .A2(_0745_));
 sg13g2_nand2_1 _3837_ (.Y(_0748_),
    .A(net712),
    .B(net636));
 sg13g2_nand2_1 _3838_ (.Y(_0749_),
    .A(net711),
    .B(net641));
 sg13g2_xor2_1 _3839_ (.B(_0748_),
    .A(_0735_),
    .X(_0750_));
 sg13g2_nand2b_1 _3840_ (.Y(_0751_),
    .B(_0750_),
    .A_N(_0749_));
 sg13g2_o21ai_1 _3841_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0735_),
    .A2(_0748_));
 sg13g2_xnor2_1 _3842_ (.Y(_0753_),
    .A(_0741_),
    .B(_0744_));
 sg13g2_xnor2_1 _3843_ (.Y(_0754_),
    .A(_0742_),
    .B(_0744_));
 sg13g2_nand2_1 _3844_ (.Y(_0755_),
    .A(net737),
    .B(net618));
 sg13g2_inv_1 _3845_ (.Y(_0756_),
    .A(_0755_));
 sg13g2_nand4_1 _3846_ (.B(net733),
    .C(net618),
    .A(net738),
    .Y(_0757_),
    .D(net615));
 sg13g2_inv_1 _3847_ (.Y(_0758_),
    .A(_0757_));
 sg13g2_a22oi_1 _3848_ (.Y(_0759_),
    .B1(net615),
    .B2(net738),
    .A2(net618),
    .A1(net733));
 sg13g2_nor2_1 _3849_ (.A(_0758_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_xnor2_1 _3850_ (.Y(_0761_),
    .A(_0749_),
    .B(_0750_));
 sg13g2_o21ai_1 _3851_ (.B1(_0729_),
    .Y(_0762_),
    .A1(_0727_),
    .A2(_0730_));
 sg13g2_nand2_1 _3852_ (.Y(_0763_),
    .A(net719),
    .B(net632));
 sg13g2_and4_1 _3853_ (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .B(net723),
    .C(net625),
    .D(net619),
    .X(_0764_));
 sg13g2_nand4_1 _3854_ (.B(net723),
    .C(net625),
    .A(net728),
    .Y(_0765_),
    .D(net619));
 sg13g2_a22oi_1 _3855_ (.Y(_0766_),
    .B1(net623),
    .B2(net728),
    .A2(net625),
    .A1(net726));
 sg13g2_or3_1 _3856_ (.A(_0763_),
    .B(_0764_),
    .C(_0766_),
    .X(_0767_));
 sg13g2_o21ai_1 _3857_ (.B1(_0763_),
    .Y(_0768_),
    .A1(_0764_),
    .A2(_0766_));
 sg13g2_nand3_1 _3858_ (.B(_0767_),
    .C(_0768_),
    .A(_0762_),
    .Y(_0769_));
 sg13g2_a21o_1 _3859_ (.A2(_0768_),
    .A1(_0767_),
    .B1(_0762_),
    .X(_0770_));
 sg13g2_a21o_1 _3860_ (.A2(_0770_),
    .A1(_0769_),
    .B1(_0761_),
    .X(_0771_));
 sg13g2_nand3_1 _3861_ (.B(_0769_),
    .C(_0770_),
    .A(_0761_),
    .Y(_0772_));
 sg13g2_nand3_1 _3862_ (.B(_0771_),
    .C(_0772_),
    .A(_0760_),
    .Y(_0773_));
 sg13g2_a21o_1 _3863_ (.A2(_0772_),
    .A1(_0771_),
    .B1(_0760_),
    .X(_0774_));
 sg13g2_nand2_1 _3864_ (.Y(_0775_),
    .A(_0773_),
    .B(_0774_));
 sg13g2_nand4_1 _3865_ (.B(_0756_),
    .C(_0773_),
    .A(_0753_),
    .Y(_0776_),
    .D(_0774_));
 sg13g2_nand2_1 _3866_ (.Y(_0777_),
    .A(_0769_),
    .B(_0772_));
 sg13g2_nor2b_1 _3867_ (.A(_0776_),
    .B_N(_0777_),
    .Y(_0778_));
 sg13g2_xnor2_1 _3868_ (.Y(_0779_),
    .A(_0776_),
    .B(_0777_));
 sg13g2_xnor2_1 _3869_ (.Y(_0780_),
    .A(_0752_),
    .B(_0779_));
 sg13g2_nand2_1 _3870_ (.Y(_0781_),
    .A(net762),
    .B(net641));
 sg13g2_nand2_1 _3871_ (.Y(_0782_),
    .A(net711),
    .B(net634));
 sg13g2_and4_1 _3872_ (.A(net712),
    .B(net711),
    .C(net637),
    .D(net635),
    .X(_0783_));
 sg13g2_a22oi_1 _3873_ (.Y(_0784_),
    .B1(net635),
    .B2(net715),
    .A2(net637),
    .A1(net711));
 sg13g2_nor3_1 _3874_ (.A(_0781_),
    .B(_0783_),
    .C(_0784_),
    .Y(_0785_));
 sg13g2_o21ai_1 _3875_ (.B1(_0781_),
    .Y(_0786_),
    .A1(_0783_),
    .A2(_0784_));
 sg13g2_nor2b_1 _3876_ (.A(_0785_),
    .B_N(_0786_),
    .Y(_0787_));
 sg13g2_o21ai_1 _3877_ (.B1(_0765_),
    .Y(_0788_),
    .A1(_0763_),
    .A2(_0766_));
 sg13g2_nand2_1 _3878_ (.Y(_0789_),
    .A(net718),
    .B(net632));
 sg13g2_nand2_1 _3879_ (.Y(_0790_),
    .A(net719),
    .B(net622));
 sg13g2_and4_1 _3880_ (.A(net726),
    .B(net722),
    .C(net625),
    .D(net619),
    .X(_0791_));
 sg13g2_a22oi_1 _3881_ (.Y(_0792_),
    .B1(net623),
    .B2(net723),
    .A2(net625),
    .A1(net722));
 sg13g2_or3_1 _3882_ (.A(_0789_),
    .B(_0791_),
    .C(_0792_),
    .X(_0793_));
 sg13g2_o21ai_1 _3883_ (.B1(_0789_),
    .Y(_0794_),
    .A1(_0791_),
    .A2(_0792_));
 sg13g2_nand3_1 _3884_ (.B(_0793_),
    .C(_0794_),
    .A(_0788_),
    .Y(_0795_));
 sg13g2_a21o_1 _3885_ (.A2(_0794_),
    .A1(_0793_),
    .B1(_0788_),
    .X(_0796_));
 sg13g2_a21o_1 _3886_ (.A2(_0796_),
    .A1(_0795_),
    .B1(_0787_),
    .X(_0797_));
 sg13g2_nand3_1 _3887_ (.B(_0795_),
    .C(_0796_),
    .A(_0787_),
    .Y(_0798_));
 sg13g2_nand2_1 _3888_ (.Y(_0799_),
    .A(net728),
    .B(net618));
 sg13g2_and4_1 _3889_ (.A(net738),
    .B(net733),
    .C(net615),
    .D(net708),
    .X(_0800_));
 sg13g2_a22oi_1 _3890_ (.Y(_0801_),
    .B1(net708),
    .B2(net738),
    .A2(net615),
    .A1(net733));
 sg13g2_nor2_1 _3891_ (.A(_0800_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_nor3_1 _3892_ (.A(_0799_),
    .B(_0800_),
    .C(_0801_),
    .Y(_0803_));
 sg13g2_xnor2_1 _3893_ (.Y(_0804_),
    .A(_0799_),
    .B(_0802_));
 sg13g2_nand2_1 _3894_ (.Y(_0805_),
    .A(_0758_),
    .B(_0804_));
 sg13g2_xnor2_1 _3895_ (.Y(_0806_),
    .A(_0757_),
    .B(_0804_));
 sg13g2_and3_1 _3896_ (.X(_0807_),
    .A(_0797_),
    .B(_0798_),
    .C(_0806_));
 sg13g2_nand3_1 _3897_ (.B(_0798_),
    .C(_0806_),
    .A(_0797_),
    .Y(_0808_));
 sg13g2_a21oi_1 _3898_ (.A1(_0797_),
    .A2(_0798_),
    .Y(_0809_),
    .B1(_0806_));
 sg13g2_nor2_1 _3899_ (.A(_0807_),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_nor3_1 _3900_ (.A(_0773_),
    .B(_0807_),
    .C(_0809_),
    .Y(_0811_));
 sg13g2_xor2_1 _3901_ (.B(_0810_),
    .A(_0773_),
    .X(_0812_));
 sg13g2_nor2_1 _3902_ (.A(_0780_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_xnor2_1 _3903_ (.Y(_0814_),
    .A(_0780_),
    .B(_0812_));
 sg13g2_o21ai_1 _3904_ (.B1(_0775_),
    .Y(_0815_),
    .A1(_0754_),
    .A2(_0755_));
 sg13g2_nand2_1 _3905_ (.Y(_0816_),
    .A(_0776_),
    .B(_0815_));
 sg13g2_or3_1 _3906_ (.A(_0733_),
    .B(_0745_),
    .C(_0746_),
    .X(_0817_));
 sg13g2_and2_1 _3907_ (.A(_0747_),
    .B(_0817_),
    .X(_0818_));
 sg13g2_nand2b_1 _3908_ (.Y(_0819_),
    .B(_0818_),
    .A_N(_0816_));
 sg13g2_xor2_1 _3909_ (.B(_0819_),
    .A(_0814_),
    .X(_0820_));
 sg13g2_xnor2_1 _3910_ (.Y(_0821_),
    .A(_0747_),
    .B(_0820_));
 sg13g2_xor2_1 _3911_ (.B(_0818_),
    .A(_0816_),
    .X(_0822_));
 sg13g2_xnor2_1 _3912_ (.Y(_0823_),
    .A(_0754_),
    .B(_0756_));
 sg13g2_nand2_2 _3913_ (.Y(_0824_),
    .A(net737),
    .B(net629));
 sg13g2_nand4_1 _3914_ (.B(net732),
    .C(net629),
    .A(net737),
    .Y(_0825_),
    .D(net624));
 sg13g2_inv_1 _3915_ (.Y(_0826_),
    .A(_0825_));
 sg13g2_o21ai_1 _3916_ (.B1(_0723_),
    .Y(_0827_),
    .A1(_0721_),
    .A2(_0724_));
 sg13g2_nand2b_1 _3917_ (.Y(_0828_),
    .B(_0827_),
    .A_N(_0725_));
 sg13g2_nor2_1 _3918_ (.A(_0825_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_xnor2_1 _3919_ (.Y(_0830_),
    .A(_0826_),
    .B(_0828_));
 sg13g2_nand2_1 _3920_ (.Y(_0831_),
    .A(net718),
    .B(net640));
 sg13g2_nand2_1 _3921_ (.Y(_0832_),
    .A(net723),
    .B(net636));
 sg13g2_nand2_1 _3922_ (.Y(_0833_),
    .A(net723),
    .B(net633));
 sg13g2_xor2_1 _3923_ (.B(_0833_),
    .A(_0736_),
    .X(_0834_));
 sg13g2_nand2b_1 _3924_ (.Y(_0835_),
    .B(_0834_),
    .A_N(_0831_));
 sg13g2_xnor2_1 _3925_ (.Y(_0836_),
    .A(_0831_),
    .B(_0834_));
 sg13g2_and2_1 _3926_ (.A(_0830_),
    .B(_0836_),
    .X(_0837_));
 sg13g2_o21ai_1 _3927_ (.B1(_0835_),
    .Y(_0838_),
    .A1(_0736_),
    .A2(_0833_));
 sg13g2_o21ai_1 _3928_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_0829_),
    .A2(_0837_));
 sg13g2_or3_1 _3929_ (.A(_0829_),
    .B(_0837_),
    .C(_0838_),
    .X(_0840_));
 sg13g2_and2_1 _3930_ (.A(_0839_),
    .B(_0840_),
    .X(_0841_));
 sg13g2_nand2_1 _3931_ (.Y(_0842_),
    .A(_0823_),
    .B(_0841_));
 sg13g2_xnor2_1 _3932_ (.Y(_0843_),
    .A(_0822_),
    .B(_0842_));
 sg13g2_or2_1 _3933_ (.X(_0844_),
    .B(_0839_),
    .A(_0822_));
 sg13g2_a21oi_2 _3934_ (.B1(_0822_),
    .Y(_0845_),
    .A2(_0842_),
    .A1(_0839_));
 sg13g2_nand2_1 _3935_ (.Y(_0846_),
    .A(_0821_),
    .B(_0845_));
 sg13g2_xnor2_1 _3936_ (.Y(_0847_),
    .A(_0821_),
    .B(_0845_));
 sg13g2_nand2_1 _3937_ (.Y(_0848_),
    .A(_0839_),
    .B(_0843_));
 sg13g2_nand2_1 _3938_ (.Y(_0849_),
    .A(net719),
    .B(net640));
 sg13g2_nand2_2 _3939_ (.Y(_0850_),
    .A(net727),
    .B(net636));
 sg13g2_and2_1 _3940_ (.A(net727),
    .B(net633),
    .X(_0851_));
 sg13g2_xnor2_1 _3941_ (.Y(_0852_),
    .A(_0832_),
    .B(_0851_));
 sg13g2_nand2b_1 _3942_ (.Y(_0853_),
    .B(_0852_),
    .A_N(_0849_));
 sg13g2_xnor2_1 _3943_ (.Y(_0854_),
    .A(_0849_),
    .B(_0852_));
 sg13g2_a22oi_1 _3944_ (.Y(_0855_),
    .B1(net624),
    .B2(net737),
    .A2(net629),
    .A1(net732));
 sg13g2_nor2_1 _3945_ (.A(_0826_),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_nand2_1 _3946_ (.Y(_0857_),
    .A(_0854_),
    .B(_0856_));
 sg13g2_o21ai_1 _3947_ (.B1(_0853_),
    .Y(_0858_),
    .A1(_0833_),
    .A2(_0850_));
 sg13g2_nand2b_1 _3948_ (.Y(_0859_),
    .B(_0858_),
    .A_N(_0857_));
 sg13g2_xor2_1 _3949_ (.B(_0858_),
    .A(_0857_),
    .X(_0860_));
 sg13g2_xnor2_1 _3950_ (.Y(_0861_),
    .A(_0830_),
    .B(_0836_));
 sg13g2_nor2_1 _3951_ (.A(_0860_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_xor2_1 _3952_ (.B(_0841_),
    .A(_0823_),
    .X(_0863_));
 sg13g2_nand2_1 _3953_ (.Y(_0864_),
    .A(_0862_),
    .B(_0863_));
 sg13g2_and2_1 _3954_ (.A(net732),
    .B(net636),
    .X(_0865_));
 sg13g2_nand2_1 _3955_ (.Y(_0866_),
    .A(net732),
    .B(net633));
 sg13g2_nand2_1 _3956_ (.Y(_0867_),
    .A(_0850_),
    .B(_0866_));
 sg13g2_xnor2_1 _3957_ (.Y(_0868_),
    .A(_0850_),
    .B(_0866_));
 sg13g2_nor2_1 _3958_ (.A(_2220_),
    .B(_2227_),
    .Y(_0869_));
 sg13g2_xor2_1 _3959_ (.B(_0869_),
    .A(_0868_),
    .X(_0870_));
 sg13g2_a22oi_1 _3960_ (.Y(_0871_),
    .B1(_0867_),
    .B2(_0869_),
    .A2(_0865_),
    .A1(_0851_));
 sg13g2_or3_1 _3961_ (.A(_0824_),
    .B(_0870_),
    .C(_0871_),
    .X(_0872_));
 sg13g2_inv_1 _3962_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_o21ai_1 _3963_ (.B1(_0871_),
    .Y(_0874_),
    .A1(_0824_),
    .A2(_0870_));
 sg13g2_nand2_1 _3964_ (.Y(_0875_),
    .A(_0872_),
    .B(_0874_));
 sg13g2_xnor2_1 _3965_ (.Y(_0876_),
    .A(_0854_),
    .B(_0856_));
 sg13g2_and4_1 _3966_ (.A(net737),
    .B(net640),
    .C(_0865_),
    .D(_0868_),
    .X(_0877_));
 sg13g2_a21oi_1 _3967_ (.A1(net727),
    .A2(net640),
    .Y(_0878_),
    .B1(_0865_));
 sg13g2_nand2_1 _3968_ (.Y(_0879_),
    .A(net737),
    .B(net633));
 sg13g2_nand3_1 _3969_ (.B(net640),
    .C(_0865_),
    .A(net727),
    .Y(_0880_));
 sg13g2_a21oi_1 _3970_ (.A1(_0879_),
    .A2(_0880_),
    .Y(_0881_),
    .B1(_0878_));
 sg13g2_nand2_1 _3971_ (.Y(_0882_),
    .A(_0877_),
    .B(_0881_));
 sg13g2_xor2_1 _3972_ (.B(_0870_),
    .A(_0824_),
    .X(_0883_));
 sg13g2_o21ai_1 _3973_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0877_),
    .A2(_0881_));
 sg13g2_a22oi_1 _3974_ (.Y(_0885_),
    .B1(_0882_),
    .B2(_0884_),
    .A2(_0876_),
    .A1(_0875_));
 sg13g2_o21ai_1 _3975_ (.B1(_0872_),
    .Y(_0886_),
    .A1(_0875_),
    .A2(_0876_));
 sg13g2_nand2_1 _3976_ (.Y(_0887_),
    .A(_0860_),
    .B(_0861_));
 sg13g2_o21ai_1 _3977_ (.B1(_0887_),
    .Y(_0888_),
    .A1(_0885_),
    .A2(_0886_));
 sg13g2_nor2_1 _3978_ (.A(_0862_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_a21oi_1 _3979_ (.A1(_0873_),
    .A2(_0885_),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_nor2_1 _3980_ (.A(_0862_),
    .B(_0863_),
    .Y(_0891_));
 sg13g2_o21ai_1 _3981_ (.B1(_0891_),
    .Y(_0892_),
    .A1(_0859_),
    .A2(_0890_));
 sg13g2_nand3_1 _3982_ (.B(_0864_),
    .C(_0890_),
    .A(_0859_),
    .Y(_0893_));
 sg13g2_nand4_1 _3983_ (.B(_0848_),
    .C(_0892_),
    .A(_0844_),
    .Y(_0894_),
    .D(_0893_));
 sg13g2_xor2_1 _3984_ (.B(_0894_),
    .A(_0847_),
    .X(_0895_));
 sg13g2_o21ai_1 _3985_ (.B1(net792),
    .Y(_0896_),
    .A1(net609),
    .A2(_0895_));
 sg13g2_a21oi_1 _3986_ (.A1(net609),
    .A2(_2202_),
    .Y(_0173_),
    .B1(_0896_));
 sg13g2_a21oi_2 _3987_ (.B1(_0814_),
    .Y(_0897_),
    .A2(_0819_),
    .A1(_0747_));
 sg13g2_a21o_1 _3988_ (.A2(_0779_),
    .A1(_0752_),
    .B1(_0778_),
    .X(_0898_));
 sg13g2_or2_1 _3989_ (.X(_0899_),
    .B(_0785_),
    .A(_0783_));
 sg13g2_nand2_1 _3990_ (.Y(_0900_),
    .A(_0795_),
    .B(_0798_));
 sg13g2_xor2_1 _3991_ (.B(_0900_),
    .A(_0811_),
    .X(_0901_));
 sg13g2_and2_1 _3992_ (.A(_0899_),
    .B(_0901_),
    .X(_0902_));
 sg13g2_xnor2_1 _3993_ (.Y(_0903_),
    .A(_0899_),
    .B(_0901_));
 sg13g2_nand2_2 _3994_ (.Y(_0904_),
    .A(net739),
    .B(net702));
 sg13g2_nor2_1 _3995_ (.A(_0800_),
    .B(_0803_),
    .Y(_0905_));
 sg13g2_nand2_1 _3996_ (.Y(_0906_),
    .A(net725),
    .B(net617));
 sg13g2_nand2_1 _3997_ (.Y(_0907_),
    .A(net729),
    .B(net704));
 sg13g2_and4_1 _3998_ (.A(net735),
    .B(net729),
    .C(net611),
    .D(net704),
    .X(_0908_));
 sg13g2_a22oi_1 _3999_ (.Y(_0909_),
    .B1(net704),
    .B2(net735),
    .A2(net611),
    .A1(net729));
 sg13g2_nor2_1 _4000_ (.A(_0908_),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_nor3_1 _4001_ (.A(_0906_),
    .B(_0908_),
    .C(_0909_),
    .Y(_0911_));
 sg13g2_xnor2_1 _4002_ (.Y(_0912_),
    .A(_0906_),
    .B(_0910_));
 sg13g2_nand2b_1 _4003_ (.Y(_0913_),
    .B(_0912_),
    .A_N(_0905_));
 sg13g2_xnor2_1 _4004_ (.Y(_0914_),
    .A(_0905_),
    .B(_0912_));
 sg13g2_nor2b_1 _4005_ (.A(_0805_),
    .B_N(_0914_),
    .Y(_0915_));
 sg13g2_xnor2_1 _4006_ (.Y(_0916_),
    .A(_0805_),
    .B(_0914_));
 sg13g2_nand2_1 _4007_ (.Y(_0917_),
    .A(net758),
    .B(net641));
 sg13g2_nand2_1 _4008_ (.Y(_0918_),
    .A(net762),
    .B(net634));
 sg13g2_nand2_1 _4009_ (.Y(_0919_),
    .A(net762),
    .B(net637));
 sg13g2_xor2_1 _4010_ (.B(_0919_),
    .A(_0782_),
    .X(_0920_));
 sg13g2_nand2b_1 _4011_ (.Y(_0921_),
    .B(_0920_),
    .A_N(_0917_));
 sg13g2_xor2_1 _4012_ (.B(_0920_),
    .A(_0917_),
    .X(_0922_));
 sg13g2_nand2b_2 _4013_ (.Y(_0923_),
    .B(_0793_),
    .A_N(_0791_));
 sg13g2_nand2_1 _4014_ (.Y(_0924_),
    .A(net712),
    .B(net631));
 sg13g2_nand2_1 _4015_ (.Y(_0925_),
    .A(net717),
    .B(net622));
 sg13g2_nand2_2 _4016_ (.Y(_0926_),
    .A(net717),
    .B(net628));
 sg13g2_or2_1 _4017_ (.X(_0927_),
    .B(_0926_),
    .A(_0790_));
 sg13g2_and2_1 _4018_ (.A(_0790_),
    .B(_0926_),
    .X(_0928_));
 sg13g2_xor2_1 _4019_ (.B(_0926_),
    .A(_0790_),
    .X(_0929_));
 sg13g2_xnor2_1 _4020_ (.Y(_0930_),
    .A(_0924_),
    .B(_0929_));
 sg13g2_nand2_1 _4021_ (.Y(_0931_),
    .A(_0923_),
    .B(_0930_));
 sg13g2_xnor2_1 _4022_ (.Y(_0932_),
    .A(_0923_),
    .B(_0930_));
 sg13g2_xor2_1 _4023_ (.B(_0932_),
    .A(_0922_),
    .X(_0933_));
 sg13g2_xnor2_1 _4024_ (.Y(_0934_),
    .A(_0916_),
    .B(_0933_));
 sg13g2_nor2_1 _4025_ (.A(_0808_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_xnor2_1 _4026_ (.Y(_0936_),
    .A(_0808_),
    .B(_0934_));
 sg13g2_or2_1 _4027_ (.X(_0937_),
    .B(_0936_),
    .A(_0904_));
 sg13g2_xor2_1 _4028_ (.B(_0936_),
    .A(_0904_),
    .X(_0938_));
 sg13g2_nor2b_1 _4029_ (.A(_0903_),
    .B_N(_0938_),
    .Y(_0939_));
 sg13g2_xnor2_1 _4030_ (.Y(_0940_),
    .A(_0903_),
    .B(_0938_));
 sg13g2_xnor2_1 _4031_ (.Y(_0941_),
    .A(_0813_),
    .B(_0940_));
 sg13g2_nor2b_1 _4032_ (.A(_0941_),
    .B_N(_0898_),
    .Y(_0942_));
 sg13g2_xnor2_1 _4033_ (.Y(_0943_),
    .A(_0898_),
    .B(_0941_));
 sg13g2_nor2_1 _4034_ (.A(_0897_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_inv_1 _4035_ (.Y(_0945_),
    .A(_0944_));
 sg13g2_xor2_1 _4036_ (.B(_0943_),
    .A(_0897_),
    .X(_0946_));
 sg13g2_o21ai_1 _4037_ (.B1(_0846_),
    .Y(_0947_),
    .A1(_0847_),
    .A2(_0894_));
 sg13g2_xnor2_1 _4038_ (.Y(_0948_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_o21ai_1 _4039_ (.B1(net792),
    .Y(_0949_),
    .A1(net674),
    .A2(net260));
 sg13g2_a21oi_1 _4040_ (.A1(net674),
    .A2(_0948_),
    .Y(_0174_),
    .B1(net261));
 sg13g2_a21oi_1 _4041_ (.A1(_0813_),
    .A2(_0940_),
    .Y(_0950_),
    .B1(_0942_));
 sg13g2_a21o_1 _4042_ (.A2(_0900_),
    .A1(_0811_),
    .B1(_0902_),
    .X(_0951_));
 sg13g2_o21ai_1 _4043_ (.B1(_0921_),
    .Y(_0952_),
    .A1(_0782_),
    .A2(_0919_));
 sg13g2_o21ai_1 _4044_ (.B1(_0931_),
    .Y(_0953_),
    .A1(_0922_),
    .A2(_0932_));
 sg13g2_xor2_1 _4045_ (.B(_0953_),
    .A(_0935_),
    .X(_0954_));
 sg13g2_and2_1 _4046_ (.A(_0952_),
    .B(_0954_),
    .X(_0955_));
 sg13g2_xnor2_1 _4047_ (.Y(_0956_),
    .A(_0952_),
    .B(_0954_));
 sg13g2_nand2_2 _4048_ (.Y(_0957_),
    .A(net735),
    .B(net699));
 sg13g2_nor2_2 _4049_ (.A(_0904_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_a22oi_1 _4050_ (.Y(_0959_),
    .B1(net700),
    .B2(net738),
    .A2(net702),
    .A1(net733));
 sg13g2_nor2_1 _4051_ (.A(_0958_),
    .B(_0959_),
    .Y(_0960_));
 sg13g2_nor2_1 _4052_ (.A(_0908_),
    .B(_0911_),
    .Y(_0961_));
 sg13g2_nand2_1 _4053_ (.Y(_0962_),
    .A(net720),
    .B(net617));
 sg13g2_nand2_1 _4054_ (.Y(_0963_),
    .A(net724),
    .B(net704));
 sg13g2_nand2_1 _4055_ (.Y(_0964_),
    .A(net725),
    .B(net611));
 sg13g2_or2_1 _4056_ (.X(_0965_),
    .B(_0964_),
    .A(_0907_));
 sg13g2_xor2_1 _4057_ (.B(_0964_),
    .A(_0907_),
    .X(_0966_));
 sg13g2_nand2b_1 _4058_ (.Y(_0967_),
    .B(_0966_),
    .A_N(_0962_));
 sg13g2_xnor2_1 _4059_ (.Y(_0968_),
    .A(_0962_),
    .B(_0966_));
 sg13g2_nand2b_1 _4060_ (.Y(_0969_),
    .B(_0968_),
    .A_N(_0961_));
 sg13g2_inv_1 _4061_ (.Y(_0970_),
    .A(_0969_));
 sg13g2_xnor2_1 _4062_ (.Y(_0971_),
    .A(_0961_),
    .B(_0968_));
 sg13g2_nor2b_1 _4063_ (.A(_0913_),
    .B_N(_0971_),
    .Y(_0972_));
 sg13g2_xnor2_1 _4064_ (.Y(_0973_),
    .A(_0913_),
    .B(_0971_));
 sg13g2_nand2_1 _4065_ (.Y(_0974_),
    .A(net755),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[23] ));
 sg13g2_nand2_1 _4066_ (.Y(_0975_),
    .A(net758),
    .B(net634));
 sg13g2_nand2_1 _4067_ (.Y(_0976_),
    .A(net758),
    .B(net638));
 sg13g2_xor2_1 _4068_ (.B(_0976_),
    .A(_0918_),
    .X(_0977_));
 sg13g2_nand2b_1 _4069_ (.Y(_0978_),
    .B(_0977_),
    .A_N(_0974_));
 sg13g2_xnor2_1 _4070_ (.Y(_0979_),
    .A(_0974_),
    .B(_0977_));
 sg13g2_inv_1 _4071_ (.Y(_0980_),
    .A(_0979_));
 sg13g2_o21ai_1 _4072_ (.B1(_0927_),
    .Y(_0981_),
    .A1(_0924_),
    .A2(_0928_));
 sg13g2_nand2_1 _4073_ (.Y(_0982_),
    .A(net710),
    .B(net631));
 sg13g2_nand2_2 _4074_ (.Y(_0983_),
    .A(net714),
    .B(net622));
 sg13g2_nand2_1 _4075_ (.Y(_0984_),
    .A(net714),
    .B(net628));
 sg13g2_or2_1 _4076_ (.X(_0985_),
    .B(_0983_),
    .A(_0926_));
 sg13g2_xnor2_1 _4077_ (.Y(_0986_),
    .A(_0925_),
    .B(_0984_));
 sg13g2_xor2_1 _4078_ (.B(_0986_),
    .A(_0982_),
    .X(_0987_));
 sg13g2_nand2_1 _4079_ (.Y(_0988_),
    .A(_0981_),
    .B(_0987_));
 sg13g2_xnor2_1 _4080_ (.Y(_0989_),
    .A(_0981_),
    .B(_0987_));
 sg13g2_xnor2_1 _4081_ (.Y(_0990_),
    .A(_0979_),
    .B(_0989_));
 sg13g2_xnor2_1 _4082_ (.Y(_0991_),
    .A(_0973_),
    .B(_0990_));
 sg13g2_a21oi_1 _4083_ (.A1(_0916_),
    .A2(_0933_),
    .Y(_0992_),
    .B1(_0915_));
 sg13g2_nor2_1 _4084_ (.A(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_xnor2_1 _4085_ (.Y(_0994_),
    .A(_0991_),
    .B(_0992_));
 sg13g2_or3_1 _4086_ (.A(_0958_),
    .B(_0959_),
    .C(_0994_),
    .X(_0995_));
 sg13g2_xor2_1 _4087_ (.B(_0994_),
    .A(_0960_),
    .X(_0996_));
 sg13g2_nor2_1 _4088_ (.A(_0937_),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_xor2_1 _4089_ (.B(_0996_),
    .A(_0937_),
    .X(_0998_));
 sg13g2_nor2b_1 _4090_ (.A(_0956_),
    .B_N(_0998_),
    .Y(_0999_));
 sg13g2_xnor2_1 _4091_ (.Y(_1000_),
    .A(_0956_),
    .B(_0998_));
 sg13g2_xnor2_1 _4092_ (.Y(_1001_),
    .A(_0939_),
    .B(_1000_));
 sg13g2_nor2b_1 _4093_ (.A(_1001_),
    .B_N(_0951_),
    .Y(_1002_));
 sg13g2_xor2_1 _4094_ (.B(_1001_),
    .A(_0951_),
    .X(_1003_));
 sg13g2_nor2_1 _4095_ (.A(_0950_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_xor2_1 _4096_ (.B(_1003_),
    .A(_0950_),
    .X(_1005_));
 sg13g2_a22oi_1 _4097_ (.Y(_1006_),
    .B1(_0897_),
    .B2(_0943_),
    .A2(_0845_),
    .A1(_0821_));
 sg13g2_o21ai_1 _4098_ (.B1(_1006_),
    .Y(_1007_),
    .A1(_0847_),
    .A2(_0894_));
 sg13g2_a21oi_1 _4099_ (.A1(_0945_),
    .A2(_1007_),
    .Y(_1008_),
    .B1(_1005_));
 sg13g2_and3_1 _4100_ (.X(_1009_),
    .A(_0945_),
    .B(_1005_),
    .C(_1007_));
 sg13g2_or2_1 _4101_ (.X(_1010_),
    .B(_1009_),
    .A(_1008_));
 sg13g2_o21ai_1 _4102_ (.B1(net793),
    .Y(_1011_),
    .A1(net674),
    .A2(net218));
 sg13g2_a21oi_1 _4103_ (.A1(net674),
    .A2(_1010_),
    .Y(_0175_),
    .B1(net219));
 sg13g2_a21oi_1 _4104_ (.A1(_0939_),
    .A2(_1000_),
    .Y(_1012_),
    .B1(_1002_));
 sg13g2_a21oi_1 _4105_ (.A1(_0935_),
    .A2(_0953_),
    .Y(_1013_),
    .B1(_0955_));
 sg13g2_nor2_1 _4106_ (.A(_0997_),
    .B(_0999_),
    .Y(_1014_));
 sg13g2_o21ai_1 _4107_ (.B1(_0978_),
    .Y(_1015_),
    .A1(_0918_),
    .A2(_0976_));
 sg13g2_o21ai_1 _4108_ (.B1(_0988_),
    .Y(_1016_),
    .A1(_0980_),
    .A2(_0989_));
 sg13g2_xor2_1 _4109_ (.B(_1016_),
    .A(_0993_),
    .X(_1017_));
 sg13g2_and2_1 _4110_ (.A(_1015_),
    .B(_1017_),
    .X(_1018_));
 sg13g2_xnor2_1 _4111_ (.Y(_1019_),
    .A(_1015_),
    .B(_1017_));
 sg13g2_inv_1 _4112_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_nand2_1 _4113_ (.Y(_1021_),
    .A(net729),
    .B(net702));
 sg13g2_nand2_1 _4114_ (.Y(_1022_),
    .A(net739),
    .B(net696));
 sg13g2_or2_1 _4115_ (.X(_1023_),
    .B(_1022_),
    .A(_0957_));
 sg13g2_and2_1 _4116_ (.A(_0957_),
    .B(_1022_),
    .X(_1024_));
 sg13g2_xor2_1 _4117_ (.B(_1022_),
    .A(_0957_),
    .X(_1025_));
 sg13g2_xnor2_1 _4118_ (.Y(_1026_),
    .A(_1021_),
    .B(_1025_));
 sg13g2_inv_1 _4119_ (.Y(_1027_),
    .A(_1026_));
 sg13g2_and2_1 _4120_ (.A(_0965_),
    .B(_0967_),
    .X(_1028_));
 sg13g2_nand2_1 _4121_ (.Y(_1029_),
    .A(net717),
    .B(net617));
 sg13g2_nand2_1 _4122_ (.Y(_1030_),
    .A(net720),
    .B(net611));
 sg13g2_or2_1 _4123_ (.X(_1031_),
    .B(_1030_),
    .A(_0963_));
 sg13g2_xnor2_1 _4124_ (.Y(_1032_),
    .A(_0963_),
    .B(_1030_));
 sg13g2_xor2_1 _4125_ (.B(_1032_),
    .A(_1029_),
    .X(_1033_));
 sg13g2_nand2_1 _4126_ (.Y(_1034_),
    .A(_0958_),
    .B(_1033_));
 sg13g2_nor2_1 _4127_ (.A(_0958_),
    .B(_1033_),
    .Y(_1035_));
 sg13g2_xor2_1 _4128_ (.B(_1033_),
    .A(_0958_),
    .X(_1036_));
 sg13g2_xnor2_1 _4129_ (.Y(_1037_),
    .A(_1028_),
    .B(_1036_));
 sg13g2_nand2_1 _4130_ (.Y(_1038_),
    .A(_0970_),
    .B(_1037_));
 sg13g2_xnor2_1 _4131_ (.Y(_1039_),
    .A(_0970_),
    .B(_1037_));
 sg13g2_nand2_1 _4132_ (.Y(_1040_),
    .A(net751),
    .B(net641));
 sg13g2_nand2_1 _4133_ (.Y(_1041_),
    .A(net755),
    .B(net635));
 sg13g2_nand2_1 _4134_ (.Y(_1042_),
    .A(net755),
    .B(net638));
 sg13g2_xor2_1 _4135_ (.B(_1042_),
    .A(_0975_),
    .X(_1043_));
 sg13g2_nand2b_1 _4136_ (.Y(_1044_),
    .B(_1043_),
    .A_N(_1040_));
 sg13g2_xnor2_1 _4137_ (.Y(_1045_),
    .A(_1040_),
    .B(_1043_));
 sg13g2_inv_1 _4138_ (.Y(_1046_),
    .A(_1045_));
 sg13g2_o21ai_1 _4139_ (.B1(_0985_),
    .Y(_1047_),
    .A1(_0982_),
    .A2(_0986_));
 sg13g2_nand2_1 _4140_ (.Y(_1048_),
    .A(net760),
    .B(net631));
 sg13g2_nand2_1 _4141_ (.Y(_1049_),
    .A(net710),
    .B(net621));
 sg13g2_nand2_1 _4142_ (.Y(_1050_),
    .A(net710),
    .B(net628));
 sg13g2_xor2_1 _4143_ (.B(_1050_),
    .A(_0983_),
    .X(_1051_));
 sg13g2_nand2b_1 _4144_ (.Y(_1052_),
    .B(_1051_),
    .A_N(_1048_));
 sg13g2_xnor2_1 _4145_ (.Y(_1053_),
    .A(_1048_),
    .B(_1051_));
 sg13g2_nand2_1 _4146_ (.Y(_1054_),
    .A(_1047_),
    .B(_1053_));
 sg13g2_xnor2_1 _4147_ (.Y(_1055_),
    .A(_1047_),
    .B(_1053_));
 sg13g2_xnor2_1 _4148_ (.Y(_1056_),
    .A(_1046_),
    .B(_1055_));
 sg13g2_xnor2_1 _4149_ (.Y(_1057_),
    .A(_1039_),
    .B(_1056_));
 sg13g2_a21oi_1 _4150_ (.A1(_0973_),
    .A2(_0990_),
    .Y(_1058_),
    .B1(_0972_));
 sg13g2_nor2_1 _4151_ (.A(_1057_),
    .B(_1058_),
    .Y(_1059_));
 sg13g2_xnor2_1 _4152_ (.Y(_1060_),
    .A(_1057_),
    .B(_1058_));
 sg13g2_or2_1 _4153_ (.X(_1061_),
    .B(_1060_),
    .A(_1027_));
 sg13g2_xnor2_1 _4154_ (.Y(_1062_),
    .A(_1027_),
    .B(_1060_));
 sg13g2_nor2_1 _4155_ (.A(_0995_),
    .B(_1062_),
    .Y(_1063_));
 sg13g2_xor2_1 _4156_ (.B(_1062_),
    .A(_0995_),
    .X(_1064_));
 sg13g2_xnor2_1 _4157_ (.Y(_1065_),
    .A(_1019_),
    .B(_1064_));
 sg13g2_nand2b_1 _4158_ (.Y(_1066_),
    .B(_1065_),
    .A_N(_1014_));
 sg13g2_nor2b_1 _4159_ (.A(_1065_),
    .B_N(_1014_),
    .Y(_1067_));
 sg13g2_xnor2_1 _4160_ (.Y(_1068_),
    .A(_1014_),
    .B(_1065_));
 sg13g2_xnor2_1 _4161_ (.Y(_1069_),
    .A(_1013_),
    .B(_1068_));
 sg13g2_nand2b_1 _4162_ (.Y(_1070_),
    .B(_1069_),
    .A_N(_1012_));
 sg13g2_xnor2_1 _4163_ (.Y(_1071_),
    .A(_1012_),
    .B(_1069_));
 sg13g2_nor3_1 _4164_ (.A(_1004_),
    .B(_1009_),
    .C(_1071_),
    .Y(_1072_));
 sg13g2_o21ai_1 _4165_ (.B1(_1071_),
    .Y(_1073_),
    .A1(_1004_),
    .A2(_1009_));
 sg13g2_nor2b_2 _4166_ (.A(_1072_),
    .B_N(_1073_),
    .Y(_1074_));
 sg13g2_o21ai_1 _4167_ (.B1(net793),
    .Y(_1075_),
    .A1(net609),
    .A2(_1074_));
 sg13g2_a21oi_1 _4168_ (.A1(net609),
    .A2(_2201_),
    .Y(_0176_),
    .B1(_1075_));
 sg13g2_nand2_1 _4169_ (.Y(_1076_),
    .A(_1070_),
    .B(_1073_));
 sg13g2_a21o_1 _4170_ (.A2(_1016_),
    .A1(_0993_),
    .B1(_1018_),
    .X(_1077_));
 sg13g2_a21oi_1 _4171_ (.A1(_1020_),
    .A2(_1064_),
    .Y(_1078_),
    .B1(_1063_));
 sg13g2_o21ai_1 _4172_ (.B1(_1044_),
    .Y(_1079_),
    .A1(_0975_),
    .A2(_1042_));
 sg13g2_o21ai_1 _4173_ (.B1(_1054_),
    .Y(_1080_),
    .A1(_1046_),
    .A2(_1055_));
 sg13g2_xor2_1 _4174_ (.B(_1080_),
    .A(_1059_),
    .X(_1081_));
 sg13g2_and2_1 _4175_ (.A(_1079_),
    .B(_1081_),
    .X(_1082_));
 sg13g2_xor2_1 _4176_ (.B(_1081_),
    .A(_1079_),
    .X(_1083_));
 sg13g2_nand2_2 _4177_ (.Y(_1084_),
    .A(net739),
    .B(net692));
 sg13g2_nand2_1 _4178_ (.Y(_1085_),
    .A(net724),
    .B(net701));
 sg13g2_nand2_1 _4179_ (.Y(_1086_),
    .A(net730),
    .B(net694));
 sg13g2_nor2_1 _4180_ (.A(_0957_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_nand4_1 _4181_ (.B(net730),
    .C(net699),
    .A(net735),
    .Y(_1088_),
    .D(net695));
 sg13g2_a22oi_1 _4182_ (.Y(_1089_),
    .B1(net695),
    .B2(net735),
    .A2(net699),
    .A1(net730));
 sg13g2_nor2_1 _4183_ (.A(_1087_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_xnor2_1 _4184_ (.Y(_1091_),
    .A(_1085_),
    .B(_1090_));
 sg13g2_nand2b_1 _4185_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_1084_));
 sg13g2_xnor2_1 _4186_ (.Y(_1093_),
    .A(_1084_),
    .B(_1091_));
 sg13g2_o21ai_1 _4187_ (.B1(_1034_),
    .Y(_1094_),
    .A1(_1028_),
    .A2(_1035_));
 sg13g2_o21ai_1 _4188_ (.B1(_1031_),
    .Y(_1095_),
    .A1(_1029_),
    .A2(_1032_));
 sg13g2_o21ai_1 _4189_ (.B1(_1023_),
    .Y(_1096_),
    .A1(_1021_),
    .A2(_1024_));
 sg13g2_nand2_1 _4190_ (.Y(_1097_),
    .A(net714),
    .B(net616));
 sg13g2_and4_1 _4191_ (.A(net720),
    .B(net716),
    .C(net612),
    .D(net704),
    .X(_1098_));
 sg13g2_nand4_1 _4192_ (.B(net716),
    .C(net612),
    .A(net721),
    .Y(_1099_),
    .D(net705));
 sg13g2_a22oi_1 _4193_ (.Y(_1100_),
    .B1(net705),
    .B2(net721),
    .A2(net612),
    .A1(net716));
 sg13g2_nor3_1 _4194_ (.A(_1097_),
    .B(_1098_),
    .C(_1100_),
    .Y(_1101_));
 sg13g2_o21ai_1 _4195_ (.B1(_1097_),
    .Y(_1102_),
    .A1(_1098_),
    .A2(_1100_));
 sg13g2_nor2b_1 _4196_ (.A(_1101_),
    .B_N(_1102_),
    .Y(_1103_));
 sg13g2_and2_1 _4197_ (.A(_1096_),
    .B(_1103_),
    .X(_1104_));
 sg13g2_xor2_1 _4198_ (.B(_1103_),
    .A(_1096_),
    .X(_1105_));
 sg13g2_xnor2_1 _4199_ (.Y(_1106_),
    .A(_1095_),
    .B(_1105_));
 sg13g2_nand2b_1 _4200_ (.Y(_1107_),
    .B(_1094_),
    .A_N(_1106_));
 sg13g2_xor2_1 _4201_ (.B(_1106_),
    .A(_1094_),
    .X(_1108_));
 sg13g2_nand2_1 _4202_ (.Y(_1109_),
    .A(net749),
    .B(net641));
 sg13g2_nand2_1 _4203_ (.Y(_1110_),
    .A(net751),
    .B(net635));
 sg13g2_nand2_1 _4204_ (.Y(_1111_),
    .A(net751),
    .B(net638));
 sg13g2_xor2_1 _4205_ (.B(_1111_),
    .A(_1041_),
    .X(_1112_));
 sg13g2_nand2b_1 _4206_ (.Y(_1113_),
    .B(_1112_),
    .A_N(_1109_));
 sg13g2_xnor2_1 _4207_ (.Y(_1114_),
    .A(_1109_),
    .B(_1112_));
 sg13g2_inv_1 _4208_ (.Y(_1115_),
    .A(_1114_));
 sg13g2_o21ai_1 _4209_ (.B1(_1052_),
    .Y(_1116_),
    .A1(_0983_),
    .A2(_1050_));
 sg13g2_nand2_1 _4210_ (.Y(_1117_),
    .A(net758),
    .B(net630));
 sg13g2_nand2_1 _4211_ (.Y(_1118_),
    .A(net760),
    .B(net621));
 sg13g2_nand2_1 _4212_ (.Y(_1119_),
    .A(net760),
    .B(net628));
 sg13g2_xor2_1 _4213_ (.B(_1119_),
    .A(_1049_),
    .X(_1120_));
 sg13g2_nand2b_1 _4214_ (.Y(_1121_),
    .B(_1120_),
    .A_N(_1117_));
 sg13g2_xnor2_1 _4215_ (.Y(_1122_),
    .A(_1117_),
    .B(_1120_));
 sg13g2_nand2_1 _4216_ (.Y(_1123_),
    .A(_1116_),
    .B(_1122_));
 sg13g2_xnor2_1 _4217_ (.Y(_1124_),
    .A(_1116_),
    .B(_1122_));
 sg13g2_xnor2_1 _4218_ (.Y(_1125_),
    .A(_1115_),
    .B(_1124_));
 sg13g2_xor2_1 _4219_ (.B(_1125_),
    .A(_1108_),
    .X(_1126_));
 sg13g2_o21ai_1 _4220_ (.B1(_1038_),
    .Y(_1127_),
    .A1(_1039_),
    .A2(_1056_));
 sg13g2_nand2_1 _4221_ (.Y(_1128_),
    .A(_1126_),
    .B(_1127_));
 sg13g2_xor2_1 _4222_ (.B(_1127_),
    .A(_1126_),
    .X(_1129_));
 sg13g2_nand2_1 _4223_ (.Y(_1130_),
    .A(_1093_),
    .B(_1129_));
 sg13g2_xnor2_1 _4224_ (.Y(_1131_),
    .A(_1093_),
    .B(_1129_));
 sg13g2_nor2_1 _4225_ (.A(_1061_),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_xor2_1 _4226_ (.B(_1131_),
    .A(_1061_),
    .X(_1133_));
 sg13g2_xor2_1 _4227_ (.B(_1133_),
    .A(_1083_),
    .X(_1134_));
 sg13g2_nor2b_1 _4228_ (.A(_1078_),
    .B_N(_1134_),
    .Y(_1135_));
 sg13g2_xnor2_1 _4229_ (.Y(_1136_),
    .A(_1078_),
    .B(_1134_));
 sg13g2_xnor2_1 _4230_ (.Y(_1137_),
    .A(_1077_),
    .B(_1136_));
 sg13g2_o21ai_1 _4231_ (.B1(_1066_),
    .Y(_1138_),
    .A1(_1013_),
    .A2(_1067_));
 sg13g2_nor2b_1 _4232_ (.A(_1137_),
    .B_N(_1138_),
    .Y(_1139_));
 sg13g2_xnor2_1 _4233_ (.Y(_1140_),
    .A(_1137_),
    .B(_1138_));
 sg13g2_xnor2_1 _4234_ (.Y(_1141_),
    .A(_1076_),
    .B(_1140_));
 sg13g2_o21ai_1 _4235_ (.B1(net792),
    .Y(_1142_),
    .A1(net674),
    .A2(net223));
 sg13g2_a21oi_1 _4236_ (.A1(net674),
    .A2(_1141_),
    .Y(_0177_),
    .B1(net224));
 sg13g2_a21oi_1 _4237_ (.A1(_1077_),
    .A2(_1136_),
    .Y(_1143_),
    .B1(_1135_));
 sg13g2_a21o_1 _4238_ (.A2(_1080_),
    .A1(_1059_),
    .B1(_1082_),
    .X(_1144_));
 sg13g2_a21oi_1 _4239_ (.A1(_1083_),
    .A2(_1133_),
    .Y(_1145_),
    .B1(_1132_));
 sg13g2_o21ai_1 _4240_ (.B1(_1113_),
    .Y(_1146_),
    .A1(_1041_),
    .A2(_1111_));
 sg13g2_inv_1 _4241_ (.Y(_1147_),
    .A(_1146_));
 sg13g2_o21ai_1 _4242_ (.B1(_1123_),
    .Y(_1148_),
    .A1(_1115_),
    .A2(_1124_));
 sg13g2_nand3_1 _4243_ (.B(_1127_),
    .C(_1148_),
    .A(_1126_),
    .Y(_1149_));
 sg13g2_xor2_1 _4244_ (.B(_1148_),
    .A(_1128_),
    .X(_1150_));
 sg13g2_xnor2_1 _4245_ (.Y(_1151_),
    .A(_1147_),
    .B(_1150_));
 sg13g2_nand2_2 _4246_ (.Y(_1152_),
    .A(net735),
    .B(net691));
 sg13g2_or2_1 _4247_ (.X(_1153_),
    .B(_1152_),
    .A(_1084_));
 sg13g2_inv_1 _4248_ (.Y(_1154_),
    .A(_1153_));
 sg13g2_a22oi_1 _4249_ (.Y(_1155_),
    .B1(net691),
    .B2(net739),
    .A2(net692),
    .A1(net735));
 sg13g2_nor2_1 _4250_ (.A(_1154_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_nand2_1 _4251_ (.Y(_1157_),
    .A(net721),
    .B(net701));
 sg13g2_nand2_1 _4252_ (.Y(_1158_),
    .A(net724),
    .B(net698));
 sg13g2_nand4_1 _4253_ (.B(net724),
    .C(net698),
    .A(net730),
    .Y(_1159_),
    .D(net694));
 sg13g2_a22oi_1 _4254_ (.Y(_1160_),
    .B1(net694),
    .B2(net730),
    .A2(net698),
    .A1(net724));
 sg13g2_xor2_1 _4255_ (.B(_1158_),
    .A(_1086_),
    .X(_1161_));
 sg13g2_xnor2_1 _4256_ (.Y(_1162_),
    .A(_1157_),
    .B(_1161_));
 sg13g2_nand2_1 _4257_ (.Y(_1163_),
    .A(_1156_),
    .B(_1162_));
 sg13g2_xnor2_1 _4258_ (.Y(_1164_),
    .A(_1156_),
    .B(_1162_));
 sg13g2_nor2_1 _4259_ (.A(_1092_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_xor2_1 _4260_ (.B(_1164_),
    .A(_1092_),
    .X(_1166_));
 sg13g2_a21o_1 _4261_ (.A2(_1105_),
    .A1(_1095_),
    .B1(_1104_),
    .X(_1167_));
 sg13g2_o21ai_1 _4262_ (.B1(_1099_),
    .Y(_1168_),
    .A1(_1097_),
    .A2(_1100_));
 sg13g2_inv_1 _4263_ (.Y(_1169_),
    .A(_1168_));
 sg13g2_o21ai_1 _4264_ (.B1(_1088_),
    .Y(_1170_),
    .A1(_1085_),
    .A2(_1089_));
 sg13g2_nand2_1 _4265_ (.Y(_1171_),
    .A(net709),
    .B(net616));
 sg13g2_and4_1 _4266_ (.A(net716),
    .B(net713),
    .C(net612),
    .D(net705),
    .X(_1172_));
 sg13g2_a22oi_1 _4267_ (.Y(_1173_),
    .B1(net705),
    .B2(net716),
    .A2(net612),
    .A1(net713));
 sg13g2_or3_1 _4268_ (.A(_1171_),
    .B(_1172_),
    .C(_1173_),
    .X(_1174_));
 sg13g2_o21ai_1 _4269_ (.B1(_1171_),
    .Y(_1175_),
    .A1(_1172_),
    .A2(_1173_));
 sg13g2_and3_1 _4270_ (.X(_1176_),
    .A(_1170_),
    .B(_1174_),
    .C(_1175_));
 sg13g2_nand3_1 _4271_ (.B(_1174_),
    .C(_1175_),
    .A(_1170_),
    .Y(_1177_));
 sg13g2_a21oi_1 _4272_ (.A1(_1174_),
    .A2(_1175_),
    .Y(_1178_),
    .B1(_1170_));
 sg13g2_nor2_1 _4273_ (.A(_1176_),
    .B(_1178_),
    .Y(_1179_));
 sg13g2_xnor2_1 _4274_ (.Y(_1180_),
    .A(_1168_),
    .B(_1179_));
 sg13g2_nand2b_1 _4275_ (.Y(_1181_),
    .B(_1167_),
    .A_N(_1180_));
 sg13g2_xor2_1 _4276_ (.B(_1180_),
    .A(_1167_),
    .X(_1182_));
 sg13g2_nand2_1 _4277_ (.Y(_1183_),
    .A(net747),
    .B(net641));
 sg13g2_nand2_1 _4278_ (.Y(_1184_),
    .A(net750),
    .B(net635));
 sg13g2_nand2_1 _4279_ (.Y(_1185_),
    .A(net749),
    .B(net638));
 sg13g2_xor2_1 _4280_ (.B(_1185_),
    .A(_1110_),
    .X(_1186_));
 sg13g2_nand2b_1 _4281_ (.Y(_1187_),
    .B(_1186_),
    .A_N(_1183_));
 sg13g2_xnor2_1 _4282_ (.Y(_1188_),
    .A(_1183_),
    .B(_1186_));
 sg13g2_inv_1 _4283_ (.Y(_1189_),
    .A(_1188_));
 sg13g2_o21ai_1 _4284_ (.B1(_1121_),
    .Y(_1190_),
    .A1(_1049_),
    .A2(_1119_));
 sg13g2_nand2_1 _4285_ (.Y(_1191_),
    .A(net754),
    .B(net630));
 sg13g2_nand2_1 _4286_ (.Y(_1192_),
    .A(net757),
    .B(net626));
 sg13g2_or2_1 _4287_ (.X(_1193_),
    .B(_1192_),
    .A(_1118_));
 sg13g2_and2_1 _4288_ (.A(_1118_),
    .B(_1192_),
    .X(_1194_));
 sg13g2_xor2_1 _4289_ (.B(_1192_),
    .A(_1118_),
    .X(_1195_));
 sg13g2_xnor2_1 _4290_ (.Y(_1196_),
    .A(_1191_),
    .B(_1195_));
 sg13g2_nand2_1 _4291_ (.Y(_1197_),
    .A(_1190_),
    .B(_1196_));
 sg13g2_xnor2_1 _4292_ (.Y(_1198_),
    .A(_1190_),
    .B(_1196_));
 sg13g2_xnor2_1 _4293_ (.Y(_1199_),
    .A(_1189_),
    .B(_1198_));
 sg13g2_xor2_1 _4294_ (.B(_1199_),
    .A(_1182_),
    .X(_1200_));
 sg13g2_o21ai_1 _4295_ (.B1(_1107_),
    .Y(_1201_),
    .A1(_1108_),
    .A2(_1125_));
 sg13g2_nand2_1 _4296_ (.Y(_1202_),
    .A(_1200_),
    .B(_1201_));
 sg13g2_xor2_1 _4297_ (.B(_1201_),
    .A(_1200_),
    .X(_1203_));
 sg13g2_and2_1 _4298_ (.A(_1166_),
    .B(_1203_),
    .X(_1204_));
 sg13g2_xnor2_1 _4299_ (.Y(_1205_),
    .A(_1166_),
    .B(_1203_));
 sg13g2_or2_1 _4300_ (.X(_1206_),
    .B(_1205_),
    .A(_1130_));
 sg13g2_xnor2_1 _4301_ (.Y(_1207_),
    .A(_1130_),
    .B(_1205_));
 sg13g2_xor2_1 _4302_ (.B(_1207_),
    .A(_1151_),
    .X(_1208_));
 sg13g2_nor2b_1 _4303_ (.A(_1145_),
    .B_N(_1208_),
    .Y(_1209_));
 sg13g2_xnor2_1 _4304_ (.Y(_1210_),
    .A(_1145_),
    .B(_1208_));
 sg13g2_xnor2_1 _4305_ (.Y(_1211_),
    .A(_1144_),
    .B(_1210_));
 sg13g2_nand2_1 _4306_ (.Y(_1212_),
    .A(_1143_),
    .B(_1211_));
 sg13g2_nor2_1 _4307_ (.A(_1143_),
    .B(_1211_),
    .Y(_1213_));
 sg13g2_xor2_1 _4308_ (.B(_1211_),
    .A(_1143_),
    .X(_1214_));
 sg13g2_a21oi_1 _4309_ (.A1(_1076_),
    .A2(_1140_),
    .Y(_1215_),
    .B1(_1139_));
 sg13g2_xnor2_1 _4310_ (.Y(_1216_),
    .A(_1214_),
    .B(_1215_));
 sg13g2_o21ai_1 _4311_ (.B1(net793),
    .Y(_1217_),
    .A1(net609),
    .A2(_1216_));
 sg13g2_a21oi_1 _4312_ (.A1(net609),
    .A2(_2200_),
    .Y(_0178_),
    .B1(_1217_));
 sg13g2_o21ai_1 _4313_ (.B1(_1149_),
    .Y(_1218_),
    .A1(_1147_),
    .A2(_1150_));
 sg13g2_inv_1 _4314_ (.Y(_1219_),
    .A(_1218_));
 sg13g2_o21ai_1 _4315_ (.B1(_1206_),
    .Y(_1220_),
    .A1(_1151_),
    .A2(_1207_));
 sg13g2_o21ai_1 _4316_ (.B1(_1187_),
    .Y(_1221_),
    .A1(_1110_),
    .A2(_1185_));
 sg13g2_inv_1 _4317_ (.Y(_1222_),
    .A(_1221_));
 sg13g2_o21ai_1 _4318_ (.B1(_1197_),
    .Y(_1223_),
    .A1(_1189_),
    .A2(_1198_));
 sg13g2_nand3_1 _4319_ (.B(_1201_),
    .C(_1223_),
    .A(_1200_),
    .Y(_1224_));
 sg13g2_xor2_1 _4320_ (.B(_1223_),
    .A(_1202_),
    .X(_1225_));
 sg13g2_xnor2_1 _4321_ (.Y(_1226_),
    .A(_1221_),
    .B(_1225_));
 sg13g2_nand2_1 _4322_ (.Y(_1227_),
    .A(net716),
    .B(net701));
 sg13g2_nand2_2 _4323_ (.Y(_1228_),
    .A(net721),
    .B(net694));
 sg13g2_nor2_1 _4324_ (.A(_1158_),
    .B(_1228_),
    .Y(_1229_));
 sg13g2_or2_1 _4325_ (.X(_1230_),
    .B(_1228_),
    .A(_1158_));
 sg13g2_a22oi_1 _4326_ (.Y(_1231_),
    .B1(net694),
    .B2(net724),
    .A2(net698),
    .A1(net721));
 sg13g2_nor3_1 _4327_ (.A(_1227_),
    .B(_1229_),
    .C(_1231_),
    .Y(_1232_));
 sg13g2_o21ai_1 _4328_ (.B1(_1227_),
    .Y(_1233_),
    .A1(_1229_),
    .A2(_1231_));
 sg13g2_nor2b_1 _4329_ (.A(_1232_),
    .B_N(_1233_),
    .Y(_1234_));
 sg13g2_nand2_1 _4330_ (.Y(_1235_),
    .A(net730),
    .B(net692));
 sg13g2_nand2_1 _4331_ (.Y(_1236_),
    .A(net735),
    .B(net688));
 sg13g2_nand2_1 _4332_ (.Y(_1237_),
    .A(net739),
    .B(net688));
 sg13g2_xor2_1 _4333_ (.B(_1237_),
    .A(_1152_),
    .X(_1238_));
 sg13g2_nand2b_1 _4334_ (.Y(_1239_),
    .B(_1238_),
    .A_N(_1235_));
 sg13g2_xnor2_1 _4335_ (.Y(_1240_),
    .A(_1235_),
    .B(_1238_));
 sg13g2_xnor2_1 _4336_ (.Y(_1241_),
    .A(_1153_),
    .B(_1240_));
 sg13g2_and2_1 _4337_ (.A(_1234_),
    .B(_1241_),
    .X(_1242_));
 sg13g2_xnor2_1 _4338_ (.Y(_1243_),
    .A(_1234_),
    .B(_1241_));
 sg13g2_nor2_1 _4339_ (.A(_1163_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_xnor2_1 _4340_ (.Y(_1245_),
    .A(_1163_),
    .B(_1243_));
 sg13g2_o21ai_1 _4341_ (.B1(_1181_),
    .Y(_1246_),
    .A1(_1182_),
    .A2(_1199_));
 sg13g2_o21ai_1 _4342_ (.B1(_1177_),
    .Y(_1247_),
    .A1(_1169_),
    .A2(_1178_));
 sg13g2_nand2b_1 _4343_ (.Y(_1248_),
    .B(_1174_),
    .A_N(_1172_));
 sg13g2_o21ai_1 _4344_ (.B1(_1159_),
    .Y(_1249_),
    .A1(_1157_),
    .A2(_1160_));
 sg13g2_nand2_1 _4345_ (.Y(_1250_),
    .A(net761),
    .B(net616));
 sg13g2_nand2_1 _4346_ (.Y(_1251_),
    .A(net709),
    .B(net706));
 sg13g2_and4_1 _4347_ (.A(net713),
    .B(net709),
    .C(net612),
    .D(net705),
    .X(_1252_));
 sg13g2_a22oi_1 _4348_ (.Y(_1253_),
    .B1(net705),
    .B2(net713),
    .A2(net612),
    .A1(net709));
 sg13g2_or3_1 _4349_ (.A(_1250_),
    .B(_1252_),
    .C(_1253_),
    .X(_1254_));
 sg13g2_o21ai_1 _4350_ (.B1(_1250_),
    .Y(_1255_),
    .A1(_1252_),
    .A2(_1253_));
 sg13g2_nand3_1 _4351_ (.B(_1254_),
    .C(_1255_),
    .A(_1249_),
    .Y(_1256_));
 sg13g2_a21o_1 _4352_ (.A2(_1255_),
    .A1(_1254_),
    .B1(_1249_),
    .X(_1257_));
 sg13g2_nand3_1 _4353_ (.B(_1256_),
    .C(_1257_),
    .A(_1248_),
    .Y(_1258_));
 sg13g2_a21o_1 _4354_ (.A2(_1257_),
    .A1(_1256_),
    .B1(_1248_),
    .X(_1259_));
 sg13g2_nand3_1 _4355_ (.B(_1258_),
    .C(_1259_),
    .A(_1247_),
    .Y(_1260_));
 sg13g2_a21o_1 _4356_ (.A2(_1259_),
    .A1(_1258_),
    .B1(_1247_),
    .X(_1261_));
 sg13g2_nand2_1 _4357_ (.Y(_1262_),
    .A(net745),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[23] ));
 sg13g2_nand2_1 _4358_ (.Y(_1263_),
    .A(net747),
    .B(net634));
 sg13g2_nand2_1 _4359_ (.Y(_1264_),
    .A(net748),
    .B(net639));
 sg13g2_xor2_1 _4360_ (.B(_1264_),
    .A(_1184_),
    .X(_1265_));
 sg13g2_nand2b_1 _4361_ (.Y(_1266_),
    .B(_1265_),
    .A_N(_1262_));
 sg13g2_xnor2_1 _4362_ (.Y(_1267_),
    .A(_1262_),
    .B(_1265_));
 sg13g2_inv_1 _4363_ (.Y(_1268_),
    .A(_1267_));
 sg13g2_o21ai_1 _4364_ (.B1(_1193_),
    .Y(_1269_),
    .A1(_1191_),
    .A2(_1194_));
 sg13g2_nand2_1 _4365_ (.Y(_1270_),
    .A(net751),
    .B(net630));
 sg13g2_nand2_1 _4366_ (.Y(_1271_),
    .A(net754),
    .B(net620));
 sg13g2_and4_1 _4367_ (.A(net757),
    .B(net754),
    .C(net626),
    .D(net621),
    .X(_1272_));
 sg13g2_a22oi_1 _4368_ (.Y(_1273_),
    .B1(net621),
    .B2(net757),
    .A2(net626),
    .A1(net754));
 sg13g2_nor3_1 _4369_ (.A(_1270_),
    .B(_1272_),
    .C(_1273_),
    .Y(_1274_));
 sg13g2_o21ai_1 _4370_ (.B1(_1270_),
    .Y(_1275_),
    .A1(_1272_),
    .A2(_1273_));
 sg13g2_nor2b_1 _4371_ (.A(_1274_),
    .B_N(_1275_),
    .Y(_1276_));
 sg13g2_nand2_1 _4372_ (.Y(_1277_),
    .A(_1269_),
    .B(_1276_));
 sg13g2_xnor2_1 _4373_ (.Y(_1278_),
    .A(_1269_),
    .B(_1276_));
 sg13g2_xnor2_1 _4374_ (.Y(_1279_),
    .A(_1267_),
    .B(_1278_));
 sg13g2_nand3_1 _4375_ (.B(_1261_),
    .C(_1279_),
    .A(_1260_),
    .Y(_1280_));
 sg13g2_a21o_1 _4376_ (.A2(_1261_),
    .A1(_1260_),
    .B1(_1279_),
    .X(_1281_));
 sg13g2_nand3_1 _4377_ (.B(_1280_),
    .C(_1281_),
    .A(_1165_),
    .Y(_1282_));
 sg13g2_a21o_1 _4378_ (.A2(_1281_),
    .A1(_1280_),
    .B1(_1165_),
    .X(_1283_));
 sg13g2_a21oi_1 _4379_ (.A1(_1282_),
    .A2(_1283_),
    .Y(_1284_),
    .B1(_1246_));
 sg13g2_and3_1 _4380_ (.X(_1285_),
    .A(_1246_),
    .B(_1282_),
    .C(_1283_));
 sg13g2_nand3_1 _4381_ (.B(_1282_),
    .C(_1283_),
    .A(_1246_),
    .Y(_1286_));
 sg13g2_nor3_1 _4382_ (.A(_1245_),
    .B(_1284_),
    .C(_1285_),
    .Y(_1287_));
 sg13g2_or3_1 _4383_ (.A(_1245_),
    .B(_1284_),
    .C(_1285_),
    .X(_1288_));
 sg13g2_o21ai_1 _4384_ (.B1(_1245_),
    .Y(_1289_),
    .A1(_1284_),
    .A2(_1285_));
 sg13g2_nand3_1 _4385_ (.B(_1288_),
    .C(_1289_),
    .A(_1204_),
    .Y(_1290_));
 sg13g2_a21o_1 _4386_ (.A2(_1289_),
    .A1(_1288_),
    .B1(_1204_),
    .X(_1291_));
 sg13g2_nand3_1 _4387_ (.B(_1290_),
    .C(_1291_),
    .A(_1226_),
    .Y(_1292_));
 sg13g2_a21o_1 _4388_ (.A2(_1291_),
    .A1(_1290_),
    .B1(_1226_),
    .X(_1293_));
 sg13g2_nand3_1 _4389_ (.B(_1292_),
    .C(_1293_),
    .A(_1220_),
    .Y(_1294_));
 sg13g2_a21oi_1 _4390_ (.A1(_1292_),
    .A2(_1293_),
    .Y(_1295_),
    .B1(_1220_));
 sg13g2_a21o_1 _4391_ (.A2(_1293_),
    .A1(_1292_),
    .B1(_1220_),
    .X(_1296_));
 sg13g2_a21oi_1 _4392_ (.A1(_1294_),
    .A2(_1296_),
    .Y(_1297_),
    .B1(_1218_));
 sg13g2_nand3_1 _4393_ (.B(_1294_),
    .C(_1296_),
    .A(_1218_),
    .Y(_1298_));
 sg13g2_nand2b_1 _4394_ (.Y(_1299_),
    .B(_1298_),
    .A_N(_1297_));
 sg13g2_a21o_1 _4395_ (.A2(_1210_),
    .A1(_1144_),
    .B1(_1209_),
    .X(_1300_));
 sg13g2_nand3b_1 _4396_ (.B(_1298_),
    .C(_1300_),
    .Y(_1301_),
    .A_N(_1297_));
 sg13g2_xnor2_1 _4397_ (.Y(_1302_),
    .A(_1299_),
    .B(_1300_));
 sg13g2_nand2_1 _4398_ (.Y(_1303_),
    .A(_1140_),
    .B(_1214_));
 sg13g2_a21oi_1 _4399_ (.A1(_1070_),
    .A2(_1073_),
    .Y(_1304_),
    .B1(_1303_));
 sg13g2_a21o_1 _4400_ (.A2(_1073_),
    .A1(_1070_),
    .B1(_1303_),
    .X(_1305_));
 sg13g2_a21o_1 _4401_ (.A2(_1212_),
    .A1(_1139_),
    .B1(_1213_),
    .X(_1306_));
 sg13g2_o21ai_1 _4402_ (.B1(_1302_),
    .Y(_1307_),
    .A1(_1304_),
    .A2(_1306_));
 sg13g2_or3_1 _4403_ (.A(_1302_),
    .B(_1304_),
    .C(_1306_),
    .X(_1308_));
 sg13g2_and2_1 _4404_ (.A(_1307_),
    .B(_1308_),
    .X(_1309_));
 sg13g2_o21ai_1 _4405_ (.B1(net793),
    .Y(_1310_),
    .A1(net610),
    .A2(_1309_));
 sg13g2_a21oi_1 _4406_ (.A1(net609),
    .A2(_2199_),
    .Y(_0179_),
    .B1(_1310_));
 sg13g2_nand2_1 _4407_ (.Y(_1311_),
    .A(_1301_),
    .B(_1307_));
 sg13g2_o21ai_1 _4408_ (.B1(_1294_),
    .Y(_1312_),
    .A1(_1219_),
    .A2(_1295_));
 sg13g2_inv_1 _4409_ (.Y(_1313_),
    .A(_1312_));
 sg13g2_o21ai_1 _4410_ (.B1(_1224_),
    .Y(_1314_),
    .A1(_1222_),
    .A2(_1225_));
 sg13g2_nand2_1 _4411_ (.Y(_1315_),
    .A(_1290_),
    .B(_1292_));
 sg13g2_o21ai_1 _4412_ (.B1(_1266_),
    .Y(_1316_),
    .A1(_1184_),
    .A2(_1264_));
 sg13g2_and2_1 _4413_ (.A(_1282_),
    .B(_1286_),
    .X(_1317_));
 sg13g2_o21ai_1 _4414_ (.B1(_1277_),
    .Y(_1318_),
    .A1(_1268_),
    .A2(_1278_));
 sg13g2_inv_1 _4415_ (.Y(_1319_),
    .A(_1318_));
 sg13g2_xnor2_1 _4416_ (.Y(_1320_),
    .A(_1317_),
    .B(_1319_));
 sg13g2_nand2b_1 _4417_ (.Y(_1321_),
    .B(_1316_),
    .A_N(_1320_));
 sg13g2_xor2_1 _4418_ (.B(_1320_),
    .A(_1316_),
    .X(_1322_));
 sg13g2_nand2_1 _4419_ (.Y(_1323_),
    .A(_1260_),
    .B(_1280_));
 sg13g2_nand2_1 _4420_ (.Y(_1324_),
    .A(_1256_),
    .B(_1258_));
 sg13g2_nand2b_1 _4421_ (.Y(_1325_),
    .B(_1254_),
    .A_N(_1252_));
 sg13g2_o21ai_1 _4422_ (.B1(_1230_),
    .Y(_1326_),
    .A1(_1227_),
    .A2(_1231_));
 sg13g2_nand2_1 _4423_ (.Y(_1327_),
    .A(net757),
    .B(net616));
 sg13g2_nand2_1 _4424_ (.Y(_1328_),
    .A(net761),
    .B(net706));
 sg13g2_nand2_1 _4425_ (.Y(_1329_),
    .A(net761),
    .B(net613));
 sg13g2_or2_1 _4426_ (.X(_1330_),
    .B(_1329_),
    .A(_1251_));
 sg13g2_xnor2_1 _4427_ (.Y(_1331_),
    .A(_1251_),
    .B(_1329_));
 sg13g2_xor2_1 _4428_ (.B(_1331_),
    .A(_1327_),
    .X(_1332_));
 sg13g2_xnor2_1 _4429_ (.Y(_1333_),
    .A(_1326_),
    .B(_1332_));
 sg13g2_nor2b_1 _4430_ (.A(_1333_),
    .B_N(_1325_),
    .Y(_1334_));
 sg13g2_xnor2_1 _4431_ (.Y(_1335_),
    .A(_1325_),
    .B(_1333_));
 sg13g2_nand2_1 _4432_ (.Y(_1336_),
    .A(_1324_),
    .B(_1335_));
 sg13g2_xnor2_1 _4433_ (.Y(_1337_),
    .A(_1324_),
    .B(_1335_));
 sg13g2_nand2_2 _4434_ (.Y(_1338_),
    .A(net742),
    .B(net641));
 sg13g2_nand2_2 _4435_ (.Y(_1339_),
    .A(net745),
    .B(net638));
 sg13g2_xor2_1 _4436_ (.B(_1339_),
    .A(_1263_),
    .X(_1340_));
 sg13g2_nand2b_1 _4437_ (.Y(_1341_),
    .B(_1340_),
    .A_N(_1338_));
 sg13g2_xnor2_1 _4438_ (.Y(_1342_),
    .A(_1338_),
    .B(_1340_));
 sg13g2_inv_1 _4439_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_or2_1 _4440_ (.X(_1344_),
    .B(_1274_),
    .A(_1272_));
 sg13g2_nand2_1 _4441_ (.Y(_1345_),
    .A(net750),
    .B(net630));
 sg13g2_nand2_1 _4442_ (.Y(_1346_),
    .A(net752),
    .B(net620));
 sg13g2_nand2_1 _4443_ (.Y(_1347_),
    .A(net752),
    .B(net626));
 sg13g2_xor2_1 _4444_ (.B(_1347_),
    .A(_1271_),
    .X(_1348_));
 sg13g2_nand2b_1 _4445_ (.Y(_1349_),
    .B(_1348_),
    .A_N(_1345_));
 sg13g2_xnor2_1 _4446_ (.Y(_1350_),
    .A(_1345_),
    .B(_1348_));
 sg13g2_nand2_1 _4447_ (.Y(_1351_),
    .A(_1344_),
    .B(_1350_));
 sg13g2_xnor2_1 _4448_ (.Y(_1352_),
    .A(_1344_),
    .B(_1350_));
 sg13g2_xnor2_1 _4449_ (.Y(_1353_),
    .A(_1343_),
    .B(_1352_));
 sg13g2_xor2_1 _4450_ (.B(_1353_),
    .A(_1337_),
    .X(_1354_));
 sg13g2_and2_1 _4451_ (.A(_1244_),
    .B(_1354_),
    .X(_1355_));
 sg13g2_xor2_1 _4452_ (.B(_1354_),
    .A(_1244_),
    .X(_1356_));
 sg13g2_xnor2_1 _4453_ (.Y(_1357_),
    .A(_1323_),
    .B(_1356_));
 sg13g2_nand2_2 _4454_ (.Y(_1358_),
    .A(net739),
    .B(net686));
 sg13g2_inv_4 _4455_ (.A(_1358_),
    .Y(_1359_));
 sg13g2_a21oi_1 _4456_ (.A1(_1154_),
    .A2(_1240_),
    .Y(_1360_),
    .B1(_1242_));
 sg13g2_o21ai_1 _4457_ (.B1(_1239_),
    .Y(_1361_),
    .A1(_1152_),
    .A2(_1237_));
 sg13g2_nand2_1 _4458_ (.Y(_1362_),
    .A(net724),
    .B(net693));
 sg13g2_nand2_2 _4459_ (.Y(_1363_),
    .A(net731),
    .B(net689));
 sg13g2_nand2_1 _4460_ (.Y(_1364_),
    .A(net730),
    .B(net691));
 sg13g2_xor2_1 _4461_ (.B(_1364_),
    .A(_1236_),
    .X(_1365_));
 sg13g2_nand2b_1 _4462_ (.Y(_1366_),
    .B(_1365_),
    .A_N(_1362_));
 sg13g2_xnor2_1 _4463_ (.Y(_1367_),
    .A(_1362_),
    .B(_1365_));
 sg13g2_and2_1 _4464_ (.A(_1361_),
    .B(_1367_),
    .X(_1368_));
 sg13g2_xnor2_1 _4465_ (.Y(_1369_),
    .A(_1361_),
    .B(_1367_));
 sg13g2_nand2_1 _4466_ (.Y(_1370_),
    .A(net713),
    .B(net701));
 sg13g2_nand2_1 _4467_ (.Y(_1371_),
    .A(net716),
    .B(net694));
 sg13g2_nand2_1 _4468_ (.Y(_1372_),
    .A(net716),
    .B(net698));
 sg13g2_xor2_1 _4469_ (.B(_1372_),
    .A(_1228_),
    .X(_1373_));
 sg13g2_nand2b_1 _4470_ (.Y(_1374_),
    .B(_1373_),
    .A_N(_1370_));
 sg13g2_xnor2_1 _4471_ (.Y(_1375_),
    .A(_1370_),
    .B(_1373_));
 sg13g2_nor2b_1 _4472_ (.A(_1369_),
    .B_N(_1375_),
    .Y(_1376_));
 sg13g2_xnor2_1 _4473_ (.Y(_1377_),
    .A(_1369_),
    .B(_1375_));
 sg13g2_nand2b_1 _4474_ (.Y(_1378_),
    .B(_1377_),
    .A_N(_1360_));
 sg13g2_xnor2_1 _4475_ (.Y(_1379_),
    .A(_1360_),
    .B(_1377_));
 sg13g2_and2_1 _4476_ (.A(_1359_),
    .B(_1379_),
    .X(_1380_));
 sg13g2_xnor2_1 _4477_ (.Y(_1381_),
    .A(_1358_),
    .B(_1379_));
 sg13g2_nor2b_1 _4478_ (.A(_1357_),
    .B_N(_1381_),
    .Y(_1382_));
 sg13g2_xnor2_1 _4479_ (.Y(_1383_),
    .A(_1357_),
    .B(_1381_));
 sg13g2_nand2_1 _4480_ (.Y(_1384_),
    .A(_1287_),
    .B(_1383_));
 sg13g2_xnor2_1 _4481_ (.Y(_1385_),
    .A(_1287_),
    .B(_1383_));
 sg13g2_xor2_1 _4482_ (.B(_1385_),
    .A(_1322_),
    .X(_1386_));
 sg13g2_xnor2_1 _4483_ (.Y(_1387_),
    .A(_1315_),
    .B(_1386_));
 sg13g2_nor2b_1 _4484_ (.A(_1387_),
    .B_N(_1314_),
    .Y(_1388_));
 sg13g2_xor2_1 _4485_ (.B(_1387_),
    .A(_1314_),
    .X(_1389_));
 sg13g2_nand2_1 _4486_ (.Y(_1390_),
    .A(_1313_),
    .B(_1389_));
 sg13g2_xnor2_1 _4487_ (.Y(_1391_),
    .A(_1312_),
    .B(_1389_));
 sg13g2_xnor2_1 _4488_ (.Y(_1392_),
    .A(_1311_),
    .B(_1391_));
 sg13g2_o21ai_1 _4489_ (.B1(net796),
    .Y(_1393_),
    .A1(net673),
    .A2(net245));
 sg13g2_a21oi_1 _4490_ (.A1(net673),
    .A2(_1392_),
    .Y(_0180_),
    .B1(net246));
 sg13g2_o21ai_1 _4491_ (.B1(_1321_),
    .Y(_1394_),
    .A1(_1317_),
    .A2(_1319_));
 sg13g2_o21ai_1 _4492_ (.B1(_1384_),
    .Y(_1395_),
    .A1(_1322_),
    .A2(_1385_));
 sg13g2_o21ai_1 _4493_ (.B1(_1341_),
    .Y(_1396_),
    .A1(_1263_),
    .A2(_1339_));
 sg13g2_inv_1 _4494_ (.Y(_1397_),
    .A(_1396_));
 sg13g2_a21oi_1 _4495_ (.A1(_1323_),
    .A2(_1356_),
    .Y(_1398_),
    .B1(_1355_));
 sg13g2_o21ai_1 _4496_ (.B1(_1351_),
    .Y(_1399_),
    .A1(_1343_),
    .A2(_1352_));
 sg13g2_nand2b_1 _4497_ (.Y(_1400_),
    .B(_1399_),
    .A_N(_1398_));
 sg13g2_xor2_1 _4498_ (.B(_1399_),
    .A(_1398_),
    .X(_1401_));
 sg13g2_xnor2_1 _4499_ (.Y(_1402_),
    .A(_1397_),
    .B(_1401_));
 sg13g2_nor2_2 _4500_ (.A(_2219_),
    .B(_2233_),
    .Y(_1403_));
 sg13g2_nand2_2 _4501_ (.Y(_1404_),
    .A(net736),
    .B(_1359_));
 sg13g2_o21ai_1 _4502_ (.B1(_1404_),
    .Y(_1405_),
    .A1(_1359_),
    .A2(_1403_));
 sg13g2_o21ai_1 _4503_ (.B1(_1366_),
    .Y(_1406_),
    .A1(_1152_),
    .A2(_1363_));
 sg13g2_nand2_1 _4504_ (.Y(_1407_),
    .A(net720),
    .B(net692));
 sg13g2_nand2_1 _4505_ (.Y(_1408_),
    .A(net725),
    .B(net689));
 sg13g2_nand2_1 _4506_ (.Y(_1409_),
    .A(net724),
    .B(net691));
 sg13g2_xor2_1 _4507_ (.B(_1409_),
    .A(_1363_),
    .X(_1410_));
 sg13g2_nand2b_1 _4508_ (.Y(_1411_),
    .B(_1410_),
    .A_N(_1407_));
 sg13g2_xnor2_1 _4509_ (.Y(_1412_),
    .A(_1407_),
    .B(_1410_));
 sg13g2_and2_1 _4510_ (.A(_1406_),
    .B(_1412_),
    .X(_1413_));
 sg13g2_xnor2_1 _4511_ (.Y(_1414_),
    .A(_1406_),
    .B(_1412_));
 sg13g2_nand2_1 _4512_ (.Y(_1415_),
    .A(net709),
    .B(net701));
 sg13g2_nand2_1 _4513_ (.Y(_1416_),
    .A(net715),
    .B(net694));
 sg13g2_nand2_1 _4514_ (.Y(_1417_),
    .A(net713),
    .B(net698));
 sg13g2_xor2_1 _4515_ (.B(_1417_),
    .A(_1371_),
    .X(_1418_));
 sg13g2_nand2b_1 _4516_ (.Y(_1419_),
    .B(_1418_),
    .A_N(_1415_));
 sg13g2_xnor2_1 _4517_ (.Y(_1420_),
    .A(_1415_),
    .B(_1418_));
 sg13g2_nor2b_1 _4518_ (.A(_1414_),
    .B_N(_1420_),
    .Y(_1421_));
 sg13g2_xnor2_1 _4519_ (.Y(_1422_),
    .A(_1414_),
    .B(_1420_));
 sg13g2_o21ai_1 _4520_ (.B1(_1422_),
    .Y(_1423_),
    .A1(_1368_),
    .A2(_1376_));
 sg13g2_or3_1 _4521_ (.A(_1368_),
    .B(_1376_),
    .C(_1422_),
    .X(_1424_));
 sg13g2_and2_1 _4522_ (.A(_1423_),
    .B(_1424_),
    .X(_1425_));
 sg13g2_nor2b_1 _4523_ (.A(net556),
    .B_N(_1425_),
    .Y(_1426_));
 sg13g2_xnor2_1 _4524_ (.Y(_1427_),
    .A(net556),
    .B(_1425_));
 sg13g2_nand2_1 _4525_ (.Y(_1428_),
    .A(_1380_),
    .B(_1427_));
 sg13g2_xnor2_1 _4526_ (.Y(_1429_),
    .A(_1380_),
    .B(_1427_));
 sg13g2_o21ai_1 _4527_ (.B1(_1336_),
    .Y(_1430_),
    .A1(_1337_),
    .A2(_1353_));
 sg13g2_a21o_1 _4528_ (.A2(_1332_),
    .A1(_1326_),
    .B1(_1334_),
    .X(_1431_));
 sg13g2_o21ai_1 _4529_ (.B1(_1330_),
    .Y(_1432_),
    .A1(_1327_),
    .A2(_1331_));
 sg13g2_o21ai_1 _4530_ (.B1(_1374_),
    .Y(_1433_),
    .A1(_1228_),
    .A2(_1372_));
 sg13g2_nand2_1 _4531_ (.Y(_1434_),
    .A(net754),
    .B(net617));
 sg13g2_nand2_1 _4532_ (.Y(_1435_),
    .A(net757),
    .B(net706));
 sg13g2_nand2_1 _4533_ (.Y(_1436_),
    .A(net757),
    .B(net613));
 sg13g2_or2_1 _4534_ (.X(_1437_),
    .B(_1435_),
    .A(_1329_));
 sg13g2_xnor2_1 _4535_ (.Y(_1438_),
    .A(_1328_),
    .B(_1436_));
 sg13g2_xor2_1 _4536_ (.B(_1438_),
    .A(_1434_),
    .X(_1439_));
 sg13g2_xnor2_1 _4537_ (.Y(_1440_),
    .A(_1433_),
    .B(_1439_));
 sg13g2_nor2b_1 _4538_ (.A(_1440_),
    .B_N(_1432_),
    .Y(_1441_));
 sg13g2_xnor2_1 _4539_ (.Y(_1442_),
    .A(_1432_),
    .B(_1440_));
 sg13g2_nand2_1 _4540_ (.Y(_1443_),
    .A(_1431_),
    .B(_1442_));
 sg13g2_xnor2_1 _4541_ (.Y(_1444_),
    .A(_1431_),
    .B(_1442_));
 sg13g2_nor3_1 _4542_ (.A(_2226_),
    .B(_2228_),
    .C(_1339_),
    .Y(_1445_));
 sg13g2_a22oi_1 _4543_ (.Y(_1446_),
    .B1(net634),
    .B2(net745),
    .A2(net638),
    .A1(net742));
 sg13g2_nor3_1 _4544_ (.A(_1338_),
    .B(_1445_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_o21ai_1 _4545_ (.B1(_1338_),
    .Y(_1448_),
    .A1(_1445_),
    .A2(_1446_));
 sg13g2_nor2b_1 _4546_ (.A(_1447_),
    .B_N(_1448_),
    .Y(_1449_));
 sg13g2_inv_1 _4547_ (.Y(_1450_),
    .A(_1449_));
 sg13g2_o21ai_1 _4548_ (.B1(_1349_),
    .Y(_1451_),
    .A1(_1271_),
    .A2(_1347_));
 sg13g2_nand2_1 _4549_ (.Y(_1452_),
    .A(net748),
    .B(net631));
 sg13g2_nand2_2 _4550_ (.Y(_1453_),
    .A(net749),
    .B(net620));
 sg13g2_nand2_1 _4551_ (.Y(_1454_),
    .A(net749),
    .B(net627));
 sg13g2_xor2_1 _4552_ (.B(_1454_),
    .A(_1346_),
    .X(_1455_));
 sg13g2_nand2b_1 _4553_ (.Y(_1456_),
    .B(_1455_),
    .A_N(_1452_));
 sg13g2_xnor2_1 _4554_ (.Y(_1457_),
    .A(_1452_),
    .B(_1455_));
 sg13g2_nand2_1 _4555_ (.Y(_1458_),
    .A(_1451_),
    .B(_1457_));
 sg13g2_xnor2_1 _4556_ (.Y(_1459_),
    .A(_1451_),
    .B(_1457_));
 sg13g2_xnor2_1 _4557_ (.Y(_1460_),
    .A(_1450_),
    .B(_1459_));
 sg13g2_xor2_1 _4558_ (.B(_1460_),
    .A(_1444_),
    .X(_1461_));
 sg13g2_nor2b_1 _4559_ (.A(_1378_),
    .B_N(_1461_),
    .Y(_1462_));
 sg13g2_xnor2_1 _4560_ (.Y(_1463_),
    .A(_1378_),
    .B(_1461_));
 sg13g2_xnor2_1 _4561_ (.Y(_1464_),
    .A(_1430_),
    .B(_1463_));
 sg13g2_xor2_1 _4562_ (.B(_1464_),
    .A(_1429_),
    .X(_1465_));
 sg13g2_nand2_1 _4563_ (.Y(_1466_),
    .A(_1382_),
    .B(_1465_));
 sg13g2_xnor2_1 _4564_ (.Y(_1467_),
    .A(_1382_),
    .B(_1465_));
 sg13g2_xor2_1 _4565_ (.B(_1467_),
    .A(_1402_),
    .X(_1468_));
 sg13g2_xnor2_1 _4566_ (.Y(_1469_),
    .A(_1395_),
    .B(_1468_));
 sg13g2_nor2b_1 _4567_ (.A(_1469_),
    .B_N(_1394_),
    .Y(_1470_));
 sg13g2_xor2_1 _4568_ (.B(_1469_),
    .A(_1394_),
    .X(_1471_));
 sg13g2_a21o_1 _4569_ (.A2(_1386_),
    .A1(_1315_),
    .B1(_1388_),
    .X(_1472_));
 sg13g2_nor2b_1 _4570_ (.A(_1471_),
    .B_N(_1472_),
    .Y(_1473_));
 sg13g2_xor2_1 _4571_ (.B(_1472_),
    .A(_1471_),
    .X(_1474_));
 sg13g2_o21ai_1 _4572_ (.B1(_1301_),
    .Y(_1475_),
    .A1(_1313_),
    .A2(_1389_));
 sg13g2_nand2_1 _4573_ (.Y(_1476_),
    .A(_1390_),
    .B(_1475_));
 sg13g2_a21oi_1 _4574_ (.A1(_1390_),
    .A2(_1475_),
    .Y(_1477_),
    .B1(_1306_));
 sg13g2_nand2_1 _4575_ (.Y(_1478_),
    .A(_1302_),
    .B(_1391_));
 sg13g2_a22oi_1 _4576_ (.Y(_1479_),
    .B1(_1478_),
    .B2(_1476_),
    .A2(_1477_),
    .A1(_1305_));
 sg13g2_a221oi_1 _4577_ (.B2(_1476_),
    .C1(_1474_),
    .B1(_1478_),
    .A1(_1305_),
    .Y(_1480_),
    .A2(_1477_));
 sg13g2_xnor2_1 _4578_ (.Y(_1481_),
    .A(_1474_),
    .B(_1479_));
 sg13g2_o21ai_1 _4579_ (.B1(net793),
    .Y(_1482_),
    .A1(net610),
    .A2(_1481_));
 sg13g2_a21oi_1 _4580_ (.A1(net610),
    .A2(_2198_),
    .Y(_0181_),
    .B1(_1482_));
 sg13g2_nor2_1 _4581_ (.A(_1473_),
    .B(_1480_),
    .Y(_1483_));
 sg13g2_a21o_1 _4582_ (.A2(_1468_),
    .A1(_1395_),
    .B1(_1470_),
    .X(_1484_));
 sg13g2_o21ai_1 _4583_ (.B1(_1400_),
    .Y(_1485_),
    .A1(_1397_),
    .A2(_1401_));
 sg13g2_o21ai_1 _4584_ (.B1(_1466_),
    .Y(_1486_),
    .A1(_1402_),
    .A2(_1467_));
 sg13g2_or2_1 _4585_ (.X(_1487_),
    .B(_1447_),
    .A(_1445_));
 sg13g2_a21oi_1 _4586_ (.A1(_1430_),
    .A2(_1463_),
    .Y(_1488_),
    .B1(_1462_));
 sg13g2_o21ai_1 _4587_ (.B1(_1458_),
    .Y(_1489_),
    .A1(_1450_),
    .A2(_1459_));
 sg13g2_nor2b_1 _4588_ (.A(_1488_),
    .B_N(_1489_),
    .Y(_1490_));
 sg13g2_xor2_1 _4589_ (.B(_1489_),
    .A(_1488_),
    .X(_1491_));
 sg13g2_nor2b_1 _4590_ (.A(_1491_),
    .B_N(_1487_),
    .Y(_1492_));
 sg13g2_xor2_1 _4591_ (.B(_1491_),
    .A(_1487_),
    .X(_1493_));
 sg13g2_o21ai_1 _4592_ (.B1(_1428_),
    .Y(_1494_),
    .A1(_1429_),
    .A2(_1464_));
 sg13g2_nand2_2 _4593_ (.Y(_1495_),
    .A(net729),
    .B(net686));
 sg13g2_nand2_1 _4594_ (.Y(_1496_),
    .A(net729),
    .B(_1403_));
 sg13g2_nand3_1 _4595_ (.B(_1359_),
    .C(_1403_),
    .A(net730),
    .Y(_1497_));
 sg13g2_nor2_1 _4596_ (.A(net556),
    .B(_1495_),
    .Y(_1498_));
 sg13g2_xor2_1 _4597_ (.B(_1495_),
    .A(net556),
    .X(_1499_));
 sg13g2_mux2_1 _4598_ (.A0(_1495_),
    .A1(_1499_),
    .S(_1404_),
    .X(_1500_));
 sg13g2_o21ai_1 _4599_ (.B1(_1411_),
    .Y(_1501_),
    .A1(_1363_),
    .A2(_1409_));
 sg13g2_nand2_1 _4600_ (.Y(_1502_),
    .A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .B(net692));
 sg13g2_nand2_1 _4601_ (.Y(_1503_),
    .A(net720),
    .B(net689));
 sg13g2_nand2_1 _4602_ (.Y(_1504_),
    .A(net721),
    .B(net690));
 sg13g2_xor2_1 _4603_ (.B(_1504_),
    .A(_1408_),
    .X(_1505_));
 sg13g2_nand2b_1 _4604_ (.Y(_1506_),
    .B(_1505_),
    .A_N(_1502_));
 sg13g2_xnor2_1 _4605_ (.Y(_1507_),
    .A(_1502_),
    .B(_1505_));
 sg13g2_nand2_1 _4606_ (.Y(_1508_),
    .A(_1501_),
    .B(_1507_));
 sg13g2_xnor2_1 _4607_ (.Y(_1509_),
    .A(_1501_),
    .B(_1507_));
 sg13g2_nand2_1 _4608_ (.Y(_1510_),
    .A(net761),
    .B(net701));
 sg13g2_nand2_1 _4609_ (.Y(_1511_),
    .A(net709),
    .B(net695));
 sg13g2_nand2_1 _4610_ (.Y(_1512_),
    .A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .B(net698));
 sg13g2_xor2_1 _4611_ (.B(_1512_),
    .A(_1416_),
    .X(_1513_));
 sg13g2_nand2b_1 _4612_ (.Y(_1514_),
    .B(_1513_),
    .A_N(_1510_));
 sg13g2_xnor2_1 _4613_ (.Y(_1515_),
    .A(_1510_),
    .B(_1513_));
 sg13g2_nand2b_1 _4614_ (.Y(_1516_),
    .B(_1515_),
    .A_N(_1509_));
 sg13g2_xnor2_1 _4615_ (.Y(_1517_),
    .A(_1509_),
    .B(_1515_));
 sg13g2_o21ai_1 _4616_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_1413_),
    .A2(_1421_));
 sg13g2_or3_1 _4617_ (.A(_1413_),
    .B(_1421_),
    .C(_1517_),
    .X(_1519_));
 sg13g2_and2_1 _4618_ (.A(_1518_),
    .B(_1519_),
    .X(_1520_));
 sg13g2_and2_1 _4619_ (.A(_1500_),
    .B(_1520_),
    .X(_1521_));
 sg13g2_xnor2_1 _4620_ (.Y(_1522_),
    .A(_1500_),
    .B(_1520_));
 sg13g2_inv_1 _4621_ (.Y(_1523_),
    .A(_1522_));
 sg13g2_nand2_1 _4622_ (.Y(_1524_),
    .A(_1426_),
    .B(_1523_));
 sg13g2_xor2_1 _4623_ (.B(_1522_),
    .A(_1426_),
    .X(_1525_));
 sg13g2_o21ai_1 _4624_ (.B1(_1443_),
    .Y(_1526_),
    .A1(_1444_),
    .A2(_1460_));
 sg13g2_o21ai_1 _4625_ (.B1(net742),
    .Y(_1527_),
    .A1(net638),
    .A2(net634));
 sg13g2_nand3_1 _4626_ (.B(net638),
    .C(net634),
    .A(net742),
    .Y(_1528_));
 sg13g2_nand2b_1 _4627_ (.Y(_1529_),
    .B(_1528_),
    .A_N(_1527_));
 sg13g2_xor2_1 _4628_ (.B(_1529_),
    .A(_1338_),
    .X(_1530_));
 sg13g2_xnor2_1 _4629_ (.Y(_1531_),
    .A(_1338_),
    .B(_1529_));
 sg13g2_o21ai_1 _4630_ (.B1(_1456_),
    .Y(_1532_),
    .A1(_1346_),
    .A2(_1454_));
 sg13g2_nand2_1 _4631_ (.Y(_1533_),
    .A(net745),
    .B(net630));
 sg13g2_nand2_2 _4632_ (.Y(_1534_),
    .A(net747),
    .B(net626));
 sg13g2_xor2_1 _4633_ (.B(_1534_),
    .A(_1453_),
    .X(_1535_));
 sg13g2_nand2b_1 _4634_ (.Y(_1536_),
    .B(_1535_),
    .A_N(_1533_));
 sg13g2_xnor2_1 _4635_ (.Y(_1537_),
    .A(_1533_),
    .B(_1535_));
 sg13g2_nand2_1 _4636_ (.Y(_1538_),
    .A(_1532_),
    .B(_1537_));
 sg13g2_xnor2_1 _4637_ (.Y(_1539_),
    .A(_1532_),
    .B(_1537_));
 sg13g2_xnor2_1 _4638_ (.Y(_1540_),
    .A(_1531_),
    .B(_1539_));
 sg13g2_a21o_1 _4639_ (.A2(_1439_),
    .A1(_1433_),
    .B1(_1441_),
    .X(_1541_));
 sg13g2_o21ai_1 _4640_ (.B1(_1437_),
    .Y(_1542_),
    .A1(_1434_),
    .A2(_1438_));
 sg13g2_o21ai_1 _4641_ (.B1(_1419_),
    .Y(_1543_),
    .A1(_1371_),
    .A2(_1417_));
 sg13g2_nand2_1 _4642_ (.Y(_1544_),
    .A(net752),
    .B(net616));
 sg13g2_nand2_1 _4643_ (.Y(_1545_),
    .A(net754),
    .B(net705));
 sg13g2_nand2_1 _4644_ (.Y(_1546_),
    .A(net755),
    .B(net613));
 sg13g2_or2_1 _4645_ (.X(_1547_),
    .B(_1545_),
    .A(_1436_));
 sg13g2_xnor2_1 _4646_ (.Y(_1548_),
    .A(_1435_),
    .B(_1546_));
 sg13g2_xor2_1 _4647_ (.B(_1548_),
    .A(_1544_),
    .X(_1549_));
 sg13g2_xnor2_1 _4648_ (.Y(_1550_),
    .A(_1543_),
    .B(_1549_));
 sg13g2_nor2b_1 _4649_ (.A(_1550_),
    .B_N(_1542_),
    .Y(_1551_));
 sg13g2_xnor2_1 _4650_ (.Y(_1552_),
    .A(_1542_),
    .B(_1550_));
 sg13g2_nand2_1 _4651_ (.Y(_1553_),
    .A(_1541_),
    .B(_1552_));
 sg13g2_xnor2_1 _4652_ (.Y(_1554_),
    .A(_1541_),
    .B(_1552_));
 sg13g2_xor2_1 _4653_ (.B(_1554_),
    .A(_1540_),
    .X(_1555_));
 sg13g2_nor2b_1 _4654_ (.A(_1423_),
    .B_N(_1555_),
    .Y(_1556_));
 sg13g2_xnor2_1 _4655_ (.Y(_1557_),
    .A(_1423_),
    .B(_1555_));
 sg13g2_and2_1 _4656_ (.A(_1526_),
    .B(_1557_),
    .X(_1558_));
 sg13g2_xnor2_1 _4657_ (.Y(_1559_),
    .A(_1526_),
    .B(_1557_));
 sg13g2_xor2_1 _4658_ (.B(_1559_),
    .A(_1525_),
    .X(_1560_));
 sg13g2_xnor2_1 _4659_ (.Y(_1561_),
    .A(_1494_),
    .B(_1560_));
 sg13g2_nor2_1 _4660_ (.A(_1493_),
    .B(_1561_),
    .Y(_1562_));
 sg13g2_xor2_1 _4661_ (.B(_1561_),
    .A(_1493_),
    .X(_1563_));
 sg13g2_xnor2_1 _4662_ (.Y(_1564_),
    .A(_1486_),
    .B(_1563_));
 sg13g2_nor2b_1 _4663_ (.A(_1564_),
    .B_N(_1485_),
    .Y(_1565_));
 sg13g2_xor2_1 _4664_ (.B(_1564_),
    .A(_1485_),
    .X(_1566_));
 sg13g2_nor2b_1 _4665_ (.A(_1566_),
    .B_N(_1484_),
    .Y(_1567_));
 sg13g2_nor2b_2 _4666_ (.A(_1484_),
    .B_N(_1566_),
    .Y(_1568_));
 sg13g2_nor2_1 _4667_ (.A(_1567_),
    .B(_1568_),
    .Y(_1569_));
 sg13g2_xnor2_1 _4668_ (.Y(_1570_),
    .A(_1483_),
    .B(_1569_));
 sg13g2_o21ai_1 _4669_ (.B1(net793),
    .Y(_1571_),
    .A1(net610),
    .A2(_1570_));
 sg13g2_a21oi_1 _4670_ (.A1(net609),
    .A2(_2197_),
    .Y(_0182_),
    .B1(_1571_));
 sg13g2_nor2_2 _4671_ (.A(_1490_),
    .B(_1492_),
    .Y(_1572_));
 sg13g2_a21oi_2 _4672_ (.B1(_1562_),
    .Y(_1573_),
    .A2(_1560_),
    .A1(_1494_));
 sg13g2_o21ai_1 _4673_ (.B1(_1524_),
    .Y(_1574_),
    .A1(_1525_),
    .A2(_1559_));
 sg13g2_a21oi_2 _4674_ (.B1(_1498_),
    .Y(_1575_),
    .A2(_1359_),
    .A1(net736));
 sg13g2_nor2_2 _4675_ (.A(_2220_),
    .B(_2233_),
    .Y(_1576_));
 sg13g2_nand2_1 _4676_ (.Y(_1577_),
    .A(net725),
    .B(net686));
 sg13g2_o21ai_1 _4677_ (.B1(net687),
    .Y(_1578_),
    .A1(net736),
    .A2(net729));
 sg13g2_a21oi_1 _4678_ (.A1(net731),
    .A2(_1403_),
    .Y(_1579_),
    .B1(_1578_));
 sg13g2_xnor2_1 _4679_ (.Y(_1580_),
    .A(_1577_),
    .B(_1579_));
 sg13g2_nand2b_1 _4680_ (.Y(_1581_),
    .B(_1580_),
    .A_N(_1575_));
 sg13g2_xnor2_1 _4681_ (.Y(_1582_),
    .A(_1575_),
    .B(_1580_));
 sg13g2_and2_1 _4682_ (.A(_1359_),
    .B(_1582_),
    .X(_1583_));
 sg13g2_xnor2_1 _4683_ (.Y(_1584_),
    .A(_1359_),
    .B(_1582_));
 sg13g2_nand2_1 _4684_ (.Y(_1585_),
    .A(_1508_),
    .B(_1516_));
 sg13g2_nand2_2 _4685_ (.Y(_1586_),
    .A(net759),
    .B(net702));
 sg13g2_nand2_1 _4686_ (.Y(_1587_),
    .A(net760),
    .B(net694));
 sg13g2_nand2_1 _4687_ (.Y(_1588_),
    .A(net761),
    .B(net699));
 sg13g2_xor2_1 _4688_ (.B(_1588_),
    .A(_1511_),
    .X(_1589_));
 sg13g2_nand2b_1 _4689_ (.Y(_1590_),
    .B(_1589_),
    .A_N(_1586_));
 sg13g2_xnor2_1 _4690_ (.Y(_1591_),
    .A(_1586_),
    .B(_1589_));
 sg13g2_inv_1 _4691_ (.Y(_1592_),
    .A(_1591_));
 sg13g2_o21ai_1 _4692_ (.B1(_1506_),
    .Y(_1593_),
    .A1(_1408_),
    .A2(_1504_));
 sg13g2_nand2_1 _4693_ (.Y(_1594_),
    .A(net713),
    .B(net692));
 sg13g2_nand2_2 _4694_ (.Y(_1595_),
    .A(net717),
    .B(net690));
 sg13g2_xor2_1 _4695_ (.B(_1595_),
    .A(_1503_),
    .X(_1596_));
 sg13g2_nand2b_1 _4696_ (.Y(_1597_),
    .B(_1596_),
    .A_N(_1594_));
 sg13g2_xnor2_1 _4697_ (.Y(_1598_),
    .A(_1594_),
    .B(_1596_));
 sg13g2_nand2_1 _4698_ (.Y(_1599_),
    .A(_1593_),
    .B(_1598_));
 sg13g2_xnor2_1 _4699_ (.Y(_1600_),
    .A(_1593_),
    .B(_1598_));
 sg13g2_xnor2_1 _4700_ (.Y(_1601_),
    .A(_1592_),
    .B(_1600_));
 sg13g2_nor2_1 _4701_ (.A(_1497_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_xor2_1 _4702_ (.B(_1601_),
    .A(_1497_),
    .X(_1603_));
 sg13g2_xnor2_1 _4703_ (.Y(_1604_),
    .A(_1585_),
    .B(_1603_));
 sg13g2_nor2_1 _4704_ (.A(_1584_),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_xnor2_1 _4705_ (.Y(_1606_),
    .A(_1584_),
    .B(_1604_));
 sg13g2_inv_1 _4706_ (.Y(_1607_),
    .A(_1606_));
 sg13g2_xor2_1 _4707_ (.B(_1606_),
    .A(_1521_),
    .X(_1608_));
 sg13g2_o21ai_1 _4708_ (.B1(_1553_),
    .Y(_1609_),
    .A1(_1540_),
    .A2(_1554_));
 sg13g2_o21ai_1 _4709_ (.B1(_1536_),
    .Y(_1610_),
    .A1(_1453_),
    .A2(_1534_));
 sg13g2_nand2_2 _4710_ (.Y(_1611_),
    .A(net742),
    .B(net630));
 sg13g2_nor3_1 _4711_ (.A(_2225_),
    .B(_2230_),
    .C(_1534_),
    .Y(_1612_));
 sg13g2_a22oi_1 _4712_ (.Y(_1613_),
    .B1(net620),
    .B2(net747),
    .A2(net626),
    .A1(net746));
 sg13g2_nor3_1 _4713_ (.A(_1611_),
    .B(_1612_),
    .C(_1613_),
    .Y(_1614_));
 sg13g2_o21ai_1 _4714_ (.B1(_1611_),
    .Y(_1615_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_nor2b_2 _4715_ (.A(_1614_),
    .B_N(_1615_),
    .Y(_1616_));
 sg13g2_nand2_1 _4716_ (.Y(_1617_),
    .A(_1610_),
    .B(_1616_));
 sg13g2_xnor2_1 _4717_ (.Y(_1618_),
    .A(_1610_),
    .B(_1616_));
 sg13g2_xnor2_1 _4718_ (.Y(_1619_),
    .A(_1531_),
    .B(_1618_));
 sg13g2_a21o_1 _4719_ (.A2(_1549_),
    .A1(_1543_),
    .B1(_1551_),
    .X(_1620_));
 sg13g2_o21ai_1 _4720_ (.B1(_1547_),
    .Y(_1621_),
    .A1(_1544_),
    .A2(_1548_));
 sg13g2_o21ai_1 _4721_ (.B1(_1514_),
    .Y(_1622_),
    .A1(_1416_),
    .A2(_1512_));
 sg13g2_nand2_1 _4722_ (.Y(_1623_),
    .A(net749),
    .B(net616));
 sg13g2_nand2_1 _4723_ (.Y(_1624_),
    .A(net752),
    .B(net705));
 sg13g2_nand2_1 _4724_ (.Y(_1625_),
    .A(net752),
    .B(net612));
 sg13g2_or2_1 _4725_ (.X(_1626_),
    .B(_1624_),
    .A(_1546_));
 sg13g2_xnor2_1 _4726_ (.Y(_1627_),
    .A(_1545_),
    .B(_1625_));
 sg13g2_xor2_1 _4727_ (.B(_1627_),
    .A(_1623_),
    .X(_1628_));
 sg13g2_xnor2_1 _4728_ (.Y(_1629_),
    .A(_1622_),
    .B(_1628_));
 sg13g2_nor2b_1 _4729_ (.A(_1629_),
    .B_N(_1621_),
    .Y(_1630_));
 sg13g2_xnor2_1 _4730_ (.Y(_1631_),
    .A(_1621_),
    .B(_1629_));
 sg13g2_nand2_1 _4731_ (.Y(_1632_),
    .A(_1620_),
    .B(_1631_));
 sg13g2_xnor2_1 _4732_ (.Y(_1633_),
    .A(_1620_),
    .B(_1631_));
 sg13g2_xor2_1 _4733_ (.B(_1633_),
    .A(_1619_),
    .X(_1634_));
 sg13g2_nor2b_1 _4734_ (.A(_1518_),
    .B_N(_1634_),
    .Y(_1635_));
 sg13g2_xnor2_1 _4735_ (.Y(_1636_),
    .A(_1518_),
    .B(_1634_));
 sg13g2_and2_1 _4736_ (.A(_1609_),
    .B(_1636_),
    .X(_1637_));
 sg13g2_xnor2_1 _4737_ (.Y(_1638_),
    .A(_1609_),
    .B(_1636_));
 sg13g2_nor2_1 _4738_ (.A(_1608_),
    .B(_1638_),
    .Y(_1639_));
 sg13g2_xor2_1 _4739_ (.B(_1638_),
    .A(_1608_),
    .X(_1640_));
 sg13g2_and2_1 _4740_ (.A(_1574_),
    .B(_1640_),
    .X(_1641_));
 sg13g2_or2_1 _4741_ (.X(_1642_),
    .B(_1640_),
    .A(_1574_));
 sg13g2_nand2b_1 _4742_ (.Y(_1643_),
    .B(_1642_),
    .A_N(_1641_));
 sg13g2_o21ai_1 _4743_ (.B1(_1528_),
    .Y(_1644_),
    .A1(_1338_),
    .A2(_1527_));
 sg13g2_inv_2 _4744_ (.Y(_1645_),
    .A(_1644_));
 sg13g2_o21ai_1 _4745_ (.B1(_1538_),
    .Y(_1646_),
    .A1(_1531_),
    .A2(_1539_));
 sg13g2_o21ai_1 _4746_ (.B1(_1646_),
    .Y(_1647_),
    .A1(_1556_),
    .A2(_1558_));
 sg13g2_or3_1 _4747_ (.A(_1556_),
    .B(_1558_),
    .C(_1646_),
    .X(_1648_));
 sg13g2_nand2_1 _4748_ (.Y(_1649_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_xnor2_1 _4749_ (.Y(_1650_),
    .A(_1644_),
    .B(_1649_));
 sg13g2_xnor2_1 _4750_ (.Y(_1651_),
    .A(_1643_),
    .B(_1650_));
 sg13g2_nand2b_1 _4751_ (.Y(_1652_),
    .B(_1651_),
    .A_N(_1573_));
 sg13g2_nor2b_1 _4752_ (.A(_1651_),
    .B_N(_1573_),
    .Y(_1653_));
 sg13g2_xor2_1 _4753_ (.B(_1651_),
    .A(_1573_),
    .X(_1654_));
 sg13g2_xnor2_1 _4754_ (.Y(_1655_),
    .A(_1572_),
    .B(_1654_));
 sg13g2_a21o_2 _4755_ (.A2(_1563_),
    .A1(_1486_),
    .B1(_1565_),
    .X(_1656_));
 sg13g2_nor2b_1 _4756_ (.A(_1655_),
    .B_N(_1656_),
    .Y(_1657_));
 sg13g2_nand2b_1 _4757_ (.Y(_1658_),
    .B(_1656_),
    .A_N(_1655_));
 sg13g2_xnor2_1 _4758_ (.Y(_1659_),
    .A(_1655_),
    .B(_1656_));
 sg13g2_or3_1 _4759_ (.A(_1473_),
    .B(_1480_),
    .C(_1567_),
    .X(_1660_));
 sg13g2_nand2b_1 _4760_ (.Y(_1661_),
    .B(_1660_),
    .A_N(_1568_));
 sg13g2_nand3b_1 _4761_ (.B(_1659_),
    .C(_1660_),
    .Y(_1662_),
    .A_N(_1568_));
 sg13g2_xnor2_1 _4762_ (.Y(_1663_),
    .A(_1659_),
    .B(_1661_));
 sg13g2_o21ai_1 _4763_ (.B1(net793),
    .Y(_1664_),
    .A1(net610),
    .A2(_1663_));
 sg13g2_a21oi_1 _4764_ (.A1(net610),
    .A2(_2196_),
    .Y(_0183_),
    .B1(_1664_));
 sg13g2_o21ai_1 _4765_ (.B1(_1652_),
    .Y(_1665_),
    .A1(_1572_),
    .A2(_1653_));
 sg13g2_o21ai_1 _4766_ (.B1(_1647_),
    .Y(_1666_),
    .A1(_1645_),
    .A2(_1649_));
 sg13g2_a21oi_1 _4767_ (.A1(_1642_),
    .A2(_1650_),
    .Y(_1667_),
    .B1(_1641_));
 sg13g2_a21oi_1 _4768_ (.A1(_1521_),
    .A2(_1607_),
    .Y(_1668_),
    .B1(_1639_));
 sg13g2_mux2_1 _4769_ (.A0(_2220_),
    .A1(_1576_),
    .S(_1495_),
    .X(_1669_));
 sg13g2_nor2_2 _4770_ (.A(_2221_),
    .B(_2233_),
    .Y(_1670_));
 sg13g2_xor2_1 _4771_ (.B(_1670_),
    .A(_1669_),
    .X(_1671_));
 sg13g2_o21ai_1 _4772_ (.B1(_1496_),
    .Y(_1672_),
    .A1(_1577_),
    .A2(_1578_));
 sg13g2_nand2_1 _4773_ (.Y(_1673_),
    .A(_1671_),
    .B(_1672_));
 sg13g2_xor2_1 _4774_ (.B(_1672_),
    .A(_1671_),
    .X(_1674_));
 sg13g2_inv_1 _4775_ (.Y(_1675_),
    .A(_1674_));
 sg13g2_xnor2_1 _4776_ (.Y(_1676_),
    .A(_1405_),
    .B(_1674_));
 sg13g2_nand2_1 _4777_ (.Y(_1677_),
    .A(_1583_),
    .B(_1676_));
 sg13g2_xnor2_1 _4778_ (.Y(_1678_),
    .A(_1583_),
    .B(_1676_));
 sg13g2_o21ai_1 _4779_ (.B1(_1599_),
    .Y(_1679_),
    .A1(_1592_),
    .A2(_1600_));
 sg13g2_nand2_1 _4780_ (.Y(_1680_),
    .A(net754),
    .B(net701));
 sg13g2_nand2_1 _4781_ (.Y(_1681_),
    .A(net757),
    .B(net695));
 sg13g2_nand2_1 _4782_ (.Y(_1682_),
    .A(net757),
    .B(net698));
 sg13g2_xor2_1 _4783_ (.B(_1682_),
    .A(_1587_),
    .X(_1683_));
 sg13g2_nand2b_1 _4784_ (.Y(_1684_),
    .B(_1683_),
    .A_N(_1680_));
 sg13g2_xor2_1 _4785_ (.B(_1683_),
    .A(_1680_),
    .X(_1685_));
 sg13g2_o21ai_1 _4786_ (.B1(_1597_),
    .Y(_1686_),
    .A1(_1503_),
    .A2(_1595_));
 sg13g2_nand2_1 _4787_ (.Y(_1687_),
    .A(net709),
    .B(net692));
 sg13g2_nand2_2 _4788_ (.Y(_1688_),
    .A(net715),
    .B(net689));
 sg13g2_nor2_1 _4789_ (.A(_1595_),
    .B(_1688_),
    .Y(_1689_));
 sg13g2_or2_1 _4790_ (.X(_1690_),
    .B(_1688_),
    .A(_1595_));
 sg13g2_a22oi_1 _4791_ (.Y(_1691_),
    .B1(net689),
    .B2(net717),
    .A2(net691),
    .A1(net713));
 sg13g2_or2_1 _4792_ (.X(_1692_),
    .B(_1691_),
    .A(_1689_));
 sg13g2_xor2_1 _4793_ (.B(_1692_),
    .A(_1687_),
    .X(_1693_));
 sg13g2_nand2_1 _4794_ (.Y(_1694_),
    .A(_1686_),
    .B(_1693_));
 sg13g2_xnor2_1 _4795_ (.Y(_1695_),
    .A(_1686_),
    .B(_1693_));
 sg13g2_xnor2_1 _4796_ (.Y(_1696_),
    .A(_1685_),
    .B(_1695_));
 sg13g2_nor2_1 _4797_ (.A(_1581_),
    .B(_1696_),
    .Y(_1697_));
 sg13g2_xor2_1 _4798_ (.B(_1696_),
    .A(_1581_),
    .X(_1698_));
 sg13g2_xnor2_1 _4799_ (.Y(_1699_),
    .A(_1679_),
    .B(_1698_));
 sg13g2_xor2_1 _4800_ (.B(_1699_),
    .A(_1678_),
    .X(_1700_));
 sg13g2_xnor2_1 _4801_ (.Y(_1701_),
    .A(_1605_),
    .B(_1700_));
 sg13g2_o21ai_1 _4802_ (.B1(_1632_),
    .Y(_1702_),
    .A1(_1619_),
    .A2(_1633_));
 sg13g2_a21oi_1 _4803_ (.A1(_1585_),
    .A2(_1603_),
    .Y(_1703_),
    .B1(_1602_));
 sg13g2_a21o_1 _4804_ (.A2(_1628_),
    .A1(_1622_),
    .B1(_1630_),
    .X(_1704_));
 sg13g2_o21ai_1 _4805_ (.B1(_1626_),
    .Y(_1705_),
    .A1(_1623_),
    .A2(_1627_));
 sg13g2_o21ai_1 _4806_ (.B1(_1590_),
    .Y(_1706_),
    .A1(_1511_),
    .A2(_1588_));
 sg13g2_nand2_1 _4807_ (.Y(_1707_),
    .A(net747),
    .B(net616));
 sg13g2_nand2_1 _4808_ (.Y(_1708_),
    .A(net749),
    .B(net706));
 sg13g2_nand2_1 _4809_ (.Y(_1709_),
    .A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .B(net613));
 sg13g2_or2_1 _4810_ (.X(_1710_),
    .B(_1708_),
    .A(_1625_));
 sg13g2_xnor2_1 _4811_ (.Y(_1711_),
    .A(_1624_),
    .B(_1709_));
 sg13g2_xor2_1 _4812_ (.B(_1711_),
    .A(_1707_),
    .X(_1712_));
 sg13g2_xnor2_1 _4813_ (.Y(_1713_),
    .A(_1706_),
    .B(_1712_));
 sg13g2_nor2b_1 _4814_ (.A(_1713_),
    .B_N(_1705_),
    .Y(_1714_));
 sg13g2_xnor2_1 _4815_ (.Y(_1715_),
    .A(_1705_),
    .B(_1713_));
 sg13g2_nand2_1 _4816_ (.Y(_1716_),
    .A(_1704_),
    .B(_1715_));
 sg13g2_xnor2_1 _4817_ (.Y(_1717_),
    .A(_1704_),
    .B(_1715_));
 sg13g2_or2_1 _4818_ (.X(_1718_),
    .B(_1614_),
    .A(_1612_));
 sg13g2_a22oi_1 _4819_ (.Y(_1719_),
    .B1(net621),
    .B2(net746),
    .A2(net626),
    .A1(net743));
 sg13g2_nand4_1 _4820_ (.B(net743),
    .C(net626),
    .A(net746),
    .Y(_1720_),
    .D(net621));
 sg13g2_nor2b_1 _4821_ (.A(_1719_),
    .B_N(_1720_),
    .Y(_1721_));
 sg13g2_xnor2_1 _4822_ (.Y(_1722_),
    .A(_1611_),
    .B(_1721_));
 sg13g2_nand2_1 _4823_ (.Y(_1723_),
    .A(_1718_),
    .B(_1722_));
 sg13g2_xnor2_1 _4824_ (.Y(_1724_),
    .A(_1718_),
    .B(_1722_));
 sg13g2_xnor2_1 _4825_ (.Y(_1725_),
    .A(_1531_),
    .B(_1724_));
 sg13g2_xor2_1 _4826_ (.B(_1725_),
    .A(_1717_),
    .X(_1726_));
 sg13g2_nor2b_1 _4827_ (.A(_1703_),
    .B_N(_1726_),
    .Y(_1727_));
 sg13g2_xnor2_1 _4828_ (.Y(_1728_),
    .A(_1703_),
    .B(_1726_));
 sg13g2_and2_1 _4829_ (.A(_1702_),
    .B(_1728_),
    .X(_1729_));
 sg13g2_xnor2_1 _4830_ (.Y(_1730_),
    .A(_1702_),
    .B(_1728_));
 sg13g2_nor2_1 _4831_ (.A(_1701_),
    .B(_1730_),
    .Y(_1731_));
 sg13g2_xnor2_1 _4832_ (.Y(_1732_),
    .A(_1701_),
    .B(_1730_));
 sg13g2_nor2_1 _4833_ (.A(_1668_),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_xor2_1 _4834_ (.B(_1732_),
    .A(_1668_),
    .X(_1734_));
 sg13g2_o21ai_1 _4835_ (.B1(_1617_),
    .Y(_1735_),
    .A1(_1531_),
    .A2(_1618_));
 sg13g2_o21ai_1 _4836_ (.B1(_1735_),
    .Y(_1736_),
    .A1(_1635_),
    .A2(_1637_));
 sg13g2_or3_1 _4837_ (.A(_1635_),
    .B(_1637_),
    .C(_1735_),
    .X(_1737_));
 sg13g2_nand2_1 _4838_ (.Y(_1738_),
    .A(_1736_),
    .B(_1737_));
 sg13g2_xnor2_1 _4839_ (.Y(_1739_),
    .A(_1644_),
    .B(_1738_));
 sg13g2_xnor2_1 _4840_ (.Y(_1740_),
    .A(_1734_),
    .B(_1739_));
 sg13g2_xor2_1 _4841_ (.B(_1740_),
    .A(_1667_),
    .X(_1741_));
 sg13g2_nand2_1 _4842_ (.Y(_1742_),
    .A(_1666_),
    .B(_1741_));
 sg13g2_xnor2_1 _4843_ (.Y(_1743_),
    .A(_1666_),
    .B(_1741_));
 sg13g2_nand2b_1 _4844_ (.Y(_1744_),
    .B(_1743_),
    .A_N(_1665_));
 sg13g2_nor2b_1 _4845_ (.A(_1743_),
    .B_N(_1665_),
    .Y(_1745_));
 sg13g2_xor2_1 _4846_ (.B(_1743_),
    .A(_1665_),
    .X(_1746_));
 sg13g2_nand3_1 _4847_ (.B(_1662_),
    .C(_1746_),
    .A(_1658_),
    .Y(_1747_));
 sg13g2_a21o_2 _4848_ (.A2(_1662_),
    .A1(_1658_),
    .B1(_1746_),
    .X(_1748_));
 sg13g2_a21oi_1 _4849_ (.A1(_1747_),
    .A2(_1748_),
    .Y(_1749_),
    .B1(net610));
 sg13g2_o21ai_1 _4850_ (.B1(net796),
    .Y(_1750_),
    .A1(net673),
    .A2(net286));
 sg13g2_nor2_1 _4851_ (.A(_1749_),
    .B(net287),
    .Y(_0184_));
 sg13g2_o21ai_1 _4852_ (.B1(_1744_),
    .Y(_1751_),
    .A1(_1657_),
    .A2(_1745_));
 sg13g2_o21ai_1 _4853_ (.B1(_1751_),
    .Y(_1752_),
    .A1(_1662_),
    .A2(_1746_));
 sg13g2_o21ai_1 _4854_ (.B1(_1742_),
    .Y(_1753_),
    .A1(_1667_),
    .A2(_1740_));
 sg13g2_o21ai_1 _4855_ (.B1(_1736_),
    .Y(_1754_),
    .A1(_1645_),
    .A2(_1738_));
 sg13g2_a21oi_1 _4856_ (.A1(_1734_),
    .A2(_1739_),
    .Y(_1755_),
    .B1(_1733_));
 sg13g2_a21oi_1 _4857_ (.A1(_1605_),
    .A2(_1700_),
    .Y(_1756_),
    .B1(_1731_));
 sg13g2_o21ai_1 _4858_ (.B1(_1677_),
    .Y(_1757_),
    .A1(_1678_),
    .A2(_1699_));
 sg13g2_a22oi_1 _4859_ (.Y(_1758_),
    .B1(_1669_),
    .B2(_1670_),
    .A2(_1576_),
    .A1(net729));
 sg13g2_nand2_1 _4860_ (.Y(_1759_),
    .A(net720),
    .B(_1576_));
 sg13g2_o21ai_1 _4861_ (.B1(_1759_),
    .Y(_1760_),
    .A1(_1576_),
    .A2(_1670_));
 sg13g2_and2_1 _4862_ (.A(net717),
    .B(net686),
    .X(_1761_));
 sg13g2_nor2b_1 _4863_ (.A(_1760_),
    .B_N(_1761_),
    .Y(_1762_));
 sg13g2_xnor2_1 _4864_ (.Y(_1763_),
    .A(_1760_),
    .B(_1761_));
 sg13g2_nand2b_1 _4865_ (.Y(_1764_),
    .B(_1763_),
    .A_N(_1404_));
 sg13g2_xnor2_1 _4866_ (.Y(_1765_),
    .A(_1404_),
    .B(_1763_));
 sg13g2_inv_1 _4867_ (.Y(_1766_),
    .A(_1765_));
 sg13g2_xnor2_1 _4868_ (.Y(_1767_),
    .A(_1758_),
    .B(_1765_));
 sg13g2_nand2_1 _4869_ (.Y(_1768_),
    .A(_1499_),
    .B(_1767_));
 sg13g2_xnor2_1 _4870_ (.Y(_1769_),
    .A(_1499_),
    .B(_1767_));
 sg13g2_nor3_1 _4871_ (.A(net556),
    .B(_1675_),
    .C(_1769_),
    .Y(_1770_));
 sg13g2_o21ai_1 _4872_ (.B1(_1769_),
    .Y(_1771_),
    .A1(net556),
    .A2(_1675_));
 sg13g2_nand2b_1 _4873_ (.Y(_1772_),
    .B(_1771_),
    .A_N(_1770_));
 sg13g2_o21ai_1 _4874_ (.B1(_1694_),
    .Y(_1773_),
    .A1(_1685_),
    .A2(_1695_));
 sg13g2_nand2_1 _4875_ (.Y(_1774_),
    .A(net751),
    .B(net701));
 sg13g2_nand2_1 _4876_ (.Y(_1775_),
    .A(net755),
    .B(net696));
 sg13g2_nand2_1 _4877_ (.Y(_1776_),
    .A(net754),
    .B(net699));
 sg13g2_xor2_1 _4878_ (.B(_1776_),
    .A(_1681_),
    .X(_1777_));
 sg13g2_nand2b_1 _4879_ (.Y(_1778_),
    .B(_1777_),
    .A_N(_1774_));
 sg13g2_xnor2_1 _4880_ (.Y(_1779_),
    .A(_1774_),
    .B(_1777_));
 sg13g2_inv_1 _4881_ (.Y(_1780_),
    .A(_1779_));
 sg13g2_o21ai_1 _4882_ (.B1(_1690_),
    .Y(_1781_),
    .A1(_1687_),
    .A2(_1692_));
 sg13g2_nand2_1 _4883_ (.Y(_1782_),
    .A(net760),
    .B(net692));
 sg13g2_nand2_1 _4884_ (.Y(_1783_),
    .A(net710),
    .B(net688));
 sg13g2_nand2_1 _4885_ (.Y(_1784_),
    .A(net709),
    .B(net691));
 sg13g2_xor2_1 _4886_ (.B(_1784_),
    .A(_1688_),
    .X(_1785_));
 sg13g2_nand2b_1 _4887_ (.Y(_1786_),
    .B(_1785_),
    .A_N(_1782_));
 sg13g2_xnor2_1 _4888_ (.Y(_1787_),
    .A(_1782_),
    .B(_1785_));
 sg13g2_nand2_1 _4889_ (.Y(_1788_),
    .A(_1781_),
    .B(_1787_));
 sg13g2_xnor2_1 _4890_ (.Y(_1789_),
    .A(_1781_),
    .B(_1787_));
 sg13g2_xnor2_1 _4891_ (.Y(_1790_),
    .A(_1780_),
    .B(_1789_));
 sg13g2_xor2_1 _4892_ (.B(_1790_),
    .A(_1673_),
    .X(_1791_));
 sg13g2_nand2_1 _4893_ (.Y(_1792_),
    .A(_1773_),
    .B(_1791_));
 sg13g2_xnor2_1 _4894_ (.Y(_1793_),
    .A(_1773_),
    .B(_1791_));
 sg13g2_nor2_1 _4895_ (.A(_1772_),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_xor2_1 _4896_ (.B(_1793_),
    .A(_1772_),
    .X(_1795_));
 sg13g2_nand2_1 _4897_ (.Y(_1796_),
    .A(_1757_),
    .B(_1795_));
 sg13g2_xnor2_1 _4898_ (.Y(_1797_),
    .A(_1757_),
    .B(_1795_));
 sg13g2_o21ai_1 _4899_ (.B1(_1716_),
    .Y(_1798_),
    .A1(_1717_),
    .A2(_1725_));
 sg13g2_a21oi_1 _4900_ (.A1(_1679_),
    .A2(_1698_),
    .Y(_1799_),
    .B1(_1697_));
 sg13g2_o21ai_1 _4901_ (.B1(net742),
    .Y(_1800_),
    .A1(net627),
    .A2(net620));
 sg13g2_nand3_1 _4902_ (.B(net627),
    .C(net620),
    .A(net742),
    .Y(_1801_));
 sg13g2_nor2b_1 _4903_ (.A(_1800_),
    .B_N(_1801_),
    .Y(_1802_));
 sg13g2_nand2b_1 _4904_ (.Y(_1803_),
    .B(_1719_),
    .A_N(_1611_));
 sg13g2_o21ai_1 _4905_ (.B1(_1803_),
    .Y(_1804_),
    .A1(net630),
    .A2(_1720_));
 sg13g2_xnor2_1 _4906_ (.Y(_1805_),
    .A(_1802_),
    .B(_1804_));
 sg13g2_xnor2_1 _4907_ (.Y(_1806_),
    .A(_1531_),
    .B(_1805_));
 sg13g2_a21o_1 _4908_ (.A2(_1712_),
    .A1(_1706_),
    .B1(_1714_),
    .X(_1807_));
 sg13g2_o21ai_1 _4909_ (.B1(_1710_),
    .Y(_1808_),
    .A1(_1707_),
    .A2(_1711_));
 sg13g2_o21ai_1 _4910_ (.B1(_1684_),
    .Y(_1809_),
    .A1(_1587_),
    .A2(_1682_));
 sg13g2_nand2_1 _4911_ (.Y(_1810_),
    .A(net745),
    .B(net616));
 sg13g2_nand2_2 _4912_ (.Y(_1811_),
    .A(net747),
    .B(net614));
 sg13g2_or2_1 _4913_ (.X(_1812_),
    .B(_1811_),
    .A(_1708_));
 sg13g2_xnor2_1 _4914_ (.Y(_1813_),
    .A(_1708_),
    .B(_1811_));
 sg13g2_xor2_1 _4915_ (.B(_1813_),
    .A(_1810_),
    .X(_1814_));
 sg13g2_xnor2_1 _4916_ (.Y(_1815_),
    .A(_1809_),
    .B(_1814_));
 sg13g2_nor2b_1 _4917_ (.A(_1815_),
    .B_N(_1808_),
    .Y(_1816_));
 sg13g2_xnor2_1 _4918_ (.Y(_1817_),
    .A(_1808_),
    .B(_1815_));
 sg13g2_nand2_1 _4919_ (.Y(_1818_),
    .A(_1807_),
    .B(_1817_));
 sg13g2_xnor2_1 _4920_ (.Y(_1819_),
    .A(_1807_),
    .B(_1817_));
 sg13g2_xnor2_1 _4921_ (.Y(_1820_),
    .A(_1806_),
    .B(_1819_));
 sg13g2_nor2_1 _4922_ (.A(_1799_),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_xor2_1 _4923_ (.B(_1820_),
    .A(_1799_),
    .X(_1822_));
 sg13g2_xnor2_1 _4924_ (.Y(_1823_),
    .A(_1798_),
    .B(_1822_));
 sg13g2_xnor2_1 _4925_ (.Y(_1824_),
    .A(_1797_),
    .B(_1823_));
 sg13g2_nor2_1 _4926_ (.A(_1756_),
    .B(_1824_),
    .Y(_1825_));
 sg13g2_xor2_1 _4927_ (.B(_1824_),
    .A(_1756_),
    .X(_1826_));
 sg13g2_o21ai_1 _4928_ (.B1(_1723_),
    .Y(_1827_),
    .A1(_1531_),
    .A2(_1724_));
 sg13g2_o21ai_1 _4929_ (.B1(_1827_),
    .Y(_1828_),
    .A1(_1727_),
    .A2(_1729_));
 sg13g2_or3_1 _4930_ (.A(_1727_),
    .B(_1729_),
    .C(_1827_),
    .X(_1829_));
 sg13g2_nand2_1 _4931_ (.Y(_1830_),
    .A(_1828_),
    .B(_1829_));
 sg13g2_xnor2_1 _4932_ (.Y(_1831_),
    .A(_1644_),
    .B(_1830_));
 sg13g2_xnor2_1 _4933_ (.Y(_1832_),
    .A(_1826_),
    .B(_1831_));
 sg13g2_xor2_1 _4934_ (.B(_1832_),
    .A(_1755_),
    .X(_1833_));
 sg13g2_nand2_1 _4935_ (.Y(_1834_),
    .A(_1754_),
    .B(_1833_));
 sg13g2_xor2_1 _4936_ (.B(_1833_),
    .A(_1754_),
    .X(_1835_));
 sg13g2_and2_1 _4937_ (.A(_1753_),
    .B(_1835_),
    .X(_1836_));
 sg13g2_or2_1 _4938_ (.X(_1837_),
    .B(_1835_),
    .A(_1753_));
 sg13g2_nor2b_1 _4939_ (.A(_1836_),
    .B_N(_1837_),
    .Y(_1838_));
 sg13g2_xnor2_1 _4940_ (.Y(_1839_),
    .A(_1752_),
    .B(_1838_));
 sg13g2_o21ai_1 _4941_ (.B1(net793),
    .Y(_1840_),
    .A1(net672),
    .A2(net248));
 sg13g2_a21oi_1 _4942_ (.A1(net672),
    .A2(_1839_),
    .Y(_0185_),
    .B1(_1840_));
 sg13g2_a21oi_1 _4943_ (.A1(_1752_),
    .A2(_1837_),
    .Y(_1841_),
    .B1(_1836_));
 sg13g2_o21ai_1 _4944_ (.B1(_1834_),
    .Y(_1842_),
    .A1(_1755_),
    .A2(_1832_));
 sg13g2_o21ai_1 _4945_ (.B1(_1828_),
    .Y(_1843_),
    .A1(_1645_),
    .A2(_1830_));
 sg13g2_a21oi_1 _4946_ (.A1(_1826_),
    .A2(_1831_),
    .Y(_1844_),
    .B1(_1825_));
 sg13g2_o21ai_1 _4947_ (.B1(_1796_),
    .Y(_1845_),
    .A1(_1797_),
    .A2(_1823_));
 sg13g2_nor2_1 _4948_ (.A(_1770_),
    .B(_1794_),
    .Y(_1846_));
 sg13g2_nand2_1 _4949_ (.Y(_1847_),
    .A(_1359_),
    .B(_1580_));
 sg13g2_xnor2_1 _4950_ (.Y(_1848_),
    .A(_1358_),
    .B(_1580_));
 sg13g2_a21oi_1 _4951_ (.A1(net720),
    .A2(_1576_),
    .Y(_1849_),
    .B1(_1762_));
 sg13g2_nand2_1 _4952_ (.Y(_1850_),
    .A(net720),
    .B(_1761_));
 sg13g2_o21ai_1 _4953_ (.B1(_1850_),
    .Y(_1851_),
    .A1(_1670_),
    .A2(_1761_));
 sg13g2_nand2_1 _4954_ (.Y(_1852_),
    .A(net714),
    .B(net686));
 sg13g2_xor2_1 _4955_ (.B(_1852_),
    .A(_1851_),
    .X(_1853_));
 sg13g2_inv_1 _4956_ (.Y(_1854_),
    .A(_1853_));
 sg13g2_xnor2_1 _4957_ (.Y(_1855_),
    .A(_1575_),
    .B(_1853_));
 sg13g2_nand2b_1 _4958_ (.Y(_1856_),
    .B(_1855_),
    .A_N(_1849_));
 sg13g2_xor2_1 _4959_ (.B(_1855_),
    .A(_1849_),
    .X(_1857_));
 sg13g2_inv_1 _4960_ (.Y(_1858_),
    .A(_1857_));
 sg13g2_nand2_1 _4961_ (.Y(_1859_),
    .A(_1848_),
    .B(_1858_));
 sg13g2_xnor2_1 _4962_ (.Y(_1860_),
    .A(_1848_),
    .B(_1857_));
 sg13g2_nor2b_1 _4963_ (.A(_1768_),
    .B_N(_1860_),
    .Y(_1861_));
 sg13g2_xnor2_1 _4964_ (.Y(_1862_),
    .A(_1768_),
    .B(_1860_));
 sg13g2_o21ai_1 _4965_ (.B1(_1788_),
    .Y(_1863_),
    .A1(_1780_),
    .A2(_1789_));
 sg13g2_o21ai_1 _4966_ (.B1(_1764_),
    .Y(_1864_),
    .A1(_1758_),
    .A2(_1766_));
 sg13g2_nand2_1 _4967_ (.Y(_1865_),
    .A(net749),
    .B(net702));
 sg13g2_nand2_1 _4968_ (.Y(_1866_),
    .A(net751),
    .B(net696));
 sg13g2_nand2_1 _4969_ (.Y(_1867_),
    .A(net751),
    .B(net700));
 sg13g2_xor2_1 _4970_ (.B(_1867_),
    .A(_1775_),
    .X(_1868_));
 sg13g2_nand2b_1 _4971_ (.Y(_1869_),
    .B(_1868_),
    .A_N(_1865_));
 sg13g2_xnor2_1 _4972_ (.Y(_1870_),
    .A(_1865_),
    .B(_1868_));
 sg13g2_inv_1 _4973_ (.Y(_1871_),
    .A(_1870_));
 sg13g2_o21ai_1 _4974_ (.B1(_1786_),
    .Y(_1872_),
    .A1(_1688_),
    .A2(_1784_));
 sg13g2_nand2_1 _4975_ (.Y(_1873_),
    .A(net758),
    .B(net693));
 sg13g2_nand2_2 _4976_ (.Y(_1874_),
    .A(net760),
    .B(net690));
 sg13g2_xor2_1 _4977_ (.B(_1874_),
    .A(_1783_),
    .X(_1875_));
 sg13g2_nand2b_1 _4978_ (.Y(_1876_),
    .B(_1875_),
    .A_N(_1873_));
 sg13g2_xnor2_1 _4979_ (.Y(_1877_),
    .A(_1873_),
    .B(_1875_));
 sg13g2_nand2_1 _4980_ (.Y(_1878_),
    .A(_1872_),
    .B(_1877_));
 sg13g2_xnor2_1 _4981_ (.Y(_1879_),
    .A(_1872_),
    .B(_1877_));
 sg13g2_xnor2_1 _4982_ (.Y(_1880_),
    .A(_1870_),
    .B(_1879_));
 sg13g2_xnor2_1 _4983_ (.Y(_1881_),
    .A(_1864_),
    .B(_1880_));
 sg13g2_nor2b_1 _4984_ (.A(_1881_),
    .B_N(_1863_),
    .Y(_1882_));
 sg13g2_xor2_1 _4985_ (.B(_1881_),
    .A(_1863_),
    .X(_1883_));
 sg13g2_inv_1 _4986_ (.Y(_1884_),
    .A(_1883_));
 sg13g2_xor2_1 _4987_ (.B(_1883_),
    .A(_1862_),
    .X(_1885_));
 sg13g2_or2_1 _4988_ (.X(_1886_),
    .B(_1885_),
    .A(_1846_));
 sg13g2_xnor2_1 _4989_ (.Y(_1887_),
    .A(_1846_),
    .B(_1885_));
 sg13g2_o21ai_1 _4990_ (.B1(_1818_),
    .Y(_1888_),
    .A1(_1806_),
    .A2(_1819_));
 sg13g2_o21ai_1 _4991_ (.B1(_1792_),
    .Y(_1889_),
    .A1(_1673_),
    .A2(_1790_));
 sg13g2_nand4_1 _4992_ (.B(net630),
    .C(net627),
    .A(net742),
    .Y(_1890_),
    .D(net620));
 sg13g2_inv_1 _4993_ (.Y(_1891_),
    .A(_1890_));
 sg13g2_a21oi_1 _4994_ (.A1(_1611_),
    .A2(_1800_),
    .Y(_1892_),
    .B1(_1891_));
 sg13g2_xnor2_1 _4995_ (.Y(_1893_),
    .A(_1530_),
    .B(_1892_));
 sg13g2_a21o_2 _4996_ (.A2(_1814_),
    .A1(_1809_),
    .B1(_1816_),
    .X(_1894_));
 sg13g2_o21ai_1 _4997_ (.B1(_1812_),
    .Y(_1895_),
    .A1(_1810_),
    .A2(_1813_));
 sg13g2_o21ai_1 _4998_ (.B1(_1778_),
    .Y(_1896_),
    .A1(_1681_),
    .A2(_1776_));
 sg13g2_nand2_2 _4999_ (.Y(_1897_),
    .A(net743),
    .B(net617));
 sg13g2_nor3_1 _5000_ (.A(_2225_),
    .B(_2232_),
    .C(_1811_),
    .Y(_1898_));
 sg13g2_a22oi_1 _5001_ (.Y(_1899_),
    .B1(net704),
    .B2(net747),
    .A2(net611),
    .A1(net745));
 sg13g2_nor3_1 _5002_ (.A(_1897_),
    .B(_1898_),
    .C(_1899_),
    .Y(_1900_));
 sg13g2_o21ai_1 _5003_ (.B1(_1897_),
    .Y(_1901_),
    .A1(_1898_),
    .A2(_1899_));
 sg13g2_nor2b_1 _5004_ (.A(_1900_),
    .B_N(_1901_),
    .Y(_1902_));
 sg13g2_xnor2_1 _5005_ (.Y(_1903_),
    .A(_1896_),
    .B(_1902_));
 sg13g2_nor2b_1 _5006_ (.A(_1903_),
    .B_N(_1895_),
    .Y(_1904_));
 sg13g2_xor2_1 _5007_ (.B(_1903_),
    .A(_1895_),
    .X(_1905_));
 sg13g2_inv_1 _5008_ (.Y(_1906_),
    .A(_1905_));
 sg13g2_xnor2_1 _5009_ (.Y(_1907_),
    .A(_1894_),
    .B(_1906_));
 sg13g2_nor2_1 _5010_ (.A(_1893_),
    .B(_1907_),
    .Y(_1908_));
 sg13g2_xor2_1 _5011_ (.B(_1907_),
    .A(_1893_),
    .X(_1909_));
 sg13g2_xor2_1 _5012_ (.B(_1909_),
    .A(_1889_),
    .X(_1910_));
 sg13g2_and2_1 _5013_ (.A(_1888_),
    .B(_1910_),
    .X(_1911_));
 sg13g2_xnor2_1 _5014_ (.Y(_1912_),
    .A(_1888_),
    .B(_1910_));
 sg13g2_xnor2_1 _5015_ (.Y(_1913_),
    .A(_1887_),
    .B(_1912_));
 sg13g2_nor2b_1 _5016_ (.A(_1913_),
    .B_N(_1845_),
    .Y(_1914_));
 sg13g2_nand2b_1 _5017_ (.Y(_1915_),
    .B(_1913_),
    .A_N(_1845_));
 sg13g2_nand2b_1 _5018_ (.Y(_1916_),
    .B(_1915_),
    .A_N(_1914_));
 sg13g2_a21oi_1 _5019_ (.A1(_1798_),
    .A2(_1822_),
    .Y(_1917_),
    .B1(_1821_));
 sg13g2_o21ai_1 _5020_ (.B1(_1890_),
    .Y(_1918_),
    .A1(_1531_),
    .A2(_1805_));
 sg13g2_nand2b_1 _5021_ (.Y(_1919_),
    .B(_1918_),
    .A_N(_1917_));
 sg13g2_xor2_1 _5022_ (.B(_1918_),
    .A(_1917_),
    .X(_1920_));
 sg13g2_xnor2_1 _5023_ (.Y(_1921_),
    .A(_1644_),
    .B(_1920_));
 sg13g2_xnor2_1 _5024_ (.Y(_1922_),
    .A(_1916_),
    .B(_1921_));
 sg13g2_nor2b_1 _5025_ (.A(_1844_),
    .B_N(_1922_),
    .Y(_1923_));
 sg13g2_xnor2_1 _5026_ (.Y(_1924_),
    .A(_1844_),
    .B(_1922_));
 sg13g2_xor2_1 _5027_ (.B(_1924_),
    .A(_1843_),
    .X(_1925_));
 sg13g2_nand2_1 _5028_ (.Y(_1926_),
    .A(_1842_),
    .B(_1925_));
 sg13g2_xnor2_1 _5029_ (.Y(_1927_),
    .A(_1842_),
    .B(_1925_));
 sg13g2_xnor2_1 _5030_ (.Y(_1928_),
    .A(_1841_),
    .B(_1927_));
 sg13g2_o21ai_1 _5031_ (.B1(net796),
    .Y(_1929_),
    .A1(net672),
    .A2(net290));
 sg13g2_a21oi_1 _5032_ (.A1(net672),
    .A2(_1928_),
    .Y(_0186_),
    .B1(_1929_));
 sg13g2_o21ai_1 _5033_ (.B1(_1926_),
    .Y(_1930_),
    .A1(_1841_),
    .A2(_1927_));
 sg13g2_a21o_1 _5034_ (.A2(_1924_),
    .A1(_1843_),
    .B1(_1923_),
    .X(_1931_));
 sg13g2_o21ai_1 _5035_ (.B1(_1919_),
    .Y(_1932_),
    .A1(_1645_),
    .A2(_1920_));
 sg13g2_a21oi_1 _5036_ (.A1(_1915_),
    .A2(_1921_),
    .Y(_1933_),
    .B1(_1914_));
 sg13g2_a21oi_1 _5037_ (.A1(_1889_),
    .A2(_1909_),
    .Y(_1934_),
    .B1(_1911_));
 sg13g2_a21o_2 _5038_ (.A2(_1892_),
    .A1(_1530_),
    .B1(_1891_),
    .X(_1935_));
 sg13g2_nand2b_1 _5039_ (.Y(_1936_),
    .B(_1935_),
    .A_N(_1934_));
 sg13g2_xor2_1 _5040_ (.B(_1935_),
    .A(_1934_),
    .X(_1937_));
 sg13g2_xnor2_1 _5041_ (.Y(_1938_),
    .A(_1644_),
    .B(_1937_));
 sg13g2_o21ai_1 _5042_ (.B1(_1886_),
    .Y(_1939_),
    .A1(_1887_),
    .A2(_1912_));
 sg13g2_a21oi_1 _5043_ (.A1(_1894_),
    .A2(_1906_),
    .Y(_1940_),
    .B1(_1908_));
 sg13g2_a21o_1 _5044_ (.A2(_1880_),
    .A1(_1864_),
    .B1(_1882_),
    .X(_1941_));
 sg13g2_a21o_1 _5045_ (.A2(_1902_),
    .A1(_1896_),
    .B1(_1904_),
    .X(_1942_));
 sg13g2_or2_1 _5046_ (.X(_1943_),
    .B(_1900_),
    .A(_1898_));
 sg13g2_o21ai_1 _5047_ (.B1(_1869_),
    .Y(_1944_),
    .A1(_1775_),
    .A2(_1867_));
 sg13g2_and4_1 _5048_ (.A(net745),
    .B(net743),
    .C(net611),
    .D(net707),
    .X(_1945_));
 sg13g2_a22oi_1 _5049_ (.Y(_1946_),
    .B1(net704),
    .B2(net745),
    .A2(net611),
    .A1(net743));
 sg13g2_nor3_1 _5050_ (.A(_1897_),
    .B(_1945_),
    .C(_1946_),
    .Y(_1947_));
 sg13g2_o21ai_1 _5051_ (.B1(_1897_),
    .Y(_1948_),
    .A1(_1945_),
    .A2(_1946_));
 sg13g2_nor2b_1 _5052_ (.A(_1947_),
    .B_N(_1948_),
    .Y(_1949_));
 sg13g2_xnor2_1 _5053_ (.Y(_1950_),
    .A(_1944_),
    .B(_1949_));
 sg13g2_nor2b_1 _5054_ (.A(_1950_),
    .B_N(_1943_),
    .Y(_1951_));
 sg13g2_xnor2_1 _5055_ (.Y(_1952_),
    .A(_1943_),
    .B(_1950_));
 sg13g2_nand2_1 _5056_ (.Y(_1953_),
    .A(_1942_),
    .B(_1952_));
 sg13g2_xnor2_1 _5057_ (.Y(_1954_),
    .A(_1942_),
    .B(_1952_));
 sg13g2_xor2_1 _5058_ (.B(_1954_),
    .A(_1893_),
    .X(_1955_));
 sg13g2_nand2_1 _5059_ (.Y(_1956_),
    .A(_1941_),
    .B(_1955_));
 sg13g2_xnor2_1 _5060_ (.Y(_1957_),
    .A(_1941_),
    .B(_1955_));
 sg13g2_xnor2_1 _5061_ (.Y(_1958_),
    .A(_1940_),
    .B(_1957_));
 sg13g2_a21oi_1 _5062_ (.A1(_1862_),
    .A2(_1884_),
    .Y(_1959_),
    .B1(_1861_));
 sg13g2_o21ai_1 _5063_ (.B1(_1878_),
    .Y(_1960_),
    .A1(_1871_),
    .A2(_1879_));
 sg13g2_o21ai_1 _5064_ (.B1(_1856_),
    .Y(_1961_),
    .A1(_1575_),
    .A2(_1854_));
 sg13g2_nand2_1 _5065_ (.Y(_1962_),
    .A(net747),
    .B(net702));
 sg13g2_nand2_1 _5066_ (.Y(_1963_),
    .A(net750),
    .B(net697));
 sg13g2_nand2_1 _5067_ (.Y(_1964_),
    .A(net749),
    .B(net700));
 sg13g2_xor2_1 _5068_ (.B(_1964_),
    .A(_1866_),
    .X(_1965_));
 sg13g2_nand2b_1 _5069_ (.Y(_1966_),
    .B(_1965_),
    .A_N(_1962_));
 sg13g2_xnor2_1 _5070_ (.Y(_1967_),
    .A(_1962_),
    .B(_1965_));
 sg13g2_inv_1 _5071_ (.Y(_1968_),
    .A(_1967_));
 sg13g2_o21ai_1 _5072_ (.B1(_1876_),
    .Y(_1969_),
    .A1(_1783_),
    .A2(_1874_));
 sg13g2_nand2_1 _5073_ (.Y(_1970_),
    .A(net755),
    .B(net693));
 sg13g2_nand2_1 _5074_ (.Y(_1971_),
    .A(net758),
    .B(net688));
 sg13g2_nor2_1 _5075_ (.A(_1874_),
    .B(_1971_),
    .Y(_1972_));
 sg13g2_or2_1 _5076_ (.X(_1973_),
    .B(_1971_),
    .A(_1874_));
 sg13g2_a22oi_1 _5077_ (.Y(_1974_),
    .B1(net688),
    .B2(net760),
    .A2(net690),
    .A1(net758));
 sg13g2_nor2_1 _5078_ (.A(_1972_),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_xnor2_1 _5079_ (.Y(_1976_),
    .A(_1970_),
    .B(_1975_));
 sg13g2_xnor2_1 _5080_ (.Y(_1977_),
    .A(_1969_),
    .B(_1976_));
 sg13g2_nor2_1 _5081_ (.A(_1968_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_xnor2_1 _5082_ (.Y(_1979_),
    .A(_1967_),
    .B(_1977_));
 sg13g2_xnor2_1 _5083_ (.Y(_1980_),
    .A(_1961_),
    .B(_1979_));
 sg13g2_nor2b_1 _5084_ (.A(_1980_),
    .B_N(_1960_),
    .Y(_1981_));
 sg13g2_xnor2_1 _5085_ (.Y(_1982_),
    .A(_1960_),
    .B(_1980_));
 sg13g2_nor2b_1 _5086_ (.A(net556),
    .B_N(_1671_),
    .Y(_1983_));
 sg13g2_xnor2_1 _5087_ (.Y(_1984_),
    .A(net556),
    .B(_1671_));
 sg13g2_nand2b_1 _5088_ (.Y(_1985_),
    .B(_1984_),
    .A_N(_1847_));
 sg13g2_xnor2_1 _5089_ (.Y(_1986_),
    .A(_1847_),
    .B(_1984_));
 sg13g2_o21ai_1 _5090_ (.B1(_1850_),
    .Y(_1987_),
    .A1(_1851_),
    .A2(_1852_));
 sg13g2_o21ai_1 _5091_ (.B1(net686),
    .Y(_1988_),
    .A1(net717),
    .A2(net714));
 sg13g2_nand2_1 _5092_ (.Y(_1989_),
    .A(net714),
    .B(_1761_));
 sg13g2_a21oi_1 _5093_ (.A1(net714),
    .A2(_1761_),
    .Y(_1990_),
    .B1(_1988_));
 sg13g2_nand2_1 _5094_ (.Y(_1991_),
    .A(net710),
    .B(net686));
 sg13g2_xnor2_1 _5095_ (.Y(_1992_),
    .A(_1990_),
    .B(_1991_));
 sg13g2_xnor2_1 _5096_ (.Y(_1993_),
    .A(_1672_),
    .B(_1992_));
 sg13g2_nor2b_1 _5097_ (.A(_1993_),
    .B_N(_1987_),
    .Y(_1994_));
 sg13g2_xnor2_1 _5098_ (.Y(_1995_),
    .A(_1987_),
    .B(_1993_));
 sg13g2_nand2_1 _5099_ (.Y(_1996_),
    .A(_1986_),
    .B(_1995_));
 sg13g2_xnor2_1 _5100_ (.Y(_1997_),
    .A(_1986_),
    .B(_1995_));
 sg13g2_nor2_1 _5101_ (.A(_1859_),
    .B(_1997_),
    .Y(_1998_));
 sg13g2_xor2_1 _5102_ (.B(_1997_),
    .A(_1859_),
    .X(_1999_));
 sg13g2_xor2_1 _5103_ (.B(_1999_),
    .A(_1982_),
    .X(_2000_));
 sg13g2_nand2b_1 _5104_ (.Y(_2001_),
    .B(_2000_),
    .A_N(_1959_));
 sg13g2_xnor2_1 _5105_ (.Y(_2002_),
    .A(_1959_),
    .B(_2000_));
 sg13g2_nand2b_1 _5106_ (.Y(_2003_),
    .B(_2002_),
    .A_N(_1958_));
 sg13g2_xnor2_1 _5107_ (.Y(_2004_),
    .A(_1958_),
    .B(_2002_));
 sg13g2_and2_1 _5108_ (.A(_1939_),
    .B(_2004_),
    .X(_2005_));
 sg13g2_xor2_1 _5109_ (.B(_2004_),
    .A(_1939_),
    .X(_2006_));
 sg13g2_xor2_1 _5110_ (.B(_2006_),
    .A(_1938_),
    .X(_2007_));
 sg13g2_nor2b_1 _5111_ (.A(_1933_),
    .B_N(_2007_),
    .Y(_2008_));
 sg13g2_xnor2_1 _5112_ (.Y(_2009_),
    .A(_1933_),
    .B(_2007_));
 sg13g2_xor2_1 _5113_ (.B(_2009_),
    .A(_1932_),
    .X(_2010_));
 sg13g2_and2_1 _5114_ (.A(_1931_),
    .B(_2010_),
    .X(_2011_));
 sg13g2_xnor2_1 _5115_ (.Y(_2012_),
    .A(_1931_),
    .B(_2010_));
 sg13g2_inv_1 _5116_ (.Y(_2013_),
    .A(_2012_));
 sg13g2_xnor2_1 _5117_ (.Y(_2014_),
    .A(_1930_),
    .B(_2013_));
 sg13g2_inv_1 _5118_ (.Y(_2015_),
    .A(_2014_));
 sg13g2_o21ai_1 _5119_ (.B1(net795),
    .Y(_2016_),
    .A1(net672),
    .A2(net234));
 sg13g2_a21oi_1 _5120_ (.A1(net672),
    .A2(_2014_),
    .Y(_0187_),
    .B1(_2016_));
 sg13g2_a21oi_1 _5121_ (.A1(_1930_),
    .A2(_2013_),
    .Y(_2017_),
    .B1(_2011_));
 sg13g2_a21oi_1 _5122_ (.A1(_1932_),
    .A2(_2009_),
    .Y(_2018_),
    .B1(_2008_));
 sg13g2_a21oi_1 _5123_ (.A1(_1938_),
    .A2(_2006_),
    .Y(_2019_),
    .B1(_2005_));
 sg13g2_nand2_1 _5124_ (.Y(_2020_),
    .A(_2001_),
    .B(_2003_));
 sg13g2_o21ai_1 _5125_ (.B1(_1956_),
    .Y(_2021_),
    .A1(_1940_),
    .A2(_1957_));
 sg13g2_xnor2_1 _5126_ (.Y(_2022_),
    .A(_2020_),
    .B(_2021_));
 sg13g2_a21oi_1 _5127_ (.A1(_1982_),
    .A2(_1999_),
    .Y(_2023_),
    .B1(_1998_));
 sg13g2_a21oi_1 _5128_ (.A1(_1969_),
    .A2(_1976_),
    .Y(_2024_),
    .B1(_1978_));
 sg13g2_a21oi_1 _5129_ (.A1(_1672_),
    .A2(_1992_),
    .Y(_2025_),
    .B1(_1994_));
 sg13g2_nand2_1 _5130_ (.Y(_2026_),
    .A(net751),
    .B(net693));
 sg13g2_nand2_1 _5131_ (.Y(_2027_),
    .A(net748),
    .B(net700));
 sg13g2_xor2_1 _5132_ (.B(_2027_),
    .A(_1963_),
    .X(_2028_));
 sg13g2_nand2_1 _5133_ (.Y(_2029_),
    .A(net755),
    .B(net690));
 sg13g2_xor2_1 _5134_ (.B(_2029_),
    .A(_1971_),
    .X(_2030_));
 sg13g2_xnor2_1 _5135_ (.Y(_2031_),
    .A(_2028_),
    .B(_2030_));
 sg13g2_xnor2_1 _5136_ (.Y(_2032_),
    .A(_2026_),
    .B(_2031_));
 sg13g2_o21ai_1 _5137_ (.B1(_1973_),
    .Y(_2033_),
    .A1(_1970_),
    .A2(_1974_));
 sg13g2_nand2_1 _5138_ (.Y(_2034_),
    .A(net746),
    .B(net702));
 sg13g2_xnor2_1 _5139_ (.Y(_2035_),
    .A(_2033_),
    .B(_2034_));
 sg13g2_xnor2_1 _5140_ (.Y(_2036_),
    .A(_2032_),
    .B(_2035_));
 sg13g2_xnor2_1 _5141_ (.Y(_2037_),
    .A(_2025_),
    .B(_2036_));
 sg13g2_xnor2_1 _5142_ (.Y(_2038_),
    .A(_2024_),
    .B(_2037_));
 sg13g2_nor2_1 _5143_ (.A(_1945_),
    .B(_1947_),
    .Y(_2039_));
 sg13g2_o21ai_1 _5144_ (.B1(_1966_),
    .Y(_2040_),
    .A1(_1866_),
    .A2(_1964_));
 sg13g2_a21oi_1 _5145_ (.A1(_1944_),
    .A2(_1949_),
    .Y(_2041_),
    .B1(_1951_));
 sg13g2_xor2_1 _5146_ (.B(net704),
    .A(net611),
    .X(_2042_));
 sg13g2_a21oi_1 _5147_ (.A1(net617),
    .A2(_2042_),
    .Y(_2043_),
    .B1(_2226_));
 sg13g2_o21ai_1 _5148_ (.B1(_2043_),
    .Y(_2044_),
    .A1(net617),
    .A2(_2042_));
 sg13g2_xnor2_1 _5149_ (.Y(_2045_),
    .A(_2040_),
    .B(_2044_));
 sg13g2_xnor2_1 _5150_ (.Y(_2046_),
    .A(_2039_),
    .B(_2045_));
 sg13g2_xnor2_1 _5151_ (.Y(_2047_),
    .A(_2041_),
    .B(_2046_));
 sg13g2_xnor2_1 _5152_ (.Y(_2048_),
    .A(_1893_),
    .B(_2047_));
 sg13g2_xnor2_1 _5153_ (.Y(_2049_),
    .A(_1644_),
    .B(_1935_));
 sg13g2_and2_1 _5154_ (.A(_1985_),
    .B(_1996_),
    .X(_2050_));
 sg13g2_xnor2_1 _5155_ (.Y(_2051_),
    .A(_1758_),
    .B(_1983_));
 sg13g2_o21ai_1 _5156_ (.B1(_1989_),
    .Y(_2052_),
    .A1(_1988_),
    .A2(_1991_));
 sg13g2_xor2_1 _5157_ (.B(net760),
    .A(net714),
    .X(_2053_));
 sg13g2_o21ai_1 _5158_ (.B1(net686),
    .Y(_2054_),
    .A1(net710),
    .A2(_2053_));
 sg13g2_a21oi_1 _5159_ (.A1(net710),
    .A2(_2053_),
    .Y(_2055_),
    .B1(_2054_));
 sg13g2_xor2_1 _5160_ (.B(_2055_),
    .A(_2052_),
    .X(_2056_));
 sg13g2_xnor2_1 _5161_ (.Y(_2057_),
    .A(_2051_),
    .B(_2056_));
 sg13g2_xnor2_1 _5162_ (.Y(_2058_),
    .A(_1500_),
    .B(_1763_));
 sg13g2_xnor2_1 _5163_ (.Y(_2059_),
    .A(_2057_),
    .B(_2058_));
 sg13g2_xnor2_1 _5164_ (.Y(_2060_),
    .A(_2050_),
    .B(_2059_));
 sg13g2_o21ai_1 _5165_ (.B1(_1953_),
    .Y(_2061_),
    .A1(_1893_),
    .A2(_1954_));
 sg13g2_a21oi_1 _5166_ (.A1(_1961_),
    .A2(_1979_),
    .Y(_2062_),
    .B1(_1981_));
 sg13g2_xnor2_1 _5167_ (.Y(_2063_),
    .A(_2048_),
    .B(_2062_));
 sg13g2_xnor2_1 _5168_ (.Y(_2064_),
    .A(_2038_),
    .B(_2060_));
 sg13g2_xnor2_1 _5169_ (.Y(_2065_),
    .A(_2061_),
    .B(_2064_));
 sg13g2_xnor2_1 _5170_ (.Y(_2066_),
    .A(_2023_),
    .B(_2063_));
 sg13g2_xnor2_1 _5171_ (.Y(_2067_),
    .A(_2065_),
    .B(_2066_));
 sg13g2_xnor2_1 _5172_ (.Y(_2068_),
    .A(_2049_),
    .B(_2067_));
 sg13g2_xnor2_1 _5173_ (.Y(_2069_),
    .A(_2022_),
    .B(_2068_));
 sg13g2_o21ai_1 _5174_ (.B1(_1936_),
    .Y(_2070_),
    .A1(_1645_),
    .A2(_1937_));
 sg13g2_xnor2_1 _5175_ (.Y(_2071_),
    .A(_2019_),
    .B(_2070_));
 sg13g2_xnor2_1 _5176_ (.Y(_2072_),
    .A(_2069_),
    .B(_2071_));
 sg13g2_xnor2_1 _5177_ (.Y(_2073_),
    .A(_2018_),
    .B(_2072_));
 sg13g2_xnor2_1 _5178_ (.Y(_2074_),
    .A(_2017_),
    .B(_2073_));
 sg13g2_o21ai_1 _5179_ (.B1(net795),
    .Y(_2075_),
    .A1(net265),
    .A2(net672));
 sg13g2_a21oi_1 _5180_ (.A1(net673),
    .A2(_2074_),
    .Y(_0188_),
    .B1(_2075_));
 sg13g2_nor2_1 _5181_ (.A(net670),
    .B(mac_en_clear),
    .Y(_2076_));
 sg13g2_nand2_2 _5182_ (.Y(_2077_),
    .A(net294),
    .B(_0895_));
 sg13g2_inv_1 _5183_ (.Y(_2078_),
    .A(_2077_));
 sg13g2_o21ai_1 _5184_ (.B1(net670),
    .Y(_2079_),
    .A1(net294),
    .A2(_0895_));
 sg13g2_inv_1 _5185_ (.Y(_2080_),
    .A(_2079_));
 sg13g2_a22oi_1 _5186_ (.Y(_2081_),
    .B1(_2077_),
    .B2(_2080_),
    .A2(net594),
    .A1(net294));
 sg13g2_nor2_1 _5187_ (.A(net772),
    .B(net295),
    .Y(_0189_));
 sg13g2_nor2b_1 _5188_ (.A(_0948_),
    .B_N(\mac_inst.accumulator[1] ),
    .Y(_2082_));
 sg13g2_nand2b_1 _5189_ (.Y(_2083_),
    .B(_0948_),
    .A_N(net252));
 sg13g2_nand2b_1 _5190_ (.Y(_2084_),
    .B(_2083_),
    .A_N(_2082_));
 sg13g2_o21ai_1 _5191_ (.B1(net670),
    .Y(_2085_),
    .A1(_2077_),
    .A2(_2084_));
 sg13g2_a21oi_1 _5192_ (.A1(_2077_),
    .A2(_2084_),
    .Y(_2086_),
    .B1(_2085_));
 sg13g2_a21oi_1 _5193_ (.A1(net252),
    .A2(net594),
    .Y(_2087_),
    .B1(_2086_));
 sg13g2_nor2_1 _5194_ (.A(net772),
    .B(net253),
    .Y(_0190_));
 sg13g2_a21oi_1 _5195_ (.A1(_2078_),
    .A2(_2083_),
    .Y(_2088_),
    .B1(_2082_));
 sg13g2_or2_1 _5196_ (.X(_2089_),
    .B(_1010_),
    .A(_2194_));
 sg13g2_xnor2_1 _5197_ (.Y(_2090_),
    .A(_2194_),
    .B(_1010_));
 sg13g2_o21ai_1 _5198_ (.B1(net670),
    .Y(_2091_),
    .A1(_2088_),
    .A2(_2090_));
 sg13g2_a21oi_1 _5199_ (.A1(_2088_),
    .A2(_2090_),
    .Y(_2092_),
    .B1(_2091_));
 sg13g2_a21oi_1 _5200_ (.A1(net202),
    .A2(net594),
    .Y(_2093_),
    .B1(_2092_));
 sg13g2_nor2_1 _5201_ (.A(net772),
    .B(net203),
    .Y(_0191_));
 sg13g2_nand2_1 _5202_ (.Y(_2094_),
    .A(net211),
    .B(net594));
 sg13g2_o21ai_1 _5203_ (.B1(_2089_),
    .Y(_2095_),
    .A1(_2088_),
    .A2(_2090_));
 sg13g2_and2_1 _5204_ (.A(\mac_inst.accumulator[3] ),
    .B(_1074_),
    .X(_2096_));
 sg13g2_xor2_1 _5205_ (.B(_1074_),
    .A(net211),
    .X(_2097_));
 sg13g2_a21oi_1 _5206_ (.A1(_2095_),
    .A2(_2097_),
    .Y(_2098_),
    .B1(_2217_));
 sg13g2_o21ai_1 _5207_ (.B1(_2098_),
    .Y(_2099_),
    .A1(_2095_),
    .A2(_2097_));
 sg13g2_a21oi_1 _5208_ (.A1(net212),
    .A2(_2099_),
    .Y(_0192_),
    .B1(net772));
 sg13g2_a21oi_1 _5209_ (.A1(_2095_),
    .A2(_2097_),
    .Y(_2100_),
    .B1(_2096_));
 sg13g2_or2_1 _5210_ (.X(_2101_),
    .B(_1141_),
    .A(_2193_));
 sg13g2_xnor2_1 _5211_ (.Y(_2102_),
    .A(_2193_),
    .B(_1141_));
 sg13g2_o21ai_1 _5212_ (.B1(net670),
    .Y(_2103_),
    .A1(_2100_),
    .A2(_2102_));
 sg13g2_a21oi_1 _5213_ (.A1(_2100_),
    .A2(_2102_),
    .Y(_2104_),
    .B1(_2103_));
 sg13g2_a21oi_1 _5214_ (.A1(net205),
    .A2(net594),
    .Y(_2105_),
    .B1(_2104_));
 sg13g2_nor2_1 _5215_ (.A(net772),
    .B(net206),
    .Y(_0193_));
 sg13g2_o21ai_1 _5216_ (.B1(_2101_),
    .Y(_2106_),
    .A1(_2100_),
    .A2(_2102_));
 sg13g2_and2_1 _5217_ (.A(\mac_inst.accumulator[5] ),
    .B(_1216_),
    .X(_2107_));
 sg13g2_xor2_1 _5218_ (.B(_1216_),
    .A(net288),
    .X(_2108_));
 sg13g2_o21ai_1 _5219_ (.B1(net670),
    .Y(_2109_),
    .A1(_2106_),
    .A2(_2108_));
 sg13g2_a21oi_1 _5220_ (.A1(_2106_),
    .A2(_2108_),
    .Y(_2110_),
    .B1(_2109_));
 sg13g2_a21oi_1 _5221_ (.A1(net288),
    .A2(net594),
    .Y(_2111_),
    .B1(_2110_));
 sg13g2_nor2_1 _5222_ (.A(net772),
    .B(net289),
    .Y(_0194_));
 sg13g2_a21oi_1 _5223_ (.A1(_2106_),
    .A2(_2108_),
    .Y(_2112_),
    .B1(_2107_));
 sg13g2_nand2_1 _5224_ (.Y(_2113_),
    .A(\mac_inst.accumulator[6] ),
    .B(_1309_));
 sg13g2_xnor2_1 _5225_ (.Y(_2114_),
    .A(net277),
    .B(_1309_));
 sg13g2_o21ai_1 _5226_ (.B1(net670),
    .Y(_2115_),
    .A1(_2112_),
    .A2(_2114_));
 sg13g2_a21oi_1 _5227_ (.A1(_2112_),
    .A2(_2114_),
    .Y(_2116_),
    .B1(_2115_));
 sg13g2_a21oi_1 _5228_ (.A1(net277),
    .A2(net594),
    .Y(_2117_),
    .B1(_2116_));
 sg13g2_nor2_1 _5229_ (.A(net771),
    .B(net278),
    .Y(_0195_));
 sg13g2_o21ai_1 _5230_ (.B1(_2113_),
    .Y(_2118_),
    .A1(_2112_),
    .A2(_2114_));
 sg13g2_nor2b_1 _5231_ (.A(_1392_),
    .B_N(net263),
    .Y(_2119_));
 sg13g2_xnor2_1 _5232_ (.Y(_2120_),
    .A(net263),
    .B(_1392_));
 sg13g2_o21ai_1 _5233_ (.B1(net671),
    .Y(_2121_),
    .A1(_2118_),
    .A2(_2120_));
 sg13g2_a21oi_1 _5234_ (.A1(_2118_),
    .A2(_2120_),
    .Y(_2122_),
    .B1(_2121_));
 sg13g2_a21oi_1 _5235_ (.A1(net263),
    .A2(net593),
    .Y(_2123_),
    .B1(_2122_));
 sg13g2_nor2_1 _5236_ (.A(net771),
    .B(net264),
    .Y(_0196_));
 sg13g2_a21oi_1 _5237_ (.A1(_2118_),
    .A2(_2120_),
    .Y(_2124_),
    .B1(_2119_));
 sg13g2_a21o_1 _5238_ (.A2(_2120_),
    .A1(_2118_),
    .B1(_2119_),
    .X(_2125_));
 sg13g2_and2_1 _5239_ (.A(\mac_inst.accumulator[8] ),
    .B(_1481_),
    .X(_2126_));
 sg13g2_xnor2_1 _5240_ (.Y(_2127_),
    .A(net316),
    .B(_1481_));
 sg13g2_nor2_1 _5241_ (.A(_2124_),
    .B(_2127_),
    .Y(_2128_));
 sg13g2_nand2_1 _5242_ (.Y(_2129_),
    .A(_2124_),
    .B(_2127_));
 sg13g2_nor2_1 _5243_ (.A(_2217_),
    .B(_2128_),
    .Y(_2130_));
 sg13g2_a22oi_1 _5244_ (.Y(_2131_),
    .B1(_2129_),
    .B2(_2130_),
    .A2(net593),
    .A1(net316));
 sg13g2_nor2_1 _5245_ (.A(net771),
    .B(_2131_),
    .Y(_0197_));
 sg13g2_nand2_1 _5246_ (.Y(_2132_),
    .A(net272),
    .B(net593));
 sg13g2_nor2_1 _5247_ (.A(_2126_),
    .B(_2128_),
    .Y(_2133_));
 sg13g2_nor2_1 _5248_ (.A(\mac_inst.accumulator[9] ),
    .B(_1570_),
    .Y(_2134_));
 sg13g2_xnor2_1 _5249_ (.Y(_2135_),
    .A(net272),
    .B(_1570_));
 sg13g2_a21oi_1 _5250_ (.A1(_2133_),
    .A2(_2135_),
    .Y(_2136_),
    .B1(_2217_));
 sg13g2_o21ai_1 _5251_ (.B1(_2136_),
    .Y(_2137_),
    .A1(_2133_),
    .A2(_2135_));
 sg13g2_a21oi_1 _5252_ (.A1(net273),
    .A2(_2137_),
    .Y(_0198_),
    .B1(net773));
 sg13g2_nand2_1 _5253_ (.Y(_2138_),
    .A(\mac_inst.accumulator[10] ),
    .B(_1663_));
 sg13g2_xnor2_1 _5254_ (.Y(_2139_),
    .A(\mac_inst.accumulator[10] ),
    .B(_1663_));
 sg13g2_or2_1 _5255_ (.X(_2140_),
    .B(_2135_),
    .A(_2127_));
 sg13g2_inv_1 _5256_ (.Y(_2141_),
    .A(_2140_));
 sg13g2_a21oi_1 _5257_ (.A1(\mac_inst.accumulator[9] ),
    .A2(_1570_),
    .Y(_2142_),
    .B1(_2126_));
 sg13g2_nor2_1 _5258_ (.A(_2134_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_a21oi_1 _5259_ (.A1(_2125_),
    .A2(_2141_),
    .Y(_2144_),
    .B1(_2143_));
 sg13g2_or2_1 _5260_ (.X(_2145_),
    .B(_2144_),
    .A(_2139_));
 sg13g2_a21oi_1 _5261_ (.A1(_2139_),
    .A2(_2144_),
    .Y(_2146_),
    .B1(_2217_));
 sg13g2_a22oi_1 _5262_ (.Y(_2147_),
    .B1(_2145_),
    .B2(_2146_),
    .A2(net593),
    .A1(net331));
 sg13g2_nor2_1 _5263_ (.A(net771),
    .B(_2147_),
    .Y(_0199_));
 sg13g2_and2_1 _5264_ (.A(_2138_),
    .B(_2145_),
    .X(_2148_));
 sg13g2_a21oi_1 _5265_ (.A1(_1747_),
    .A2(_1748_),
    .Y(_2149_),
    .B1(\mac_inst.accumulator[11] ));
 sg13g2_and3_1 _5266_ (.X(_2150_),
    .A(\mac_inst.accumulator[11] ),
    .B(_1747_),
    .C(_1748_));
 sg13g2_nand3_1 _5267_ (.B(_1747_),
    .C(_1748_),
    .A(\mac_inst.accumulator[11] ),
    .Y(_2151_));
 sg13g2_nand2b_1 _5268_ (.Y(_2152_),
    .B(_2151_),
    .A_N(_2149_));
 sg13g2_or2_1 _5269_ (.X(_2153_),
    .B(_2152_),
    .A(_2148_));
 sg13g2_a21oi_1 _5270_ (.A1(_2148_),
    .A2(_2152_),
    .Y(_2154_),
    .B1(_2217_));
 sg13g2_a22oi_1 _5271_ (.Y(_2155_),
    .B1(_2153_),
    .B2(_2154_),
    .A2(net593),
    .A1(net335));
 sg13g2_nor2_1 _5272_ (.A(net773),
    .B(_2155_),
    .Y(_0200_));
 sg13g2_nand2_1 _5273_ (.Y(_2156_),
    .A(net230),
    .B(net593));
 sg13g2_a21oi_1 _5274_ (.A1(_2138_),
    .A2(_2151_),
    .Y(_2157_),
    .B1(_2149_));
 sg13g2_nor3_1 _5275_ (.A(_2139_),
    .B(_2149_),
    .C(_2150_),
    .Y(_2158_));
 sg13g2_nor4_1 _5276_ (.A(_2139_),
    .B(_2140_),
    .C(_2149_),
    .D(_2150_),
    .Y(_2159_));
 sg13g2_a221oi_1 _5277_ (.B2(_2125_),
    .C1(_2157_),
    .B1(_2159_),
    .A1(_2143_),
    .Y(_2160_),
    .A2(_2158_));
 sg13g2_nor2_1 _5278_ (.A(_2192_),
    .B(_1839_),
    .Y(_2161_));
 sg13g2_xnor2_1 _5279_ (.Y(_2162_),
    .A(net230),
    .B(_1839_));
 sg13g2_inv_1 _5280_ (.Y(_2163_),
    .A(_2162_));
 sg13g2_nor2_1 _5281_ (.A(_2160_),
    .B(_2163_),
    .Y(_2164_));
 sg13g2_a21oi_1 _5282_ (.A1(_2160_),
    .A2(_2163_),
    .Y(_2165_),
    .B1(_2217_));
 sg13g2_nand2b_1 _5283_ (.Y(_2166_),
    .B(_2165_),
    .A_N(_2164_));
 sg13g2_a21oi_1 _5284_ (.A1(net231),
    .A2(_2166_),
    .Y(_0201_),
    .B1(net771));
 sg13g2_nor2_1 _5285_ (.A(_2191_),
    .B(_1928_),
    .Y(_2167_));
 sg13g2_nand2_1 _5286_ (.Y(_2168_),
    .A(_2191_),
    .B(_1928_));
 sg13g2_xnor2_1 _5287_ (.Y(_2169_),
    .A(_2191_),
    .B(_1928_));
 sg13g2_nor2_1 _5288_ (.A(_2161_),
    .B(_2164_),
    .Y(_2170_));
 sg13g2_or2_1 _5289_ (.X(_2171_),
    .B(_2170_),
    .A(_2169_));
 sg13g2_a21oi_1 _5290_ (.A1(_2169_),
    .A2(_2170_),
    .Y(_2172_),
    .B1(_2217_));
 sg13g2_a22oi_1 _5291_ (.Y(_2173_),
    .B1(_2171_),
    .B2(_2172_),
    .A2(net593),
    .A1(net279));
 sg13g2_nor2_1 _5292_ (.A(net771),
    .B(_2173_),
    .Y(_0202_));
 sg13g2_nand2_1 _5293_ (.Y(_2174_),
    .A(net242),
    .B(net593));
 sg13g2_nor3_1 _5294_ (.A(_2160_),
    .B(_2163_),
    .C(_2169_),
    .Y(_2175_));
 sg13g2_a21o_1 _5295_ (.A2(_2168_),
    .A1(_2161_),
    .B1(_2167_),
    .X(_2176_));
 sg13g2_nand2_1 _5296_ (.Y(_2177_),
    .A(\mac_inst.accumulator[14] ),
    .B(_2015_));
 sg13g2_xnor2_1 _5297_ (.Y(_2178_),
    .A(net242),
    .B(_2014_));
 sg13g2_o21ai_1 _5298_ (.B1(_2178_),
    .Y(_2179_),
    .A1(_2175_),
    .A2(_2176_));
 sg13g2_or3_1 _5299_ (.A(_2175_),
    .B(_2176_),
    .C(_2178_),
    .X(_2180_));
 sg13g2_nand3_1 _5300_ (.B(_2179_),
    .C(_2180_),
    .A(net671),
    .Y(_2181_));
 sg13g2_a21oi_1 _5301_ (.A1(net243),
    .A2(_2181_),
    .Y(_0203_),
    .B1(net771));
 sg13g2_nand2_1 _5302_ (.Y(_2182_),
    .A(net164),
    .B(_2076_));
 sg13g2_xor2_1 _5303_ (.B(_2074_),
    .A(net164),
    .X(_2183_));
 sg13g2_nand3_1 _5304_ (.B(_2179_),
    .C(_2183_),
    .A(_2177_),
    .Y(_2184_));
 sg13g2_a21oi_1 _5305_ (.A1(_2177_),
    .A2(_2179_),
    .Y(_2185_),
    .B1(_2183_));
 sg13g2_nand3b_1 _5306_ (.B(net671),
    .C(_2184_),
    .Y(_2186_),
    .A_N(_2185_));
 sg13g2_a21oi_1 _5307_ (.A1(net165),
    .A2(_2186_),
    .Y(_0204_),
    .B1(net771));
 sg13g2_o21ai_1 _5308_ (.B1(net794),
    .Y(_2187_),
    .A1(\mac_inst.RDY_get_multiply ),
    .A2(net672));
 sg13g2_nor2_1 _5309_ (.A(net129),
    .B(_2187_),
    .Y(_0205_));
 sg13g2_o21ai_1 _5310_ (.B1(net795),
    .Y(_2188_),
    .A1(\mac_inst.RDY_get_mac ),
    .A2(net671));
 sg13g2_nor2_1 _5311_ (.A(net131),
    .B(_2188_),
    .Y(_0206_));
 sg13g2_nor2_1 _5312_ (.A(_2308_),
    .B(_2366_),
    .Y(_0047_));
 sg13g2_dfrbpq_1 _5313_ (.RESET_B(net782),
    .D(net416),
    .Q(\byte_counter[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5314_ (.RESET_B(net782),
    .D(net413),
    .Q(\byte_counter[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5315_ (.RESET_B(net29),
    .D(_0012_),
    .Q(\cordic_inst.current_op[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5316_ (.RESET_B(net61),
    .D(_0013_),
    .Q(\cordic_inst.current_op[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5317_ (.RESET_B(net76),
    .D(_0014_),
    .Q(\cordic_inst.current_op[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5318_ (.RESET_B(net788),
    .D(_0021_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5319_ (.RESET_B(net785),
    .D(_0022_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5320_ (.RESET_B(net785),
    .D(_0023_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5321_ (.RESET_B(net785),
    .D(_0024_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5322_ (.RESET_B(net787),
    .D(_0025_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5323_ (.RESET_B(net787),
    .D(_0026_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5324_ (.RESET_B(net787),
    .D(_0027_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5325_ (.RESET_B(net785),
    .D(_0028_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5326_ (.RESET_B(net783),
    .D(net233),
    .Q(\result_reg[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5327_ (.RESET_B(net779),
    .D(net160),
    .Q(\result_reg[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5328_ (.RESET_B(net778),
    .D(net195),
    .Q(\result_reg[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5329_ (.RESET_B(net776),
    .D(net210),
    .Q(\result_reg[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5330_ (.RESET_B(net781),
    .D(net181),
    .Q(\result_reg[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5331_ (.RESET_B(net779),
    .D(net229),
    .Q(\result_reg[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5332_ (.RESET_B(net777),
    .D(net199),
    .Q(\result_reg[6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5333_ (.RESET_B(net782),
    .D(net175),
    .Q(\result_reg[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5334_ (.RESET_B(net781),
    .D(net216),
    .Q(\result_reg[8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5335_ (.RESET_B(net779),
    .D(net197),
    .Q(\result_reg[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5336_ (.RESET_B(net777),
    .D(_0041_),
    .Q(\result_reg[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5337_ (.RESET_B(net776),
    .D(net158),
    .Q(\result_reg[11] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5338_ (.RESET_B(net781),
    .D(net187),
    .Q(\result_reg[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5339_ (.RESET_B(net776),
    .D(net185),
    .Q(\result_reg[13] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5340_ (.RESET_B(net777),
    .D(net179),
    .Q(\result_reg[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5341_ (.RESET_B(net782),
    .D(net239),
    .Q(\result_reg[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5342_ (.RESET_B(net75),
    .D(_0047_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5343_ (.RESET_B(net74),
    .D(_0000_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5344_ (.RESET_B(net73),
    .D(_0051_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5345_ (.RESET_B(net72),
    .D(_0052_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5346_ (.RESET_B(net71),
    .D(_0053_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5347_ (.RESET_B(net70),
    .D(_0054_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5348_ (.RESET_B(net781),
    .D(_0055_),
    .Q(uo_out[0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5349_ (.RESET_B(net779),
    .D(_0056_),
    .Q(uo_out[1]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5350_ (.RESET_B(net777),
    .D(_0057_),
    .Q(uo_out[2]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _5351_ (.RESET_B(net779),
    .D(_0058_),
    .Q(uo_out[3]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5352_ (.RESET_B(net781),
    .D(_0059_),
    .Q(uo_out[4]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5353_ (.RESET_B(net779),
    .D(_0060_),
    .Q(uo_out[5]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5354_ (.RESET_B(net778),
    .D(_0061_),
    .Q(uo_out[6]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5355_ (.RESET_B(net782),
    .D(net301),
    .Q(uo_out[7]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5356_ (.RESET_B(net791),
    .D(net333),
    .Q(\state[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5357_ (.RESET_B(net791),
    .D(_0064_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5358_ (.RESET_B(net791),
    .D(_0065_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5359_ (.RESET_B(net790),
    .D(_0066_),
    .Q(\cmd_reg[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5360_ (.RESET_B(net790),
    .D(_0067_),
    .Q(\cmd_reg[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5361_ (.RESET_B(net794),
    .D(_0068_),
    .Q(\cmd_reg[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5362_ (.RESET_B(net790),
    .D(_0069_),
    .Q(\cmd_reg[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5363_ (.RESET_B(net794),
    .D(net259),
    .Q(\cmd_reg[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5364_ (.RESET_B(net795),
    .D(_0071_),
    .Q(\cmd_reg[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5365_ (.RESET_B(net794),
    .D(net177),
    .Q(\cmd_reg[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5366_ (.RESET_B(net790),
    .D(_0073_),
    .Q(\cmd_reg[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5367_ (.RESET_B(net786),
    .D(_0074_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5368_ (.RESET_B(net789),
    .D(_0075_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5369_ (.RESET_B(net789),
    .D(_0076_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5370_ (.RESET_B(net785),
    .D(_0077_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5371_ (.RESET_B(net787),
    .D(_0078_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5372_ (.RESET_B(net789),
    .D(_0079_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5373_ (.RESET_B(net789),
    .D(_0080_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _5374_ (.RESET_B(net786),
    .D(_0081_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5375_ (.RESET_B(net788),
    .D(_0082_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[31] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5376_ (.RESET_B(net788),
    .D(_0083_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5377_ (.RESET_B(net788),
    .D(_0084_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5378_ (.RESET_B(net786),
    .D(_0085_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5379_ (.RESET_B(net789),
    .D(_0086_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5380_ (.RESET_B(net789),
    .D(_0087_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5381_ (.RESET_B(net789),
    .D(_0088_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5382_ (.RESET_B(net785),
    .D(_0089_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5383_ (.RESET_B(net777),
    .D(net257),
    .Q(\result_reg[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5384_ (.RESET_B(net777),
    .D(net237),
    .Q(\result_reg[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5385_ (.RESET_B(net778),
    .D(net222),
    .Q(\result_reg[18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5386_ (.RESET_B(net776),
    .D(net183),
    .Q(\result_reg[19] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5387_ (.RESET_B(net780),
    .D(net214),
    .Q(\result_reg[20] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5388_ (.RESET_B(net779),
    .D(net173),
    .Q(\result_reg[21] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5389_ (.RESET_B(net777),
    .D(net241),
    .Q(\result_reg[22] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5390_ (.RESET_B(net781),
    .D(net189),
    .Q(\result_reg[23] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5391_ (.RESET_B(net781),
    .D(net149),
    .Q(\result_reg[24] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5392_ (.RESET_B(net780),
    .D(net191),
    .Q(\result_reg[25] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5393_ (.RESET_B(net778),
    .D(net193),
    .Q(\result_reg[26] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5394_ (.RESET_B(net776),
    .D(net227),
    .Q(\result_reg[27] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5395_ (.RESET_B(net780),
    .D(net163),
    .Q(\result_reg[28] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5396_ (.RESET_B(net779),
    .D(net208),
    .Q(\result_reg[29] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5397_ (.RESET_B(net777),
    .D(net201),
    .Q(\result_reg[30] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5398_ (.RESET_B(net782),
    .D(net171),
    .Q(\result_reg[31] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5399_ (.RESET_B(net791),
    .D(net9),
    .Q(wr_prev),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5400_ (.RESET_B(net781),
    .D(net10),
    .Q(rd_prev),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5401_ (.RESET_B(net792),
    .D(_0005_),
    .Q(cordic_en_sin_cos),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5402_ (.RESET_B(net792),
    .D(net137),
    .Q(cordic_en_atan2),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5403_ (.RESET_B(net792),
    .D(_0006_),
    .Q(cordic_en_sqrt),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5404_ (.RESET_B(net791),
    .D(_0003_),
    .Q(cordic_en_get_sin_cos),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5405_ (.RESET_B(net790),
    .D(_0002_),
    .Q(cordic_en_get_atan2),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5406_ (.RESET_B(net790),
    .D(_0004_),
    .Q(cordic_en_get_sqrt),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5407_ (.RESET_B(net790),
    .D(net134),
    .Q(mac_en_multiply),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5408_ (.RESET_B(net794),
    .D(_0009_),
    .Q(mac_en_get_multiply),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5409_ (.RESET_B(net794),
    .D(net140),
    .Q(mac_en_mac),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5410_ (.RESET_B(net794),
    .D(_0008_),
    .Q(mac_en_get_mac),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5411_ (.RESET_B(net794),
    .D(_0007_),
    .Q(mac_en_clear),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5412_ (.RESET_B(net69),
    .D(net305),
    .Q(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5413_ (.RESET_B(net67),
    .D(_0107_),
    .Q(cordic_busy),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5414_ (.RESET_B(net65),
    .D(_0108_),
    .Q(\cordic_inst.cordic_state[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5415_ (.RESET_B(net63),
    .D(_0109_),
    .Q(\cordic_inst.cordic_state[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5416_ (.RESET_B(net60),
    .D(_0110_),
    .Q(\cordic_inst.cordic_state[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5417_ (.RESET_B(net58),
    .D(_0111_),
    .Q(\cordic_inst.cordic_state[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5418_ (.RESET_B(net56),
    .D(_0112_),
    .Q(\cordic_inst.cordic_state[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5419_ (.RESET_B(net54),
    .D(_0113_),
    .Q(\cordic_atan2_result[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5420_ (.RESET_B(net52),
    .D(_0114_),
    .Q(\cordic_atan2_result[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5421_ (.RESET_B(net50),
    .D(_0115_),
    .Q(\cordic_atan2_result[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5422_ (.RESET_B(net48),
    .D(_0116_),
    .Q(\cordic_atan2_result[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5423_ (.RESET_B(net46),
    .D(_0117_),
    .Q(\cordic_atan2_result[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5424_ (.RESET_B(net45),
    .D(_0118_),
    .Q(\cordic_atan2_result[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5425_ (.RESET_B(net43),
    .D(_0119_),
    .Q(\cordic_atan2_result[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5426_ (.RESET_B(net41),
    .D(_0120_),
    .Q(\cordic_atan2_result[7] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5427_ (.RESET_B(net39),
    .D(_0121_),
    .Q(\cordic_atan2_result[8] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5428_ (.RESET_B(net38),
    .D(_0122_),
    .Q(\cordic_atan2_result[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5429_ (.RESET_B(net37),
    .D(net340),
    .Q(\cordic_atan2_result[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5430_ (.RESET_B(net36),
    .D(_0124_),
    .Q(\cordic_atan2_result[11] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5431_ (.RESET_B(net35),
    .D(_0125_),
    .Q(\cordic_atan2_result[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5432_ (.RESET_B(net34),
    .D(_0126_),
    .Q(\cordic_atan2_result[13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5433_ (.RESET_B(net33),
    .D(_0127_),
    .Q(\cordic_atan2_result[14] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5434_ (.RESET_B(net32),
    .D(_0128_),
    .Q(\cordic_atan2_result[15] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5435_ (.RESET_B(net31),
    .D(_0129_),
    .Q(\cordic_inst.cordic_state[23] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5436_ (.RESET_B(net28),
    .D(_0130_),
    .Q(\cordic_inst.cordic_state[24] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5437_ (.RESET_B(net128),
    .D(_0131_),
    .Q(\cordic_inst.cordic_state[25] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5438_ (.RESET_B(net126),
    .D(_0132_),
    .Q(\cordic_inst.cordic_state[26] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5439_ (.RESET_B(net124),
    .D(_0133_),
    .Q(\cordic_inst.cordic_state[27] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5440_ (.RESET_B(net122),
    .D(net360),
    .Q(\cordic_inst.cordic_state[28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5441_ (.RESET_B(net121),
    .D(net373),
    .Q(\cordic_inst.cordic_state[29] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5442_ (.RESET_B(net119),
    .D(_0136_),
    .Q(\cordic_inst.cordic_state[30] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _5443_ (.RESET_B(net117),
    .D(_0137_),
    .Q(\cordic_inst.cordic_state[31] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _5444_ (.RESET_B(net115),
    .D(_0138_),
    .Q(\cordic_inst.cordic_state[32] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5445_ (.RESET_B(net113),
    .D(_0139_),
    .Q(\cordic_inst.cordic_state[33] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _5446_ (.RESET_B(net111),
    .D(_0140_),
    .Q(\cordic_inst.cordic_state[34] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5447_ (.RESET_B(net109),
    .D(_0141_),
    .Q(\cordic_inst.cordic_state[35] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5448_ (.RESET_B(net107),
    .D(_0142_),
    .Q(\cordic_inst.cordic_state[36] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5449_ (.RESET_B(net105),
    .D(_0143_),
    .Q(\cordic_inst.cordic_state[37] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5450_ (.RESET_B(net103),
    .D(net346),
    .Q(\cordic_inst.cordic_state[38] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5451_ (.RESET_B(net101),
    .D(_0145_),
    .Q(\cordic_inst.cordic_state[39] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5452_ (.RESET_B(net99),
    .D(_0146_),
    .Q(\cordic_inst.cordic_state[40] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5453_ (.RESET_B(net97),
    .D(_0147_),
    .Q(\cordic_inst.cordic_state[41] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5454_ (.RESET_B(net95),
    .D(_0148_),
    .Q(\cordic_inst.cordic_state[42] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5455_ (.RESET_B(net93),
    .D(_0149_),
    .Q(\cordic_inst.cordic_state[43] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5456_ (.RESET_B(net91),
    .D(_0150_),
    .Q(\cordic_inst.cordic_state[44] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5457_ (.RESET_B(net89),
    .D(_0151_),
    .Q(\cordic_inst.cordic_state[45] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5458_ (.RESET_B(net87),
    .D(_0152_),
    .Q(\cordic_inst.cordic_state[46] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5459_ (.RESET_B(net85),
    .D(_0153_),
    .Q(\cordic_inst.cordic_state[47] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _5460_ (.RESET_B(net83),
    .D(_0154_),
    .Q(\cordic_inst.cordic_state[48] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _5461_ (.RESET_B(net81),
    .D(_0155_),
    .Q(\cordic_inst.cordic_state[49] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5462_ (.RESET_B(net79),
    .D(_0156_),
    .Q(\cordic_inst.cordic_state[50] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5463_ (.RESET_B(net77),
    .D(net350),
    .Q(\cordic_inst.cordic_state[51] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5464_ (.RESET_B(net66),
    .D(net357),
    .Q(\cordic_inst.cordic_state[52] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5465_ (.RESET_B(net62),
    .D(net354),
    .Q(\cordic_inst.cordic_state[53] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5466_ (.RESET_B(net57),
    .D(_0160_),
    .Q(\cordic_inst.cordic_state[54] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5467_ (.RESET_B(net53),
    .D(_0161_),
    .Q(\cordic_inst.operation_pending ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5468_ (.RESET_B(net49),
    .D(net169),
    .Q(\cordic_inst.result_ready ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5469_ (.RESET_B(net791),
    .D(_0018_),
    .Q(_0017_),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5470_ (.RESET_B(net790),
    .D(net251),
    .Q(\exec_phase[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5471_ (.RESET_B(net791),
    .D(_0016_),
    .Q(\exec_phase[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5472_ (.RESET_B(net42),
    .D(_0163_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5473_ (.RESET_B(net40),
    .D(_0164_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_6_TO_3_0_201_1_119_2_63_ETC__q3[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5474_ (.RESET_B(net786),
    .D(_0165_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[23] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5475_ (.RESET_B(net788),
    .D(_0166_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[24] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5476_ (.RESET_B(net788),
    .D(_0167_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[25] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5477_ (.RESET_B(net785),
    .D(_0168_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[26] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5478_ (.RESET_B(net787),
    .D(_0169_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[27] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5479_ (.RESET_B(net789),
    .D(_0170_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[28] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5480_ (.RESET_B(net788),
    .D(_0171_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[29] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5481_ (.RESET_B(net785),
    .D(_0172_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[30] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5482_ (.RESET_B(net30),
    .D(_0173_),
    .Q(\mac_inst.get_multiply[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5483_ (.RESET_B(net127),
    .D(net262),
    .Q(\mac_inst.get_multiply[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5484_ (.RESET_B(net123),
    .D(net220),
    .Q(\mac_inst.get_multiply[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5485_ (.RESET_B(net120),
    .D(_0176_),
    .Q(\mac_inst.get_multiply[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5486_ (.RESET_B(net116),
    .D(net225),
    .Q(\mac_inst.get_multiply[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5487_ (.RESET_B(net112),
    .D(_0178_),
    .Q(\mac_inst.get_multiply[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5488_ (.RESET_B(net108),
    .D(_0179_),
    .Q(\mac_inst.get_multiply[6] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5489_ (.RESET_B(net104),
    .D(net247),
    .Q(\mac_inst.get_multiply[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5490_ (.RESET_B(net100),
    .D(_0181_),
    .Q(\mac_inst.get_multiply[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5491_ (.RESET_B(net96),
    .D(_0182_),
    .Q(\mac_inst.get_multiply[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5492_ (.RESET_B(net92),
    .D(_0183_),
    .Q(\mac_inst.get_multiply[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5493_ (.RESET_B(net88),
    .D(_0184_),
    .Q(\mac_inst.get_multiply[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5494_ (.RESET_B(net84),
    .D(net249),
    .Q(\mac_inst.get_multiply[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5495_ (.RESET_B(net80),
    .D(net291),
    .Q(\mac_inst.get_multiply[13] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5496_ (.RESET_B(net68),
    .D(net235),
    .Q(\mac_inst.get_multiply[14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5497_ (.RESET_B(net59),
    .D(net266),
    .Q(\mac_inst.get_multiply[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5498_ (.RESET_B(net51),
    .D(_0189_),
    .Q(\mac_inst.accumulator[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5499_ (.RESET_B(net44),
    .D(_0190_),
    .Q(\mac_inst.accumulator[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5500_ (.RESET_B(net125),
    .D(_0191_),
    .Q(\mac_inst.accumulator[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5501_ (.RESET_B(net118),
    .D(_0192_),
    .Q(\mac_inst.accumulator[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5502_ (.RESET_B(net110),
    .D(_0193_),
    .Q(\mac_inst.accumulator[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5503_ (.RESET_B(net102),
    .D(_0194_),
    .Q(\mac_inst.accumulator[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5504_ (.RESET_B(net94),
    .D(_0195_),
    .Q(\mac_inst.accumulator[6] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _5505_ (.RESET_B(net86),
    .D(_0196_),
    .Q(\mac_inst.accumulator[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5506_ (.RESET_B(net78),
    .D(_0197_),
    .Q(\mac_inst.accumulator[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5507_ (.RESET_B(net55),
    .D(net274),
    .Q(\mac_inst.accumulator[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5508_ (.RESET_B(net27),
    .D(_0199_),
    .Q(\mac_inst.accumulator[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5509_ (.RESET_B(net114),
    .D(_0200_),
    .Q(\mac_inst.accumulator[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5510_ (.RESET_B(net98),
    .D(_0201_),
    .Q(\mac_inst.accumulator[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5511_ (.RESET_B(net82),
    .D(_0202_),
    .Q(\mac_inst.accumulator[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5512_ (.RESET_B(net47),
    .D(net244),
    .Q(\mac_inst.accumulator[14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5513_ (.RESET_B(net106),
    .D(net166),
    .Q(\mac_inst.accumulator[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5514_ (.RESET_B(net64),
    .D(net130),
    .Q(\mac_inst.RDY_get_multiply ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5515_ (.RESET_B(net90),
    .D(net132),
    .Q(\mac_inst.RDY_get_mac ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_tiehi _5436__28 (.L_HI(net28));
 sg13g2_tiehi _5315__29 (.L_HI(net29));
 sg13g2_tiehi _5482__30 (.L_HI(net30));
 sg13g2_tiehi _5435__31 (.L_HI(net31));
 sg13g2_tiehi _5434__32 (.L_HI(net32));
 sg13g2_tiehi _5433__33 (.L_HI(net33));
 sg13g2_tiehi _5432__34 (.L_HI(net34));
 sg13g2_tiehi _5431__35 (.L_HI(net35));
 sg13g2_tiehi _5430__36 (.L_HI(net36));
 sg13g2_tiehi _5429__37 (.L_HI(net37));
 sg13g2_tiehi _5428__38 (.L_HI(net38));
 sg13g2_tiehi _5427__39 (.L_HI(net39));
 sg13g2_tiehi _5473__40 (.L_HI(net40));
 sg13g2_tiehi _5426__41 (.L_HI(net41));
 sg13g2_tiehi _5472__42 (.L_HI(net42));
 sg13g2_tiehi _5425__43 (.L_HI(net43));
 sg13g2_tiehi _5499__44 (.L_HI(net44));
 sg13g2_tiehi _5424__45 (.L_HI(net45));
 sg13g2_tiehi _5423__46 (.L_HI(net46));
 sg13g2_tiehi _5512__47 (.L_HI(net47));
 sg13g2_tiehi _5422__48 (.L_HI(net48));
 sg13g2_tiehi _5468__49 (.L_HI(net49));
 sg13g2_tiehi _5421__50 (.L_HI(net50));
 sg13g2_tiehi _5498__51 (.L_HI(net51));
 sg13g2_tiehi _5420__52 (.L_HI(net52));
 sg13g2_tiehi _5467__53 (.L_HI(net53));
 sg13g2_tiehi _5419__54 (.L_HI(net54));
 sg13g2_tiehi _5507__55 (.L_HI(net55));
 sg13g2_tiehi _5418__56 (.L_HI(net56));
 sg13g2_tiehi _5466__57 (.L_HI(net57));
 sg13g2_tiehi _5417__58 (.L_HI(net58));
 sg13g2_tiehi _5497__59 (.L_HI(net59));
 sg13g2_tiehi _5416__60 (.L_HI(net60));
 sg13g2_tiehi _5316__61 (.L_HI(net61));
 sg13g2_tiehi _5465__62 (.L_HI(net62));
 sg13g2_tiehi _5415__63 (.L_HI(net63));
 sg13g2_tiehi _5514__64 (.L_HI(net64));
 sg13g2_tiehi _5414__65 (.L_HI(net65));
 sg13g2_tiehi _5464__66 (.L_HI(net66));
 sg13g2_tiehi _5413__67 (.L_HI(net67));
 sg13g2_tiehi _5496__68 (.L_HI(net68));
 sg13g2_tiehi _5412__69 (.L_HI(net69));
 sg13g2_tiehi _5347__70 (.L_HI(net70));
 sg13g2_tiehi _5346__71 (.L_HI(net71));
 sg13g2_tiehi _5345__72 (.L_HI(net72));
 sg13g2_tiehi _5344__73 (.L_HI(net73));
 sg13g2_tiehi _5343__74 (.L_HI(net74));
 sg13g2_tiehi _5342__75 (.L_HI(net75));
 sg13g2_tiehi _5317__76 (.L_HI(net76));
 sg13g2_tiehi _5463__77 (.L_HI(net77));
 sg13g2_tiehi _5506__78 (.L_HI(net78));
 sg13g2_tiehi _5462__79 (.L_HI(net79));
 sg13g2_tiehi _5495__80 (.L_HI(net80));
 sg13g2_tiehi _5461__81 (.L_HI(net81));
 sg13g2_tiehi _5511__82 (.L_HI(net82));
 sg13g2_tiehi _5460__83 (.L_HI(net83));
 sg13g2_tiehi _5494__84 (.L_HI(net84));
 sg13g2_tiehi _5459__85 (.L_HI(net85));
 sg13g2_tiehi _5505__86 (.L_HI(net86));
 sg13g2_tiehi _5458__87 (.L_HI(net87));
 sg13g2_tiehi _5493__88 (.L_HI(net88));
 sg13g2_tiehi _5457__89 (.L_HI(net89));
 sg13g2_tiehi _5515__90 (.L_HI(net90));
 sg13g2_tiehi _5456__91 (.L_HI(net91));
 sg13g2_tiehi _5492__92 (.L_HI(net92));
 sg13g2_tiehi _5455__93 (.L_HI(net93));
 sg13g2_tiehi _5504__94 (.L_HI(net94));
 sg13g2_tiehi _5454__95 (.L_HI(net95));
 sg13g2_tiehi _5491__96 (.L_HI(net96));
 sg13g2_tiehi _5453__97 (.L_HI(net97));
 sg13g2_tiehi _5510__98 (.L_HI(net98));
 sg13g2_tiehi _5452__99 (.L_HI(net99));
 sg13g2_tiehi _5490__100 (.L_HI(net100));
 sg13g2_tiehi _5451__101 (.L_HI(net101));
 sg13g2_tiehi _5503__102 (.L_HI(net102));
 sg13g2_tiehi _5450__103 (.L_HI(net103));
 sg13g2_tiehi _5489__104 (.L_HI(net104));
 sg13g2_tiehi _5449__105 (.L_HI(net105));
 sg13g2_tiehi _5513__106 (.L_HI(net106));
 sg13g2_tiehi _5448__107 (.L_HI(net107));
 sg13g2_tiehi _5488__108 (.L_HI(net108));
 sg13g2_tiehi _5447__109 (.L_HI(net109));
 sg13g2_tiehi _5502__110 (.L_HI(net110));
 sg13g2_tiehi _5446__111 (.L_HI(net111));
 sg13g2_tiehi _5487__112 (.L_HI(net112));
 sg13g2_tiehi _5445__113 (.L_HI(net113));
 sg13g2_tiehi _5509__114 (.L_HI(net114));
 sg13g2_tiehi _5444__115 (.L_HI(net115));
 sg13g2_tiehi _5486__116 (.L_HI(net116));
 sg13g2_tiehi _5443__117 (.L_HI(net117));
 sg13g2_tiehi _5501__118 (.L_HI(net118));
 sg13g2_tiehi _5442__119 (.L_HI(net119));
 sg13g2_tiehi _5485__120 (.L_HI(net120));
 sg13g2_tiehi _5441__121 (.L_HI(net121));
 sg13g2_tiehi _5440__122 (.L_HI(net122));
 sg13g2_tiehi _5484__123 (.L_HI(net123));
 sg13g2_tiehi _5439__124 (.L_HI(net124));
 sg13g2_tiehi _5500__125 (.L_HI(net125));
 sg13g2_tiehi _5438__126 (.L_HI(net126));
 sg13g2_tiehi _5483__127 (.L_HI(net127));
 sg13g2_tiehi _5437__128 (.L_HI(net128));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_herald_12 (.L_LO(net12));
 sg13g2_tielo tt_um_herald_13 (.L_LO(net13));
 sg13g2_tielo tt_um_herald_14 (.L_LO(net14));
 sg13g2_tielo tt_um_herald_15 (.L_LO(net15));
 sg13g2_tielo tt_um_herald_16 (.L_LO(net16));
 sg13g2_tielo tt_um_herald_17 (.L_LO(net17));
 sg13g2_tielo tt_um_herald_18 (.L_LO(net18));
 sg13g2_tielo tt_um_herald_19 (.L_LO(net19));
 sg13g2_tielo tt_um_herald_20 (.L_LO(net20));
 sg13g2_tielo tt_um_herald_21 (.L_LO(net21));
 sg13g2_tielo tt_um_herald_22 (.L_LO(net22));
 sg13g2_tielo tt_um_herald_23 (.L_LO(net23));
 sg13g2_tielo tt_um_herald_24 (.L_LO(net24));
 sg13g2_tielo tt_um_herald_25 (.L_LO(net25));
 sg13g2_tielo tt_um_herald_26 (.L_LO(net26));
 sg13g2_tiehi _5508__27 (.L_HI(net27));
 sg13g2_buf_8 fanout542 (.A(net544),
    .X(net542));
 sg13g2_buf_1 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(_2566_),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(net547),
    .X(net545));
 sg13g2_buf_1 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(_2376_),
    .X(net547));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_8 fanout550 (.A(_2475_),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(_2466_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_2466_),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_8 fanout555 (.A(_2250_),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(_1405_),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(_2496_),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(net561),
    .X(net559));
 sg13g2_buf_1 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_8 fanout562 (.A(_2495_),
    .X(net562));
 sg13g2_buf_8 fanout563 (.A(net565),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(_2278_),
    .X(net565));
 sg13g2_buf_8 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(_2276_),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(_2273_),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(net573),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(net573),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_2248_),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(_0715_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_0715_),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(_2481_),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(_2472_),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(_2299_),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net583),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_2299_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(_2291_),
    .X(net584));
 sg13g2_buf_8 fanout585 (.A(_2300_),
    .X(net585));
 sg13g2_buf_1 fanout586 (.A(_2300_),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(_2300_),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(_2289_),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(_2289_),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(_2237_),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(_2076_),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(_0243_),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(_0243_),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(_0235_),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(_2283_),
    .X(net600));
 sg13g2_buf_8 fanout601 (.A(net603),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(_2280_),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(_2216_),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(_2211_),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(_2211_),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_2210_),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(_2195_),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(_2195_),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(net614),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_1 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(net375),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(net365),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net623),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(net621),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[28] ),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(net418),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(net628),
    .X(net626));
 sg13g2_buf_1 fanout627 (.A(net628),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[27] ),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(net632),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net409),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net635),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net414),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net639),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(net639),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net417),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net420),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(net133),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net645),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(net388),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(\cordic_inst.cordic_state[38] ),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net401),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(net404),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(net400),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net654),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(net397),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(\cordic_inst.cordic_state[5] ),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(\cordic_inst.cordic_state[4] ),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(\cordic_inst.cordic_state[4] ),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(net669),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_1 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(\cordic_inst.cordic_state[3] ),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(mac_en_mac),
    .X(net671));
 sg13g2_buf_8 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_8 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(mac_en_multiply),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(cordic_en_sqrt),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net680),
    .X(net677));
 sg13g2_buf_8 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(cordic_en_sqrt),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(cordic_en_atan2),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(cordic_en_sin_cos),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net369),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(net395),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(net396),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(net384),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net381),
    .X(net697));
 sg13g2_buf_8 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net386),
    .X(net700));
 sg13g2_buf_8 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(net366),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net707),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(net707),
    .X(net705));
 sg13g2_buf_1 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(net393),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(net710),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(net403),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(net715),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(net715),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(net419),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(net717),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(net398),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net722),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(net722),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net407),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net726),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(net411),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(net402),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(net731),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net736),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(net410),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_8 fanout739 (.A(net408),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(net135),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net298),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(net387),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(net385),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_8 fanout748 (.A(net377),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net399),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(net753),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net376),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(net370),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(net378),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net760));
 sg13g2_buf_1 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net394),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net764),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net412),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net415),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(_2215_),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(_2215_),
    .X(net770));
 sg13g2_buf_8 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(_2215_),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(net798),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net798),
    .X(net775));
 sg13g2_buf_8 fanout776 (.A(net784),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net780),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net780),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net784),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net783),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net798),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net786),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net797),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net797),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net797),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net797),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net796),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(rst_n),
    .X(net798));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_tielo tt_um_herald_11 (.L_LO(net11));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_0_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_9_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_17_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(mac_en_get_multiply),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0205_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold3 (.A(mac_en_get_mac),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0206_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0017_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0011_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cmd_reg[0] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold8 (.A(_2249_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0001_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cmd_reg[3] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold11 (.A(_2241_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0010_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac_inst.get_multiply[3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac_inst.get_multiply[0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cordic_inst.operation_pending ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0713_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mac_inst.get_multiply[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mac_inst.get_multiply[8] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold19 (.A(\result_reg[24] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold20 (.A(_2476_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0098_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac_inst.get_multiply[10] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac_inst.get_multiply[6] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cordic_inst.current_op[2] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold25 (.A(_2286_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mac_inst.get_multiply[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cordic_inst.current_op[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold28 (.A(_2315_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold29 (.A(\result_reg[11] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0042_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold31 (.A(\result_reg[1] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0032_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold33 (.A(\result_reg[28] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold34 (.A(_2477_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0102_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac_inst.accumulator[15] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2182_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0204_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold39 (.A(cordic_en_get_sin_cos),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0714_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0162_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold42 (.A(\result_reg[31] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0105_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold44 (.A(\result_reg[21] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0095_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold46 (.A(\result_reg[7] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0038_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cmd_reg[6] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0072_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold50 (.A(\result_reg[14] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0045_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold52 (.A(\result_reg[4] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0035_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold54 (.A(\result_reg[19] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0093_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold56 (.A(\result_reg[13] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0044_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold58 (.A(\result_reg[12] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0043_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold60 (.A(\result_reg[23] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0097_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold62 (.A(\result_reg[25] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0099_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold64 (.A(\result_reg[26] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0100_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold66 (.A(\result_reg[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0033_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold68 (.A(\result_reg[9] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0040_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold70 (.A(\result_reg[6] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0037_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold72 (.A(\result_reg[30] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0104_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mac_inst.accumulator[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold75 (.A(_2093_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold76 (.A(\result_reg[10] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mac_inst.accumulator[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold78 (.A(_2105_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold79 (.A(\result_reg[29] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0103_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold81 (.A(\result_reg[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0034_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mac_inst.accumulator[3] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold84 (.A(_2094_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold85 (.A(\result_reg[20] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0094_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold87 (.A(\result_reg[8] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0039_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cmd_reg[7] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mac_inst.get_multiply[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold91 (.A(_1011_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0175_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold93 (.A(\result_reg[18] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0092_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac_inst.get_multiply[4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold96 (.A(_1142_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0177_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold98 (.A(\result_reg[27] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0101_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold100 (.A(\result_reg[5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0036_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac_inst.accumulator[12] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold103 (.A(_2156_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold104 (.A(\result_reg[0] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0031_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mac_inst.get_multiply[14] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0187_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold108 (.A(\result_reg[17] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0091_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold110 (.A(\result_reg[15] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0046_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold112 (.A(\result_reg[22] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0096_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mac_inst.accumulator[14] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold115 (.A(_2174_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0203_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac_inst.get_multiply[7] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold118 (.A(_1393_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0180_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac_inst.get_multiply[12] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0185_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold122 (.A(\exec_phase[1] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0015_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mac_inst.accumulator[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold125 (.A(_2087_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold126 (.A(\exec_phase[2] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold127 (.A(_2321_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold128 (.A(\result_reg[16] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0090_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cmd_reg[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0070_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac_inst.get_multiply[1] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0949_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0174_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac_inst.accumulator[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold136 (.A(_2123_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mac_inst.get_multiply[15] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0188_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold139 (.A(uo_out[3]),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold140 (.A(_2440_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold141 (.A(uo_out[0]),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold142 (.A(_2434_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cmd_reg[5] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mac_inst.accumulator[9] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold145 (.A(_2132_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0198_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold147 (.A(uo_out[4]),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2442_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mac_inst.accumulator[6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold150 (.A(_2117_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac_inst.accumulator[13] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold152 (.A(uo_out[2]),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold153 (.A(_2438_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold154 (.A(uo_out[1]),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold155 (.A(_2436_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold156 (.A(uo_out[5]),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold157 (.A(_2444_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mac_inst.get_multiply[11] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold159 (.A(_1750_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac_inst.accumulator[5] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2111_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mac_inst.get_multiply[13] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0186_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cordic_atan2_result[9] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold165 (.A(_2581_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mac_inst.accumulator[0] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold167 (.A(_2081_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cordic_inst.cordic_state[0] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold169 (.A(_2480_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold170 (.A(\state[2] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold171 (.A(uo_out[7]),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold172 (.A(_2452_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0062_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cordic_atan2_result[1] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold175 (.A(_2505_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0106_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cordic_atan2_result[11] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold179 (.A(_2595_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cordic_atan2_result[7] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cordic_atan2_result[3] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cordic_inst.current_op[0] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold183 (.A(_2319_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold184 (.A(uo_out[6]),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold185 (.A(_2446_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cordic_inst.cordic_state[41] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold187 (.A(wr_prev),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mac_inst.accumulator[8] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cmd_reg[1] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cordic_atan2_result[12] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold191 (.A(_2604_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cmd_reg[2] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cordic_atan2_result[14] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0221_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold195 (.A(\cordic_atan2_result[13] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0213_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cordic_inst.cordic_state[40] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cordic_atan2_result[5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cordic_atan2_result[6] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cordic_atan2_result[0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2485_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cordic_atan2_result[2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac_inst.accumulator[10] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold204 (.A(\state[0] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0063_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cordic_atan2_result[4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mac_inst.accumulator[11] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cordic_inst.cordic_state[42] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold209 (.A(\cordic_atan2_result[8] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold210 (.A(_2574_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cordic_atan2_result[10] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0123_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold213 (.A(\cordic_inst.cordic_state[45] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cordic_atan2_result[15] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0228_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold216 (.A(\state[1] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold217 (.A(\cordic_inst.cordic_state[38] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0144_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cordic_inst.cordic_state[43] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cordic_inst.cordic_state[39] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cordic_inst.cordic_state[51] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0157_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cordic_inst.cordic_state[46] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0619_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cordic_inst.cordic_state[53] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0159_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cordic_inst.cordic_state[23] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold228 (.A(\cordic_inst.cordic_state[52] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0158_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold230 (.A(\cordic_inst.cordic_state[44] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cordic_inst.cordic_state[28] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0134_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cordic_inst.cordic_state[48] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0643_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold235 (.A(\cordic_inst.cordic_state[26] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cordic_inst.cordic_state[24] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold237 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[29] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cordic_inst.cordic_state[50] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0665_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cordic_inst.cordic_state[36] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cordic_inst.cordic_state[29] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0135_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cordic_inst.cordic_state[47] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold247 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[30] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold248 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold251 (.A(\state[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold252 (.A(_2261_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold254 (.A(cordic_busy),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cordic_inst.cordic_state[30] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold257 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cordic_inst.cordic_state[54] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold261 (.A(\cordic_inst.cordic_state[37] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cordic_inst.cordic_state[49] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cordic_inst.cordic_state[27] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold264 (.A(\cordic_inst.cordic_state[25] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[31] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold267 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold269 (.A(\cordic_inst.cordic_state[6] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold271 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cordic_inst.cordic_state[32] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold273 (.A(\cordic_inst.cordic_state[34] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold275 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cordic_inst.cordic_state[33] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold277 (.A(\cordic_inst.cordic_state[35] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cordic_inst.cordic_state[31] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold279 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold281 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[26] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold284 (.A(\byte_counter[1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0020_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold286 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[25] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold287 (.A(\byte_counter[0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0019_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[24] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[27] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[23] ),
    .X(net420));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_4 FILLER_24_581 ();
 sg13g2_fill_1 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_591 ();
 sg13g2_fill_1 FILLER_24_598 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_4 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_506 ();
 sg13g2_decap_8 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_531 ();
 sg13g2_decap_8 FILLER_25_538 ();
 sg13g2_decap_8 FILLER_25_545 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_4 FILLER_25_559 ();
 sg13g2_decap_4 FILLER_25_574 ();
 sg13g2_fill_2 FILLER_25_586 ();
 sg13g2_fill_2 FILLER_25_600 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_fill_1 FILLER_25_629 ();
 sg13g2_fill_2 FILLER_25_638 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_657 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_685 ();
 sg13g2_decap_8 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_8 FILLER_25_706 ();
 sg13g2_decap_8 FILLER_25_713 ();
 sg13g2_decap_8 FILLER_25_720 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_decap_8 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_decap_8 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_762 ();
 sg13g2_decap_8 FILLER_25_769 ();
 sg13g2_decap_8 FILLER_25_776 ();
 sg13g2_decap_8 FILLER_25_783 ();
 sg13g2_decap_8 FILLER_25_790 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_decap_8 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_846 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_4 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_457 ();
 sg13g2_decap_8 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_471 ();
 sg13g2_fill_1 FILLER_26_473 ();
 sg13g2_decap_8 FILLER_26_484 ();
 sg13g2_fill_2 FILLER_26_491 ();
 sg13g2_decap_4 FILLER_26_530 ();
 sg13g2_fill_2 FILLER_26_534 ();
 sg13g2_decap_4 FILLER_26_549 ();
 sg13g2_fill_1 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_578 ();
 sg13g2_decap_8 FILLER_26_585 ();
 sg13g2_decap_4 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_596 ();
 sg13g2_decap_8 FILLER_26_618 ();
 sg13g2_decap_4 FILLER_26_625 ();
 sg13g2_fill_2 FILLER_26_629 ();
 sg13g2_fill_2 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_666 ();
 sg13g2_decap_8 FILLER_26_673 ();
 sg13g2_fill_2 FILLER_26_680 ();
 sg13g2_fill_1 FILLER_26_682 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_fill_2 FILLER_27_441 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_fill_2 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_472 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_4 FILLER_27_511 ();
 sg13g2_fill_2 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_551 ();
 sg13g2_decap_4 FILLER_27_558 ();
 sg13g2_fill_2 FILLER_27_562 ();
 sg13g2_fill_2 FILLER_27_569 ();
 sg13g2_decap_8 FILLER_27_587 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_4 FILLER_27_619 ();
 sg13g2_fill_2 FILLER_27_623 ();
 sg13g2_fill_2 FILLER_27_633 ();
 sg13g2_fill_1 FILLER_27_635 ();
 sg13g2_decap_8 FILLER_27_645 ();
 sg13g2_fill_2 FILLER_27_652 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_fill_2 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_696 ();
 sg13g2_decap_8 FILLER_27_703 ();
 sg13g2_fill_1 FILLER_27_710 ();
 sg13g2_fill_2 FILLER_27_715 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_decap_8 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_738 ();
 sg13g2_decap_8 FILLER_27_745 ();
 sg13g2_decap_8 FILLER_27_752 ();
 sg13g2_decap_8 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_766 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_decap_8 FILLER_27_780 ();
 sg13g2_decap_8 FILLER_27_787 ();
 sg13g2_decap_8 FILLER_27_794 ();
 sg13g2_decap_8 FILLER_27_801 ();
 sg13g2_decap_8 FILLER_27_808 ();
 sg13g2_decap_8 FILLER_27_815 ();
 sg13g2_decap_8 FILLER_27_822 ();
 sg13g2_decap_8 FILLER_27_829 ();
 sg13g2_decap_8 FILLER_27_836 ();
 sg13g2_decap_8 FILLER_27_843 ();
 sg13g2_decap_8 FILLER_27_850 ();
 sg13g2_decap_4 FILLER_27_857 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_4 FILLER_28_410 ();
 sg13g2_fill_2 FILLER_28_414 ();
 sg13g2_fill_2 FILLER_28_420 ();
 sg13g2_fill_1 FILLER_28_422 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_fill_2 FILLER_28_441 ();
 sg13g2_decap_4 FILLER_28_461 ();
 sg13g2_fill_2 FILLER_28_478 ();
 sg13g2_fill_1 FILLER_28_480 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_fill_1 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_fill_1 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_4 FILLER_28_533 ();
 sg13g2_fill_2 FILLER_28_545 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_decap_4 FILLER_28_554 ();
 sg13g2_fill_1 FILLER_28_558 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_4 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_621 ();
 sg13g2_fill_2 FILLER_28_625 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_fill_2 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_fill_2 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_29_409 ();
 sg13g2_decap_8 FILLER_29_436 ();
 sg13g2_decap_4 FILLER_29_443 ();
 sg13g2_fill_2 FILLER_29_447 ();
 sg13g2_decap_4 FILLER_29_457 ();
 sg13g2_fill_1 FILLER_29_461 ();
 sg13g2_fill_1 FILLER_29_467 ();
 sg13g2_decap_8 FILLER_29_485 ();
 sg13g2_fill_1 FILLER_29_492 ();
 sg13g2_fill_1 FILLER_29_512 ();
 sg13g2_fill_2 FILLER_29_540 ();
 sg13g2_decap_4 FILLER_29_577 ();
 sg13g2_fill_1 FILLER_29_581 ();
 sg13g2_fill_2 FILLER_29_598 ();
 sg13g2_decap_4 FILLER_29_613 ();
 sg13g2_fill_2 FILLER_29_637 ();
 sg13g2_fill_2 FILLER_29_652 ();
 sg13g2_fill_1 FILLER_29_654 ();
 sg13g2_decap_4 FILLER_29_684 ();
 sg13g2_fill_1 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_fill_2 FILLER_29_709 ();
 sg13g2_fill_1 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_4 FILLER_29_741 ();
 sg13g2_fill_1 FILLER_29_745 ();
 sg13g2_fill_2 FILLER_29_759 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_fill_1 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_801 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_4 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_400 ();
 sg13g2_fill_1 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_415 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_2 FILLER_30_429 ();
 sg13g2_decap_4 FILLER_30_468 ();
 sg13g2_decap_4 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_504 ();
 sg13g2_fill_1 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_512 ();
 sg13g2_fill_1 FILLER_30_519 ();
 sg13g2_decap_8 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_fill_2 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_4 FILLER_30_581 ();
 sg13g2_fill_2 FILLER_30_585 ();
 sg13g2_decap_8 FILLER_30_607 ();
 sg13g2_decap_8 FILLER_30_614 ();
 sg13g2_decap_8 FILLER_30_621 ();
 sg13g2_decap_4 FILLER_30_633 ();
 sg13g2_fill_2 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_4 FILLER_30_658 ();
 sg13g2_fill_2 FILLER_30_662 ();
 sg13g2_fill_2 FILLER_30_669 ();
 sg13g2_decap_4 FILLER_30_675 ();
 sg13g2_fill_2 FILLER_30_679 ();
 sg13g2_fill_1 FILLER_30_712 ();
 sg13g2_fill_2 FILLER_30_726 ();
 sg13g2_fill_1 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_741 ();
 sg13g2_decap_4 FILLER_30_748 ();
 sg13g2_fill_2 FILLER_30_752 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_fill_2 FILLER_30_767 ();
 sg13g2_fill_2 FILLER_30_786 ();
 sg13g2_fill_1 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_820 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_decap_8 FILLER_30_834 ();
 sg13g2_decap_8 FILLER_30_841 ();
 sg13g2_decap_8 FILLER_30_848 ();
 sg13g2_decap_8 FILLER_30_855 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_decap_4 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_fill_2 FILLER_31_423 ();
 sg13g2_fill_2 FILLER_31_433 ();
 sg13g2_decap_8 FILLER_31_444 ();
 sg13g2_decap_8 FILLER_31_451 ();
 sg13g2_decap_8 FILLER_31_458 ();
 sg13g2_decap_4 FILLER_31_465 ();
 sg13g2_fill_2 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_501 ();
 sg13g2_decap_8 FILLER_31_515 ();
 sg13g2_fill_2 FILLER_31_522 ();
 sg13g2_fill_1 FILLER_31_524 ();
 sg13g2_decap_4 FILLER_31_538 ();
 sg13g2_fill_1 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_579 ();
 sg13g2_decap_4 FILLER_31_586 ();
 sg13g2_fill_1 FILLER_31_590 ();
 sg13g2_fill_2 FILLER_31_596 ();
 sg13g2_fill_1 FILLER_31_598 ();
 sg13g2_decap_8 FILLER_31_612 ();
 sg13g2_fill_1 FILLER_31_619 ();
 sg13g2_decap_8 FILLER_31_629 ();
 sg13g2_fill_2 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_decap_4 FILLER_31_692 ();
 sg13g2_fill_1 FILLER_31_696 ();
 sg13g2_decap_8 FILLER_31_702 ();
 sg13g2_decap_8 FILLER_31_709 ();
 sg13g2_decap_8 FILLER_31_716 ();
 sg13g2_fill_1 FILLER_31_723 ();
 sg13g2_fill_1 FILLER_31_731 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_790 ();
 sg13g2_fill_1 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_fill_2 FILLER_31_809 ();
 sg13g2_fill_2 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_396 ();
 sg13g2_fill_1 FILLER_32_400 ();
 sg13g2_fill_1 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_32_436 ();
 sg13g2_decap_8 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_450 ();
 sg13g2_fill_1 FILLER_32_472 ();
 sg13g2_fill_2 FILLER_32_478 ();
 sg13g2_fill_1 FILLER_32_480 ();
 sg13g2_decap_8 FILLER_32_486 ();
 sg13g2_decap_4 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_497 ();
 sg13g2_fill_1 FILLER_32_507 ();
 sg13g2_decap_8 FILLER_32_513 ();
 sg13g2_decap_4 FILLER_32_520 ();
 sg13g2_fill_1 FILLER_32_524 ();
 sg13g2_decap_8 FILLER_32_538 ();
 sg13g2_decap_8 FILLER_32_545 ();
 sg13g2_fill_1 FILLER_32_552 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_fill_1 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_608 ();
 sg13g2_fill_2 FILLER_32_615 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_decap_8 FILLER_32_635 ();
 sg13g2_decap_8 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_fill_1 FILLER_32_680 ();
 sg13g2_decap_4 FILLER_32_693 ();
 sg13g2_decap_4 FILLER_32_714 ();
 sg13g2_fill_1 FILLER_32_730 ();
 sg13g2_decap_4 FILLER_32_743 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_fill_2 FILLER_32_752 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_fill_1 FILLER_32_777 ();
 sg13g2_fill_2 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_784 ();
 sg13g2_fill_1 FILLER_32_794 ();
 sg13g2_fill_2 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_842 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_4 FILLER_32_856 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_293 ();
 sg13g2_decap_4 FILLER_33_300 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_383 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_438 ();
 sg13g2_decap_8 FILLER_33_460 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_524 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_decap_8 FILLER_33_555 ();
 sg13g2_decap_8 FILLER_33_577 ();
 sg13g2_fill_1 FILLER_33_584 ();
 sg13g2_decap_4 FILLER_33_610 ();
 sg13g2_fill_1 FILLER_33_614 ();
 sg13g2_decap_8 FILLER_33_638 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_647 ();
 sg13g2_decap_8 FILLER_33_656 ();
 sg13g2_decap_8 FILLER_33_663 ();
 sg13g2_fill_2 FILLER_33_678 ();
 sg13g2_fill_1 FILLER_33_680 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_4 FILLER_33_706 ();
 sg13g2_fill_1 FILLER_33_710 ();
 sg13g2_fill_1 FILLER_33_715 ();
 sg13g2_fill_2 FILLER_33_724 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_fill_1 FILLER_33_758 ();
 sg13g2_fill_1 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_fill_2 FILLER_33_816 ();
 sg13g2_fill_1 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_419 ();
 sg13g2_decap_4 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_438 ();
 sg13g2_fill_1 FILLER_34_450 ();
 sg13g2_fill_1 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_fill_1 FILLER_34_488 ();
 sg13g2_decap_4 FILLER_34_528 ();
 sg13g2_fill_2 FILLER_34_532 ();
 sg13g2_fill_2 FILLER_34_541 ();
 sg13g2_decap_8 FILLER_34_548 ();
 sg13g2_decap_8 FILLER_34_555 ();
 sg13g2_decap_4 FILLER_34_562 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_fill_2 FILLER_34_573 ();
 sg13g2_fill_1 FILLER_34_575 ();
 sg13g2_fill_2 FILLER_34_598 ();
 sg13g2_decap_8 FILLER_34_605 ();
 sg13g2_fill_2 FILLER_34_612 ();
 sg13g2_decap_4 FILLER_34_635 ();
 sg13g2_fill_1 FILLER_34_657 ();
 sg13g2_decap_8 FILLER_34_678 ();
 sg13g2_decap_4 FILLER_34_685 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_decap_8 FILLER_34_737 ();
 sg13g2_fill_1 FILLER_34_744 ();
 sg13g2_decap_4 FILLER_34_749 ();
 sg13g2_fill_2 FILLER_34_753 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_4 FILLER_34_786 ();
 sg13g2_fill_2 FILLER_34_790 ();
 sg13g2_fill_1 FILLER_34_798 ();
 sg13g2_fill_2 FILLER_34_814 ();
 sg13g2_fill_1 FILLER_34_816 ();
 sg13g2_fill_2 FILLER_34_829 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_fill_2 FILLER_35_462 ();
 sg13g2_decap_4 FILLER_35_474 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_fill_2 FILLER_35_504 ();
 sg13g2_fill_1 FILLER_35_514 ();
 sg13g2_decap_8 FILLER_35_527 ();
 sg13g2_fill_2 FILLER_35_558 ();
 sg13g2_fill_1 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_decap_8 FILLER_35_598 ();
 sg13g2_decap_8 FILLER_35_605 ();
 sg13g2_decap_4 FILLER_35_633 ();
 sg13g2_fill_1 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_fill_2 FILLER_35_694 ();
 sg13g2_fill_1 FILLER_35_696 ();
 sg13g2_decap_8 FILLER_35_702 ();
 sg13g2_decap_8 FILLER_35_709 ();
 sg13g2_decap_8 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_723 ();
 sg13g2_fill_2 FILLER_35_730 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_4 FILLER_35_764 ();
 sg13g2_decap_4 FILLER_35_776 ();
 sg13g2_fill_2 FILLER_35_780 ();
 sg13g2_decap_4 FILLER_35_790 ();
 sg13g2_fill_1 FILLER_35_794 ();
 sg13g2_fill_2 FILLER_35_801 ();
 sg13g2_fill_1 FILLER_35_803 ();
 sg13g2_decap_4 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_4 FILLER_35_857 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_8 FILLER_36_404 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_36_430 ();
 sg13g2_decap_8 FILLER_36_444 ();
 sg13g2_decap_4 FILLER_36_451 ();
 sg13g2_decap_8 FILLER_36_470 ();
 sg13g2_decap_4 FILLER_36_477 ();
 sg13g2_fill_2 FILLER_36_499 ();
 sg13g2_decap_8 FILLER_36_505 ();
 sg13g2_decap_4 FILLER_36_512 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_4 FILLER_36_539 ();
 sg13g2_fill_2 FILLER_36_543 ();
 sg13g2_fill_2 FILLER_36_549 ();
 sg13g2_decap_8 FILLER_36_561 ();
 sg13g2_fill_1 FILLER_36_568 ();
 sg13g2_decap_8 FILLER_36_577 ();
 sg13g2_fill_2 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_601 ();
 sg13g2_decap_8 FILLER_36_608 ();
 sg13g2_fill_1 FILLER_36_615 ();
 sg13g2_fill_2 FILLER_36_634 ();
 sg13g2_fill_1 FILLER_36_640 ();
 sg13g2_decap_4 FILLER_36_653 ();
 sg13g2_fill_2 FILLER_36_657 ();
 sg13g2_decap_4 FILLER_36_684 ();
 sg13g2_fill_1 FILLER_36_706 ();
 sg13g2_decap_4 FILLER_36_717 ();
 sg13g2_fill_1 FILLER_36_721 ();
 sg13g2_fill_1 FILLER_36_725 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_749 ();
 sg13g2_decap_4 FILLER_36_754 ();
 sg13g2_fill_1 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_fill_1 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_4 FILLER_36_835 ();
 sg13g2_fill_2 FILLER_36_839 ();
 sg13g2_decap_8 FILLER_36_846 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_decap_4 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_decap_4 FILLER_37_310 ();
 sg13g2_decap_4 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_decap_4 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_fill_2 FILLER_37_376 ();
 sg13g2_fill_1 FILLER_37_378 ();
 sg13g2_decap_4 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_426 ();
 sg13g2_decap_4 FILLER_37_433 ();
 sg13g2_fill_2 FILLER_37_437 ();
 sg13g2_decap_4 FILLER_37_443 ();
 sg13g2_fill_2 FILLER_37_447 ();
 sg13g2_decap_4 FILLER_37_472 ();
 sg13g2_fill_2 FILLER_37_476 ();
 sg13g2_fill_2 FILLER_37_482 ();
 sg13g2_fill_1 FILLER_37_496 ();
 sg13g2_fill_1 FILLER_37_532 ();
 sg13g2_fill_2 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_568 ();
 sg13g2_decap_4 FILLER_37_601 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_decap_4 FILLER_37_625 ();
 sg13g2_fill_2 FILLER_37_640 ();
 sg13g2_decap_8 FILLER_37_649 ();
 sg13g2_decap_8 FILLER_37_656 ();
 sg13g2_decap_4 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_689 ();
 sg13g2_decap_8 FILLER_37_708 ();
 sg13g2_decap_8 FILLER_37_737 ();
 sg13g2_fill_2 FILLER_37_744 ();
 sg13g2_decap_8 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_766 ();
 sg13g2_fill_1 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_780 ();
 sg13g2_fill_1 FILLER_37_782 ();
 sg13g2_fill_1 FILLER_37_786 ();
 sg13g2_fill_1 FILLER_37_792 ();
 sg13g2_fill_2 FILLER_37_806 ();
 sg13g2_fill_1 FILLER_37_808 ();
 sg13g2_decap_4 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_73 ();
 sg13g2_decap_8 FILLER_38_80 ();
 sg13g2_decap_4 FILLER_38_87 ();
 sg13g2_fill_1 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_131 ();
 sg13g2_fill_2 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_4 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_4 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_409 ();
 sg13g2_fill_2 FILLER_38_423 ();
 sg13g2_decap_8 FILLER_38_439 ();
 sg13g2_fill_1 FILLER_38_446 ();
 sg13g2_fill_1 FILLER_38_486 ();
 sg13g2_decap_8 FILLER_38_501 ();
 sg13g2_fill_2 FILLER_38_508 ();
 sg13g2_fill_1 FILLER_38_510 ();
 sg13g2_decap_4 FILLER_38_528 ();
 sg13g2_fill_2 FILLER_38_532 ();
 sg13g2_fill_1 FILLER_38_547 ();
 sg13g2_fill_1 FILLER_38_552 ();
 sg13g2_decap_8 FILLER_38_562 ();
 sg13g2_decap_8 FILLER_38_569 ();
 sg13g2_fill_2 FILLER_38_576 ();
 sg13g2_fill_1 FILLER_38_578 ();
 sg13g2_fill_2 FILLER_38_592 ();
 sg13g2_fill_1 FILLER_38_594 ();
 sg13g2_fill_2 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_618 ();
 sg13g2_fill_2 FILLER_38_625 ();
 sg13g2_decap_8 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_655 ();
 sg13g2_decap_4 FILLER_38_662 ();
 sg13g2_fill_1 FILLER_38_666 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_fill_2 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_fill_2 FILLER_38_725 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_739 ();
 sg13g2_decap_4 FILLER_38_769 ();
 sg13g2_fill_1 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_fill_2 FILLER_38_794 ();
 sg13g2_fill_1 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_4 FILLER_38_816 ();
 sg13g2_fill_2 FILLER_38_820 ();
 sg13g2_fill_1 FILLER_38_826 ();
 sg13g2_decap_4 FILLER_38_840 ();
 sg13g2_fill_1 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_853 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_fill_2 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_4 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_fill_2 FILLER_39_145 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_fill_2 FILLER_39_180 ();
 sg13g2_fill_2 FILLER_39_187 ();
 sg13g2_fill_1 FILLER_39_197 ();
 sg13g2_fill_2 FILLER_39_212 ();
 sg13g2_decap_4 FILLER_39_224 ();
 sg13g2_fill_2 FILLER_39_228 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_2 FILLER_39_273 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_326 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_346 ();
 sg13g2_decap_8 FILLER_39_353 ();
 sg13g2_fill_2 FILLER_39_360 ();
 sg13g2_decap_4 FILLER_39_428 ();
 sg13g2_fill_2 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_493 ();
 sg13g2_fill_2 FILLER_39_551 ();
 sg13g2_decap_4 FILLER_39_569 ();
 sg13g2_fill_2 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_579 ();
 sg13g2_decap_4 FILLER_39_594 ();
 sg13g2_decap_4 FILLER_39_603 ();
 sg13g2_decap_8 FILLER_39_617 ();
 sg13g2_fill_2 FILLER_39_624 ();
 sg13g2_fill_1 FILLER_39_626 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_decap_8 FILLER_39_649 ();
 sg13g2_decap_4 FILLER_39_688 ();
 sg13g2_fill_1 FILLER_39_692 ();
 sg13g2_decap_4 FILLER_39_718 ();
 sg13g2_fill_1 FILLER_39_744 ();
 sg13g2_decap_8 FILLER_39_762 ();
 sg13g2_decap_4 FILLER_39_769 ();
 sg13g2_fill_1 FILLER_39_790 ();
 sg13g2_fill_2 FILLER_39_799 ();
 sg13g2_decap_4 FILLER_39_823 ();
 sg13g2_fill_1 FILLER_39_840 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_4 FILLER_40_25 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_2 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_57 ();
 sg13g2_decap_4 FILLER_40_64 ();
 sg13g2_fill_2 FILLER_40_68 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_81 ();
 sg13g2_fill_2 FILLER_40_107 ();
 sg13g2_decap_4 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_152 ();
 sg13g2_decap_4 FILLER_40_163 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_fill_2 FILLER_40_184 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_decap_4 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_239 ();
 sg13g2_decap_4 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_249 ();
 sg13g2_fill_2 FILLER_40_270 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_348 ();
 sg13g2_decap_8 FILLER_40_353 ();
 sg13g2_decap_8 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_fill_1 FILLER_40_465 ();
 sg13g2_fill_2 FILLER_40_488 ();
 sg13g2_fill_1 FILLER_40_495 ();
 sg13g2_decap_8 FILLER_40_499 ();
 sg13g2_decap_8 FILLER_40_506 ();
 sg13g2_fill_2 FILLER_40_513 ();
 sg13g2_fill_1 FILLER_40_515 ();
 sg13g2_decap_8 FILLER_40_529 ();
 sg13g2_decap_4 FILLER_40_536 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_554 ();
 sg13g2_fill_2 FILLER_40_564 ();
 sg13g2_fill_1 FILLER_40_570 ();
 sg13g2_fill_2 FILLER_40_584 ();
 sg13g2_fill_2 FILLER_40_590 ();
 sg13g2_decap_4 FILLER_40_602 ();
 sg13g2_fill_2 FILLER_40_614 ();
 sg13g2_fill_1 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_fill_1 FILLER_40_637 ();
 sg13g2_fill_1 FILLER_40_644 ();
 sg13g2_fill_2 FILLER_40_661 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_fill_2 FILLER_40_683 ();
 sg13g2_fill_1 FILLER_40_685 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_fill_2 FILLER_40_719 ();
 sg13g2_fill_1 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_739 ();
 sg13g2_decap_4 FILLER_40_746 ();
 sg13g2_fill_1 FILLER_40_750 ();
 sg13g2_fill_1 FILLER_40_759 ();
 sg13g2_fill_2 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_decap_4 FILLER_40_794 ();
 sg13g2_fill_1 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_fill_2 FILLER_40_814 ();
 sg13g2_fill_1 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_829 ();
 sg13g2_decap_4 FILLER_40_836 ();
 sg13g2_fill_2 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_850 ();
 sg13g2_decap_4 FILLER_40_857 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_11 ();
 sg13g2_fill_2 FILLER_41_76 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_128 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_142 ();
 sg13g2_decap_8 FILLER_41_148 ();
 sg13g2_fill_2 FILLER_41_155 ();
 sg13g2_decap_8 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_169 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_fill_2 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_decap_4 FILLER_41_183 ();
 sg13g2_fill_2 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_229 ();
 sg13g2_fill_1 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_240 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_fill_2 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_270 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_decap_4 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_359 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_fill_2 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_425 ();
 sg13g2_fill_2 FILLER_41_439 ();
 sg13g2_fill_2 FILLER_41_495 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_fill_2 FILLER_41_571 ();
 sg13g2_decap_4 FILLER_41_582 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_decap_8 FILLER_41_596 ();
 sg13g2_fill_1 FILLER_41_603 ();
 sg13g2_decap_4 FILLER_41_618 ();
 sg13g2_decap_4 FILLER_41_651 ();
 sg13g2_fill_1 FILLER_41_655 ();
 sg13g2_decap_4 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_673 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_687 ();
 sg13g2_decap_4 FILLER_41_693 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_decap_8 FILLER_41_706 ();
 sg13g2_decap_4 FILLER_41_743 ();
 sg13g2_decap_4 FILLER_41_764 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_4 FILLER_41_800 ();
 sg13g2_decap_4 FILLER_41_809 ();
 sg13g2_fill_1 FILLER_41_813 ();
 sg13g2_fill_2 FILLER_41_823 ();
 sg13g2_fill_2 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_859 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_fill_2 FILLER_42_84 ();
 sg13g2_fill_1 FILLER_42_86 ();
 sg13g2_fill_1 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_122 ();
 sg13g2_fill_1 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_177 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_191 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_decap_4 FILLER_42_230 ();
 sg13g2_fill_2 FILLER_42_234 ();
 sg13g2_decap_4 FILLER_42_250 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_fill_1 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_272 ();
 sg13g2_decap_8 FILLER_42_279 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_312 ();
 sg13g2_decap_4 FILLER_42_378 ();
 sg13g2_fill_2 FILLER_42_410 ();
 sg13g2_fill_1 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_450 ();
 sg13g2_decap_4 FILLER_42_457 ();
 sg13g2_fill_2 FILLER_42_461 ();
 sg13g2_decap_8 FILLER_42_498 ();
 sg13g2_decap_8 FILLER_42_505 ();
 sg13g2_decap_4 FILLER_42_512 ();
 sg13g2_fill_2 FILLER_42_516 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_fill_1 FILLER_42_559 ();
 sg13g2_decap_4 FILLER_42_581 ();
 sg13g2_fill_2 FILLER_42_585 ();
 sg13g2_decap_4 FILLER_42_591 ();
 sg13g2_fill_1 FILLER_42_595 ();
 sg13g2_fill_1 FILLER_42_604 ();
 sg13g2_decap_8 FILLER_42_620 ();
 sg13g2_decap_8 FILLER_42_627 ();
 sg13g2_decap_8 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_641 ();
 sg13g2_fill_2 FILLER_42_658 ();
 sg13g2_fill_1 FILLER_42_660 ();
 sg13g2_fill_2 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_fill_1 FILLER_42_710 ();
 sg13g2_decap_8 FILLER_42_715 ();
 sg13g2_decap_4 FILLER_42_739 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_fill_1 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_787 ();
 sg13g2_decap_4 FILLER_42_794 ();
 sg13g2_fill_2 FILLER_42_807 ();
 sg13g2_fill_1 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_835 ();
 sg13g2_fill_1 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_855 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_2 FILLER_43_66 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_decap_8 FILLER_43_86 ();
 sg13g2_decap_8 FILLER_43_93 ();
 sg13g2_fill_2 FILLER_43_100 ();
 sg13g2_fill_1 FILLER_43_102 ();
 sg13g2_decap_4 FILLER_43_124 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_146 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_decap_8 FILLER_43_199 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_222 ();
 sg13g2_decap_4 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_233 ();
 sg13g2_decap_8 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_247 ();
 sg13g2_fill_2 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_decap_4 FILLER_43_307 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_2 FILLER_43_349 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_decap_8 FILLER_43_411 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_425 ();
 sg13g2_fill_1 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_fill_2 FILLER_43_466 ();
 sg13g2_decap_8 FILLER_43_503 ();
 sg13g2_decap_4 FILLER_43_510 ();
 sg13g2_fill_1 FILLER_43_514 ();
 sg13g2_fill_2 FILLER_43_549 ();
 sg13g2_fill_1 FILLER_43_551 ();
 sg13g2_decap_4 FILLER_43_564 ();
 sg13g2_fill_2 FILLER_43_568 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_4 FILLER_43_581 ();
 sg13g2_fill_1 FILLER_43_589 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_4 FILLER_43_602 ();
 sg13g2_decap_4 FILLER_43_610 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_636 ();
 sg13g2_fill_2 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_655 ();
 sg13g2_decap_4 FILLER_43_662 ();
 sg13g2_fill_1 FILLER_43_666 ();
 sg13g2_decap_8 FILLER_43_675 ();
 sg13g2_fill_2 FILLER_43_686 ();
 sg13g2_fill_2 FILLER_43_701 ();
 sg13g2_decap_8 FILLER_43_720 ();
 sg13g2_fill_1 FILLER_43_727 ();
 sg13g2_decap_8 FILLER_43_733 ();
 sg13g2_fill_2 FILLER_43_740 ();
 sg13g2_fill_1 FILLER_43_742 ();
 sg13g2_fill_1 FILLER_43_751 ();
 sg13g2_decap_8 FILLER_43_757 ();
 sg13g2_decap_8 FILLER_43_764 ();
 sg13g2_decap_8 FILLER_43_786 ();
 sg13g2_fill_1 FILLER_43_793 ();
 sg13g2_decap_4 FILLER_43_827 ();
 sg13g2_fill_2 FILLER_43_831 ();
 sg13g2_decap_4 FILLER_43_856 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_13 ();
 sg13g2_decap_8 FILLER_44_20 ();
 sg13g2_fill_2 FILLER_44_61 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_fill_2 FILLER_44_105 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_142 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_fill_2 FILLER_44_163 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_4 FILLER_44_225 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_242 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_fill_2 FILLER_44_272 ();
 sg13g2_fill_1 FILLER_44_274 ();
 sg13g2_fill_2 FILLER_44_280 ();
 sg13g2_fill_2 FILLER_44_288 ();
 sg13g2_fill_2 FILLER_44_366 ();
 sg13g2_fill_1 FILLER_44_368 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_fill_2 FILLER_44_393 ();
 sg13g2_decap_4 FILLER_44_432 ();
 sg13g2_fill_1 FILLER_44_436 ();
 sg13g2_fill_1 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_532 ();
 sg13g2_fill_1 FILLER_44_534 ();
 sg13g2_fill_1 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_548 ();
 sg13g2_fill_1 FILLER_44_555 ();
 sg13g2_decap_4 FILLER_44_601 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_625 ();
 sg13g2_fill_1 FILLER_44_632 ();
 sg13g2_decap_8 FILLER_44_646 ();
 sg13g2_fill_1 FILLER_44_653 ();
 sg13g2_fill_2 FILLER_44_667 ();
 sg13g2_decap_8 FILLER_44_685 ();
 sg13g2_decap_8 FILLER_44_692 ();
 sg13g2_decap_8 FILLER_44_717 ();
 sg13g2_decap_4 FILLER_44_724 ();
 sg13g2_fill_1 FILLER_44_728 ();
 sg13g2_decap_4 FILLER_44_737 ();
 sg13g2_fill_1 FILLER_44_741 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_4 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_fill_1 FILLER_44_802 ();
 sg13g2_decap_4 FILLER_44_808 ();
 sg13g2_fill_1 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_818 ();
 sg13g2_decap_4 FILLER_44_825 ();
 sg13g2_fill_2 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_857 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_decap_4 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_31 ();
 sg13g2_decap_8 FILLER_45_74 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_fill_2 FILLER_45_88 ();
 sg13g2_decap_4 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_decap_4 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_170 ();
 sg13g2_decap_8 FILLER_45_188 ();
 sg13g2_decap_8 FILLER_45_195 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_fill_1 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_257 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_decap_4 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_343 ();
 sg13g2_fill_1 FILLER_45_363 ();
 sg13g2_decap_4 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_377 ();
 sg13g2_decap_8 FILLER_45_447 ();
 sg13g2_fill_2 FILLER_45_454 ();
 sg13g2_decap_8 FILLER_45_482 ();
 sg13g2_decap_4 FILLER_45_503 ();
 sg13g2_fill_2 FILLER_45_507 ();
 sg13g2_fill_2 FILLER_45_535 ();
 sg13g2_fill_2 FILLER_45_557 ();
 sg13g2_decap_4 FILLER_45_567 ();
 sg13g2_decap_4 FILLER_45_574 ();
 sg13g2_decap_4 FILLER_45_583 ();
 sg13g2_fill_1 FILLER_45_587 ();
 sg13g2_decap_8 FILLER_45_593 ();
 sg13g2_fill_1 FILLER_45_600 ();
 sg13g2_fill_2 FILLER_45_609 ();
 sg13g2_fill_1 FILLER_45_611 ();
 sg13g2_decap_8 FILLER_45_620 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_decap_8 FILLER_45_643 ();
 sg13g2_fill_1 FILLER_45_650 ();
 sg13g2_decap_4 FILLER_45_667 ();
 sg13g2_fill_1 FILLER_45_677 ();
 sg13g2_decap_4 FILLER_45_688 ();
 sg13g2_fill_2 FILLER_45_692 ();
 sg13g2_fill_2 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_708 ();
 sg13g2_decap_4 FILLER_45_739 ();
 sg13g2_fill_1 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_fill_2 FILLER_45_771 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_fill_2 FILLER_45_782 ();
 sg13g2_fill_1 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_790 ();
 sg13g2_fill_1 FILLER_45_797 ();
 sg13g2_fill_2 FILLER_45_806 ();
 sg13g2_decap_4 FILLER_45_824 ();
 sg13g2_decap_4 FILLER_45_840 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_1 FILLER_46_107 ();
 sg13g2_fill_2 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_fill_2 FILLER_46_186 ();
 sg13g2_decap_4 FILLER_46_204 ();
 sg13g2_fill_1 FILLER_46_208 ();
 sg13g2_fill_2 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_240 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_293 ();
 sg13g2_fill_2 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_1 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_559 ();
 sg13g2_decap_4 FILLER_46_600 ();
 sg13g2_fill_2 FILLER_46_604 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_fill_2 FILLER_46_637 ();
 sg13g2_fill_1 FILLER_46_639 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_fill_1 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_685 ();
 sg13g2_decap_4 FILLER_46_692 ();
 sg13g2_fill_2 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_713 ();
 sg13g2_decap_4 FILLER_46_720 ();
 sg13g2_fill_2 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_4 FILLER_46_745 ();
 sg13g2_decap_4 FILLER_46_752 ();
 sg13g2_decap_4 FILLER_46_764 ();
 sg13g2_fill_2 FILLER_46_768 ();
 sg13g2_fill_1 FILLER_46_778 ();
 sg13g2_decap_4 FILLER_46_795 ();
 sg13g2_fill_2 FILLER_46_799 ();
 sg13g2_decap_4 FILLER_46_806 ();
 sg13g2_fill_2 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_decap_4 FILLER_46_824 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_17 ();
 sg13g2_fill_1 FILLER_47_19 ();
 sg13g2_decap_8 FILLER_47_30 ();
 sg13g2_decap_4 FILLER_47_37 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_fill_2 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_60 ();
 sg13g2_decap_4 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_4 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_152 ();
 sg13g2_decap_4 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_fill_2 FILLER_47_180 ();
 sg13g2_decap_8 FILLER_47_194 ();
 sg13g2_decap_8 FILLER_47_201 ();
 sg13g2_decap_8 FILLER_47_208 ();
 sg13g2_decap_8 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_250 ();
 sg13g2_decap_8 FILLER_47_256 ();
 sg13g2_fill_2 FILLER_47_263 ();
 sg13g2_decap_4 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_decap_8 FILLER_47_281 ();
 sg13g2_decap_8 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_decap_4 FILLER_47_314 ();
 sg13g2_decap_8 FILLER_47_331 ();
 sg13g2_decap_8 FILLER_47_338 ();
 sg13g2_fill_2 FILLER_47_345 ();
 sg13g2_decap_4 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_359 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_fill_1 FILLER_47_385 ();
 sg13g2_fill_1 FILLER_47_435 ();
 sg13g2_fill_2 FILLER_47_449 ();
 sg13g2_fill_1 FILLER_47_451 ();
 sg13g2_decap_8 FILLER_47_505 ();
 sg13g2_decap_8 FILLER_47_512 ();
 sg13g2_decap_4 FILLER_47_519 ();
 sg13g2_decap_4 FILLER_47_529 ();
 sg13g2_fill_1 FILLER_47_533 ();
 sg13g2_decap_8 FILLER_47_557 ();
 sg13g2_decap_4 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_568 ();
 sg13g2_fill_2 FILLER_47_574 ();
 sg13g2_decap_4 FILLER_47_580 ();
 sg13g2_fill_2 FILLER_47_584 ();
 sg13g2_decap_8 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_604 ();
 sg13g2_fill_1 FILLER_47_613 ();
 sg13g2_decap_8 FILLER_47_627 ();
 sg13g2_decap_4 FILLER_47_687 ();
 sg13g2_fill_2 FILLER_47_691 ();
 sg13g2_decap_4 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_fill_1 FILLER_47_759 ();
 sg13g2_fill_2 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_792 ();
 sg13g2_decap_4 FILLER_47_799 ();
 sg13g2_fill_2 FILLER_47_808 ();
 sg13g2_fill_1 FILLER_47_815 ();
 sg13g2_decap_4 FILLER_47_836 ();
 sg13g2_fill_2 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_25 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_1 FILLER_48_55 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_decap_4 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_122 ();
 sg13g2_fill_2 FILLER_48_129 ();
 sg13g2_decap_8 FILLER_48_166 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_fill_2 FILLER_48_196 ();
 sg13g2_decap_4 FILLER_48_212 ();
 sg13g2_fill_2 FILLER_48_216 ();
 sg13g2_decap_4 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_243 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_decap_8 FILLER_48_285 ();
 sg13g2_decap_8 FILLER_48_292 ();
 sg13g2_fill_2 FILLER_48_304 ();
 sg13g2_decap_4 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_315 ();
 sg13g2_decap_4 FILLER_48_322 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_fill_1 FILLER_48_335 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_fill_2 FILLER_48_375 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_fill_2 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_391 ();
 sg13g2_fill_2 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_4 FILLER_48_420 ();
 sg13g2_fill_1 FILLER_48_481 ();
 sg13g2_decap_4 FILLER_48_501 ();
 sg13g2_fill_2 FILLER_48_505 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_8 FILLER_48_542 ();
 sg13g2_fill_2 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_580 ();
 sg13g2_fill_2 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_603 ();
 sg13g2_decap_8 FILLER_48_610 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_fill_1 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_fill_1 FILLER_48_665 ();
 sg13g2_fill_1 FILLER_48_670 ();
 sg13g2_decap_8 FILLER_48_681 ();
 sg13g2_decap_8 FILLER_48_688 ();
 sg13g2_fill_2 FILLER_48_695 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_709 ();
 sg13g2_fill_2 FILLER_48_716 ();
 sg13g2_decap_4 FILLER_48_739 ();
 sg13g2_fill_2 FILLER_48_743 ();
 sg13g2_fill_2 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_decap_8 FILLER_48_774 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_fill_2 FILLER_48_793 ();
 sg13g2_fill_1 FILLER_48_803 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_fill_2 FILLER_48_826 ();
 sg13g2_fill_2 FILLER_48_841 ();
 sg13g2_fill_1 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_36 ();
 sg13g2_fill_1 FILLER_49_38 ();
 sg13g2_decap_8 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_decap_4 FILLER_49_77 ();
 sg13g2_decap_4 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_109 ();
 sg13g2_fill_2 FILLER_49_115 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_decap_4 FILLER_49_143 ();
 sg13g2_fill_2 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_fill_2 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_fill_1 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_4 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_218 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_decap_8 FILLER_49_237 ();
 sg13g2_decap_8 FILLER_49_244 ();
 sg13g2_decap_4 FILLER_49_251 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_311 ();
 sg13g2_decap_4 FILLER_49_338 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_357 ();
 sg13g2_fill_1 FILLER_49_372 ();
 sg13g2_fill_1 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_410 ();
 sg13g2_fill_1 FILLER_49_412 ();
 sg13g2_fill_1 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_490 ();
 sg13g2_decap_4 FILLER_49_501 ();
 sg13g2_fill_2 FILLER_49_505 ();
 sg13g2_decap_8 FILLER_49_535 ();
 sg13g2_decap_4 FILLER_49_542 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_fill_2 FILLER_49_574 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_fill_2 FILLER_49_595 ();
 sg13g2_fill_2 FILLER_49_605 ();
 sg13g2_fill_2 FILLER_49_654 ();
 sg13g2_fill_1 FILLER_49_656 ();
 sg13g2_fill_2 FILLER_49_685 ();
 sg13g2_fill_1 FILLER_49_687 ();
 sg13g2_decap_8 FILLER_49_713 ();
 sg13g2_decap_4 FILLER_49_720 ();
 sg13g2_fill_1 FILLER_49_724 ();
 sg13g2_fill_2 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_740 ();
 sg13g2_fill_2 FILLER_49_747 ();
 sg13g2_fill_1 FILLER_49_749 ();
 sg13g2_fill_2 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_fill_2 FILLER_49_808 ();
 sg13g2_fill_1 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_4 FILLER_49_831 ();
 sg13g2_fill_1 FILLER_49_835 ();
 sg13g2_decap_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_22 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_fill_2 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_59 ();
 sg13g2_fill_1 FILLER_50_61 ();
 sg13g2_decap_8 FILLER_50_66 ();
 sg13g2_decap_4 FILLER_50_73 ();
 sg13g2_decap_8 FILLER_50_82 ();
 sg13g2_decap_4 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_114 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_decap_8 FILLER_50_162 ();
 sg13g2_decap_8 FILLER_50_169 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_decap_4 FILLER_50_193 ();
 sg13g2_decap_4 FILLER_50_219 ();
 sg13g2_decap_4 FILLER_50_244 ();
 sg13g2_decap_8 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_decap_4 FILLER_50_319 ();
 sg13g2_decap_8 FILLER_50_347 ();
 sg13g2_decap_4 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_4 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_fill_2 FILLER_50_441 ();
 sg13g2_fill_1 FILLER_50_443 ();
 sg13g2_fill_2 FILLER_50_466 ();
 sg13g2_fill_2 FILLER_50_534 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_2 FILLER_50_572 ();
 sg13g2_fill_2 FILLER_50_578 ();
 sg13g2_decap_8 FILLER_50_606 ();
 sg13g2_fill_2 FILLER_50_613 ();
 sg13g2_decap_8 FILLER_50_623 ();
 sg13g2_fill_2 FILLER_50_630 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_decap_8 FILLER_50_658 ();
 sg13g2_fill_2 FILLER_50_665 ();
 sg13g2_fill_1 FILLER_50_667 ();
 sg13g2_fill_2 FILLER_50_676 ();
 sg13g2_decap_8 FILLER_50_682 ();
 sg13g2_fill_2 FILLER_50_702 ();
 sg13g2_fill_1 FILLER_50_704 ();
 sg13g2_fill_1 FILLER_50_726 ();
 sg13g2_decap_8 FILLER_50_748 ();
 sg13g2_decap_4 FILLER_50_755 ();
 sg13g2_fill_1 FILLER_50_759 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_fill_1 FILLER_50_767 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_4 FILLER_50_800 ();
 sg13g2_fill_2 FILLER_50_804 ();
 sg13g2_decap_4 FILLER_50_831 ();
 sg13g2_fill_2 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_24 ();
 sg13g2_fill_2 FILLER_51_45 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_1 FILLER_51_66 ();
 sg13g2_decap_8 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_121 ();
 sg13g2_fill_2 FILLER_51_127 ();
 sg13g2_fill_1 FILLER_51_129 ();
 sg13g2_decap_8 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_fill_1 FILLER_51_156 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_fill_2 FILLER_51_181 ();
 sg13g2_fill_1 FILLER_51_183 ();
 sg13g2_fill_1 FILLER_51_192 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_223 ();
 sg13g2_decap_4 FILLER_51_240 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_decap_4 FILLER_51_269 ();
 sg13g2_decap_4 FILLER_51_281 ();
 sg13g2_decap_8 FILLER_51_289 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_fill_2 FILLER_51_331 ();
 sg13g2_fill_1 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_406 ();
 sg13g2_fill_2 FILLER_51_460 ();
 sg13g2_fill_1 FILLER_51_462 ();
 sg13g2_fill_1 FILLER_51_467 ();
 sg13g2_fill_2 FILLER_51_478 ();
 sg13g2_fill_1 FILLER_51_480 ();
 sg13g2_fill_2 FILLER_51_566 ();
 sg13g2_fill_1 FILLER_51_568 ();
 sg13g2_fill_2 FILLER_51_579 ();
 sg13g2_fill_1 FILLER_51_581 ();
 sg13g2_decap_8 FILLER_51_588 ();
 sg13g2_fill_1 FILLER_51_603 ();
 sg13g2_decap_4 FILLER_51_620 ();
 sg13g2_fill_1 FILLER_51_624 ();
 sg13g2_fill_1 FILLER_51_631 ();
 sg13g2_decap_8 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_660 ();
 sg13g2_fill_1 FILLER_51_667 ();
 sg13g2_decap_8 FILLER_51_688 ();
 sg13g2_decap_4 FILLER_51_695 ();
 sg13g2_fill_1 FILLER_51_699 ();
 sg13g2_fill_1 FILLER_51_717 ();
 sg13g2_decap_8 FILLER_51_726 ();
 sg13g2_fill_1 FILLER_51_745 ();
 sg13g2_decap_4 FILLER_51_754 ();
 sg13g2_decap_8 FILLER_51_771 ();
 sg13g2_fill_2 FILLER_51_815 ();
 sg13g2_decap_4 FILLER_51_830 ();
 sg13g2_fill_2 FILLER_51_834 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_decap_8 FILLER_51_851 ();
 sg13g2_decap_4 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_31 ();
 sg13g2_decap_8 FILLER_52_38 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_decap_4 FILLER_52_67 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_119 ();
 sg13g2_decap_4 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_2 FILLER_52_193 ();
 sg13g2_fill_1 FILLER_52_195 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_decap_8 FILLER_52_243 ();
 sg13g2_decap_8 FILLER_52_250 ();
 sg13g2_fill_1 FILLER_52_262 ();
 sg13g2_decap_8 FILLER_52_268 ();
 sg13g2_fill_2 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_364 ();
 sg13g2_decap_4 FILLER_52_391 ();
 sg13g2_fill_2 FILLER_52_413 ();
 sg13g2_fill_2 FILLER_52_424 ();
 sg13g2_fill_1 FILLER_52_426 ();
 sg13g2_fill_1 FILLER_52_467 ();
 sg13g2_decap_8 FILLER_52_481 ();
 sg13g2_decap_8 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_505 ();
 sg13g2_decap_8 FILLER_52_558 ();
 sg13g2_fill_1 FILLER_52_569 ();
 sg13g2_decap_8 FILLER_52_583 ();
 sg13g2_fill_2 FILLER_52_590 ();
 sg13g2_fill_1 FILLER_52_592 ();
 sg13g2_fill_2 FILLER_52_606 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_626 ();
 sg13g2_decap_8 FILLER_52_643 ();
 sg13g2_decap_4 FILLER_52_650 ();
 sg13g2_fill_1 FILLER_52_654 ();
 sg13g2_decap_4 FILLER_52_673 ();
 sg13g2_fill_1 FILLER_52_685 ();
 sg13g2_decap_8 FILLER_52_691 ();
 sg13g2_decap_8 FILLER_52_698 ();
 sg13g2_fill_2 FILLER_52_705 ();
 sg13g2_fill_1 FILLER_52_707 ();
 sg13g2_fill_1 FILLER_52_713 ();
 sg13g2_fill_1 FILLER_52_722 ();
 sg13g2_decap_8 FILLER_52_727 ();
 sg13g2_decap_8 FILLER_52_734 ();
 sg13g2_fill_1 FILLER_52_741 ();
 sg13g2_decap_8 FILLER_52_747 ();
 sg13g2_decap_8 FILLER_52_754 ();
 sg13g2_fill_2 FILLER_52_761 ();
 sg13g2_fill_1 FILLER_52_780 ();
 sg13g2_decap_8 FILLER_52_789 ();
 sg13g2_decap_8 FILLER_52_796 ();
 sg13g2_decap_4 FILLER_52_803 ();
 sg13g2_decap_4 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_852 ();
 sg13g2_fill_2 FILLER_52_859 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_29 ();
 sg13g2_decap_4 FILLER_53_36 ();
 sg13g2_decap_8 FILLER_53_66 ();
 sg13g2_decap_8 FILLER_53_73 ();
 sg13g2_fill_1 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_114 ();
 sg13g2_fill_2 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_decap_4 FILLER_53_144 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_decap_8 FILLER_53_172 ();
 sg13g2_decap_8 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_199 ();
 sg13g2_decap_4 FILLER_53_224 ();
 sg13g2_fill_2 FILLER_53_228 ();
 sg13g2_decap_8 FILLER_53_240 ();
 sg13g2_decap_4 FILLER_53_247 ();
 sg13g2_fill_2 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_fill_2 FILLER_53_310 ();
 sg13g2_fill_1 FILLER_53_312 ();
 sg13g2_decap_8 FILLER_53_354 ();
 sg13g2_decap_4 FILLER_53_361 ();
 sg13g2_fill_2 FILLER_53_398 ();
 sg13g2_fill_2 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_4 FILLER_53_441 ();
 sg13g2_fill_1 FILLER_53_445 ();
 sg13g2_fill_1 FILLER_53_475 ();
 sg13g2_decap_8 FILLER_53_578 ();
 sg13g2_decap_8 FILLER_53_585 ();
 sg13g2_decap_8 FILLER_53_592 ();
 sg13g2_decap_4 FILLER_53_620 ();
 sg13g2_fill_1 FILLER_53_624 ();
 sg13g2_decap_8 FILLER_53_635 ();
 sg13g2_fill_2 FILLER_53_642 ();
 sg13g2_fill_1 FILLER_53_644 ();
 sg13g2_fill_2 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_decap_4 FILLER_53_675 ();
 sg13g2_fill_2 FILLER_53_679 ();
 sg13g2_fill_1 FILLER_53_697 ();
 sg13g2_decap_4 FILLER_53_703 ();
 sg13g2_fill_2 FILLER_53_720 ();
 sg13g2_fill_1 FILLER_53_722 ();
 sg13g2_decap_8 FILLER_53_757 ();
 sg13g2_fill_1 FILLER_53_772 ();
 sg13g2_fill_1 FILLER_53_786 ();
 sg13g2_decap_8 FILLER_53_799 ();
 sg13g2_fill_1 FILLER_53_817 ();
 sg13g2_decap_4 FILLER_53_826 ();
 sg13g2_fill_1 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_12 ();
 sg13g2_decap_8 FILLER_54_19 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_57 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_decap_4 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_74 ();
 sg13g2_decap_4 FILLER_54_98 ();
 sg13g2_fill_2 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_108 ();
 sg13g2_decap_4 FILLER_54_123 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_decap_8 FILLER_54_141 ();
 sg13g2_decap_8 FILLER_54_148 ();
 sg13g2_fill_2 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_157 ();
 sg13g2_decap_4 FILLER_54_163 ();
 sg13g2_decap_8 FILLER_54_172 ();
 sg13g2_decap_4 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_192 ();
 sg13g2_fill_2 FILLER_54_199 ();
 sg13g2_fill_1 FILLER_54_201 ();
 sg13g2_decap_8 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_241 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_8 FILLER_54_264 ();
 sg13g2_decap_4 FILLER_54_271 ();
 sg13g2_decap_4 FILLER_54_281 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_decap_8 FILLER_54_291 ();
 sg13g2_fill_2 FILLER_54_298 ();
 sg13g2_fill_1 FILLER_54_300 ();
 sg13g2_fill_2 FILLER_54_327 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_decap_8 FILLER_54_353 ();
 sg13g2_decap_4 FILLER_54_360 ();
 sg13g2_fill_1 FILLER_54_364 ();
 sg13g2_fill_2 FILLER_54_379 ();
 sg13g2_fill_1 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_fill_1 FILLER_54_398 ();
 sg13g2_fill_2 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_424 ();
 sg13g2_decap_8 FILLER_54_504 ();
 sg13g2_fill_1 FILLER_54_511 ();
 sg13g2_decap_8 FILLER_54_518 ();
 sg13g2_fill_2 FILLER_54_525 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_2 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_582 ();
 sg13g2_fill_1 FILLER_54_591 ();
 sg13g2_decap_8 FILLER_54_612 ();
 sg13g2_fill_1 FILLER_54_619 ();
 sg13g2_fill_1 FILLER_54_635 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_decap_8 FILLER_54_655 ();
 sg13g2_decap_4 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_681 ();
 sg13g2_fill_2 FILLER_54_692 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_decap_8 FILLER_54_711 ();
 sg13g2_decap_4 FILLER_54_718 ();
 sg13g2_fill_1 FILLER_54_722 ();
 sg13g2_decap_8 FILLER_54_735 ();
 sg13g2_decap_4 FILLER_54_759 ();
 sg13g2_fill_1 FILLER_54_763 ();
 sg13g2_decap_8 FILLER_54_776 ();
 sg13g2_fill_2 FILLER_54_783 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_fill_2 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_807 ();
 sg13g2_decap_4 FILLER_54_813 ();
 sg13g2_fill_2 FILLER_54_817 ();
 sg13g2_decap_8 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_836 ();
 sg13g2_decap_8 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_4 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_1 FILLER_55_31 ();
 sg13g2_decap_8 FILLER_55_52 ();
 sg13g2_fill_2 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_71 ();
 sg13g2_decap_8 FILLER_55_82 ();
 sg13g2_decap_8 FILLER_55_89 ();
 sg13g2_decap_4 FILLER_55_96 ();
 sg13g2_fill_1 FILLER_55_116 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_decap_4 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_decap_8 FILLER_55_183 ();
 sg13g2_decap_4 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_199 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_216 ();
 sg13g2_decap_8 FILLER_55_223 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_decap_8 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_253 ();
 sg13g2_decap_8 FILLER_55_260 ();
 sg13g2_decap_4 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_276 ();
 sg13g2_decap_8 FILLER_55_283 ();
 sg13g2_decap_8 FILLER_55_290 ();
 sg13g2_decap_8 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_312 ();
 sg13g2_decap_8 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_326 ();
 sg13g2_decap_4 FILLER_55_359 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_fill_2 FILLER_55_373 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_decap_4 FILLER_55_402 ();
 sg13g2_decap_4 FILLER_55_438 ();
 sg13g2_fill_2 FILLER_55_464 ();
 sg13g2_fill_1 FILLER_55_466 ();
 sg13g2_decap_8 FILLER_55_480 ();
 sg13g2_fill_2 FILLER_55_497 ();
 sg13g2_fill_1 FILLER_55_499 ();
 sg13g2_fill_2 FILLER_55_554 ();
 sg13g2_fill_2 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_574 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_decap_8 FILLER_55_596 ();
 sg13g2_decap_8 FILLER_55_608 ();
 sg13g2_decap_8 FILLER_55_615 ();
 sg13g2_decap_4 FILLER_55_622 ();
 sg13g2_fill_1 FILLER_55_626 ();
 sg13g2_fill_1 FILLER_55_636 ();
 sg13g2_fill_1 FILLER_55_650 ();
 sg13g2_decap_8 FILLER_55_662 ();
 sg13g2_fill_2 FILLER_55_669 ();
 sg13g2_fill_1 FILLER_55_671 ();
 sg13g2_fill_2 FILLER_55_680 ();
 sg13g2_fill_1 FILLER_55_682 ();
 sg13g2_decap_8 FILLER_55_691 ();
 sg13g2_fill_2 FILLER_55_698 ();
 sg13g2_decap_8 FILLER_55_710 ();
 sg13g2_decap_8 FILLER_55_717 ();
 sg13g2_decap_4 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_754 ();
 sg13g2_decap_8 FILLER_55_761 ();
 sg13g2_fill_2 FILLER_55_768 ();
 sg13g2_fill_1 FILLER_55_770 ();
 sg13g2_fill_2 FILLER_55_779 ();
 sg13g2_fill_1 FILLER_55_781 ();
 sg13g2_decap_8 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_810 ();
 sg13g2_decap_4 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_4 FILLER_55_857 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_12 ();
 sg13g2_fill_2 FILLER_56_19 ();
 sg13g2_fill_1 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_40 ();
 sg13g2_fill_2 FILLER_56_50 ();
 sg13g2_fill_1 FILLER_56_52 ();
 sg13g2_fill_2 FILLER_56_88 ();
 sg13g2_fill_1 FILLER_56_90 ();
 sg13g2_decap_4 FILLER_56_106 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_fill_2 FILLER_56_122 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_decap_4 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_167 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_267 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_decap_4 FILLER_56_314 ();
 sg13g2_fill_2 FILLER_56_318 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_fill_1 FILLER_56_363 ();
 sg13g2_fill_2 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_397 ();
 sg13g2_fill_2 FILLER_56_413 ();
 sg13g2_fill_1 FILLER_56_419 ();
 sg13g2_decap_8 FILLER_56_429 ();
 sg13g2_decap_8 FILLER_56_436 ();
 sg13g2_fill_2 FILLER_56_443 ();
 sg13g2_fill_1 FILLER_56_445 ();
 sg13g2_decap_8 FILLER_56_456 ();
 sg13g2_fill_1 FILLER_56_463 ();
 sg13g2_fill_2 FILLER_56_473 ();
 sg13g2_decap_8 FILLER_56_503 ();
 sg13g2_decap_8 FILLER_56_510 ();
 sg13g2_decap_8 FILLER_56_564 ();
 sg13g2_fill_1 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_fill_2 FILLER_56_589 ();
 sg13g2_fill_1 FILLER_56_591 ();
 sg13g2_decap_4 FILLER_56_636 ();
 sg13g2_fill_2 FILLER_56_640 ();
 sg13g2_decap_8 FILLER_56_652 ();
 sg13g2_decap_4 FILLER_56_659 ();
 sg13g2_fill_1 FILLER_56_663 ();
 sg13g2_decap_4 FILLER_56_672 ();
 sg13g2_fill_2 FILLER_56_715 ();
 sg13g2_decap_8 FILLER_56_735 ();
 sg13g2_fill_2 FILLER_56_742 ();
 sg13g2_fill_1 FILLER_56_744 ();
 sg13g2_decap_8 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_765 ();
 sg13g2_decap_4 FILLER_56_788 ();
 sg13g2_fill_1 FILLER_56_796 ();
 sg13g2_decap_4 FILLER_56_809 ();
 sg13g2_fill_2 FILLER_56_813 ();
 sg13g2_decap_8 FILLER_56_837 ();
 sg13g2_decap_8 FILLER_56_844 ();
 sg13g2_decap_8 FILLER_56_851 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_37 ();
 sg13g2_fill_2 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_104 ();
 sg13g2_decap_4 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_118 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_fill_1 FILLER_57_158 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_fill_2 FILLER_57_176 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_194 ();
 sg13g2_fill_1 FILLER_57_201 ();
 sg13g2_decap_4 FILLER_57_221 ();
 sg13g2_fill_2 FILLER_57_225 ();
 sg13g2_decap_4 FILLER_57_233 ();
 sg13g2_fill_2 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_274 ();
 sg13g2_decap_4 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_311 ();
 sg13g2_fill_2 FILLER_57_358 ();
 sg13g2_fill_1 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_379 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_387 ();
 sg13g2_decap_4 FILLER_57_394 ();
 sg13g2_fill_2 FILLER_57_398 ();
 sg13g2_fill_2 FILLER_57_405 ();
 sg13g2_fill_1 FILLER_57_407 ();
 sg13g2_fill_2 FILLER_57_412 ();
 sg13g2_decap_8 FILLER_57_479 ();
 sg13g2_fill_1 FILLER_57_518 ();
 sg13g2_decap_8 FILLER_57_565 ();
 sg13g2_decap_4 FILLER_57_572 ();
 sg13g2_fill_1 FILLER_57_576 ();
 sg13g2_decap_8 FILLER_57_582 ();
 sg13g2_decap_8 FILLER_57_589 ();
 sg13g2_decap_8 FILLER_57_609 ();
 sg13g2_decap_8 FILLER_57_616 ();
 sg13g2_decap_4 FILLER_57_623 ();
 sg13g2_decap_4 FILLER_57_660 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_fill_1 FILLER_57_686 ();
 sg13g2_fill_2 FILLER_57_700 ();
 sg13g2_fill_1 FILLER_57_702 ();
 sg13g2_decap_8 FILLER_57_716 ();
 sg13g2_fill_2 FILLER_57_723 ();
 sg13g2_fill_1 FILLER_57_725 ();
 sg13g2_decap_8 FILLER_57_734 ();
 sg13g2_decap_8 FILLER_57_761 ();
 sg13g2_decap_4 FILLER_57_768 ();
 sg13g2_fill_1 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_fill_2 FILLER_57_800 ();
 sg13g2_fill_1 FILLER_57_815 ();
 sg13g2_decap_8 FILLER_57_824 ();
 sg13g2_decap_8 FILLER_57_831 ();
 sg13g2_decap_8 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_40 ();
 sg13g2_fill_2 FILLER_58_88 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_168 ();
 sg13g2_fill_1 FILLER_58_170 ();
 sg13g2_fill_2 FILLER_58_181 ();
 sg13g2_fill_1 FILLER_58_183 ();
 sg13g2_decap_8 FILLER_58_188 ();
 sg13g2_decap_8 FILLER_58_195 ();
 sg13g2_fill_2 FILLER_58_202 ();
 sg13g2_fill_2 FILLER_58_228 ();
 sg13g2_decap_8 FILLER_58_234 ();
 sg13g2_decap_8 FILLER_58_241 ();
 sg13g2_decap_8 FILLER_58_248 ();
 sg13g2_decap_4 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_265 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_fill_2 FILLER_58_313 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_fill_2 FILLER_58_361 ();
 sg13g2_fill_1 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_58_390 ();
 sg13g2_fill_1 FILLER_58_397 ();
 sg13g2_fill_1 FILLER_58_414 ();
 sg13g2_decap_8 FILLER_58_441 ();
 sg13g2_decap_4 FILLER_58_456 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_decap_4 FILLER_58_470 ();
 sg13g2_fill_2 FILLER_58_492 ();
 sg13g2_decap_4 FILLER_58_516 ();
 sg13g2_fill_2 FILLER_58_537 ();
 sg13g2_fill_2 FILLER_58_562 ();
 sg13g2_fill_1 FILLER_58_564 ();
 sg13g2_decap_8 FILLER_58_592 ();
 sg13g2_decap_4 FILLER_58_599 ();
 sg13g2_fill_1 FILLER_58_603 ();
 sg13g2_fill_2 FILLER_58_608 ();
 sg13g2_fill_1 FILLER_58_610 ();
 sg13g2_decap_8 FILLER_58_619 ();
 sg13g2_decap_8 FILLER_58_626 ();
 sg13g2_decap_8 FILLER_58_633 ();
 sg13g2_fill_2 FILLER_58_640 ();
 sg13g2_fill_1 FILLER_58_642 ();
 sg13g2_fill_1 FILLER_58_648 ();
 sg13g2_decap_8 FILLER_58_657 ();
 sg13g2_fill_2 FILLER_58_664 ();
 sg13g2_fill_1 FILLER_58_666 ();
 sg13g2_decap_8 FILLER_58_675 ();
 sg13g2_decap_4 FILLER_58_682 ();
 sg13g2_fill_2 FILLER_58_686 ();
 sg13g2_decap_8 FILLER_58_693 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_717 ();
 sg13g2_decap_8 FILLER_58_724 ();
 sg13g2_decap_8 FILLER_58_731 ();
 sg13g2_fill_1 FILLER_58_738 ();
 sg13g2_fill_2 FILLER_58_749 ();
 sg13g2_fill_1 FILLER_58_751 ();
 sg13g2_decap_4 FILLER_58_760 ();
 sg13g2_decap_8 FILLER_58_772 ();
 sg13g2_fill_2 FILLER_58_779 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_12 ();
 sg13g2_decap_8 FILLER_59_17 ();
 sg13g2_decap_8 FILLER_59_24 ();
 sg13g2_decap_8 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_38 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_107 ();
 sg13g2_decap_4 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_118 ();
 sg13g2_decap_8 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_decap_4 FILLER_59_224 ();
 sg13g2_fill_2 FILLER_59_276 ();
 sg13g2_decap_8 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_315 ();
 sg13g2_decap_4 FILLER_59_346 ();
 sg13g2_fill_1 FILLER_59_366 ();
 sg13g2_fill_1 FILLER_59_405 ();
 sg13g2_fill_2 FILLER_59_442 ();
 sg13g2_fill_1 FILLER_59_476 ();
 sg13g2_fill_2 FILLER_59_494 ();
 sg13g2_fill_1 FILLER_59_505 ();
 sg13g2_fill_2 FILLER_59_520 ();
 sg13g2_fill_2 FILLER_59_540 ();
 sg13g2_fill_2 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_583 ();
 sg13g2_fill_2 FILLER_59_593 ();
 sg13g2_decap_4 FILLER_59_631 ();
 sg13g2_fill_2 FILLER_59_635 ();
 sg13g2_decap_8 FILLER_59_657 ();
 sg13g2_fill_2 FILLER_59_664 ();
 sg13g2_decap_4 FILLER_59_697 ();
 sg13g2_fill_1 FILLER_59_709 ();
 sg13g2_fill_2 FILLER_59_731 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_fill_2 FILLER_59_756 ();
 sg13g2_decap_4 FILLER_59_778 ();
 sg13g2_fill_1 FILLER_59_782 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_4 FILLER_59_810 ();
 sg13g2_fill_2 FILLER_59_814 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_31 ();
 sg13g2_fill_1 FILLER_60_33 ();
 sg13g2_decap_4 FILLER_60_51 ();
 sg13g2_fill_2 FILLER_60_55 ();
 sg13g2_decap_4 FILLER_60_79 ();
 sg13g2_fill_2 FILLER_60_83 ();
 sg13g2_fill_2 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_103 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_fill_2 FILLER_60_147 ();
 sg13g2_fill_1 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_159 ();
 sg13g2_decap_8 FILLER_60_174 ();
 sg13g2_fill_2 FILLER_60_181 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_fill_2 FILLER_60_237 ();
 sg13g2_fill_1 FILLER_60_255 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_decap_4 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_290 ();
 sg13g2_fill_2 FILLER_60_300 ();
 sg13g2_fill_1 FILLER_60_342 ();
 sg13g2_decap_8 FILLER_60_363 ();
 sg13g2_fill_2 FILLER_60_383 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_decap_4 FILLER_60_390 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_1 FILLER_60_401 ();
 sg13g2_decap_4 FILLER_60_446 ();
 sg13g2_decap_8 FILLER_60_455 ();
 sg13g2_decap_4 FILLER_60_462 ();
 sg13g2_fill_2 FILLER_60_479 ();
 sg13g2_fill_1 FILLER_60_506 ();
 sg13g2_decap_4 FILLER_60_512 ();
 sg13g2_decap_8 FILLER_60_520 ();
 sg13g2_fill_2 FILLER_60_541 ();
 sg13g2_decap_8 FILLER_60_556 ();
 sg13g2_decap_8 FILLER_60_563 ();
 sg13g2_fill_2 FILLER_60_570 ();
 sg13g2_decap_4 FILLER_60_600 ();
 sg13g2_fill_1 FILLER_60_604 ();
 sg13g2_fill_1 FILLER_60_611 ();
 sg13g2_decap_8 FILLER_60_650 ();
 sg13g2_decap_4 FILLER_60_657 ();
 sg13g2_fill_1 FILLER_60_661 ();
 sg13g2_decap_8 FILLER_60_675 ();
 sg13g2_fill_1 FILLER_60_682 ();
 sg13g2_decap_8 FILLER_60_693 ();
 sg13g2_decap_4 FILLER_60_700 ();
 sg13g2_fill_2 FILLER_60_704 ();
 sg13g2_fill_2 FILLER_60_714 ();
 sg13g2_decap_8 FILLER_60_726 ();
 sg13g2_decap_4 FILLER_60_733 ();
 sg13g2_fill_2 FILLER_60_742 ();
 sg13g2_fill_1 FILLER_60_744 ();
 sg13g2_decap_4 FILLER_60_755 ();
 sg13g2_fill_1 FILLER_60_759 ();
 sg13g2_decap_8 FILLER_60_772 ();
 sg13g2_decap_8 FILLER_60_779 ();
 sg13g2_fill_2 FILLER_60_786 ();
 sg13g2_fill_1 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_decap_8 FILLER_60_801 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_decap_8 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_836 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_34 ();
 sg13g2_decap_8 FILLER_61_72 ();
 sg13g2_decap_8 FILLER_61_83 ();
 sg13g2_decap_4 FILLER_61_90 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_fill_2 FILLER_61_100 ();
 sg13g2_decap_8 FILLER_61_110 ();
 sg13g2_decap_8 FILLER_61_117 ();
 sg13g2_decap_4 FILLER_61_124 ();
 sg13g2_decap_8 FILLER_61_137 ();
 sg13g2_decap_4 FILLER_61_144 ();
 sg13g2_fill_2 FILLER_61_176 ();
 sg13g2_fill_1 FILLER_61_178 ();
 sg13g2_fill_2 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_300 ();
 sg13g2_decap_8 FILLER_61_307 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_fill_1 FILLER_61_321 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_379 ();
 sg13g2_decap_4 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_442 ();
 sg13g2_fill_2 FILLER_61_524 ();
 sg13g2_decap_4 FILLER_61_549 ();
 sg13g2_fill_1 FILLER_61_553 ();
 sg13g2_fill_2 FILLER_61_572 ();
 sg13g2_fill_1 FILLER_61_591 ();
 sg13g2_decap_8 FILLER_61_597 ();
 sg13g2_decap_4 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_608 ();
 sg13g2_fill_1 FILLER_61_635 ();
 sg13g2_fill_2 FILLER_61_652 ();
 sg13g2_decap_8 FILLER_61_682 ();
 sg13g2_decap_8 FILLER_61_689 ();
 sg13g2_decap_8 FILLER_61_696 ();
 sg13g2_decap_4 FILLER_61_703 ();
 sg13g2_fill_1 FILLER_61_707 ();
 sg13g2_decap_4 FILLER_61_732 ();
 sg13g2_fill_2 FILLER_61_736 ();
 sg13g2_decap_8 FILLER_61_759 ();
 sg13g2_decap_8 FILLER_61_766 ();
 sg13g2_decap_8 FILLER_61_773 ();
 sg13g2_decap_8 FILLER_61_780 ();
 sg13g2_decap_8 FILLER_61_787 ();
 sg13g2_decap_8 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_801 ();
 sg13g2_decap_8 FILLER_61_808 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_8 FILLER_61_822 ();
 sg13g2_decap_8 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_843 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_decap_4 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_decap_8 FILLER_62_17 ();
 sg13g2_decap_8 FILLER_62_24 ();
 sg13g2_fill_2 FILLER_62_31 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_decap_4 FILLER_62_60 ();
 sg13g2_fill_1 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_decap_8 FILLER_62_167 ();
 sg13g2_fill_2 FILLER_62_174 ();
 sg13g2_fill_1 FILLER_62_176 ();
 sg13g2_fill_2 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_decap_4 FILLER_62_188 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_fill_1 FILLER_62_213 ();
 sg13g2_decap_8 FILLER_62_230 ();
 sg13g2_fill_2 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_258 ();
 sg13g2_fill_2 FILLER_62_270 ();
 sg13g2_decap_4 FILLER_62_300 ();
 sg13g2_decap_8 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_328 ();
 sg13g2_decap_4 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_fill_1 FILLER_62_353 ();
 sg13g2_fill_2 FILLER_62_371 ();
 sg13g2_fill_2 FILLER_62_384 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_fill_2 FILLER_62_422 ();
 sg13g2_fill_1 FILLER_62_447 ();
 sg13g2_fill_1 FILLER_62_452 ();
 sg13g2_decap_4 FILLER_62_456 ();
 sg13g2_fill_2 FILLER_62_460 ();
 sg13g2_fill_2 FILLER_62_471 ();
 sg13g2_decap_8 FILLER_62_486 ();
 sg13g2_fill_2 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_495 ();
 sg13g2_fill_2 FILLER_62_500 ();
 sg13g2_fill_2 FILLER_62_516 ();
 sg13g2_fill_1 FILLER_62_518 ();
 sg13g2_fill_2 FILLER_62_568 ();
 sg13g2_fill_1 FILLER_62_570 ();
 sg13g2_decap_8 FILLER_62_585 ();
 sg13g2_fill_2 FILLER_62_609 ();
 sg13g2_decap_8 FILLER_62_646 ();
 sg13g2_decap_4 FILLER_62_653 ();
 sg13g2_fill_2 FILLER_62_657 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_decap_8 FILLER_62_679 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_4 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_726 ();
 sg13g2_decap_8 FILLER_62_733 ();
 sg13g2_decap_8 FILLER_62_740 ();
 sg13g2_decap_8 FILLER_62_747 ();
 sg13g2_decap_8 FILLER_62_754 ();
 sg13g2_decap_8 FILLER_62_761 ();
 sg13g2_decap_8 FILLER_62_768 ();
 sg13g2_decap_8 FILLER_62_775 ();
 sg13g2_decap_8 FILLER_62_782 ();
 sg13g2_decap_8 FILLER_62_789 ();
 sg13g2_decap_8 FILLER_62_796 ();
 sg13g2_decap_8 FILLER_62_803 ();
 sg13g2_decap_8 FILLER_62_810 ();
 sg13g2_decap_8 FILLER_62_817 ();
 sg13g2_decap_8 FILLER_62_824 ();
 sg13g2_decap_8 FILLER_62_831 ();
 sg13g2_decap_8 FILLER_62_838 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_decap_8 FILLER_62_852 ();
 sg13g2_fill_2 FILLER_62_859 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_2 FILLER_63_30 ();
 sg13g2_fill_2 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_69 ();
 sg13g2_decap_8 FILLER_63_76 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_decap_4 FILLER_63_90 ();
 sg13g2_fill_1 FILLER_63_94 ();
 sg13g2_decap_8 FILLER_63_116 ();
 sg13g2_decap_8 FILLER_63_123 ();
 sg13g2_decap_4 FILLER_63_130 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_fill_2 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_153 ();
 sg13g2_decap_8 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_1 FILLER_63_258 ();
 sg13g2_decap_4 FILLER_63_269 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_278 ();
 sg13g2_decap_8 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_decap_4 FILLER_63_363 ();
 sg13g2_fill_1 FILLER_63_367 ();
 sg13g2_decap_8 FILLER_63_373 ();
 sg13g2_fill_2 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_387 ();
 sg13g2_fill_2 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_403 ();
 sg13g2_decap_4 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_445 ();
 sg13g2_decap_4 FILLER_63_451 ();
 sg13g2_fill_2 FILLER_63_455 ();
 sg13g2_fill_2 FILLER_63_496 ();
 sg13g2_fill_2 FILLER_63_566 ();
 sg13g2_decap_4 FILLER_63_578 ();
 sg13g2_fill_2 FILLER_63_600 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_675 ();
 sg13g2_decap_8 FILLER_63_682 ();
 sg13g2_decap_8 FILLER_63_689 ();
 sg13g2_decap_8 FILLER_63_696 ();
 sg13g2_decap_8 FILLER_63_703 ();
 sg13g2_decap_8 FILLER_63_710 ();
 sg13g2_decap_8 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_724 ();
 sg13g2_decap_8 FILLER_63_731 ();
 sg13g2_decap_8 FILLER_63_738 ();
 sg13g2_decap_8 FILLER_63_745 ();
 sg13g2_decap_8 FILLER_63_752 ();
 sg13g2_decap_8 FILLER_63_759 ();
 sg13g2_decap_8 FILLER_63_766 ();
 sg13g2_decap_8 FILLER_63_773 ();
 sg13g2_decap_8 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_787 ();
 sg13g2_decap_8 FILLER_63_794 ();
 sg13g2_decap_8 FILLER_63_801 ();
 sg13g2_decap_8 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_815 ();
 sg13g2_decap_8 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_829 ();
 sg13g2_decap_8 FILLER_63_836 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_decap_8 FILLER_63_850 ();
 sg13g2_decap_4 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_56 ();
 sg13g2_fill_2 FILLER_64_71 ();
 sg13g2_decap_4 FILLER_64_82 ();
 sg13g2_fill_2 FILLER_64_86 ();
 sg13g2_decap_8 FILLER_64_92 ();
 sg13g2_decap_8 FILLER_64_104 ();
 sg13g2_fill_2 FILLER_64_111 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_decap_8 FILLER_64_118 ();
 sg13g2_decap_8 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_132 ();
 sg13g2_fill_1 FILLER_64_141 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_decap_8 FILLER_64_166 ();
 sg13g2_decap_4 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_177 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_4 FILLER_64_196 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_fill_1 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_fill_2 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_249 ();
 sg13g2_decap_4 FILLER_64_256 ();
 sg13g2_fill_1 FILLER_64_260 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_fill_1 FILLER_64_273 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_337 ();
 sg13g2_decap_8 FILLER_64_344 ();
 sg13g2_fill_1 FILLER_64_351 ();
 sg13g2_fill_2 FILLER_64_365 ();
 sg13g2_decap_4 FILLER_64_373 ();
 sg13g2_fill_1 FILLER_64_377 ();
 sg13g2_fill_2 FILLER_64_405 ();
 sg13g2_fill_1 FILLER_64_407 ();
 sg13g2_fill_2 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_430 ();
 sg13g2_fill_2 FILLER_64_440 ();
 sg13g2_decap_4 FILLER_64_479 ();
 sg13g2_fill_2 FILLER_64_491 ();
 sg13g2_fill_2 FILLER_64_497 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_decap_4 FILLER_64_513 ();
 sg13g2_fill_2 FILLER_64_517 ();
 sg13g2_fill_2 FILLER_64_552 ();
 sg13g2_fill_2 FILLER_64_581 ();
 sg13g2_fill_1 FILLER_64_583 ();
 sg13g2_fill_1 FILLER_64_612 ();
 sg13g2_decap_8 FILLER_64_621 ();
 sg13g2_fill_1 FILLER_64_636 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_fill_1 FILLER_64_657 ();
 sg13g2_decap_8 FILLER_64_671 ();
 sg13g2_decap_8 FILLER_64_678 ();
 sg13g2_decap_8 FILLER_64_685 ();
 sg13g2_decap_8 FILLER_64_692 ();
 sg13g2_decap_8 FILLER_64_699 ();
 sg13g2_decap_8 FILLER_64_706 ();
 sg13g2_decap_8 FILLER_64_713 ();
 sg13g2_decap_8 FILLER_64_720 ();
 sg13g2_decap_8 FILLER_64_727 ();
 sg13g2_decap_8 FILLER_64_734 ();
 sg13g2_decap_8 FILLER_64_741 ();
 sg13g2_decap_8 FILLER_64_748 ();
 sg13g2_decap_8 FILLER_64_755 ();
 sg13g2_decap_8 FILLER_64_762 ();
 sg13g2_decap_8 FILLER_64_769 ();
 sg13g2_decap_8 FILLER_64_776 ();
 sg13g2_decap_8 FILLER_64_783 ();
 sg13g2_decap_8 FILLER_64_790 ();
 sg13g2_decap_8 FILLER_64_797 ();
 sg13g2_decap_8 FILLER_64_804 ();
 sg13g2_decap_8 FILLER_64_811 ();
 sg13g2_decap_8 FILLER_64_818 ();
 sg13g2_decap_8 FILLER_64_825 ();
 sg13g2_decap_8 FILLER_64_832 ();
 sg13g2_decap_8 FILLER_64_839 ();
 sg13g2_decap_8 FILLER_64_846 ();
 sg13g2_decap_8 FILLER_64_853 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_decap_4 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_80 ();
 sg13g2_fill_2 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_158 ();
 sg13g2_decap_4 FILLER_65_174 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_decap_4 FILLER_65_190 ();
 sg13g2_fill_1 FILLER_65_194 ();
 sg13g2_decap_8 FILLER_65_243 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_decap_4 FILLER_65_345 ();
 sg13g2_fill_2 FILLER_65_404 ();
 sg13g2_fill_2 FILLER_65_415 ();
 sg13g2_fill_1 FILLER_65_417 ();
 sg13g2_decap_8 FILLER_65_443 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_fill_2 FILLER_65_454 ();
 sg13g2_decap_4 FILLER_65_483 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_fill_2 FILLER_65_528 ();
 sg13g2_fill_1 FILLER_65_539 ();
 sg13g2_decap_8 FILLER_65_599 ();
 sg13g2_decap_8 FILLER_65_613 ();
 sg13g2_fill_1 FILLER_65_620 ();
 sg13g2_fill_1 FILLER_65_638 ();
 sg13g2_decap_8 FILLER_65_676 ();
 sg13g2_decap_8 FILLER_65_683 ();
 sg13g2_decap_8 FILLER_65_690 ();
 sg13g2_decap_8 FILLER_65_697 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_725 ();
 sg13g2_decap_8 FILLER_65_732 ();
 sg13g2_decap_8 FILLER_65_739 ();
 sg13g2_decap_8 FILLER_65_746 ();
 sg13g2_decap_8 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_2 FILLER_66_27 ();
 sg13g2_decap_4 FILLER_66_66 ();
 sg13g2_fill_1 FILLER_66_70 ();
 sg13g2_decap_4 FILLER_66_108 ();
 sg13g2_decap_8 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_166 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_4 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_241 ();
 sg13g2_decap_8 FILLER_66_247 ();
 sg13g2_fill_1 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_2 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_66_373 ();
 sg13g2_fill_2 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_418 ();
 sg13g2_decap_4 FILLER_66_445 ();
 sg13g2_fill_1 FILLER_66_463 ();
 sg13g2_fill_2 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_508 ();
 sg13g2_fill_1 FILLER_66_515 ();
 sg13g2_fill_1 FILLER_66_562 ();
 sg13g2_fill_2 FILLER_66_595 ();
 sg13g2_fill_1 FILLER_66_597 ();
 sg13g2_decap_4 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_621 ();
 sg13g2_fill_2 FILLER_66_637 ();
 sg13g2_fill_1 FILLER_66_639 ();
 sg13g2_decap_4 FILLER_66_650 ();
 sg13g2_decap_8 FILLER_66_667 ();
 sg13g2_decap_8 FILLER_66_674 ();
 sg13g2_decap_8 FILLER_66_681 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_decap_8 FILLER_66_709 ();
 sg13g2_decap_8 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_fill_1 FILLER_67_36 ();
 sg13g2_fill_2 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_58 ();
 sg13g2_decap_4 FILLER_67_69 ();
 sg13g2_fill_2 FILLER_67_86 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_126 ();
 sg13g2_decap_4 FILLER_67_156 ();
 sg13g2_decap_8 FILLER_67_173 ();
 sg13g2_fill_1 FILLER_67_184 ();
 sg13g2_decap_8 FILLER_67_193 ();
 sg13g2_decap_8 FILLER_67_200 ();
 sg13g2_decap_4 FILLER_67_207 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_fill_1 FILLER_67_233 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_268 ();
 sg13g2_fill_2 FILLER_67_278 ();
 sg13g2_fill_1 FILLER_67_280 ();
 sg13g2_decap_4 FILLER_67_290 ();
 sg13g2_decap_8 FILLER_67_320 ();
 sg13g2_decap_4 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_345 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_decap_4 FILLER_67_385 ();
 sg13g2_decap_4 FILLER_67_436 ();
 sg13g2_fill_2 FILLER_67_453 ();
 sg13g2_fill_2 FILLER_67_506 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_527 ();
 sg13g2_decap_8 FILLER_67_554 ();
 sg13g2_fill_1 FILLER_67_568 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_fill_2 FILLER_67_602 ();
 sg13g2_fill_1 FILLER_67_604 ();
 sg13g2_decap_4 FILLER_67_612 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_631 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_644 ();
 sg13g2_fill_2 FILLER_67_649 ();
 sg13g2_decap_8 FILLER_67_660 ();
 sg13g2_decap_8 FILLER_67_667 ();
 sg13g2_decap_8 FILLER_67_674 ();
 sg13g2_decap_8 FILLER_67_681 ();
 sg13g2_decap_8 FILLER_67_688 ();
 sg13g2_decap_8 FILLER_67_695 ();
 sg13g2_decap_8 FILLER_67_702 ();
 sg13g2_decap_8 FILLER_67_709 ();
 sg13g2_decap_8 FILLER_67_716 ();
 sg13g2_decap_8 FILLER_67_723 ();
 sg13g2_decap_8 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_737 ();
 sg13g2_decap_8 FILLER_67_744 ();
 sg13g2_decap_8 FILLER_67_751 ();
 sg13g2_decap_8 FILLER_67_758 ();
 sg13g2_decap_8 FILLER_67_765 ();
 sg13g2_decap_8 FILLER_67_772 ();
 sg13g2_decap_8 FILLER_67_779 ();
 sg13g2_decap_8 FILLER_67_786 ();
 sg13g2_decap_8 FILLER_67_793 ();
 sg13g2_decap_8 FILLER_67_800 ();
 sg13g2_decap_8 FILLER_67_807 ();
 sg13g2_decap_8 FILLER_67_814 ();
 sg13g2_decap_8 FILLER_67_821 ();
 sg13g2_decap_8 FILLER_67_828 ();
 sg13g2_decap_8 FILLER_67_835 ();
 sg13g2_decap_8 FILLER_67_842 ();
 sg13g2_decap_8 FILLER_67_849 ();
 sg13g2_decap_4 FILLER_67_856 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_decap_4 FILLER_68_60 ();
 sg13g2_fill_2 FILLER_68_104 ();
 sg13g2_fill_2 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_254 ();
 sg13g2_decap_8 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_decap_8 FILLER_68_344 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_decap_8 FILLER_68_366 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_decap_4 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_426 ();
 sg13g2_decap_8 FILLER_68_433 ();
 sg13g2_decap_4 FILLER_68_440 ();
 sg13g2_decap_4 FILLER_68_471 ();
 sg13g2_fill_2 FILLER_68_511 ();
 sg13g2_fill_1 FILLER_68_513 ();
 sg13g2_decap_8 FILLER_68_527 ();
 sg13g2_fill_2 FILLER_68_547 ();
 sg13g2_fill_1 FILLER_68_566 ();
 sg13g2_decap_8 FILLER_68_631 ();
 sg13g2_fill_2 FILLER_68_638 ();
 sg13g2_decap_8 FILLER_68_668 ();
 sg13g2_decap_8 FILLER_68_675 ();
 sg13g2_decap_8 FILLER_68_682 ();
 sg13g2_decap_8 FILLER_68_689 ();
 sg13g2_decap_8 FILLER_68_696 ();
 sg13g2_decap_8 FILLER_68_703 ();
 sg13g2_decap_8 FILLER_68_710 ();
 sg13g2_decap_8 FILLER_68_717 ();
 sg13g2_decap_8 FILLER_68_724 ();
 sg13g2_decap_8 FILLER_68_731 ();
 sg13g2_decap_8 FILLER_68_738 ();
 sg13g2_decap_8 FILLER_68_745 ();
 sg13g2_decap_8 FILLER_68_752 ();
 sg13g2_decap_8 FILLER_68_759 ();
 sg13g2_decap_8 FILLER_68_766 ();
 sg13g2_decap_8 FILLER_68_773 ();
 sg13g2_decap_8 FILLER_68_780 ();
 sg13g2_decap_8 FILLER_68_787 ();
 sg13g2_decap_8 FILLER_68_794 ();
 sg13g2_decap_8 FILLER_68_801 ();
 sg13g2_decap_8 FILLER_68_808 ();
 sg13g2_decap_8 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_decap_8 FILLER_68_829 ();
 sg13g2_decap_8 FILLER_68_836 ();
 sg13g2_decap_8 FILLER_68_843 ();
 sg13g2_decap_8 FILLER_68_850 ();
 sg13g2_decap_4 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_7 ();
 sg13g2_decap_4 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_85 ();
 sg13g2_fill_2 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_118 ();
 sg13g2_fill_1 FILLER_69_120 ();
 sg13g2_fill_2 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_182 ();
 sg13g2_fill_1 FILLER_69_184 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_fill_2 FILLER_69_228 ();
 sg13g2_decap_4 FILLER_69_244 ();
 sg13g2_fill_2 FILLER_69_248 ();
 sg13g2_decap_4 FILLER_69_290 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_fill_2 FILLER_69_305 ();
 sg13g2_fill_1 FILLER_69_307 ();
 sg13g2_decap_8 FILLER_69_321 ();
 sg13g2_decap_4 FILLER_69_328 ();
 sg13g2_fill_2 FILLER_69_332 ();
 sg13g2_decap_4 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_382 ();
 sg13g2_fill_2 FILLER_69_389 ();
 sg13g2_fill_2 FILLER_69_401 ();
 sg13g2_fill_2 FILLER_69_412 ();
 sg13g2_decap_4 FILLER_69_444 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_decap_8 FILLER_69_453 ();
 sg13g2_decap_4 FILLER_69_460 ();
 sg13g2_fill_2 FILLER_69_464 ();
 sg13g2_decap_8 FILLER_69_489 ();
 sg13g2_decap_4 FILLER_69_505 ();
 sg13g2_fill_1 FILLER_69_509 ();
 sg13g2_fill_2 FILLER_69_537 ();
 sg13g2_fill_1 FILLER_69_539 ();
 sg13g2_fill_2 FILLER_69_546 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_decap_4 FILLER_69_603 ();
 sg13g2_decap_8 FILLER_69_612 ();
 sg13g2_decap_8 FILLER_69_647 ();
 sg13g2_decap_8 FILLER_69_654 ();
 sg13g2_decap_8 FILLER_69_661 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_decap_8 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_682 ();
 sg13g2_decap_8 FILLER_69_689 ();
 sg13g2_decap_8 FILLER_69_696 ();
 sg13g2_decap_8 FILLER_69_703 ();
 sg13g2_decap_8 FILLER_69_710 ();
 sg13g2_decap_8 FILLER_69_717 ();
 sg13g2_decap_8 FILLER_69_724 ();
 sg13g2_decap_8 FILLER_69_731 ();
 sg13g2_decap_8 FILLER_69_738 ();
 sg13g2_decap_8 FILLER_69_745 ();
 sg13g2_decap_8 FILLER_69_752 ();
 sg13g2_decap_8 FILLER_69_759 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_780 ();
 sg13g2_decap_8 FILLER_69_787 ();
 sg13g2_decap_8 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_801 ();
 sg13g2_decap_8 FILLER_69_808 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_4 FILLER_69_857 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_46 ();
 sg13g2_fill_2 FILLER_70_50 ();
 sg13g2_decap_8 FILLER_70_89 ();
 sg13g2_decap_4 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_157 ();
 sg13g2_fill_2 FILLER_70_171 ();
 sg13g2_fill_2 FILLER_70_186 ();
 sg13g2_fill_2 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_204 ();
 sg13g2_fill_2 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_2 FILLER_70_246 ();
 sg13g2_fill_1 FILLER_70_248 ();
 sg13g2_fill_2 FILLER_70_306 ();
 sg13g2_fill_2 FILLER_70_348 ();
 sg13g2_fill_1 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_decap_4 FILLER_70_390 ();
 sg13g2_fill_2 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_70_473 ();
 sg13g2_fill_2 FILLER_70_520 ();
 sg13g2_fill_2 FILLER_70_531 ();
 sg13g2_fill_1 FILLER_70_574 ();
 sg13g2_fill_2 FILLER_70_584 ();
 sg13g2_fill_1 FILLER_70_586 ();
 sg13g2_decap_8 FILLER_70_598 ();
 sg13g2_decap_8 FILLER_70_605 ();
 sg13g2_decap_8 FILLER_70_612 ();
 sg13g2_fill_1 FILLER_70_632 ();
 sg13g2_decap_8 FILLER_70_642 ();
 sg13g2_decap_8 FILLER_70_649 ();
 sg13g2_decap_8 FILLER_70_656 ();
 sg13g2_decap_8 FILLER_70_663 ();
 sg13g2_decap_8 FILLER_70_670 ();
 sg13g2_decap_8 FILLER_70_677 ();
 sg13g2_decap_8 FILLER_70_684 ();
 sg13g2_decap_8 FILLER_70_691 ();
 sg13g2_decap_8 FILLER_70_698 ();
 sg13g2_decap_8 FILLER_70_705 ();
 sg13g2_decap_8 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_719 ();
 sg13g2_decap_8 FILLER_70_726 ();
 sg13g2_decap_8 FILLER_70_733 ();
 sg13g2_decap_8 FILLER_70_740 ();
 sg13g2_decap_8 FILLER_70_747 ();
 sg13g2_decap_8 FILLER_70_754 ();
 sg13g2_decap_8 FILLER_70_761 ();
 sg13g2_decap_8 FILLER_70_768 ();
 sg13g2_decap_8 FILLER_70_775 ();
 sg13g2_decap_8 FILLER_70_782 ();
 sg13g2_decap_8 FILLER_70_789 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_817 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_2 FILLER_71_27 ();
 sg13g2_decap_4 FILLER_71_47 ();
 sg13g2_fill_2 FILLER_71_51 ();
 sg13g2_fill_2 FILLER_71_85 ();
 sg13g2_fill_1 FILLER_71_87 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_197 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_237 ();
 sg13g2_fill_1 FILLER_71_265 ();
 sg13g2_fill_2 FILLER_71_285 ();
 sg13g2_fill_1 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_325 ();
 sg13g2_fill_1 FILLER_71_332 ();
 sg13g2_fill_1 FILLER_71_355 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_466 ();
 sg13g2_fill_2 FILLER_71_486 ();
 sg13g2_fill_1 FILLER_71_488 ();
 sg13g2_fill_1 FILLER_71_517 ();
 sg13g2_fill_1 FILLER_71_550 ();
 sg13g2_fill_2 FILLER_71_578 ();
 sg13g2_fill_1 FILLER_71_580 ();
 sg13g2_decap_8 FILLER_71_587 ();
 sg13g2_decap_8 FILLER_71_594 ();
 sg13g2_decap_8 FILLER_71_601 ();
 sg13g2_decap_8 FILLER_71_608 ();
 sg13g2_decap_8 FILLER_71_615 ();
 sg13g2_decap_8 FILLER_71_622 ();
 sg13g2_decap_8 FILLER_71_629 ();
 sg13g2_decap_8 FILLER_71_636 ();
 sg13g2_decap_8 FILLER_71_643 ();
 sg13g2_decap_8 FILLER_71_650 ();
 sg13g2_decap_8 FILLER_71_657 ();
 sg13g2_decap_8 FILLER_71_664 ();
 sg13g2_decap_8 FILLER_71_671 ();
 sg13g2_decap_8 FILLER_71_678 ();
 sg13g2_decap_8 FILLER_71_685 ();
 sg13g2_decap_8 FILLER_71_692 ();
 sg13g2_decap_8 FILLER_71_699 ();
 sg13g2_decap_8 FILLER_71_706 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_decap_8 FILLER_71_720 ();
 sg13g2_decap_8 FILLER_71_727 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_8 FILLER_71_748 ();
 sg13g2_decap_8 FILLER_71_755 ();
 sg13g2_decap_8 FILLER_71_762 ();
 sg13g2_decap_8 FILLER_71_769 ();
 sg13g2_decap_8 FILLER_71_776 ();
 sg13g2_decap_8 FILLER_71_783 ();
 sg13g2_decap_8 FILLER_71_790 ();
 sg13g2_decap_8 FILLER_71_797 ();
 sg13g2_decap_8 FILLER_71_804 ();
 sg13g2_decap_8 FILLER_71_811 ();
 sg13g2_decap_8 FILLER_71_818 ();
 sg13g2_decap_8 FILLER_71_825 ();
 sg13g2_decap_8 FILLER_71_832 ();
 sg13g2_decap_8 FILLER_71_839 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_fill_2 FILLER_72_37 ();
 sg13g2_fill_1 FILLER_72_39 ();
 sg13g2_decap_4 FILLER_72_61 ();
 sg13g2_fill_1 FILLER_72_65 ();
 sg13g2_decap_8 FILLER_72_194 ();
 sg13g2_fill_2 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_220 ();
 sg13g2_fill_1 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_1 FILLER_72_283 ();
 sg13g2_fill_2 FILLER_72_290 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_fill_2 FILLER_72_321 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_decap_4 FILLER_72_345 ();
 sg13g2_fill_1 FILLER_72_349 ();
 sg13g2_fill_2 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_388 ();
 sg13g2_fill_1 FILLER_72_390 ();
 sg13g2_fill_2 FILLER_72_446 ();
 sg13g2_fill_2 FILLER_72_496 ();
 sg13g2_decap_8 FILLER_72_507 ();
 sg13g2_decap_4 FILLER_72_514 ();
 sg13g2_fill_2 FILLER_72_518 ();
 sg13g2_fill_2 FILLER_72_524 ();
 sg13g2_fill_1 FILLER_72_526 ();
 sg13g2_decap_8 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_583 ();
 sg13g2_decap_8 FILLER_72_590 ();
 sg13g2_decap_8 FILLER_72_597 ();
 sg13g2_decap_8 FILLER_72_604 ();
 sg13g2_decap_8 FILLER_72_611 ();
 sg13g2_decap_8 FILLER_72_618 ();
 sg13g2_decap_8 FILLER_72_625 ();
 sg13g2_decap_8 FILLER_72_632 ();
 sg13g2_decap_8 FILLER_72_639 ();
 sg13g2_decap_8 FILLER_72_646 ();
 sg13g2_decap_8 FILLER_72_653 ();
 sg13g2_decap_8 FILLER_72_660 ();
 sg13g2_decap_8 FILLER_72_667 ();
 sg13g2_decap_8 FILLER_72_674 ();
 sg13g2_decap_8 FILLER_72_681 ();
 sg13g2_decap_8 FILLER_72_688 ();
 sg13g2_decap_8 FILLER_72_695 ();
 sg13g2_decap_8 FILLER_72_702 ();
 sg13g2_decap_8 FILLER_72_709 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_decap_8 FILLER_72_723 ();
 sg13g2_decap_8 FILLER_72_730 ();
 sg13g2_decap_8 FILLER_72_737 ();
 sg13g2_decap_8 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_758 ();
 sg13g2_decap_8 FILLER_72_765 ();
 sg13g2_decap_8 FILLER_72_772 ();
 sg13g2_decap_8 FILLER_72_779 ();
 sg13g2_decap_8 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_793 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_4 FILLER_72_856 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_63 ();
 sg13g2_fill_1 FILLER_73_74 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_fill_1 FILLER_73_90 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_115 ();
 sg13g2_fill_1 FILLER_73_117 ();
 sg13g2_decap_4 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_148 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_4 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_2 FILLER_73_239 ();
 sg13g2_decap_8 FILLER_73_264 ();
 sg13g2_fill_2 FILLER_73_288 ();
 sg13g2_decap_4 FILLER_73_295 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_fill_2 FILLER_73_322 ();
 sg13g2_fill_1 FILLER_73_324 ();
 sg13g2_fill_1 FILLER_73_348 ();
 sg13g2_decap_4 FILLER_73_373 ();
 sg13g2_fill_2 FILLER_73_377 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_fill_1 FILLER_73_468 ();
 sg13g2_fill_1 FILLER_73_478 ();
 sg13g2_decap_8 FILLER_73_493 ();
 sg13g2_fill_2 FILLER_73_500 ();
 sg13g2_fill_1 FILLER_73_502 ();
 sg13g2_fill_2 FILLER_73_534 ();
 sg13g2_decap_8 FILLER_73_563 ();
 sg13g2_decap_8 FILLER_73_570 ();
 sg13g2_decap_8 FILLER_73_577 ();
 sg13g2_decap_8 FILLER_73_584 ();
 sg13g2_decap_8 FILLER_73_591 ();
 sg13g2_decap_8 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_605 ();
 sg13g2_decap_8 FILLER_73_612 ();
 sg13g2_decap_8 FILLER_73_619 ();
 sg13g2_decap_8 FILLER_73_626 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_682 ();
 sg13g2_decap_8 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_710 ();
 sg13g2_decap_8 FILLER_73_717 ();
 sg13g2_decap_8 FILLER_73_724 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_32 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_152 ();
 sg13g2_fill_2 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_262 ();
 sg13g2_decap_4 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_273 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_decap_8 FILLER_74_302 ();
 sg13g2_fill_1 FILLER_74_309 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_decap_4 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_332 ();
 sg13g2_decap_8 FILLER_74_341 ();
 sg13g2_decap_8 FILLER_74_348 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_fill_2 FILLER_74_371 ();
 sg13g2_fill_1 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_4 FILLER_74_445 ();
 sg13g2_fill_2 FILLER_74_449 ();
 sg13g2_fill_2 FILLER_74_460 ();
 sg13g2_fill_1 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_520 ();
 sg13g2_decap_8 FILLER_74_549 ();
 sg13g2_decap_8 FILLER_74_556 ();
 sg13g2_decap_8 FILLER_74_563 ();
 sg13g2_decap_8 FILLER_74_570 ();
 sg13g2_decap_8 FILLER_74_577 ();
 sg13g2_decap_8 FILLER_74_584 ();
 sg13g2_decap_8 FILLER_74_591 ();
 sg13g2_decap_8 FILLER_74_598 ();
 sg13g2_decap_8 FILLER_74_605 ();
 sg13g2_decap_8 FILLER_74_612 ();
 sg13g2_decap_8 FILLER_74_619 ();
 sg13g2_decap_8 FILLER_74_626 ();
 sg13g2_decap_8 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_640 ();
 sg13g2_decap_8 FILLER_74_647 ();
 sg13g2_decap_8 FILLER_74_654 ();
 sg13g2_decap_8 FILLER_74_661 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_decap_8 FILLER_74_675 ();
 sg13g2_decap_8 FILLER_74_682 ();
 sg13g2_decap_8 FILLER_74_689 ();
 sg13g2_decap_8 FILLER_74_696 ();
 sg13g2_decap_8 FILLER_74_703 ();
 sg13g2_decap_8 FILLER_74_710 ();
 sg13g2_decap_8 FILLER_74_717 ();
 sg13g2_decap_8 FILLER_74_724 ();
 sg13g2_decap_8 FILLER_74_731 ();
 sg13g2_decap_8 FILLER_74_738 ();
 sg13g2_decap_8 FILLER_74_745 ();
 sg13g2_decap_8 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_759 ();
 sg13g2_decap_8 FILLER_74_766 ();
 sg13g2_decap_8 FILLER_74_773 ();
 sg13g2_decap_8 FILLER_74_780 ();
 sg13g2_decap_8 FILLER_74_787 ();
 sg13g2_decap_8 FILLER_74_794 ();
 sg13g2_decap_8 FILLER_74_801 ();
 sg13g2_decap_8 FILLER_74_808 ();
 sg13g2_decap_8 FILLER_74_815 ();
 sg13g2_decap_8 FILLER_74_822 ();
 sg13g2_decap_8 FILLER_74_829 ();
 sg13g2_decap_8 FILLER_74_836 ();
 sg13g2_decap_8 FILLER_74_843 ();
 sg13g2_decap_8 FILLER_74_850 ();
 sg13g2_decap_4 FILLER_74_857 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_4 FILLER_75_27 ();
 sg13g2_fill_1 FILLER_75_31 ();
 sg13g2_fill_1 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_136 ();
 sg13g2_fill_1 FILLER_75_173 ();
 sg13g2_fill_2 FILLER_75_211 ();
 sg13g2_fill_2 FILLER_75_219 ();
 sg13g2_fill_1 FILLER_75_221 ();
 sg13g2_fill_2 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_229 ();
 sg13g2_decap_4 FILLER_75_263 ();
 sg13g2_fill_2 FILLER_75_267 ();
 sg13g2_decap_4 FILLER_75_304 ();
 sg13g2_decap_4 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_384 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_fill_2 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_417 ();
 sg13g2_decap_4 FILLER_75_423 ();
 sg13g2_fill_2 FILLER_75_427 ();
 sg13g2_decap_4 FILLER_75_456 ();
 sg13g2_decap_8 FILLER_75_487 ();
 sg13g2_decap_8 FILLER_75_494 ();
 sg13g2_decap_8 FILLER_75_501 ();
 sg13g2_decap_8 FILLER_75_508 ();
 sg13g2_decap_8 FILLER_75_515 ();
 sg13g2_decap_8 FILLER_75_522 ();
 sg13g2_decap_8 FILLER_75_529 ();
 sg13g2_decap_4 FILLER_75_536 ();
 sg13g2_fill_1 FILLER_75_540 ();
 sg13g2_decap_8 FILLER_75_545 ();
 sg13g2_decap_8 FILLER_75_552 ();
 sg13g2_decap_8 FILLER_75_559 ();
 sg13g2_decap_8 FILLER_75_566 ();
 sg13g2_decap_8 FILLER_75_573 ();
 sg13g2_decap_8 FILLER_75_580 ();
 sg13g2_decap_8 FILLER_75_587 ();
 sg13g2_decap_8 FILLER_75_594 ();
 sg13g2_decap_8 FILLER_75_601 ();
 sg13g2_decap_8 FILLER_75_608 ();
 sg13g2_decap_8 FILLER_75_615 ();
 sg13g2_decap_8 FILLER_75_622 ();
 sg13g2_decap_8 FILLER_75_629 ();
 sg13g2_decap_8 FILLER_75_636 ();
 sg13g2_decap_8 FILLER_75_643 ();
 sg13g2_decap_8 FILLER_75_650 ();
 sg13g2_decap_8 FILLER_75_657 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_692 ();
 sg13g2_decap_8 FILLER_75_699 ();
 sg13g2_decap_8 FILLER_75_706 ();
 sg13g2_decap_8 FILLER_75_713 ();
 sg13g2_decap_8 FILLER_75_720 ();
 sg13g2_decap_8 FILLER_75_727 ();
 sg13g2_decap_8 FILLER_75_734 ();
 sg13g2_decap_8 FILLER_75_741 ();
 sg13g2_decap_8 FILLER_75_748 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_decap_8 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_776 ();
 sg13g2_decap_8 FILLER_75_783 ();
 sg13g2_decap_8 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_811 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_25 ();
 sg13g2_fill_2 FILLER_76_124 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_fill_2 FILLER_76_192 ();
 sg13g2_fill_2 FILLER_76_203 ();
 sg13g2_decap_4 FILLER_76_223 ();
 sg13g2_fill_2 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_2 FILLER_76_251 ();
 sg13g2_fill_1 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_269 ();
 sg13g2_fill_1 FILLER_76_271 ();
 sg13g2_decap_8 FILLER_76_283 ();
 sg13g2_fill_1 FILLER_76_290 ();
 sg13g2_fill_1 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_318 ();
 sg13g2_decap_8 FILLER_76_363 ();
 sg13g2_fill_1 FILLER_76_370 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_398 ();
 sg13g2_decap_8 FILLER_76_405 ();
 sg13g2_decap_8 FILLER_76_412 ();
 sg13g2_decap_8 FILLER_76_435 ();
 sg13g2_decap_8 FILLER_76_442 ();
 sg13g2_decap_8 FILLER_76_449 ();
 sg13g2_decap_4 FILLER_76_456 ();
 sg13g2_decap_8 FILLER_76_473 ();
 sg13g2_decap_8 FILLER_76_480 ();
 sg13g2_decap_8 FILLER_76_487 ();
 sg13g2_decap_8 FILLER_76_494 ();
 sg13g2_decap_8 FILLER_76_501 ();
 sg13g2_decap_8 FILLER_76_508 ();
 sg13g2_decap_8 FILLER_76_515 ();
 sg13g2_decap_8 FILLER_76_522 ();
 sg13g2_decap_8 FILLER_76_529 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_8 FILLER_76_550 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_decap_8 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_8 FILLER_76_599 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_decap_8 FILLER_76_655 ();
 sg13g2_decap_8 FILLER_76_662 ();
 sg13g2_decap_8 FILLER_76_669 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_8 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_774 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_8 FILLER_76_788 ();
 sg13g2_decap_8 FILLER_76_795 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_4 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_40 ();
 sg13g2_fill_2 FILLER_77_72 ();
 sg13g2_fill_2 FILLER_77_131 ();
 sg13g2_fill_2 FILLER_77_148 ();
 sg13g2_fill_1 FILLER_77_160 ();
 sg13g2_decap_4 FILLER_77_223 ();
 sg13g2_fill_2 FILLER_77_253 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_fill_2 FILLER_77_261 ();
 sg13g2_fill_1 FILLER_77_263 ();
 sg13g2_fill_2 FILLER_77_276 ();
 sg13g2_fill_2 FILLER_77_312 ();
 sg13g2_fill_2 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_decap_8 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_77_414 ();
 sg13g2_decap_8 FILLER_77_421 ();
 sg13g2_decap_8 FILLER_77_428 ();
 sg13g2_decap_8 FILLER_77_435 ();
 sg13g2_decap_8 FILLER_77_442 ();
 sg13g2_decap_8 FILLER_77_449 ();
 sg13g2_decap_8 FILLER_77_456 ();
 sg13g2_decap_8 FILLER_77_463 ();
 sg13g2_decap_8 FILLER_77_470 ();
 sg13g2_decap_8 FILLER_77_477 ();
 sg13g2_decap_8 FILLER_77_484 ();
 sg13g2_decap_8 FILLER_77_491 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_decap_8 FILLER_77_505 ();
 sg13g2_decap_8 FILLER_77_512 ();
 sg13g2_decap_8 FILLER_77_519 ();
 sg13g2_decap_8 FILLER_77_526 ();
 sg13g2_decap_8 FILLER_77_533 ();
 sg13g2_decap_8 FILLER_77_540 ();
 sg13g2_decap_8 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_554 ();
 sg13g2_decap_8 FILLER_77_561 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_decap_8 FILLER_77_575 ();
 sg13g2_decap_8 FILLER_77_582 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_decap_8 FILLER_77_631 ();
 sg13g2_decap_8 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_722 ();
 sg13g2_decap_8 FILLER_77_729 ();
 sg13g2_decap_8 FILLER_77_736 ();
 sg13g2_decap_8 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_fill_1 FILLER_78_21 ();
 sg13g2_fill_1 FILLER_78_96 ();
 sg13g2_fill_1 FILLER_78_119 ();
 sg13g2_fill_2 FILLER_78_165 ();
 sg13g2_fill_2 FILLER_78_332 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_363 ();
 sg13g2_fill_2 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_379 ();
 sg13g2_fill_2 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_8 FILLER_78_404 ();
 sg13g2_decap_8 FILLER_78_411 ();
 sg13g2_decap_8 FILLER_78_418 ();
 sg13g2_decap_8 FILLER_78_425 ();
 sg13g2_decap_8 FILLER_78_432 ();
 sg13g2_decap_8 FILLER_78_439 ();
 sg13g2_decap_8 FILLER_78_446 ();
 sg13g2_decap_8 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_460 ();
 sg13g2_decap_8 FILLER_78_467 ();
 sg13g2_decap_8 FILLER_78_474 ();
 sg13g2_decap_8 FILLER_78_481 ();
 sg13g2_decap_8 FILLER_78_488 ();
 sg13g2_decap_8 FILLER_78_495 ();
 sg13g2_decap_8 FILLER_78_502 ();
 sg13g2_decap_8 FILLER_78_509 ();
 sg13g2_decap_8 FILLER_78_516 ();
 sg13g2_decap_8 FILLER_78_523 ();
 sg13g2_decap_8 FILLER_78_530 ();
 sg13g2_decap_8 FILLER_78_537 ();
 sg13g2_decap_8 FILLER_78_544 ();
 sg13g2_decap_8 FILLER_78_551 ();
 sg13g2_decap_8 FILLER_78_558 ();
 sg13g2_decap_8 FILLER_78_565 ();
 sg13g2_decap_8 FILLER_78_572 ();
 sg13g2_decap_8 FILLER_78_579 ();
 sg13g2_decap_8 FILLER_78_586 ();
 sg13g2_decap_8 FILLER_78_593 ();
 sg13g2_decap_8 FILLER_78_600 ();
 sg13g2_decap_8 FILLER_78_607 ();
 sg13g2_decap_8 FILLER_78_614 ();
 sg13g2_decap_8 FILLER_78_621 ();
 sg13g2_decap_8 FILLER_78_628 ();
 sg13g2_decap_8 FILLER_78_635 ();
 sg13g2_decap_8 FILLER_78_642 ();
 sg13g2_decap_8 FILLER_78_649 ();
 sg13g2_decap_8 FILLER_78_656 ();
 sg13g2_decap_8 FILLER_78_663 ();
 sg13g2_decap_8 FILLER_78_670 ();
 sg13g2_decap_8 FILLER_78_677 ();
 sg13g2_decap_8 FILLER_78_684 ();
 sg13g2_decap_8 FILLER_78_691 ();
 sg13g2_decap_8 FILLER_78_698 ();
 sg13g2_decap_8 FILLER_78_705 ();
 sg13g2_decap_8 FILLER_78_712 ();
 sg13g2_decap_8 FILLER_78_719 ();
 sg13g2_decap_8 FILLER_78_726 ();
 sg13g2_decap_8 FILLER_78_733 ();
 sg13g2_decap_8 FILLER_78_740 ();
 sg13g2_decap_8 FILLER_78_747 ();
 sg13g2_decap_8 FILLER_78_754 ();
 sg13g2_decap_8 FILLER_78_761 ();
 sg13g2_decap_8 FILLER_78_768 ();
 sg13g2_decap_8 FILLER_78_775 ();
 sg13g2_decap_8 FILLER_78_782 ();
 sg13g2_decap_8 FILLER_78_789 ();
 sg13g2_decap_8 FILLER_78_796 ();
 sg13g2_decap_8 FILLER_78_803 ();
 sg13g2_decap_8 FILLER_78_810 ();
 sg13g2_decap_8 FILLER_78_817 ();
 sg13g2_decap_8 FILLER_78_824 ();
 sg13g2_decap_8 FILLER_78_831 ();
 sg13g2_decap_8 FILLER_78_838 ();
 sg13g2_decap_8 FILLER_78_845 ();
 sg13g2_decap_8 FILLER_78_852 ();
 sg13g2_fill_2 FILLER_78_859 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_61 ();
 sg13g2_fill_2 FILLER_79_71 ();
 sg13g2_fill_2 FILLER_79_151 ();
 sg13g2_fill_2 FILLER_79_198 ();
 sg13g2_fill_1 FILLER_79_209 ();
 sg13g2_decap_4 FILLER_79_246 ();
 sg13g2_decap_8 FILLER_79_277 ();
 sg13g2_fill_1 FILLER_79_284 ();
 sg13g2_fill_2 FILLER_79_301 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_decap_8 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_79_415 ();
 sg13g2_decap_8 FILLER_79_422 ();
 sg13g2_decap_8 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_79_436 ();
 sg13g2_decap_8 FILLER_79_443 ();
 sg13g2_decap_8 FILLER_79_450 ();
 sg13g2_decap_8 FILLER_79_457 ();
 sg13g2_decap_8 FILLER_79_464 ();
 sg13g2_decap_8 FILLER_79_471 ();
 sg13g2_decap_8 FILLER_79_478 ();
 sg13g2_decap_8 FILLER_79_485 ();
 sg13g2_decap_8 FILLER_79_492 ();
 sg13g2_decap_8 FILLER_79_499 ();
 sg13g2_decap_8 FILLER_79_506 ();
 sg13g2_decap_8 FILLER_79_513 ();
 sg13g2_decap_8 FILLER_79_520 ();
 sg13g2_decap_8 FILLER_79_527 ();
 sg13g2_decap_8 FILLER_79_534 ();
 sg13g2_decap_8 FILLER_79_541 ();
 sg13g2_decap_8 FILLER_79_548 ();
 sg13g2_decap_8 FILLER_79_555 ();
 sg13g2_decap_8 FILLER_79_562 ();
 sg13g2_decap_8 FILLER_79_569 ();
 sg13g2_decap_8 FILLER_79_576 ();
 sg13g2_decap_8 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_590 ();
 sg13g2_decap_8 FILLER_79_597 ();
 sg13g2_decap_8 FILLER_79_604 ();
 sg13g2_decap_8 FILLER_79_611 ();
 sg13g2_decap_8 FILLER_79_618 ();
 sg13g2_decap_8 FILLER_79_625 ();
 sg13g2_decap_8 FILLER_79_632 ();
 sg13g2_decap_8 FILLER_79_639 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_decap_8 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_660 ();
 sg13g2_decap_8 FILLER_79_667 ();
 sg13g2_decap_8 FILLER_79_674 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_709 ();
 sg13g2_decap_8 FILLER_79_716 ();
 sg13g2_decap_8 FILLER_79_723 ();
 sg13g2_decap_8 FILLER_79_730 ();
 sg13g2_decap_8 FILLER_79_737 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_decap_8 FILLER_79_758 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_4 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_18 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_2 FILLER_80_177 ();
 sg13g2_fill_2 FILLER_80_188 ();
 sg13g2_fill_2 FILLER_80_217 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_fill_2 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_fill_2 FILLER_80_275 ();
 sg13g2_fill_2 FILLER_80_314 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_527 ();
 sg13g2_decap_8 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule
