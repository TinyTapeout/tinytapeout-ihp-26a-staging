module tt_um_vga_tetris (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire clknet_leaf_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire vga_hs;
 wire \vga_tetris._inputs_io_downButtonActive ;
 wire \vga_tetris._inputs_io_leftButtonActive ;
 wire \vga_tetris._inputs_io_rightButtonActive ;
 wire \vga_tetris._inputs_io_rotateButtonActive ;
 wire \vga_tetris._tetrisDisplay_io_boardYCoord[0] ;
 wire \vga_tetris._tetrisDisplay_io_boardYCoord[1] ;
 wire \vga_tetris._tetrisLogic_io_gameOver ;
 wire \vga_tetris._tetrisLogic_io_score_0[0] ;
 wire \vga_tetris._tetrisLogic_io_score_0[1] ;
 wire \vga_tetris._tetrisLogic_io_score_0[2] ;
 wire \vga_tetris._tetrisLogic_io_score_0[3] ;
 wire \vga_tetris._tetrisLogic_io_score_1[0] ;
 wire \vga_tetris._tetrisLogic_io_score_1[1] ;
 wire \vga_tetris._tetrisLogic_io_score_1[2] ;
 wire \vga_tetris._tetrisLogic_io_score_1[3] ;
 wire \vga_tetris._tetrisLogic_io_score_2[0] ;
 wire \vga_tetris._tetrisLogic_io_score_2[1] ;
 wire \vga_tetris._tetrisLogic_io_score_2[2] ;
 wire \vga_tetris._tetrisLogic_io_score_2[3] ;
 wire \vga_tetris._tetrisLogic_io_score_3[0] ;
 wire \vga_tetris._tetrisLogic_io_score_3[1] ;
 wire \vga_tetris._tetrisLogic_io_score_3[2] ;
 wire \vga_tetris._tetrisLogic_io_score_3[3] ;
 wire \vga_tetris._vgaController_io_pixelPosX[0] ;
 wire \vga_tetris._vgaController_io_pixelPosX[1] ;
 wire \vga_tetris._vgaController_io_pixelPosX[2] ;
 wire \vga_tetris._vgaController_io_pixelPosX[3] ;
 wire \vga_tetris._vgaController_io_pixelPosX[4] ;
 wire \vga_tetris._vgaController_io_pixelPosX[5] ;
 wire \vga_tetris._vgaController_io_pixelPosX[6] ;
 wire \vga_tetris._vgaController_io_pixelPosX[7] ;
 wire \vga_tetris._vgaController_io_pixelPosX[8] ;
 wire \vga_tetris._vgaController_io_pixelPosX[9] ;
 wire \vga_tetris._vgaController_io_pixelPosY[0] ;
 wire \vga_tetris._vgaController_io_pixelPosY[1] ;
 wire \vga_tetris._vgaController_io_pixelPosY[2] ;
 wire \vga_tetris._vgaController_io_pixelPosY[3] ;
 wire \vga_tetris._vgaController_io_pixelPosY[6] ;
 wire \vga_tetris._vgaController_io_pixelPosY[7] ;
 wire \vga_tetris._vgaController_io_pixelPosY[8] ;
 wire \vga_tetris._vgaController_io_pixelPosY[9] ;
 wire \vga_tetris._vgaController_io_vSync ;
 wire \vga_tetris.boardMem.board_0[0] ;
 wire \vga_tetris.boardMem.board_0[10] ;
 wire \vga_tetris.boardMem.board_0[11] ;
 wire \vga_tetris.boardMem.board_0[12] ;
 wire \vga_tetris.boardMem.board_0[13] ;
 wire \vga_tetris.boardMem.board_0[14] ;
 wire \vga_tetris.boardMem.board_0[15] ;
 wire \vga_tetris.boardMem.board_0[16] ;
 wire \vga_tetris.boardMem.board_0[17] ;
 wire \vga_tetris.boardMem.board_0[18] ;
 wire \vga_tetris.boardMem.board_0[19] ;
 wire \vga_tetris.boardMem.board_0[1] ;
 wire \vga_tetris.boardMem.board_0[2] ;
 wire \vga_tetris.boardMem.board_0[3] ;
 wire \vga_tetris.boardMem.board_0[4] ;
 wire \vga_tetris.boardMem.board_0[5] ;
 wire \vga_tetris.boardMem.board_0[6] ;
 wire \vga_tetris.boardMem.board_0[7] ;
 wire \vga_tetris.boardMem.board_0[8] ;
 wire \vga_tetris.boardMem.board_0[9] ;
 wire \vga_tetris.boardMem.board_10[0] ;
 wire \vga_tetris.boardMem.board_10[10] ;
 wire \vga_tetris.boardMem.board_10[11] ;
 wire \vga_tetris.boardMem.board_10[12] ;
 wire \vga_tetris.boardMem.board_10[13] ;
 wire \vga_tetris.boardMem.board_10[14] ;
 wire \vga_tetris.boardMem.board_10[15] ;
 wire \vga_tetris.boardMem.board_10[16] ;
 wire \vga_tetris.boardMem.board_10[17] ;
 wire \vga_tetris.boardMem.board_10[18] ;
 wire \vga_tetris.boardMem.board_10[19] ;
 wire \vga_tetris.boardMem.board_10[1] ;
 wire \vga_tetris.boardMem.board_10[2] ;
 wire \vga_tetris.boardMem.board_10[3] ;
 wire \vga_tetris.boardMem.board_10[4] ;
 wire \vga_tetris.boardMem.board_10[5] ;
 wire \vga_tetris.boardMem.board_10[6] ;
 wire \vga_tetris.boardMem.board_10[7] ;
 wire \vga_tetris.boardMem.board_10[8] ;
 wire \vga_tetris.boardMem.board_10[9] ;
 wire \vga_tetris.boardMem.board_11[0] ;
 wire \vga_tetris.boardMem.board_11[10] ;
 wire \vga_tetris.boardMem.board_11[11] ;
 wire \vga_tetris.boardMem.board_11[12] ;
 wire \vga_tetris.boardMem.board_11[13] ;
 wire \vga_tetris.boardMem.board_11[14] ;
 wire \vga_tetris.boardMem.board_11[15] ;
 wire \vga_tetris.boardMem.board_11[16] ;
 wire \vga_tetris.boardMem.board_11[17] ;
 wire \vga_tetris.boardMem.board_11[18] ;
 wire \vga_tetris.boardMem.board_11[19] ;
 wire \vga_tetris.boardMem.board_11[1] ;
 wire \vga_tetris.boardMem.board_11[2] ;
 wire \vga_tetris.boardMem.board_11[3] ;
 wire \vga_tetris.boardMem.board_11[4] ;
 wire \vga_tetris.boardMem.board_11[5] ;
 wire \vga_tetris.boardMem.board_11[6] ;
 wire \vga_tetris.boardMem.board_11[7] ;
 wire \vga_tetris.boardMem.board_11[8] ;
 wire \vga_tetris.boardMem.board_11[9] ;
 wire \vga_tetris.boardMem.board_12[0] ;
 wire \vga_tetris.boardMem.board_12[10] ;
 wire \vga_tetris.boardMem.board_12[11] ;
 wire \vga_tetris.boardMem.board_12[12] ;
 wire \vga_tetris.boardMem.board_12[13] ;
 wire \vga_tetris.boardMem.board_12[14] ;
 wire \vga_tetris.boardMem.board_12[15] ;
 wire \vga_tetris.boardMem.board_12[16] ;
 wire \vga_tetris.boardMem.board_12[17] ;
 wire \vga_tetris.boardMem.board_12[18] ;
 wire \vga_tetris.boardMem.board_12[19] ;
 wire \vga_tetris.boardMem.board_12[1] ;
 wire \vga_tetris.boardMem.board_12[2] ;
 wire \vga_tetris.boardMem.board_12[3] ;
 wire \vga_tetris.boardMem.board_12[4] ;
 wire \vga_tetris.boardMem.board_12[5] ;
 wire \vga_tetris.boardMem.board_12[6] ;
 wire \vga_tetris.boardMem.board_12[7] ;
 wire \vga_tetris.boardMem.board_12[8] ;
 wire \vga_tetris.boardMem.board_12[9] ;
 wire \vga_tetris.boardMem.board_13[0] ;
 wire \vga_tetris.boardMem.board_13[10] ;
 wire \vga_tetris.boardMem.board_13[11] ;
 wire \vga_tetris.boardMem.board_13[12] ;
 wire \vga_tetris.boardMem.board_13[13] ;
 wire \vga_tetris.boardMem.board_13[14] ;
 wire \vga_tetris.boardMem.board_13[15] ;
 wire \vga_tetris.boardMem.board_13[16] ;
 wire \vga_tetris.boardMem.board_13[17] ;
 wire \vga_tetris.boardMem.board_13[18] ;
 wire \vga_tetris.boardMem.board_13[19] ;
 wire \vga_tetris.boardMem.board_13[1] ;
 wire \vga_tetris.boardMem.board_13[2] ;
 wire \vga_tetris.boardMem.board_13[3] ;
 wire \vga_tetris.boardMem.board_13[4] ;
 wire \vga_tetris.boardMem.board_13[5] ;
 wire \vga_tetris.boardMem.board_13[6] ;
 wire \vga_tetris.boardMem.board_13[7] ;
 wire \vga_tetris.boardMem.board_13[8] ;
 wire \vga_tetris.boardMem.board_13[9] ;
 wire \vga_tetris.boardMem.board_14[0] ;
 wire \vga_tetris.boardMem.board_14[10] ;
 wire \vga_tetris.boardMem.board_14[11] ;
 wire \vga_tetris.boardMem.board_14[12] ;
 wire \vga_tetris.boardMem.board_14[13] ;
 wire \vga_tetris.boardMem.board_14[14] ;
 wire \vga_tetris.boardMem.board_14[15] ;
 wire \vga_tetris.boardMem.board_14[16] ;
 wire \vga_tetris.boardMem.board_14[17] ;
 wire \vga_tetris.boardMem.board_14[18] ;
 wire \vga_tetris.boardMem.board_14[19] ;
 wire \vga_tetris.boardMem.board_14[1] ;
 wire \vga_tetris.boardMem.board_14[2] ;
 wire \vga_tetris.boardMem.board_14[3] ;
 wire \vga_tetris.boardMem.board_14[4] ;
 wire \vga_tetris.boardMem.board_14[5] ;
 wire \vga_tetris.boardMem.board_14[6] ;
 wire \vga_tetris.boardMem.board_14[7] ;
 wire \vga_tetris.boardMem.board_14[8] ;
 wire \vga_tetris.boardMem.board_14[9] ;
 wire \vga_tetris.boardMem.board_15[0] ;
 wire \vga_tetris.boardMem.board_15[10] ;
 wire \vga_tetris.boardMem.board_15[11] ;
 wire \vga_tetris.boardMem.board_15[12] ;
 wire \vga_tetris.boardMem.board_15[13] ;
 wire \vga_tetris.boardMem.board_15[14] ;
 wire \vga_tetris.boardMem.board_15[15] ;
 wire \vga_tetris.boardMem.board_15[16] ;
 wire \vga_tetris.boardMem.board_15[17] ;
 wire \vga_tetris.boardMem.board_15[18] ;
 wire \vga_tetris.boardMem.board_15[19] ;
 wire \vga_tetris.boardMem.board_15[1] ;
 wire \vga_tetris.boardMem.board_15[2] ;
 wire \vga_tetris.boardMem.board_15[3] ;
 wire \vga_tetris.boardMem.board_15[4] ;
 wire \vga_tetris.boardMem.board_15[5] ;
 wire \vga_tetris.boardMem.board_15[6] ;
 wire \vga_tetris.boardMem.board_15[7] ;
 wire \vga_tetris.boardMem.board_15[8] ;
 wire \vga_tetris.boardMem.board_15[9] ;
 wire \vga_tetris.boardMem.board_16[0] ;
 wire \vga_tetris.boardMem.board_16[10] ;
 wire \vga_tetris.boardMem.board_16[11] ;
 wire \vga_tetris.boardMem.board_16[12] ;
 wire \vga_tetris.boardMem.board_16[13] ;
 wire \vga_tetris.boardMem.board_16[14] ;
 wire \vga_tetris.boardMem.board_16[15] ;
 wire \vga_tetris.boardMem.board_16[16] ;
 wire \vga_tetris.boardMem.board_16[17] ;
 wire \vga_tetris.boardMem.board_16[18] ;
 wire \vga_tetris.boardMem.board_16[19] ;
 wire \vga_tetris.boardMem.board_16[1] ;
 wire \vga_tetris.boardMem.board_16[2] ;
 wire \vga_tetris.boardMem.board_16[3] ;
 wire \vga_tetris.boardMem.board_16[4] ;
 wire \vga_tetris.boardMem.board_16[5] ;
 wire \vga_tetris.boardMem.board_16[6] ;
 wire \vga_tetris.boardMem.board_16[7] ;
 wire \vga_tetris.boardMem.board_16[8] ;
 wire \vga_tetris.boardMem.board_16[9] ;
 wire \vga_tetris.boardMem.board_17[0] ;
 wire \vga_tetris.boardMem.board_17[10] ;
 wire \vga_tetris.boardMem.board_17[11] ;
 wire \vga_tetris.boardMem.board_17[12] ;
 wire \vga_tetris.boardMem.board_17[13] ;
 wire \vga_tetris.boardMem.board_17[14] ;
 wire \vga_tetris.boardMem.board_17[15] ;
 wire \vga_tetris.boardMem.board_17[16] ;
 wire \vga_tetris.boardMem.board_17[17] ;
 wire \vga_tetris.boardMem.board_17[18] ;
 wire \vga_tetris.boardMem.board_17[19] ;
 wire \vga_tetris.boardMem.board_17[1] ;
 wire \vga_tetris.boardMem.board_17[2] ;
 wire \vga_tetris.boardMem.board_17[3] ;
 wire \vga_tetris.boardMem.board_17[4] ;
 wire \vga_tetris.boardMem.board_17[5] ;
 wire \vga_tetris.boardMem.board_17[6] ;
 wire \vga_tetris.boardMem.board_17[7] ;
 wire \vga_tetris.boardMem.board_17[8] ;
 wire \vga_tetris.boardMem.board_17[9] ;
 wire \vga_tetris.boardMem.board_18[0] ;
 wire \vga_tetris.boardMem.board_18[10] ;
 wire \vga_tetris.boardMem.board_18[11] ;
 wire \vga_tetris.boardMem.board_18[12] ;
 wire \vga_tetris.boardMem.board_18[13] ;
 wire \vga_tetris.boardMem.board_18[14] ;
 wire \vga_tetris.boardMem.board_18[15] ;
 wire \vga_tetris.boardMem.board_18[16] ;
 wire \vga_tetris.boardMem.board_18[17] ;
 wire \vga_tetris.boardMem.board_18[18] ;
 wire \vga_tetris.boardMem.board_18[19] ;
 wire \vga_tetris.boardMem.board_18[1] ;
 wire \vga_tetris.boardMem.board_18[2] ;
 wire \vga_tetris.boardMem.board_18[3] ;
 wire \vga_tetris.boardMem.board_18[4] ;
 wire \vga_tetris.boardMem.board_18[5] ;
 wire \vga_tetris.boardMem.board_18[6] ;
 wire \vga_tetris.boardMem.board_18[7] ;
 wire \vga_tetris.boardMem.board_18[8] ;
 wire \vga_tetris.boardMem.board_18[9] ;
 wire \vga_tetris.boardMem.board_19[0] ;
 wire \vga_tetris.boardMem.board_19[10] ;
 wire \vga_tetris.boardMem.board_19[11] ;
 wire \vga_tetris.boardMem.board_19[12] ;
 wire \vga_tetris.boardMem.board_19[13] ;
 wire \vga_tetris.boardMem.board_19[14] ;
 wire \vga_tetris.boardMem.board_19[15] ;
 wire \vga_tetris.boardMem.board_19[16] ;
 wire \vga_tetris.boardMem.board_19[17] ;
 wire \vga_tetris.boardMem.board_19[18] ;
 wire \vga_tetris.boardMem.board_19[19] ;
 wire \vga_tetris.boardMem.board_19[1] ;
 wire \vga_tetris.boardMem.board_19[2] ;
 wire \vga_tetris.boardMem.board_19[3] ;
 wire \vga_tetris.boardMem.board_19[4] ;
 wire \vga_tetris.boardMem.board_19[5] ;
 wire \vga_tetris.boardMem.board_19[6] ;
 wire \vga_tetris.boardMem.board_19[7] ;
 wire \vga_tetris.boardMem.board_19[8] ;
 wire \vga_tetris.boardMem.board_19[9] ;
 wire \vga_tetris.boardMem.board_1[0] ;
 wire \vga_tetris.boardMem.board_1[10] ;
 wire \vga_tetris.boardMem.board_1[11] ;
 wire \vga_tetris.boardMem.board_1[12] ;
 wire \vga_tetris.boardMem.board_1[13] ;
 wire \vga_tetris.boardMem.board_1[14] ;
 wire \vga_tetris.boardMem.board_1[15] ;
 wire \vga_tetris.boardMem.board_1[16] ;
 wire \vga_tetris.boardMem.board_1[17] ;
 wire \vga_tetris.boardMem.board_1[18] ;
 wire \vga_tetris.boardMem.board_1[19] ;
 wire \vga_tetris.boardMem.board_1[1] ;
 wire \vga_tetris.boardMem.board_1[2] ;
 wire \vga_tetris.boardMem.board_1[3] ;
 wire \vga_tetris.boardMem.board_1[4] ;
 wire \vga_tetris.boardMem.board_1[5] ;
 wire \vga_tetris.boardMem.board_1[6] ;
 wire \vga_tetris.boardMem.board_1[7] ;
 wire \vga_tetris.boardMem.board_1[8] ;
 wire \vga_tetris.boardMem.board_1[9] ;
 wire \vga_tetris.boardMem.board_2[0] ;
 wire \vga_tetris.boardMem.board_2[10] ;
 wire \vga_tetris.boardMem.board_2[11] ;
 wire \vga_tetris.boardMem.board_2[12] ;
 wire \vga_tetris.boardMem.board_2[13] ;
 wire \vga_tetris.boardMem.board_2[14] ;
 wire \vga_tetris.boardMem.board_2[15] ;
 wire \vga_tetris.boardMem.board_2[16] ;
 wire \vga_tetris.boardMem.board_2[17] ;
 wire \vga_tetris.boardMem.board_2[18] ;
 wire \vga_tetris.boardMem.board_2[19] ;
 wire \vga_tetris.boardMem.board_2[1] ;
 wire \vga_tetris.boardMem.board_2[2] ;
 wire \vga_tetris.boardMem.board_2[3] ;
 wire \vga_tetris.boardMem.board_2[4] ;
 wire \vga_tetris.boardMem.board_2[5] ;
 wire \vga_tetris.boardMem.board_2[6] ;
 wire \vga_tetris.boardMem.board_2[7] ;
 wire \vga_tetris.boardMem.board_2[8] ;
 wire \vga_tetris.boardMem.board_2[9] ;
 wire \vga_tetris.boardMem.board_3[0] ;
 wire \vga_tetris.boardMem.board_3[10] ;
 wire \vga_tetris.boardMem.board_3[11] ;
 wire \vga_tetris.boardMem.board_3[12] ;
 wire \vga_tetris.boardMem.board_3[13] ;
 wire \vga_tetris.boardMem.board_3[14] ;
 wire \vga_tetris.boardMem.board_3[15] ;
 wire \vga_tetris.boardMem.board_3[16] ;
 wire \vga_tetris.boardMem.board_3[17] ;
 wire \vga_tetris.boardMem.board_3[18] ;
 wire \vga_tetris.boardMem.board_3[19] ;
 wire \vga_tetris.boardMem.board_3[1] ;
 wire \vga_tetris.boardMem.board_3[2] ;
 wire \vga_tetris.boardMem.board_3[3] ;
 wire \vga_tetris.boardMem.board_3[4] ;
 wire \vga_tetris.boardMem.board_3[5] ;
 wire \vga_tetris.boardMem.board_3[6] ;
 wire \vga_tetris.boardMem.board_3[7] ;
 wire \vga_tetris.boardMem.board_3[8] ;
 wire \vga_tetris.boardMem.board_3[9] ;
 wire \vga_tetris.boardMem.board_4[0] ;
 wire \vga_tetris.boardMem.board_4[10] ;
 wire \vga_tetris.boardMem.board_4[11] ;
 wire \vga_tetris.boardMem.board_4[12] ;
 wire \vga_tetris.boardMem.board_4[13] ;
 wire \vga_tetris.boardMem.board_4[14] ;
 wire \vga_tetris.boardMem.board_4[15] ;
 wire \vga_tetris.boardMem.board_4[16] ;
 wire \vga_tetris.boardMem.board_4[17] ;
 wire \vga_tetris.boardMem.board_4[18] ;
 wire \vga_tetris.boardMem.board_4[19] ;
 wire \vga_tetris.boardMem.board_4[1] ;
 wire \vga_tetris.boardMem.board_4[2] ;
 wire \vga_tetris.boardMem.board_4[3] ;
 wire \vga_tetris.boardMem.board_4[4] ;
 wire \vga_tetris.boardMem.board_4[5] ;
 wire \vga_tetris.boardMem.board_4[6] ;
 wire \vga_tetris.boardMem.board_4[7] ;
 wire \vga_tetris.boardMem.board_4[8] ;
 wire \vga_tetris.boardMem.board_4[9] ;
 wire \vga_tetris.boardMem.board_5[0] ;
 wire \vga_tetris.boardMem.board_5[10] ;
 wire \vga_tetris.boardMem.board_5[11] ;
 wire \vga_tetris.boardMem.board_5[12] ;
 wire \vga_tetris.boardMem.board_5[13] ;
 wire \vga_tetris.boardMem.board_5[14] ;
 wire \vga_tetris.boardMem.board_5[15] ;
 wire \vga_tetris.boardMem.board_5[16] ;
 wire \vga_tetris.boardMem.board_5[17] ;
 wire \vga_tetris.boardMem.board_5[18] ;
 wire \vga_tetris.boardMem.board_5[19] ;
 wire \vga_tetris.boardMem.board_5[1] ;
 wire \vga_tetris.boardMem.board_5[2] ;
 wire \vga_tetris.boardMem.board_5[3] ;
 wire \vga_tetris.boardMem.board_5[4] ;
 wire \vga_tetris.boardMem.board_5[5] ;
 wire \vga_tetris.boardMem.board_5[6] ;
 wire \vga_tetris.boardMem.board_5[7] ;
 wire \vga_tetris.boardMem.board_5[8] ;
 wire \vga_tetris.boardMem.board_5[9] ;
 wire \vga_tetris.boardMem.board_6[0] ;
 wire \vga_tetris.boardMem.board_6[10] ;
 wire \vga_tetris.boardMem.board_6[11] ;
 wire \vga_tetris.boardMem.board_6[12] ;
 wire \vga_tetris.boardMem.board_6[13] ;
 wire \vga_tetris.boardMem.board_6[14] ;
 wire \vga_tetris.boardMem.board_6[15] ;
 wire \vga_tetris.boardMem.board_6[16] ;
 wire \vga_tetris.boardMem.board_6[17] ;
 wire \vga_tetris.boardMem.board_6[18] ;
 wire \vga_tetris.boardMem.board_6[19] ;
 wire \vga_tetris.boardMem.board_6[1] ;
 wire \vga_tetris.boardMem.board_6[2] ;
 wire \vga_tetris.boardMem.board_6[3] ;
 wire \vga_tetris.boardMem.board_6[4] ;
 wire \vga_tetris.boardMem.board_6[5] ;
 wire \vga_tetris.boardMem.board_6[6] ;
 wire \vga_tetris.boardMem.board_6[7] ;
 wire \vga_tetris.boardMem.board_6[8] ;
 wire \vga_tetris.boardMem.board_6[9] ;
 wire \vga_tetris.boardMem.board_7[0] ;
 wire \vga_tetris.boardMem.board_7[10] ;
 wire \vga_tetris.boardMem.board_7[11] ;
 wire \vga_tetris.boardMem.board_7[12] ;
 wire \vga_tetris.boardMem.board_7[13] ;
 wire \vga_tetris.boardMem.board_7[14] ;
 wire \vga_tetris.boardMem.board_7[15] ;
 wire \vga_tetris.boardMem.board_7[16] ;
 wire \vga_tetris.boardMem.board_7[17] ;
 wire \vga_tetris.boardMem.board_7[18] ;
 wire \vga_tetris.boardMem.board_7[19] ;
 wire \vga_tetris.boardMem.board_7[1] ;
 wire \vga_tetris.boardMem.board_7[2] ;
 wire \vga_tetris.boardMem.board_7[3] ;
 wire \vga_tetris.boardMem.board_7[4] ;
 wire \vga_tetris.boardMem.board_7[5] ;
 wire \vga_tetris.boardMem.board_7[6] ;
 wire \vga_tetris.boardMem.board_7[7] ;
 wire \vga_tetris.boardMem.board_7[8] ;
 wire \vga_tetris.boardMem.board_7[9] ;
 wire \vga_tetris.boardMem.board_8[0] ;
 wire \vga_tetris.boardMem.board_8[10] ;
 wire \vga_tetris.boardMem.board_8[11] ;
 wire \vga_tetris.boardMem.board_8[12] ;
 wire \vga_tetris.boardMem.board_8[13] ;
 wire \vga_tetris.boardMem.board_8[14] ;
 wire \vga_tetris.boardMem.board_8[15] ;
 wire \vga_tetris.boardMem.board_8[16] ;
 wire \vga_tetris.boardMem.board_8[17] ;
 wire \vga_tetris.boardMem.board_8[18] ;
 wire \vga_tetris.boardMem.board_8[19] ;
 wire \vga_tetris.boardMem.board_8[1] ;
 wire \vga_tetris.boardMem.board_8[2] ;
 wire \vga_tetris.boardMem.board_8[3] ;
 wire \vga_tetris.boardMem.board_8[4] ;
 wire \vga_tetris.boardMem.board_8[5] ;
 wire \vga_tetris.boardMem.board_8[6] ;
 wire \vga_tetris.boardMem.board_8[7] ;
 wire \vga_tetris.boardMem.board_8[8] ;
 wire \vga_tetris.boardMem.board_8[9] ;
 wire \vga_tetris.boardMem.board_9[0] ;
 wire \vga_tetris.boardMem.board_9[10] ;
 wire \vga_tetris.boardMem.board_9[11] ;
 wire \vga_tetris.boardMem.board_9[12] ;
 wire \vga_tetris.boardMem.board_9[13] ;
 wire \vga_tetris.boardMem.board_9[14] ;
 wire \vga_tetris.boardMem.board_9[15] ;
 wire \vga_tetris.boardMem.board_9[16] ;
 wire \vga_tetris.boardMem.board_9[17] ;
 wire \vga_tetris.boardMem.board_9[18] ;
 wire \vga_tetris.boardMem.board_9[19] ;
 wire \vga_tetris.boardMem.board_9[1] ;
 wire \vga_tetris.boardMem.board_9[2] ;
 wire \vga_tetris.boardMem.board_9[3] ;
 wire \vga_tetris.boardMem.board_9[4] ;
 wire \vga_tetris.boardMem.board_9[5] ;
 wire \vga_tetris.boardMem.board_9[6] ;
 wire \vga_tetris.boardMem.board_9[7] ;
 wire \vga_tetris.boardMem.board_9[8] ;
 wire \vga_tetris.boardMem.board_9[9] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[7] ;
 wire \vga_tetris.msTimer.msTimerQ[0] ;
 wire \vga_tetris.msTimer.msTimerQ[10] ;
 wire \vga_tetris.msTimer.msTimerQ[11] ;
 wire \vga_tetris.msTimer.msTimerQ[12] ;
 wire \vga_tetris.msTimer.msTimerQ[13] ;
 wire \vga_tetris.msTimer.msTimerQ[14] ;
 wire \vga_tetris.msTimer.msTimerQ[1] ;
 wire \vga_tetris.msTimer.msTimerQ[2] ;
 wire \vga_tetris.msTimer.msTimerQ[3] ;
 wire \vga_tetris.msTimer.msTimerQ[4] ;
 wire \vga_tetris.msTimer.msTimerQ[5] ;
 wire \vga_tetris.msTimer.msTimerQ[6] ;
 wire \vga_tetris.msTimer.msTimerQ[7] ;
 wire \vga_tetris.msTimer.msTimerQ[8] ;
 wire \vga_tetris.msTimer.msTimerQ[9] ;
 wire \vga_tetris.runningTetrisLogicQ ;
 wire \vga_tetris.startTetrisLogicQ ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_done ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ;
 wire \vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ;
 wire \vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ;
 wire \vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ;
 wire \vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[2] ;
 wire \vga_tetris.tetrisLogic.gameOverResetHappenedQ ;
 wire \vga_tetris.tetrisLogic.rotationQ[0] ;
 wire \vga_tetris.tetrisLogic.rotationQ[1] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[0] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[1] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[2] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[3] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[4] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[5] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ;
 wire \vga_tetris.tetrisLogic.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.stateQ[2] ;
 wire \vga_tetris.tetrisLogic.stateQ[3] ;
 wire \vga_tetris.tetrisLogic.stateQ[4] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[0] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[1] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[2] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[3] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[4] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[5] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[6] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[7] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[8] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[9] ;
 wire \vga_tetris.vgaController.verticalCounterQ[0] ;
 wire \vga_tetris.vgaController.verticalCounterQ[1] ;
 wire \vga_tetris.vgaController.verticalCounterQ[2] ;
 wire \vga_tetris.vgaController.verticalCounterQ[3] ;
 wire \vga_tetris.vgaController.verticalCounterQ[4] ;
 wire \vga_tetris.vgaController.verticalCounterQ[5] ;
 wire \vga_tetris.vgaController.verticalCounterQ[6] ;
 wire \vga_tetris.vgaController.verticalCounterQ[7] ;
 wire \vga_tetris.vgaController.verticalCounterQ[8] ;
 wire \vga_tetris.vgaController.verticalCounterQ[9] ;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;

 sg13g2_inv_2 _3575_ (.Y(_0625_),
    .A(net1657));
 sg13g2_inv_1 _3576_ (.Y(_0626_),
    .A(net1757));
 sg13g2_inv_4 _3577_ (.A(net1907),
    .Y(_0627_));
 sg13g2_inv_2 _3578_ (.Y(_0628_),
    .A(net1809));
 sg13g2_inv_4 _3579_ (.A(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .Y(_0629_));
 sg13g2_inv_1 _3580_ (.Y(_0630_),
    .A(net1853));
 sg13g2_inv_1 _3581_ (.Y(_0631_),
    .A(net1690));
 sg13g2_inv_1 _3582_ (.Y(_0632_),
    .A(net1599));
 sg13g2_inv_1 _3583_ (.Y(_0633_),
    .A(net1279));
 sg13g2_inv_1 _3584_ (.Y(_0634_),
    .A(net1384));
 sg13g2_inv_1 _3585_ (.Y(_0635_),
    .A(net1287));
 sg13g2_inv_1 _3586_ (.Y(_0636_),
    .A(net1369));
 sg13g2_inv_1 _3587_ (.Y(_0637_),
    .A(net1383));
 sg13g2_inv_1 _3588_ (.Y(_0638_),
    .A(net756));
 sg13g2_inv_1 _3589_ (.Y(_0639_),
    .A(net1302));
 sg13g2_inv_1 _3590_ (.Y(_0640_),
    .A(net821));
 sg13g2_inv_1 _3591_ (.Y(_0641_),
    .A(net818));
 sg13g2_inv_2 _3592_ (.Y(_0642_),
    .A(net1583));
 sg13g2_inv_1 _3593_ (.Y(_0643_),
    .A(net1729));
 sg13g2_inv_1 _3594_ (.Y(_0644_),
    .A(net1605));
 sg13g2_inv_1 _3595_ (.Y(_0645_),
    .A(net1688));
 sg13g2_inv_1 _3596_ (.Y(_0646_),
    .A(net1285));
 sg13g2_inv_1 _3597_ (.Y(_0647_),
    .A(net1700));
 sg13g2_inv_1 _3598_ (.Y(_0648_),
    .A(net1445));
 sg13g2_inv_1 _3599_ (.Y(_0649_),
    .A(net1631));
 sg13g2_inv_1 _3600_ (.Y(_0650_),
    .A(net1524));
 sg13g2_inv_1 _3601_ (.Y(_0651_),
    .A(net1378));
 sg13g2_inv_1 _3602_ (.Y(_0652_),
    .A(net1367));
 sg13g2_inv_1 _3603_ (.Y(_0653_),
    .A(net1410));
 sg13g2_inv_1 _3604_ (.Y(_0654_),
    .A(net1399));
 sg13g2_inv_1 _3605_ (.Y(_0655_),
    .A(net1353));
 sg13g2_inv_1 _3606_ (.Y(_0656_),
    .A(net1331));
 sg13g2_inv_1 _3607_ (.Y(_0657_),
    .A(net1618));
 sg13g2_inv_1 _3608_ (.Y(_0658_),
    .A(net1610));
 sg13g2_inv_1 _3609_ (.Y(_0659_),
    .A(net1233));
 sg13g2_inv_2 _3610_ (.Y(_0660_),
    .A(net1843));
 sg13g2_inv_2 _3611_ (.Y(_0661_),
    .A(net1236));
 sg13g2_inv_2 _3612_ (.Y(_0662_),
    .A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ));
 sg13g2_inv_1 _3613_ (.Y(_0663_),
    .A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ));
 sg13g2_inv_2 _3614_ (.Y(_0664_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ));
 sg13g2_inv_2 _3615_ (.Y(_0665_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ));
 sg13g2_inv_2 _3616_ (.Y(_0666_),
    .A(net1376));
 sg13g2_inv_1 _3617_ (.Y(_0667_),
    .A(net1242));
 sg13g2_inv_2 _3618_ (.Y(_0668_),
    .A(\vga_tetris.tetrisLogic.stateQ[0] ));
 sg13g2_inv_1 _3619_ (.Y(_0669_),
    .A(net1811));
 sg13g2_inv_2 _3620_ (.Y(_0670_),
    .A(net1827));
 sg13g2_inv_1 _3621_ (.Y(_0671_),
    .A(net1896));
 sg13g2_inv_1 _3622_ (.Y(_0672_),
    .A(net1206));
 sg13g2_inv_1 _3623_ (.Y(_0673_),
    .A(net1501));
 sg13g2_inv_1 _3624_ (.Y(_0674_),
    .A(net1537));
 sg13g2_inv_1 _3625_ (.Y(_0675_),
    .A(net1594));
 sg13g2_inv_1 _3626_ (.Y(_0676_),
    .A(net1407));
 sg13g2_inv_1 _3627_ (.Y(_0677_),
    .A(\vga_tetris.boardMem.board_0[4] ));
 sg13g2_inv_1 _3628_ (.Y(_0678_),
    .A(\vga_tetris.boardMem.board_0[5] ));
 sg13g2_inv_1 _3629_ (.Y(_0679_),
    .A(\vga_tetris.boardMem.board_0[6] ));
 sg13g2_inv_1 _3630_ (.Y(_0680_),
    .A(\vga_tetris.boardMem.board_0[7] ));
 sg13g2_inv_1 _3631_ (.Y(_0681_),
    .A(net1527));
 sg13g2_inv_1 _3632_ (.Y(_0682_),
    .A(net1489));
 sg13g2_inv_1 _3633_ (.Y(_0683_),
    .A(net1920));
 sg13g2_inv_1 _3634_ (.Y(_0684_),
    .A(\vga_tetris.boardMem.board_0[11] ));
 sg13g2_inv_1 _3635_ (.Y(_0685_),
    .A(\vga_tetris.boardMem.board_0[12] ));
 sg13g2_inv_1 _3636_ (.Y(_0686_),
    .A(net1546));
 sg13g2_inv_1 _3637_ (.Y(_0687_),
    .A(net1539));
 sg13g2_inv_1 _3638_ (.Y(_0688_),
    .A(net1421));
 sg13g2_inv_1 _3639_ (.Y(_0689_),
    .A(\vga_tetris.boardMem.board_0[16] ));
 sg13g2_inv_1 _3640_ (.Y(_0690_),
    .A(\vga_tetris.boardMem.board_0[17] ));
 sg13g2_inv_1 _3641_ (.Y(_0691_),
    .A(\vga_tetris.boardMem.board_0[18] ));
 sg13g2_inv_1 _3642_ (.Y(_0692_),
    .A(\vga_tetris.boardMem.board_0[19] ));
 sg13g2_inv_1 _3643_ (.Y(_0693_),
    .A(\vga_tetris.msTimer.msTimerQ[2] ));
 sg13g2_inv_1 _3644_ (.Y(_0694_),
    .A(\vga_tetris.msTimer.msTimerQ[5] ));
 sg13g2_inv_1 _3645_ (.Y(_0695_),
    .A(net1871));
 sg13g2_inv_1 _3646_ (.Y(_0696_),
    .A(\vga_tetris.inputs.buttonTimerQ_2[3] ));
 sg13g2_inv_1 _3647_ (.Y(_0697_),
    .A(\vga_tetris.inputs.buttonTimerQ_2[2] ));
 sg13g2_inv_1 _3648_ (.Y(_0698_),
    .A(net1635));
 sg13g2_inv_2 _3649_ (.Y(_0699_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ));
 sg13g2_inv_4 _3650_ (.A(net1239),
    .Y(_0700_));
 sg13g2_inv_2 _3651_ (.Y(_0701_),
    .A(net1231));
 sg13g2_inv_1 _3652_ (.Y(_0702_),
    .A(net1692));
 sg13g2_inv_1 _3653_ (.Y(_0703_),
    .A(net1260));
 sg13g2_inv_1 _3654_ (.Y(_0704_),
    .A(net1798));
 sg13g2_inv_1 _3655_ (.Y(_0705_),
    .A(net1867));
 sg13g2_inv_1 _3656_ (.Y(_0706_),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ));
 sg13g2_inv_1 _3657_ (.Y(_0707_),
    .A(\vga_tetris._tetrisLogic_io_score_3[1] ));
 sg13g2_inv_1 _3658_ (.Y(_0708_),
    .A(net1453));
 sg13g2_inv_1 _3659_ (.Y(_0709_),
    .A(net1784));
 sg13g2_inv_1 _3660_ (.Y(_0710_),
    .A(net1404));
 sg13g2_inv_1 _3661_ (.Y(_0711_),
    .A(net1773));
 sg13g2_inv_1 _3662_ (.Y(_0712_),
    .A(net1858));
 sg13g2_inv_1 _3663_ (.Y(_0713_),
    .A(net1791));
 sg13g2_inv_2 _3664_ (.Y(_0714_),
    .A(net1762));
 sg13g2_or2_1 _3665_ (.X(_0715_),
    .B(net1208),
    .A(\vga_tetris._vgaController_io_pixelPosY[7] ));
 sg13g2_nand2_2 _3666_ (.Y(_0716_),
    .A(net1757),
    .B(net1208));
 sg13g2_a21o_1 _3667_ (.A2(_0716_),
    .A1(_0715_),
    .B1(net1205),
    .X(_0717_));
 sg13g2_nor2b_2 _3668_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .Y(_0718_));
 sg13g2_nor2b_2 _3669_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B_N(_0718_),
    .Y(_0719_));
 sg13g2_nand2b_2 _3670_ (.Y(_0720_),
    .B(_0718_),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ));
 sg13g2_nor2b_2 _3671_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .Y(_0721_));
 sg13g2_inv_2 _3672_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_and2_1 _3673_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0721_),
    .X(_0723_));
 sg13g2_nand2_2 _3674_ (.Y(_0724_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0721_));
 sg13g2_nor2_1 _3675_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_a21oi_1 _3676_ (.A1(_0670_),
    .A2(_0724_),
    .Y(_0726_),
    .B1(_0725_));
 sg13g2_nor2b_1 _3677_ (.A(net1233),
    .B_N(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0727_));
 sg13g2_nand3b_1 _3678_ (.B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .C(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0728_),
    .A_N(net1233));
 sg13g2_nand2_2 _3679_ (.Y(_0729_),
    .A(net1241),
    .B(_0668_));
 sg13g2_nor2_1 _3680_ (.A(_0728_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_or2_1 _3681_ (.X(_0731_),
    .B(_0729_),
    .A(_0728_));
 sg13g2_a21oi_1 _3682_ (.A1(_0643_),
    .A2(net1193),
    .Y(_0732_),
    .B1(net1180));
 sg13g2_o21ai_1 _3683_ (.B1(_0732_),
    .Y(_0733_),
    .A1(net1193),
    .A2(_0726_));
 sg13g2_inv_1 _3684_ (.Y(_0734_),
    .A(_0733_));
 sg13g2_nor2_2 _3685_ (.A(net1241),
    .B(\vga_tetris.tetrisLogic.stateQ[0] ),
    .Y(_0735_));
 sg13g2_nor2_1 _3686_ (.A(\vga_tetris.tetrisLogic.stateQ[2] ),
    .B(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0736_));
 sg13g2_nand2_1 _3687_ (.Y(_0737_),
    .A(net1234),
    .B(_0736_));
 sg13g2_nand3_1 _3688_ (.B(_0735_),
    .C(_0736_),
    .A(net1233),
    .Y(_0738_));
 sg13g2_nor2b_2 _3689_ (.A(net1796),
    .B_N(_0727_),
    .Y(_0739_));
 sg13g2_nand2b_2 _3690_ (.Y(_0740_),
    .B(_0727_),
    .A_N(\vga_tetris.tetrisLogic.stateQ[2] ));
 sg13g2_nor2b_2 _3691_ (.A(net1241),
    .B_N(\vga_tetris.tetrisLogic.stateQ[0] ),
    .Y(_0741_));
 sg13g2_and2_1 _3692_ (.A(_0739_),
    .B(_0741_),
    .X(_0742_));
 sg13g2_nor2b_1 _3693_ (.A(\vga_tetris.tetrisLogic.stateQ[3] ),
    .B_N(\vga_tetris.tetrisLogic.stateQ[2] ),
    .Y(_0743_));
 sg13g2_nand2b_1 _3694_ (.Y(_0744_),
    .B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .A_N(\vga_tetris.tetrisLogic.stateQ[3] ));
 sg13g2_nor2_2 _3695_ (.A(net1233),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_nand3_1 _3696_ (.B(net1241),
    .C(_0743_),
    .A(_0659_),
    .Y(_0746_));
 sg13g2_a22oi_1 _3697_ (.Y(_0747_),
    .B1(_0745_),
    .B2(net1242),
    .A2(_0739_),
    .A1(_0735_));
 sg13g2_nand3_1 _3698_ (.B(_0736_),
    .C(_0741_),
    .A(net1233),
    .Y(_0748_));
 sg13g2_nand2_2 _3699_ (.Y(_0749_),
    .A(net1241),
    .B(\vga_tetris.tetrisLogic.stateQ[0] ));
 sg13g2_o21ai_1 _3700_ (.B1(_0748_),
    .Y(_0750_),
    .A1(_0740_),
    .A2(_0749_));
 sg13g2_and4_1 _3701_ (.A(_0738_),
    .B(_0740_),
    .C(_0746_),
    .D(_0748_),
    .X(_0751_));
 sg13g2_nor4_2 _3702_ (.A(net1233),
    .B(net1242),
    .C(\vga_tetris.tetrisLogic.stateQ[0] ),
    .Y(_0752_),
    .D(_0744_));
 sg13g2_nand3_1 _3703_ (.B(_0735_),
    .C(_0743_),
    .A(_0659_),
    .Y(_0753_));
 sg13g2_nor2_2 _3704_ (.A(net1242),
    .B(_0728_),
    .Y(_0754_));
 sg13g2_nand2b_1 _3705_ (.Y(_0755_),
    .B(_0667_),
    .A_N(_0728_));
 sg13g2_nor2_1 _3706_ (.A(_0752_),
    .B(_0754_),
    .Y(_0756_));
 sg13g2_nand3_1 _3707_ (.B(_0753_),
    .C(_0755_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .Y(_0757_));
 sg13g2_o21ai_1 _3708_ (.B1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .Y(_0758_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_o21ai_1 _3709_ (.B1(_0758_),
    .Y(_0759_),
    .A1(_0751_),
    .A2(_0757_));
 sg13g2_and2_1 _3710_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0759_),
    .X(_0760_));
 sg13g2_nand3_1 _3711_ (.B(_0753_),
    .C(_0755_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .Y(_0761_));
 sg13g2_o21ai_1 _3712_ (.B1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .Y(_0762_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_o21ai_1 _3713_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0751_),
    .A2(_0761_));
 sg13g2_and2_1 _3714_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .B(_0763_),
    .X(_0764_));
 sg13g2_xor2_1 _3715_ (.B(_0759_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .X(_0765_));
 sg13g2_a21oi_1 _3716_ (.A1(_0764_),
    .A2(_0765_),
    .Y(_0766_),
    .B1(_0760_));
 sg13g2_o21ai_1 _3717_ (.B1(_0664_),
    .Y(_0767_),
    .A1(_0665_),
    .A2(_0766_));
 sg13g2_nand3b_1 _3718_ (.B(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .C(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .Y(_0768_),
    .A_N(_0766_));
 sg13g2_and3_1 _3719_ (.X(_0769_),
    .A(net1180),
    .B(_0767_),
    .C(_0768_));
 sg13g2_nand3_1 _3720_ (.B(_0767_),
    .C(_0768_),
    .A(net1180),
    .Y(_0770_));
 sg13g2_mux2_1 _3721_ (.A0(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .S(net1188),
    .X(_0771_));
 sg13g2_o21ai_1 _3722_ (.B1(_0730_),
    .Y(_0772_),
    .A1(_0642_),
    .A2(net1190));
 sg13g2_a21oi_1 _3723_ (.A1(net1189),
    .A2(_0771_),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_xor2_1 _3724_ (.B(_0768_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .X(_0774_));
 sg13g2_a21oi_2 _3725_ (.B1(_0773_),
    .Y(_0775_),
    .A2(_0774_),
    .A1(net1180));
 sg13g2_a21o_2 _3726_ (.A2(_0774_),
    .A1(net1180),
    .B1(_0773_),
    .X(_0776_));
 sg13g2_xnor2_1 _3727_ (.Y(_0777_),
    .A(_0665_),
    .B(_0766_));
 sg13g2_a21oi_1 _3728_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .A2(net1193),
    .Y(_0778_),
    .B1(net1180));
 sg13g2_mux2_1 _3729_ (.A0(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .S(net1188),
    .X(_0779_));
 sg13g2_nand2_1 _3730_ (.Y(_0780_),
    .A(net1190),
    .B(_0779_));
 sg13g2_a22oi_1 _3731_ (.Y(_0781_),
    .B1(_0778_),
    .B2(_0780_),
    .A2(_0777_),
    .A1(net1180));
 sg13g2_nor3_2 _3732_ (.A(_0734_),
    .B(_0769_),
    .C(_0781_),
    .Y(_0782_));
 sg13g2_nand3b_1 _3733_ (.B(_0770_),
    .C(_0733_),
    .Y(_0783_),
    .A_N(_0781_));
 sg13g2_nand2_1 _3734_ (.Y(_0784_),
    .A(_0775_),
    .B(_0783_));
 sg13g2_a21oi_1 _3735_ (.A1(_0733_),
    .A2(_0770_),
    .Y(_0785_),
    .B1(_0775_));
 sg13g2_nor3_1 _3736_ (.A(_0664_),
    .B(_0776_),
    .C(_0782_),
    .Y(_0786_));
 sg13g2_or2_1 _3737_ (.X(_0787_),
    .B(_0786_),
    .A(_0785_));
 sg13g2_o21ai_1 _3738_ (.B1(net1205),
    .Y(_0788_),
    .A1(_0785_),
    .A2(_0786_));
 sg13g2_nand3_1 _3739_ (.B(_0715_),
    .C(_0716_),
    .A(net1201),
    .Y(_0789_));
 sg13g2_or3_1 _3740_ (.A(net1202),
    .B(_0785_),
    .C(_0786_),
    .X(_0790_));
 sg13g2_nand3_1 _3741_ (.B(_0775_),
    .C(_0783_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .Y(_0791_));
 sg13g2_nand2_2 _3742_ (.Y(_0792_),
    .A(_0776_),
    .B(_0781_));
 sg13g2_nand2_2 _3743_ (.Y(_0793_),
    .A(_0791_),
    .B(_0792_));
 sg13g2_nand3_1 _3744_ (.B(_0791_),
    .C(_0792_),
    .A(net1205),
    .Y(_0794_));
 sg13g2_nand2_1 _3745_ (.Y(_0795_),
    .A(net1208),
    .B(net1201));
 sg13g2_or2_1 _3746_ (.X(_0796_),
    .B(net1205),
    .A(\vga_tetris._vgaController_io_pixelPosY[6] ));
 sg13g2_a21o_1 _3747_ (.A2(_0792_),
    .A1(_0791_),
    .B1(net1202),
    .X(_0797_));
 sg13g2_a22oi_1 _3748_ (.Y(_0798_),
    .B1(_0796_),
    .B2(_0797_),
    .A2(_0788_),
    .A1(_0717_));
 sg13g2_o21ai_1 _3749_ (.B1(_0775_),
    .Y(_0799_),
    .A1(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .A2(_0782_));
 sg13g2_nand2_1 _3750_ (.Y(_0800_),
    .A(net1206),
    .B(_0799_));
 sg13g2_nor2_1 _3751_ (.A(net1207),
    .B(_0715_),
    .Y(_0801_));
 sg13g2_a21oi_1 _3752_ (.A1(net1207),
    .A2(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_xor2_1 _3753_ (.B(_0715_),
    .A(net1207),
    .X(_0803_));
 sg13g2_and2_1 _3754_ (.A(net1201),
    .B(_0803_),
    .X(_0804_));
 sg13g2_nand2_1 _3755_ (.Y(_0805_),
    .A(net1201),
    .B(_0803_));
 sg13g2_a21oi_2 _3756_ (.B1(_0804_),
    .Y(_0806_),
    .A2(_0799_),
    .A1(net1205));
 sg13g2_a21o_1 _3757_ (.A2(_0799_),
    .A1(net1206),
    .B1(_0804_),
    .X(_0807_));
 sg13g2_xnor2_1 _3758_ (.Y(_0808_),
    .A(_0666_),
    .B(_0763_));
 sg13g2_a21oi_1 _3759_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .A2(net1193),
    .Y(_0809_),
    .B1(net1180));
 sg13g2_nand2_1 _3760_ (.Y(_0810_),
    .A(_0671_),
    .B(net1188));
 sg13g2_o21ai_1 _3761_ (.B1(_0810_),
    .Y(_0811_),
    .A1(net1229),
    .A2(net1188));
 sg13g2_o21ai_1 _3762_ (.B1(_0809_),
    .Y(_0812_),
    .A1(net1193),
    .A2(_0811_));
 sg13g2_o21ai_1 _3763_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0730_),
    .A2(_0808_));
 sg13g2_nor3_2 _3764_ (.A(_0666_),
    .B(_0776_),
    .C(_0782_),
    .Y(_0814_));
 sg13g2_a21oi_2 _3765_ (.B1(_0813_),
    .Y(_0815_),
    .A2(_0783_),
    .A1(_0775_));
 sg13g2_or2_1 _3766_ (.X(_0816_),
    .B(_0815_),
    .A(_0814_));
 sg13g2_o21ai_1 _3767_ (.B1(net1205),
    .Y(_0817_),
    .A1(_0814_),
    .A2(_0815_));
 sg13g2_nand2_2 _3768_ (.Y(_0818_),
    .A(\vga_tetris._tetrisDisplay_io_boardYCoord[0] ),
    .B(net1201));
 sg13g2_or3_1 _3769_ (.A(net1201),
    .B(_0814_),
    .C(_0815_),
    .X(_0819_));
 sg13g2_nand2_1 _3770_ (.Y(_0820_),
    .A(_0627_),
    .B(net1201));
 sg13g2_nor2_1 _3771_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .B(_0724_),
    .Y(_0821_));
 sg13g2_o21ai_1 _3772_ (.B1(net1190),
    .Y(_0822_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .A2(_0723_));
 sg13g2_a21oi_1 _3773_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .A2(net1193),
    .Y(_0823_),
    .B1(net1181));
 sg13g2_o21ai_1 _3774_ (.B1(_0823_),
    .Y(_0824_),
    .A1(_0821_),
    .A2(_0822_));
 sg13g2_xor2_1 _3775_ (.B(_0765_),
    .A(_0764_),
    .X(_0825_));
 sg13g2_o21ai_1 _3776_ (.B1(_0824_),
    .Y(_0826_),
    .A1(_0730_),
    .A2(_0825_));
 sg13g2_inv_1 _3777_ (.Y(_0827_),
    .A(_0826_));
 sg13g2_nor3_2 _3778_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0776_),
    .C(_0782_),
    .Y(_0828_));
 sg13g2_a21oi_2 _3779_ (.B1(_0827_),
    .Y(_0829_),
    .A2(_0783_),
    .A1(_0775_));
 sg13g2_nor2_1 _3780_ (.A(_0828_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_o21ai_1 _3781_ (.B1(net1205),
    .Y(_0831_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_or2_1 _3782_ (.X(_0832_),
    .B(net1205),
    .A(net1210));
 sg13g2_nand2_2 _3783_ (.Y(_0833_),
    .A(net1210),
    .B(net1201));
 sg13g2_or3_1 _3784_ (.A(net1202),
    .B(_0828_),
    .C(_0829_),
    .X(_0834_));
 sg13g2_nand2_1 _3785_ (.Y(_0835_),
    .A(_0833_),
    .B(_0834_));
 sg13g2_a22oi_1 _3786_ (.Y(_0836_),
    .B1(_0833_),
    .B2(_0834_),
    .A2(_0818_),
    .A1(_0817_));
 sg13g2_a221oi_1 _3787_ (.B2(_0834_),
    .C1(_0806_),
    .B1(_0833_),
    .A1(_0817_),
    .Y(_0837_),
    .A2(_0818_));
 sg13g2_and2_1 _3788_ (.A(net1079),
    .B(net1072),
    .X(_0838_));
 sg13g2_a22oi_1 _3789_ (.Y(_0839_),
    .B1(_0831_),
    .B2(_0832_),
    .A2(_0818_),
    .A1(_0817_));
 sg13g2_a22oi_1 _3790_ (.Y(_0840_),
    .B1(_0794_),
    .B2(_0795_),
    .A2(_0790_),
    .A1(_0789_));
 sg13g2_a221oi_1 _3791_ (.B2(_0795_),
    .C1(_0807_),
    .B1(_0794_),
    .A1(_0789_),
    .Y(_0841_),
    .A2(_0790_));
 sg13g2_and2_1 _3792_ (.A(_0839_),
    .B(net1058),
    .X(_0842_));
 sg13g2_a22oi_1 _3793_ (.Y(_0843_),
    .B1(net1021),
    .B2(\vga_tetris.boardMem.board_17[12] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[12] ));
 sg13g2_a221oi_1 _3794_ (.B2(_0832_),
    .C1(_0806_),
    .B1(_0831_),
    .A1(_0817_),
    .Y(_0844_),
    .A2(_0818_));
 sg13g2_and2_1 _3795_ (.A(net1064),
    .B(net1054),
    .X(_0845_));
 sg13g2_a22oi_1 _3796_ (.Y(_0846_),
    .B1(_0796_),
    .B2(_0797_),
    .A2(_0790_),
    .A1(_0789_));
 sg13g2_and2_1 _3797_ (.A(net1055),
    .B(net1049),
    .X(_0847_));
 sg13g2_a22oi_1 _3798_ (.Y(_0848_),
    .B1(_0831_),
    .B2(_0832_),
    .A2(_0820_),
    .A1(_0819_));
 sg13g2_nand4_1 _3799_ (.B(_0818_),
    .C(_0833_),
    .A(_0817_),
    .Y(_0849_),
    .D(_0834_));
 sg13g2_a221oi_1 _3800_ (.B2(_0832_),
    .C1(_0806_),
    .B1(_0831_),
    .A1(_0819_),
    .Y(_0850_),
    .A2(_0820_));
 sg13g2_and2_1 _3801_ (.A(net1077),
    .B(net1041),
    .X(_0851_));
 sg13g2_and2_1 _3802_ (.A(net1058),
    .B(net1043),
    .X(_0852_));
 sg13g2_a22oi_1 _3803_ (.Y(_0853_),
    .B1(_0833_),
    .B2(_0834_),
    .A2(_0820_),
    .A1(_0819_));
 sg13g2_a221oi_1 _3804_ (.B2(_0834_),
    .C1(_0806_),
    .B1(_0833_),
    .A1(_0819_),
    .Y(_0854_),
    .A2(_0820_));
 sg13g2_and2_1 _3805_ (.A(net1050),
    .B(net1036),
    .X(_0855_));
 sg13g2_and2_1 _3806_ (.A(net1077),
    .B(net1036),
    .X(_0856_));
 sg13g2_a22oi_1 _3807_ (.Y(_0857_),
    .B1(_0794_),
    .B2(_0795_),
    .A2(_0788_),
    .A1(_0717_));
 sg13g2_and2_1 _3808_ (.A(net1055),
    .B(net1031),
    .X(_0858_));
 sg13g2_and2_1 _3809_ (.A(net1041),
    .B(net1031),
    .X(_0859_));
 sg13g2_nand2_1 _3810_ (.Y(_0860_),
    .A(\vga_tetris.boardMem.board_8[12] ),
    .B(net1005));
 sg13g2_and2_1 _3811_ (.A(net1071),
    .B(net1031),
    .X(_0861_));
 sg13g2_and2_1 _3812_ (.A(net1037),
    .B(net1031),
    .X(_0862_));
 sg13g2_and2_1 _3813_ (.A(net1059),
    .B(_0853_),
    .X(_0863_));
 sg13g2_and2_1 _3814_ (.A(net1071),
    .B(net1050),
    .X(_0864_));
 sg13g2_a22oi_1 _3815_ (.Y(_0865_),
    .B1(net997),
    .B2(\vga_tetris.boardMem.board_7[12] ),
    .A2(net1000),
    .A1(\vga_tetris.boardMem.board_18[12] ));
 sg13g2_and2_1 _3816_ (.A(net1050),
    .B(net1041),
    .X(_0866_));
 sg13g2_and2_1 _3817_ (.A(net1078),
    .B(net1055),
    .X(_0867_));
 sg13g2_and2_1 _3818_ (.A(net1071),
    .B(net1064),
    .X(_0868_));
 sg13g2_a221oi_1 _3819_ (.B2(net1079),
    .C1(net1065),
    .B1(_0849_),
    .A1(_0800_),
    .Y(_0869_),
    .A2(_0805_));
 sg13g2_and2_1 _3820_ (.A(net1064),
    .B(net1037),
    .X(_0870_));
 sg13g2_nor2_2 _3821_ (.A(net1009),
    .B(net993),
    .Y(_0871_));
 sg13g2_and3_1 _3822_ (.X(_0872_),
    .A(_0807_),
    .B(_0835_),
    .C(net1065));
 sg13g2_a21o_1 _3823_ (.A2(net1056),
    .A1(net1065),
    .B1(net1061),
    .X(_0873_));
 sg13g2_nor4_2 _3824_ (.A(net1023),
    .B(_0869_),
    .C(_0872_),
    .Y(_0874_),
    .D(_0873_));
 sg13g2_and2_1 _3825_ (.A(_0871_),
    .B(net985),
    .X(_0875_));
 sg13g2_nand2_2 _3826_ (.Y(_0876_),
    .A(net986),
    .B(net985));
 sg13g2_and2_1 _3827_ (.A(_0836_),
    .B(net1058),
    .X(_0877_));
 sg13g2_a22oi_1 _3828_ (.Y(_0878_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[12] ),
    .A2(net1015),
    .A1(\vga_tetris.boardMem.board_12[12] ));
 sg13g2_a22oi_1 _3829_ (.Y(_0879_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[12] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[12] ));
 sg13g2_nand2_1 _3830_ (.Y(_0880_),
    .A(_0860_),
    .B(_0879_));
 sg13g2_a22oi_1 _3831_ (.Y(_0881_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[12] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_10[12] ));
 sg13g2_a22oi_1 _3832_ (.Y(_0882_),
    .B1(net1007),
    .B2(\vga_tetris.boardMem.board_9[12] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[12] ));
 sg13g2_a22oi_1 _3833_ (.Y(_0883_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[12] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[12] ));
 sg13g2_nand4_1 _3834_ (.B(_0865_),
    .C(_0882_),
    .A(_0843_),
    .Y(_0884_),
    .D(_0883_));
 sg13g2_a22oi_1 _3835_ (.Y(_0885_),
    .B1(net1011),
    .B2(\vga_tetris.boardMem.board_6[12] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[12] ));
 sg13g2_a22oi_1 _3836_ (.Y(_0886_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[12] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[12] ));
 sg13g2_nand4_1 _3837_ (.B(_0881_),
    .C(_0885_),
    .A(_0878_),
    .Y(_0887_),
    .D(_0886_));
 sg13g2_or4_1 _3838_ (.A(net844),
    .B(_0880_),
    .C(_0884_),
    .D(_0887_),
    .X(_0888_));
 sg13g2_nand2b_2 _3839_ (.Y(_0889_),
    .B(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .A_N(net744));
 sg13g2_or2_1 _3840_ (.X(_0890_),
    .B(net1196),
    .A(net1174));
 sg13g2_nor2_2 _3841_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0722_),
    .Y(_0891_));
 sg13g2_nor2b_1 _3842_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .Y(_0892_));
 sg13g2_nor2b_2 _3843_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .B_N(_0892_),
    .Y(_0893_));
 sg13g2_inv_1 _3844_ (.Y(_0894_),
    .A(_0893_));
 sg13g2_o21ai_1 _3845_ (.B1(net1174),
    .Y(_0895_),
    .A1(_0891_),
    .A2(_0893_));
 sg13g2_nand4_1 _3846_ (.B(_0751_),
    .C(_0890_),
    .A(net1206),
    .Y(_0896_),
    .D(_0895_));
 sg13g2_nand2_1 _3847_ (.Y(_0897_),
    .A(_0628_),
    .B(\vga_tetris._vgaController_io_pixelPosX[8] ));
 sg13g2_a21oi_1 _3848_ (.A1(net1218),
    .A2(net1219),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nand2_1 _3849_ (.Y(_0899_),
    .A(net1218),
    .B(net1220));
 sg13g2_nand2_1 _3850_ (.Y(_0900_),
    .A(_0898_),
    .B(_0899_));
 sg13g2_nor2_1 _3851_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_and2_1 _3852_ (.A(_0802_),
    .B(_0901_),
    .X(_0902_));
 sg13g2_inv_1 _3853_ (.Y(_0903_),
    .A(_0902_));
 sg13g2_nand2_2 _3854_ (.Y(_0904_),
    .A(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .B(net1224));
 sg13g2_and3_2 _3855_ (.X(_0905_),
    .A(net1225),
    .B(net1788),
    .C(net1782));
 sg13g2_and2_1 _3856_ (.A(net1819),
    .B(_0905_),
    .X(_0906_));
 sg13g2_nand2_1 _3857_ (.Y(_0907_),
    .A(net1819),
    .B(_0905_));
 sg13g2_nand2_1 _3858_ (.Y(_0908_),
    .A(net1821),
    .B(net1619));
 sg13g2_nand2_1 _3859_ (.Y(_0909_),
    .A(net1213),
    .B(net1216));
 sg13g2_nand3_1 _3860_ (.B(net1821),
    .C(net1619),
    .A(net1217),
    .Y(_0910_));
 sg13g2_nor2_2 _3861_ (.A(_0908_),
    .B(_0909_),
    .Y(_0911_));
 sg13g2_nor4_1 _3862_ (.A(net1215),
    .B(net1217),
    .C(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .D(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .Y(_0912_));
 sg13g2_nor4_2 _3863_ (.A(_0903_),
    .B(_0906_),
    .C(_0911_),
    .Y(_0913_),
    .D(_0912_));
 sg13g2_o21ai_1 _3864_ (.B1(_0896_),
    .Y(_0914_),
    .A1(net1206),
    .A2(_0913_));
 sg13g2_a21oi_1 _3865_ (.A1(_0685_),
    .A2(net844),
    .Y(_0915_),
    .B1(net1085));
 sg13g2_and2_1 _3866_ (.A(_0888_),
    .B(_0915_),
    .X(_0916_));
 sg13g2_nor2_2 _3867_ (.A(net1218),
    .B(_0629_),
    .Y(_0917_));
 sg13g2_nor2b_2 _3868_ (.A(net1223),
    .B_N(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .Y(_0918_));
 sg13g2_nand3_1 _3869_ (.B(_0917_),
    .C(_0918_),
    .A(_0916_),
    .Y(_0919_));
 sg13g2_nor2_2 _3870_ (.A(net1218),
    .B(net1219),
    .Y(_0920_));
 sg13g2_nand2b_1 _3871_ (.Y(_0921_),
    .B(net1223),
    .A_N(net1220));
 sg13g2_nand3b_1 _3872_ (.B(net1223),
    .C(_0920_),
    .Y(_0922_),
    .A_N(\vga_tetris._vgaController_io_pixelPosX[5] ));
 sg13g2_a22oi_1 _3873_ (.Y(_0923_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_18[2] ),
    .A2(net1007),
    .A1(\vga_tetris.boardMem.board_9[2] ));
 sg13g2_a22oi_1 _3874_ (.Y(_0924_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[2] ),
    .A2(net1005),
    .A1(\vga_tetris.boardMem.board_8[2] ));
 sg13g2_nand2_1 _3875_ (.Y(_0925_),
    .A(\vga_tetris.boardMem.board_11[2] ),
    .B(net1003));
 sg13g2_a22oi_1 _3876_ (.Y(_0926_),
    .B1(net1017),
    .B2(\vga_tetris.boardMem.board_5[2] ),
    .A2(net1020),
    .A1(\vga_tetris.boardMem.board_1[2] ));
 sg13g2_a22oi_1 _3877_ (.Y(_0927_),
    .B1(net1001),
    .B2(\vga_tetris.boardMem.board_10[2] ),
    .A2(net1015),
    .A1(\vga_tetris.boardMem.board_12[2] ));
 sg13g2_nand2_1 _3878_ (.Y(_0928_),
    .A(_0925_),
    .B(_0926_));
 sg13g2_a22oi_1 _3879_ (.Y(_0929_),
    .B1(net1009),
    .B2(\vga_tetris.boardMem.board_14[2] ),
    .A2(net1011),
    .A1(\vga_tetris.boardMem.board_6[2] ));
 sg13g2_a22oi_1 _3880_ (.Y(_0930_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[2] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[2] ));
 sg13g2_a22oi_1 _3881_ (.Y(_0931_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[2] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[2] ));
 sg13g2_a22oi_1 _3882_ (.Y(_0932_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[2] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_2[2] ));
 sg13g2_nand4_1 _3883_ (.B(_0930_),
    .C(_0931_),
    .A(_0929_),
    .Y(_0933_),
    .D(_0932_));
 sg13g2_a22oi_1 _3884_ (.Y(_0934_),
    .B1(net997),
    .B2(\vga_tetris.boardMem.board_7[2] ),
    .A2(net1021),
    .A1(\vga_tetris.boardMem.board_17[2] ));
 sg13g2_nand4_1 _3885_ (.B(_0924_),
    .C(_0927_),
    .A(_0923_),
    .Y(_0935_),
    .D(_0934_));
 sg13g2_or4_1 _3886_ (.A(net845),
    .B(_0928_),
    .C(_0933_),
    .D(_0935_),
    .X(_0936_));
 sg13g2_a21oi_1 _3887_ (.A1(_0675_),
    .A2(net845),
    .Y(_0937_),
    .B1(net1084));
 sg13g2_nand2_2 _3888_ (.Y(_0938_),
    .A(_0936_),
    .B(_0937_));
 sg13g2_nor2_1 _3889_ (.A(_0922_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_nand3_1 _3890_ (.B(net1073),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_14[6] ),
    .Y(_0940_));
 sg13g2_nand3_1 _3891_ (.B(net1044),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_6[6] ),
    .Y(_0941_));
 sg13g2_nand3_1 _3892_ (.B(_0839_),
    .C(net1057),
    .A(\vga_tetris.boardMem.board_17[6] ),
    .Y(_0942_));
 sg13g2_nand3_1 _3893_ (.B(net1062),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_2[6] ),
    .Y(_0943_));
 sg13g2_nand3_1 _3894_ (.B(net1070),
    .C(net1064),
    .A(\vga_tetris.boardMem.board_3[6] ),
    .Y(_0944_));
 sg13g2_nand3_1 _3895_ (.B(net1077),
    .C(net1054),
    .A(\vga_tetris.boardMem.board_13[6] ),
    .Y(_0945_));
 sg13g2_nand3_1 _3896_ (.B(net1073),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_12[6] ),
    .Y(_0946_));
 sg13g2_nand3_1 _3897_ (.B(net1064),
    .C(net1054),
    .A(\vga_tetris.boardMem.board_1[6] ),
    .Y(_0947_));
 sg13g2_nand3_1 _3898_ (.B(net1073),
    .C(net1066),
    .A(\vga_tetris.boardMem.board_15[6] ),
    .Y(_0948_));
 sg13g2_nand3_1 _3899_ (.B(net1057),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[6] ),
    .Y(_0949_));
 sg13g2_nand3_1 _3900_ (.B(net1051),
    .C(net1044),
    .A(\vga_tetris.boardMem.board_5[6] ),
    .Y(_0950_));
 sg13g2_nand3_1 _3901_ (.B(net1051),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_9[6] ),
    .Y(_0951_));
 sg13g2_nand3_1 _3902_ (.B(net1040),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_8[6] ),
    .Y(_0952_));
 sg13g2_nand3_1 _3903_ (.B(_0836_),
    .C(net1057),
    .A(\vga_tetris.boardMem.board_19[6] ),
    .Y(_0953_));
 sg13g2_nand3_1 _3904_ (.B(net1066),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_11[6] ),
    .Y(_0954_));
 sg13g2_nand3_1 _3905_ (.B(net1032),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_10[6] ),
    .Y(_0955_));
 sg13g2_nand3_1 _3906_ (.B(net1058),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[6] ),
    .Y(_0956_));
 sg13g2_nand3_1 _3907_ (.B(net1066),
    .C(net1044),
    .A(\vga_tetris.boardMem.board_7[6] ),
    .Y(_0957_));
 sg13g2_nand3_1 _3908_ (.B(net1044),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_4[6] ),
    .Y(_0958_));
 sg13g2_nand4_1 _3909_ (.B(_0945_),
    .C(_0947_),
    .A(_0944_),
    .Y(_0959_),
    .D(_0956_));
 sg13g2_a21oi_1 _3910_ (.A1(net986),
    .A2(net985),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_nand4_1 _3911_ (.B(_0946_),
    .C(_0948_),
    .A(_0940_),
    .Y(_0961_),
    .D(_0957_));
 sg13g2_nand4_1 _3912_ (.B(_0950_),
    .C(_0952_),
    .A(_0942_),
    .Y(_0962_),
    .D(_0953_));
 sg13g2_nand3_1 _3913_ (.B(_0949_),
    .C(_0955_),
    .A(_0943_),
    .Y(_0963_));
 sg13g2_nand4_1 _3914_ (.B(_0951_),
    .C(_0954_),
    .A(_0941_),
    .Y(_0964_),
    .D(_0958_));
 sg13g2_nor4_2 _3915_ (.A(_0961_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0965_),
    .D(_0964_));
 sg13g2_a221oi_1 _3916_ (.B2(_0965_),
    .C1(net1083),
    .B1(_0960_),
    .A1(_0679_),
    .Y(_0966_),
    .A2(net843));
 sg13g2_and2_1 _3917_ (.A(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .B(net1223),
    .X(_0967_));
 sg13g2_nand3_1 _3918_ (.B(_0966_),
    .C(_0967_),
    .A(_0920_),
    .Y(_0968_));
 sg13g2_nand2_2 _3919_ (.Y(_0969_),
    .A(_0917_),
    .B(_0967_));
 sg13g2_nand2_1 _3920_ (.Y(_0970_),
    .A(\vga_tetris.boardMem.board_18[14] ),
    .B(net999));
 sg13g2_a22oi_1 _3921_ (.Y(_0971_),
    .B1(net1015),
    .B2(\vga_tetris.boardMem.board_12[14] ),
    .A2(net1021),
    .A1(\vga_tetris.boardMem.board_17[14] ));
 sg13g2_a22oi_1 _3922_ (.Y(_0972_),
    .B1(net1007),
    .B2(\vga_tetris.boardMem.board_9[14] ),
    .A2(net1020),
    .A1(\vga_tetris.boardMem.board_1[14] ));
 sg13g2_a22oi_1 _3923_ (.Y(_0973_),
    .B1(net1005),
    .B2(\vga_tetris.boardMem.board_8[14] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[14] ));
 sg13g2_a22oi_1 _3924_ (.Y(_0974_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[14] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_10[14] ));
 sg13g2_a22oi_1 _3925_ (.Y(_0975_),
    .B1(net1003),
    .B2(\vga_tetris.boardMem.board_11[14] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[14] ));
 sg13g2_a22oi_1 _3926_ (.Y(_0976_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[14] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_7[14] ));
 sg13g2_a22oi_1 _3927_ (.Y(_0977_),
    .B1(net1017),
    .B2(\vga_tetris.boardMem.board_5[14] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[14] ));
 sg13g2_nand4_1 _3928_ (.B(_0975_),
    .C(_0976_),
    .A(_0974_),
    .Y(_0978_),
    .D(_0977_));
 sg13g2_nand2_1 _3929_ (.Y(_0979_),
    .A(_0970_),
    .B(_0973_));
 sg13g2_a22oi_1 _3930_ (.Y(_0980_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[14] ),
    .A2(net1011),
    .A1(\vga_tetris.boardMem.board_6[14] ));
 sg13g2_a22oi_1 _3931_ (.Y(_0981_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[14] ),
    .A2(net993),
    .A1(\vga_tetris.boardMem.board_13[14] ));
 sg13g2_nand4_1 _3932_ (.B(_0972_),
    .C(_0980_),
    .A(_0971_),
    .Y(_0982_),
    .D(_0981_));
 sg13g2_or4_1 _3933_ (.A(net845),
    .B(_0978_),
    .C(_0979_),
    .D(_0982_),
    .X(_0983_));
 sg13g2_a21oi_1 _3934_ (.A1(_0687_),
    .A2(net845),
    .Y(_0984_),
    .B1(net1084));
 sg13g2_nand2_2 _3935_ (.Y(_0985_),
    .A(_0983_),
    .B(_0984_));
 sg13g2_nor2_1 _3936_ (.A(net1220),
    .B(net1223),
    .Y(_0986_));
 sg13g2_and2_1 _3937_ (.A(_0920_),
    .B(_0986_),
    .X(_0987_));
 sg13g2_a22oi_1 _3938_ (.Y(_0988_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[0] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[0] ));
 sg13g2_nand2_1 _3939_ (.Y(_0989_),
    .A(\vga_tetris.boardMem.board_12[0] ),
    .B(net1015));
 sg13g2_a22oi_1 _3940_ (.Y(_0990_),
    .B1(net1001),
    .B2(\vga_tetris.boardMem.board_10[0] ),
    .A2(net1007),
    .A1(\vga_tetris.boardMem.board_9[0] ));
 sg13g2_a22oi_1 _3941_ (.Y(_0991_),
    .B1(net997),
    .B2(\vga_tetris.boardMem.board_7[0] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_18[0] ));
 sg13g2_nand2_1 _3942_ (.Y(_0992_),
    .A(_0989_),
    .B(_0991_));
 sg13g2_a22oi_1 _3943_ (.Y(_0993_),
    .B1(net1005),
    .B2(\vga_tetris.boardMem.board_8[0] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[0] ));
 sg13g2_a22oi_1 _3944_ (.Y(_0994_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[0] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[0] ));
 sg13g2_a22oi_1 _3945_ (.Y(_0995_),
    .B1(net1011),
    .B2(\vga_tetris.boardMem.board_6[0] ),
    .A2(net1021),
    .A1(\vga_tetris.boardMem.board_17[0] ));
 sg13g2_a22oi_1 _3946_ (.Y(_0996_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[0] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[0] ));
 sg13g2_nand4_1 _3947_ (.B(_0994_),
    .C(_0995_),
    .A(_0988_),
    .Y(_0997_),
    .D(_0996_));
 sg13g2_a22oi_1 _3948_ (.Y(_0998_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[0] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[0] ));
 sg13g2_a22oi_1 _3949_ (.Y(_0999_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[0] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[0] ));
 sg13g2_nand4_1 _3950_ (.B(_0993_),
    .C(_0998_),
    .A(_0990_),
    .Y(_1000_),
    .D(_0999_));
 sg13g2_or4_1 _3951_ (.A(net846),
    .B(_0992_),
    .C(_0997_),
    .D(_1000_),
    .X(_1001_));
 sg13g2_a21oi_2 _3952_ (.B1(net1084),
    .Y(_1002_),
    .A2(net846),
    .A1(_0673_));
 sg13g2_nand2_1 _3953_ (.Y(_1003_),
    .A(_1001_),
    .B(_1002_));
 sg13g2_nand3_1 _3954_ (.B(_1001_),
    .C(_1002_),
    .A(_0987_),
    .Y(_1004_));
 sg13g2_nand3_1 _3955_ (.B(_0836_),
    .C(net1060),
    .A(\vga_tetris.boardMem.board_19[10] ),
    .Y(_1005_));
 sg13g2_nand3_1 _3956_ (.B(net1060),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[10] ),
    .Y(_1006_));
 sg13g2_nand3_1 _3957_ (.B(net1039),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_8[10] ),
    .Y(_1007_));
 sg13g2_nand3_1 _3958_ (.B(net1034),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_10[10] ),
    .Y(_1008_));
 sg13g2_nand3_1 _3959_ (.B(net1067),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_7[10] ),
    .Y(_1009_));
 sg13g2_nand3_1 _3960_ (.B(net1053),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_9[10] ),
    .Y(_1010_));
 sg13g2_nand3_1 _3961_ (.B(net1061),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[10] ),
    .Y(_1011_));
 sg13g2_nand3_1 _3962_ (.B(net1075),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_14[10] ),
    .Y(_1012_));
 sg13g2_nand3_1 _3963_ (.B(net1052),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_5[10] ),
    .Y(_1013_));
 sg13g2_nand3_1 _3964_ (.B(_0839_),
    .C(net1060),
    .A(\vga_tetris.boardMem.board_17[10] ),
    .Y(_1014_));
 sg13g2_nand3_1 _3965_ (.B(net1067),
    .C(net1063),
    .A(\vga_tetris.boardMem.board_3[10] ),
    .Y(_1015_));
 sg13g2_nand3_1 _3966_ (.B(net1063),
    .C(net1035),
    .A(\vga_tetris.boardMem.board_2[10] ),
    .Y(_1016_));
 sg13g2_nand3_1 _3967_ (.B(net1067),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_11[10] ),
    .Y(_1017_));
 sg13g2_nand3_1 _3968_ (.B(net1075),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_12[10] ),
    .Y(_1018_));
 sg13g2_nand3_1 _3969_ (.B(net1076),
    .C(net1052),
    .A(\vga_tetris.boardMem.board_13[10] ),
    .Y(_1019_));
 sg13g2_nand3_1 _3970_ (.B(net1076),
    .C(net1068),
    .A(\vga_tetris.boardMem.board_15[10] ),
    .Y(_1020_));
 sg13g2_nand3_1 _3971_ (.B(net1047),
    .C(net1042),
    .A(\vga_tetris.boardMem.board_4[10] ),
    .Y(_1021_));
 sg13g2_nand3_1 _3972_ (.B(net1063),
    .C(net1052),
    .A(\vga_tetris.boardMem.board_1[10] ),
    .Y(_1022_));
 sg13g2_nand3_1 _3973_ (.B(net1047),
    .C(net1035),
    .A(\vga_tetris.boardMem.board_6[10] ),
    .Y(_1023_));
 sg13g2_nand4_1 _3974_ (.B(_1011_),
    .C(_1021_),
    .A(_1010_),
    .Y(_1024_),
    .D(_1023_));
 sg13g2_a21oi_1 _3975_ (.A1(net986),
    .A2(net985),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_nand4_1 _3976_ (.B(_1009_),
    .C(_1015_),
    .A(_1005_),
    .Y(_1026_),
    .D(_1022_));
 sg13g2_nand4_1 _3977_ (.B(_1013_),
    .C(_1017_),
    .A(_1007_),
    .Y(_1027_),
    .D(_1019_));
 sg13g2_nand3_1 _3978_ (.B(_1012_),
    .C(_1016_),
    .A(_1008_),
    .Y(_1028_));
 sg13g2_nand4_1 _3979_ (.B(_1014_),
    .C(_1018_),
    .A(_1006_),
    .Y(_1029_),
    .D(_1020_));
 sg13g2_nor4_1 _3980_ (.A(_1026_),
    .B(_1027_),
    .C(_1028_),
    .D(_1029_),
    .Y(_1030_));
 sg13g2_a221oi_1 _3981_ (.B2(_1030_),
    .C1(net1083),
    .B1(_1025_),
    .A1(_0683_),
    .Y(_1031_),
    .A2(net843));
 sg13g2_nor3_1 _3982_ (.A(net1218),
    .B(_0629_),
    .C(_0921_),
    .Y(_1032_));
 sg13g2_a22oi_1 _3983_ (.Y(_1033_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[8] ),
    .A2(net1005),
    .A1(\vga_tetris.boardMem.board_8[8] ));
 sg13g2_nand2_1 _3984_ (.Y(_1034_),
    .A(\vga_tetris.boardMem.board_7[8] ),
    .B(net997));
 sg13g2_a22oi_1 _3985_ (.Y(_1035_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[8] ),
    .A2(net1011),
    .A1(\vga_tetris.boardMem.board_6[8] ));
 sg13g2_a22oi_1 _3986_ (.Y(_1036_),
    .B1(net1015),
    .B2(\vga_tetris.boardMem.board_12[8] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[8] ));
 sg13g2_a22oi_1 _3987_ (.Y(_1037_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[8] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_10[8] ));
 sg13g2_a22oi_1 _3988_ (.Y(_1038_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[8] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[8] ));
 sg13g2_nand2_1 _3989_ (.Y(_1039_),
    .A(_1034_),
    .B(_1038_));
 sg13g2_a22oi_1 _3990_ (.Y(_1040_),
    .B1(net1022),
    .B2(\vga_tetris.boardMem.board_17[8] ),
    .A2(net1024),
    .A1(\vga_tetris.boardMem.board_15[8] ));
 sg13g2_a22oi_1 _3991_ (.Y(_1041_),
    .B1(net1003),
    .B2(\vga_tetris.boardMem.board_11[8] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[8] ));
 sg13g2_a22oi_1 _3992_ (.Y(_1042_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[8] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_18[8] ));
 sg13g2_a22oi_1 _3993_ (.Y(_1043_),
    .B1(net1007),
    .B2(\vga_tetris.boardMem.board_9[8] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[8] ));
 sg13g2_nand4_1 _3994_ (.B(_1041_),
    .C(_1042_),
    .A(_1040_),
    .Y(_1044_),
    .D(_1043_));
 sg13g2_nand4_1 _3995_ (.B(_1035_),
    .C(_1036_),
    .A(_1033_),
    .Y(_1045_),
    .D(_1037_));
 sg13g2_or4_1 _3996_ (.A(net846),
    .B(_1039_),
    .C(_1044_),
    .D(_1045_),
    .X(_1046_));
 sg13g2_a21oi_1 _3997_ (.A1(_0681_),
    .A2(net846),
    .Y(_1047_),
    .B1(net1084));
 sg13g2_nand2_2 _3998_ (.Y(_1048_),
    .A(_1046_),
    .B(_1047_));
 sg13g2_nand2_1 _3999_ (.Y(_1049_),
    .A(_0917_),
    .B(_0986_));
 sg13g2_nand3_1 _4000_ (.B(net1063),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_2[18] ),
    .Y(_1050_));
 sg13g2_nand3_1 _4001_ (.B(net1075),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_12[18] ),
    .Y(_1051_));
 sg13g2_nand3_1 _4002_ (.B(net1075),
    .C(net1052),
    .A(\vga_tetris.boardMem.board_13[18] ),
    .Y(_1052_));
 sg13g2_nand3_1 _4003_ (.B(net1067),
    .C(net1063),
    .A(\vga_tetris.boardMem.board_3[18] ),
    .Y(_1053_));
 sg13g2_nand3_1 _4004_ (.B(net1052),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_5[18] ),
    .Y(_1054_));
 sg13g2_nand3_1 _4005_ (.B(net1061),
    .C(_0848_),
    .A(\vga_tetris.boardMem.board_16[18] ),
    .Y(_1055_));
 sg13g2_nand3_1 _4006_ (.B(net1039),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_8[18] ),
    .Y(_1056_));
 sg13g2_nand3_1 _4007_ (.B(net1053),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_9[18] ),
    .Y(_1057_));
 sg13g2_nand3_1 _4008_ (.B(_0839_),
    .C(net1060),
    .A(\vga_tetris.boardMem.board_17[18] ),
    .Y(_1058_));
 sg13g2_nand3_1 _4009_ (.B(net1060),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[18] ),
    .Y(_1059_));
 sg13g2_nand3_1 _4010_ (.B(net1068),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_11[18] ),
    .Y(_1060_));
 sg13g2_nand3_1 _4011_ (.B(net1075),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_14[18] ),
    .Y(_1061_));
 sg13g2_nand3_1 _4012_ (.B(net1068),
    .C(net1047),
    .A(\vga_tetris.boardMem.board_7[18] ),
    .Y(_1062_));
 sg13g2_nand3_1 _4013_ (.B(net1047),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_4[18] ),
    .Y(_1063_));
 sg13g2_nand3_1 _4014_ (.B(net1046),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_6[18] ),
    .Y(_1064_));
 sg13g2_nand3_1 _4015_ (.B(net1075),
    .C(net1067),
    .A(\vga_tetris.boardMem.board_15[18] ),
    .Y(_1065_));
 sg13g2_nand3_1 _4016_ (.B(_0836_),
    .C(net1061),
    .A(\vga_tetris.boardMem.board_19[18] ),
    .Y(_1066_));
 sg13g2_nand3_1 _4017_ (.B(net1035),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_10[18] ),
    .Y(_1067_));
 sg13g2_nand3_1 _4018_ (.B(net1063),
    .C(net1052),
    .A(\vga_tetris.boardMem.board_1[18] ),
    .Y(_1068_));
 sg13g2_nand4_1 _4019_ (.B(_1057_),
    .C(_1060_),
    .A(_1056_),
    .Y(_1069_),
    .D(_1067_));
 sg13g2_a21oi_1 _4020_ (.A1(net986),
    .A2(net985),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_nand4_1 _4021_ (.B(_1054_),
    .C(_1055_),
    .A(_1050_),
    .Y(_1071_),
    .D(_1066_));
 sg13g2_nand4_1 _4022_ (.B(_1059_),
    .C(_1062_),
    .A(_1058_),
    .Y(_1072_),
    .D(_1063_));
 sg13g2_nand3_1 _4023_ (.B(_1061_),
    .C(_1065_),
    .A(_1053_),
    .Y(_1073_));
 sg13g2_nand4_1 _4024_ (.B(_1052_),
    .C(_1064_),
    .A(_1051_),
    .Y(_1074_),
    .D(_1068_));
 sg13g2_nor4_1 _4025_ (.A(_1071_),
    .B(_1072_),
    .C(_1073_),
    .D(_1074_),
    .Y(_1075_));
 sg13g2_a221oi_1 _4026_ (.B2(_1075_),
    .C1(net1083),
    .B1(_1070_),
    .A1(_0691_),
    .Y(_1076_),
    .A2(net843));
 sg13g2_nor2b_1 _4027_ (.A(net1219),
    .B_N(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .Y(_1077_));
 sg13g2_nand2_1 _4028_ (.Y(_1078_),
    .A(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .B(_0629_));
 sg13g2_nor2_1 _4029_ (.A(_0921_),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_nand2_1 _4030_ (.Y(_1080_),
    .A(_1076_),
    .B(_1079_));
 sg13g2_a22oi_1 _4031_ (.Y(_1081_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_19[16] ),
    .A2(net1012),
    .A1(\vga_tetris.boardMem.board_6[16] ));
 sg13g2_a22oi_1 _4032_ (.Y(_1082_),
    .B1(net1002),
    .B2(\vga_tetris.boardMem.board_10[16] ),
    .A2(net1014),
    .A1(\vga_tetris.boardMem.board_16[16] ));
 sg13g2_a22oi_1 _4033_ (.Y(_1083_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[16] ),
    .A2(net1018),
    .A1(\vga_tetris.boardMem.board_5[16] ));
 sg13g2_a22oi_1 _4034_ (.Y(_1084_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[16] ),
    .A2(net1015),
    .A1(\vga_tetris.boardMem.board_12[16] ));
 sg13g2_nand4_1 _4035_ (.B(_1082_),
    .C(_1083_),
    .A(_1081_),
    .Y(_1085_),
    .D(_1084_));
 sg13g2_a22oi_1 _4036_ (.Y(_1086_),
    .B1(net1006),
    .B2(\vga_tetris.boardMem.board_8[16] ),
    .A2(net1008),
    .A1(\vga_tetris.boardMem.board_9[16] ));
 sg13g2_a22oi_1 _4037_ (.Y(_1087_),
    .B1(net994),
    .B2(\vga_tetris.boardMem.board_13[16] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[16] ));
 sg13g2_a22oi_1 _4038_ (.Y(_1088_),
    .B1(net990),
    .B2(\vga_tetris.boardMem.board_2[16] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_7[16] ));
 sg13g2_a22oi_1 _4039_ (.Y(_1089_),
    .B1(net1019),
    .B2(\vga_tetris.boardMem.board_1[16] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[16] ));
 sg13g2_and4_1 _4040_ (.A(_1086_),
    .B(_1087_),
    .C(_1088_),
    .D(_1089_),
    .X(_1090_));
 sg13g2_nand2_1 _4041_ (.Y(_1091_),
    .A(\vga_tetris.boardMem.board_17[16] ),
    .B(net1021));
 sg13g2_a22oi_1 _4042_ (.Y(_1092_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_18[16] ),
    .A2(net1010),
    .A1(\vga_tetris.boardMem.board_14[16] ));
 sg13g2_nand4_1 _4043_ (.B(_1090_),
    .C(_1091_),
    .A(_0876_),
    .Y(_1093_),
    .D(_1092_));
 sg13g2_a21oi_1 _4044_ (.A1(_0689_),
    .A2(net845),
    .Y(_1094_),
    .B1(net1084));
 sg13g2_o21ai_1 _4045_ (.B1(_1094_),
    .Y(_1095_),
    .A1(_1085_),
    .A2(_1093_));
 sg13g2_nand2_1 _4046_ (.Y(_1096_),
    .A(_0986_),
    .B(_1077_));
 sg13g2_nand3_1 _4047_ (.B(net1065),
    .C(net1038),
    .A(\vga_tetris.boardMem.board_2[4] ),
    .Y(_1097_));
 sg13g2_nand3_1 _4048_ (.B(net1078),
    .C(net1036),
    .A(\vga_tetris.boardMem.board_14[4] ),
    .Y(_1098_));
 sg13g2_nand3_1 _4049_ (.B(net1079),
    .C(net1056),
    .A(\vga_tetris.boardMem.board_13[4] ),
    .Y(_1099_));
 sg13g2_nand3_1 _4050_ (.B(_0836_),
    .C(net1058),
    .A(\vga_tetris.boardMem.board_19[4] ),
    .Y(_1100_));
 sg13g2_nand3_1 _4051_ (.B(net1071),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_11[4] ),
    .Y(_1101_));
 sg13g2_nand3_1 _4052_ (.B(net1061),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[4] ),
    .Y(_1102_));
 sg13g2_nand3_1 _4053_ (.B(net1054),
    .C(net1049),
    .A(\vga_tetris.boardMem.board_5[4] ),
    .Y(_1103_));
 sg13g2_nand3_1 _4054_ (.B(net1064),
    .C(net1054),
    .A(\vga_tetris.boardMem.board_1[4] ),
    .Y(_1104_));
 sg13g2_nand3_1 _4055_ (.B(net1050),
    .C(net1037),
    .A(\vga_tetris.boardMem.board_6[4] ),
    .Y(_1105_));
 sg13g2_nand3_1 _4056_ (.B(net1061),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[4] ),
    .Y(_1106_));
 sg13g2_nand3_1 _4057_ (.B(net1078),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_12[4] ),
    .Y(_1107_));
 sg13g2_nand3_1 _4058_ (.B(net1049),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_4[4] ),
    .Y(_1108_));
 sg13g2_nand3_1 _4059_ (.B(net1077),
    .C(net1070),
    .A(\vga_tetris.boardMem.board_15[4] ),
    .Y(_1109_));
 sg13g2_nand3_1 _4060_ (.B(net1036),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_10[4] ),
    .Y(_1110_));
 sg13g2_nand3_1 _4061_ (.B(net1070),
    .C(net1065),
    .A(\vga_tetris.boardMem.board_3[4] ),
    .Y(_1111_));
 sg13g2_nand3_1 _4062_ (.B(net1055),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_9[4] ),
    .Y(_1112_));
 sg13g2_nand3_1 _4063_ (.B(net1042),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_8[4] ),
    .Y(_1113_));
 sg13g2_nand3_1 _4064_ (.B(net1070),
    .C(net1049),
    .A(\vga_tetris.boardMem.board_7[4] ),
    .Y(_1114_));
 sg13g2_nand3_1 _4065_ (.B(_0839_),
    .C(net1058),
    .A(\vga_tetris.boardMem.board_17[4] ),
    .Y(_1115_));
 sg13g2_nand4_1 _4066_ (.B(_1099_),
    .C(_1102_),
    .A(_1097_),
    .Y(_1116_),
    .D(_1106_));
 sg13g2_a21oi_1 _4067_ (.A1(net986),
    .A2(_0874_),
    .Y(_1117_),
    .B1(_1116_));
 sg13g2_nand4_1 _4068_ (.B(_1107_),
    .C(_1109_),
    .A(_1103_),
    .Y(_1118_),
    .D(_1112_));
 sg13g2_nand4_1 _4069_ (.B(_1105_),
    .C(_1111_),
    .A(_1101_),
    .Y(_1119_),
    .D(_1113_));
 sg13g2_nand3_1 _4070_ (.B(_1104_),
    .C(_1115_),
    .A(_1100_),
    .Y(_1120_));
 sg13g2_nand4_1 _4071_ (.B(_1108_),
    .C(_1110_),
    .A(_1098_),
    .Y(_1121_),
    .D(_1114_));
 sg13g2_nor4_1 _4072_ (.A(_1118_),
    .B(_1119_),
    .C(_1120_),
    .D(_1121_),
    .Y(_1122_));
 sg13g2_a221oi_1 _4073_ (.B2(_1122_),
    .C1(net1083),
    .B1(_1117_),
    .A1(_0677_),
    .Y(_1123_),
    .A2(net843));
 sg13g2_nand3_1 _4074_ (.B(_0920_),
    .C(_1123_),
    .A(_0918_),
    .Y(_1124_));
 sg13g2_o21ai_1 _4075_ (.B1(_0968_),
    .Y(_1125_),
    .A1(_1048_),
    .A2(_1049_));
 sg13g2_o21ai_1 _4076_ (.B1(_1004_),
    .Y(_1126_),
    .A1(_1095_),
    .A2(_1096_));
 sg13g2_a21oi_1 _4077_ (.A1(_1031_),
    .A2(_1032_),
    .Y(_1127_),
    .B1(_0939_));
 sg13g2_nand3_1 _4078_ (.B(_1124_),
    .C(_1127_),
    .A(_0919_),
    .Y(_1128_));
 sg13g2_o21ai_1 _4079_ (.B1(_1080_),
    .Y(_1129_),
    .A1(_0969_),
    .A2(_0985_));
 sg13g2_nor4_2 _4080_ (.A(_1125_),
    .B(_1126_),
    .C(_1128_),
    .Y(_1130_),
    .D(_1129_));
 sg13g2_nand4_1 _4081_ (.B(net1833),
    .C(net1863),
    .A(net1690),
    .Y(_1131_),
    .D(\vga_tetris.vgaController.verticalCounterQ[5] ));
 sg13g2_inv_1 _4082_ (.Y(_1132_),
    .A(net1864));
 sg13g2_nand2_1 _4083_ (.Y(_1133_),
    .A(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[9] ));
 sg13g2_a21oi_1 _4084_ (.A1(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .A2(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .Y(_1134_),
    .B1(\vga_tetris.vgaController.verticalCounterQ[9] ));
 sg13g2_nand4_1 _4085_ (.B(_1131_),
    .C(_1133_),
    .A(net1259),
    .Y(_1135_),
    .D(_1134_));
 sg13g2_inv_1 _4086_ (.Y(_1136_),
    .A(_1135_));
 sg13g2_nand2_1 _4087_ (.Y(_1137_),
    .A(_0913_),
    .B(_1136_));
 sg13g2_nor2_1 _4088_ (.A(_1130_),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_nor2_1 _4089_ (.A(net1809),
    .B(net1776),
    .Y(_1139_));
 sg13g2_nor2_1 _4090_ (.A(net1209),
    .B(net1211),
    .Y(_1140_));
 sg13g2_nand2_1 _4091_ (.Y(_1141_),
    .A(_0912_),
    .B(_1140_));
 sg13g2_nand3_1 _4092_ (.B(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .C(_1141_),
    .A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .Y(_1142_));
 sg13g2_and4_1 _4093_ (.A(_0625_),
    .B(net1207),
    .C(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .D(net1208),
    .X(_1143_));
 sg13g2_inv_1 _4094_ (.Y(_1144_),
    .A(_1143_));
 sg13g2_nor4_1 _4095_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(_0801_),
    .C(_0897_),
    .D(_1143_),
    .Y(_1145_));
 sg13g2_a22oi_1 _4096_ (.Y(_1146_),
    .B1(_1142_),
    .B2(_1145_),
    .A2(_1139_),
    .A1(_0987_));
 sg13g2_or2_1 _4097_ (.X(_1147_),
    .B(net1224),
    .A(\vga_tetris._vgaController_io_pixelPosX[3] ));
 sg13g2_a21oi_1 _4098_ (.A1(_0918_),
    .A2(_1077_),
    .Y(_1148_),
    .B1(_0987_));
 sg13g2_nor4_1 _4099_ (.A(\vga_tetris._vgaController_io_pixelPosX[1] ),
    .B(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .C(net1194),
    .D(_1148_),
    .Y(_1149_));
 sg13g2_nor2b_1 _4100_ (.A(_1146_),
    .B_N(_1149_),
    .Y(_1150_));
 sg13g2_nand2_1 _4101_ (.Y(_1151_),
    .A(_0625_),
    .B(_0801_));
 sg13g2_nor2_1 _4102_ (.A(net1207),
    .B(_0626_),
    .Y(_1152_));
 sg13g2_a21oi_1 _4103_ (.A1(net1207),
    .A2(net1208),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_nand3_1 _4104_ (.B(_0901_),
    .C(_1153_),
    .A(_0715_),
    .Y(_1154_));
 sg13g2_a21oi_1 _4105_ (.A1(_1151_),
    .A2(_1154_),
    .Y(_1155_),
    .B1(_1141_));
 sg13g2_nand2_1 _4106_ (.Y(_1156_),
    .A(net1212),
    .B(_0911_));
 sg13g2_nor3_1 _4107_ (.A(net1209),
    .B(_1144_),
    .C(_1156_),
    .Y(_1157_));
 sg13g2_nor4_1 _4108_ (.A(_0628_),
    .B(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .C(_0907_),
    .D(_0969_),
    .Y(_1158_));
 sg13g2_nor4_1 _4109_ (.A(_1150_),
    .B(_1155_),
    .C(_1157_),
    .D(_1158_),
    .Y(_1159_));
 sg13g2_inv_2 _4110_ (.Y(_1160_),
    .A(_1159_));
 sg13g2_nor2_1 _4111_ (.A(net1221),
    .B(net1194),
    .Y(_1161_));
 sg13g2_o21ai_1 _4112_ (.B1(net1220),
    .Y(_1162_),
    .A1(net1222),
    .A2(net1194));
 sg13g2_xor2_1 _4113_ (.B(_1161_),
    .A(net1220),
    .X(_1163_));
 sg13g2_a21oi_1 _4114_ (.A1(net1215),
    .A2(net1216),
    .Y(_1164_),
    .B1(net1211));
 sg13g2_nand2b_1 _4115_ (.Y(_1165_),
    .B(net1209),
    .A_N(_1164_));
 sg13g2_nand2_1 _4116_ (.Y(_1166_),
    .A(_0909_),
    .B(_1140_));
 sg13g2_and2_1 _4117_ (.A(_1165_),
    .B(_1166_),
    .X(_1167_));
 sg13g2_nand2b_1 _4118_ (.Y(_1168_),
    .B(_1167_),
    .A_N(net1216));
 sg13g2_nand2b_1 _4119_ (.Y(_1169_),
    .B(_0627_),
    .A_N(_1168_));
 sg13g2_or2_1 _4120_ (.X(_1170_),
    .B(_1168_),
    .A(net1214));
 sg13g2_nor2_2 _4121_ (.A(net1214),
    .B(_1169_),
    .Y(_1171_));
 sg13g2_nand2_1 _4122_ (.Y(_1172_),
    .A(_0627_),
    .B(net1216));
 sg13g2_a21oi_1 _4123_ (.A1(net1213),
    .A2(_1172_),
    .Y(_1173_),
    .B1(_1165_));
 sg13g2_nor3_1 _4124_ (.A(_0904_),
    .B(_1171_),
    .C(_1173_),
    .Y(_1174_));
 sg13g2_xor2_1 _4125_ (.B(_1147_),
    .A(net1221),
    .X(_1175_));
 sg13g2_xnor2_1 _4126_ (.Y(_1176_),
    .A(net1221),
    .B(net1194));
 sg13g2_nor2b_1 _4127_ (.A(net1213),
    .B_N(net1216),
    .Y(_1177_));
 sg13g2_nand2b_2 _4128_ (.Y(_1178_),
    .B(net1217),
    .A_N(net1213));
 sg13g2_and2_1 _4129_ (.A(net1209),
    .B(net1212),
    .X(_1179_));
 sg13g2_nand2_1 _4130_ (.Y(_1180_),
    .A(net1209),
    .B(net1211));
 sg13g2_a21oi_1 _4131_ (.A1(_1177_),
    .A2(_1179_),
    .Y(_1181_),
    .B1(net1224));
 sg13g2_nand2_2 _4132_ (.Y(_1182_),
    .A(_1173_),
    .B(_1178_));
 sg13g2_a21oi_1 _4133_ (.A1(net1224),
    .A2(_1182_),
    .Y(_1183_),
    .B1(_1181_));
 sg13g2_a21o_1 _4134_ (.A2(_1178_),
    .A1(net1211),
    .B1(_1164_),
    .X(_1184_));
 sg13g2_nand2_1 _4135_ (.Y(_1185_),
    .A(_1167_),
    .B(_1184_));
 sg13g2_and2_1 _4136_ (.A(_0904_),
    .B(net1194),
    .X(_1186_));
 sg13g2_nand2_2 _4137_ (.Y(_1187_),
    .A(_0904_),
    .B(net1194));
 sg13g2_nor2_1 _4138_ (.A(_1183_),
    .B(_1187_),
    .Y(_1188_));
 sg13g2_a21oi_1 _4139_ (.A1(_1185_),
    .A2(_1188_),
    .Y(_1189_),
    .B1(_1174_));
 sg13g2_xnor2_1 _4140_ (.Y(_1190_),
    .A(net1219),
    .B(_1162_));
 sg13g2_nand2b_1 _4141_ (.Y(_1191_),
    .B(_1184_),
    .A_N(_1167_));
 sg13g2_nand2_1 _4142_ (.Y(_1192_),
    .A(_1167_),
    .B(_1178_));
 sg13g2_a21oi_1 _4143_ (.A1(_1191_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(_0904_));
 sg13g2_xnor2_1 _4144_ (.Y(_1194_),
    .A(net1211),
    .B(net1216));
 sg13g2_o21ai_1 _4145_ (.B1(_1167_),
    .Y(_1195_),
    .A1(net1213),
    .A2(_1194_));
 sg13g2_a21oi_1 _4146_ (.A1(_1191_),
    .A2(_1195_),
    .Y(_1196_),
    .B1(net1225));
 sg13g2_or2_1 _4147_ (.X(_1197_),
    .B(_1196_),
    .A(_1193_));
 sg13g2_a21oi_1 _4148_ (.A1(_1171_),
    .A2(_1186_),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_o21ai_1 _4149_ (.B1(_1190_),
    .Y(_1199_),
    .A1(_1175_),
    .A2(_1198_));
 sg13g2_a21oi_1 _4150_ (.A1(_1175_),
    .A2(_1189_),
    .Y(_1200_),
    .B1(_1199_));
 sg13g2_o21ai_1 _4151_ (.B1(_1168_),
    .Y(_1201_),
    .A1(net1214),
    .A2(_1180_));
 sg13g2_nand2_1 _4152_ (.Y(_1202_),
    .A(net1221),
    .B(_1186_));
 sg13g2_nor2_1 _4153_ (.A(net1224),
    .B(_1182_),
    .Y(_1203_));
 sg13g2_o21ai_1 _4154_ (.B1(net1194),
    .Y(_1204_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_o21ai_1 _4155_ (.B1(net1209),
    .Y(_1205_),
    .A1(net1213),
    .A2(net1216));
 sg13g2_a21oi_1 _4156_ (.A1(net1213),
    .A2(net1216),
    .Y(_1206_),
    .B1(_1140_));
 sg13g2_nand2_1 _4157_ (.Y(_1207_),
    .A(net1221),
    .B(net1224));
 sg13g2_a21oi_1 _4158_ (.A1(_1205_),
    .A2(_1206_),
    .Y(_1208_),
    .B1(_1207_));
 sg13g2_nor2_1 _4159_ (.A(_1186_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_o21ai_1 _4160_ (.B1(_1209_),
    .Y(_1210_),
    .A1(_1171_),
    .A2(_1176_));
 sg13g2_nor2_1 _4161_ (.A(net1221),
    .B(_1187_),
    .Y(_1211_));
 sg13g2_nand3_1 _4162_ (.B(_1169_),
    .C(_1182_),
    .A(net1224),
    .Y(_1212_));
 sg13g2_a22oi_1 _4163_ (.Y(_1213_),
    .B1(_1211_),
    .B2(_1212_),
    .A2(_1204_),
    .A1(_1201_));
 sg13g2_a21oi_1 _4164_ (.A1(_1210_),
    .A2(_1213_),
    .Y(_1214_),
    .B1(_1190_));
 sg13g2_a22oi_1 _4165_ (.Y(_1215_),
    .B1(_1181_),
    .B2(_1185_),
    .A2(_1170_),
    .A1(net1225));
 sg13g2_nor2_1 _4166_ (.A(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_o21ai_1 _4167_ (.B1(_1176_),
    .Y(_1217_),
    .A1(_1174_),
    .A2(_1216_));
 sg13g2_nor2_1 _4168_ (.A(net1224),
    .B(_1177_),
    .Y(_1218_));
 sg13g2_nand3_1 _4169_ (.B(_1167_),
    .C(_1172_),
    .A(_0909_),
    .Y(_1219_));
 sg13g2_nand2_1 _4170_ (.Y(_1220_),
    .A(_1182_),
    .B(_1219_));
 sg13g2_o21ai_1 _4171_ (.B1(_1220_),
    .Y(_1221_),
    .A1(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .A2(_1218_));
 sg13g2_a21oi_1 _4172_ (.A1(_1171_),
    .A2(_1186_),
    .Y(_1222_),
    .B1(_1176_));
 sg13g2_nand2_1 _4173_ (.Y(_1223_),
    .A(_1163_),
    .B(_1190_));
 sg13g2_a21oi_1 _4174_ (.A1(_1221_),
    .A2(_1222_),
    .Y(_1224_),
    .B1(_1223_));
 sg13g2_nor3_1 _4175_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(net1207),
    .C(_0716_),
    .Y(_1225_));
 sg13g2_nand2_1 _4176_ (.Y(_1226_),
    .A(net1213),
    .B(_1179_));
 sg13g2_nand4_1 _4177_ (.B(_1166_),
    .C(_1225_),
    .A(net1228),
    .Y(_1227_),
    .D(_1226_));
 sg13g2_nor4_1 _4178_ (.A(_0900_),
    .B(_1135_),
    .C(_1214_),
    .D(_1227_),
    .Y(_1228_));
 sg13g2_o21ai_1 _4179_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_1163_),
    .A2(_1200_));
 sg13g2_a21oi_1 _4180_ (.A1(_1217_),
    .A2(_1224_),
    .Y(_1230_),
    .B1(_1229_));
 sg13g2_nor2_1 _4181_ (.A(_1160_),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_nor2_1 _4182_ (.A(_1135_),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_nor2b_1 _4183_ (.A(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .B_N(net1215),
    .Y(_1233_));
 sg13g2_nand2b_1 _4184_ (.Y(_1234_),
    .B(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .A_N(net1215));
 sg13g2_nor2b_1 _4185_ (.A(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .B_N(net1217),
    .Y(_1235_));
 sg13g2_a21oi_1 _4186_ (.A1(_1234_),
    .A2(_1235_),
    .Y(_1236_),
    .B1(_1233_));
 sg13g2_nand2_1 _4187_ (.Y(_1237_),
    .A(_1194_),
    .B(_1236_));
 sg13g2_nand2_1 _4188_ (.Y(_1238_),
    .A(_1172_),
    .B(_1237_));
 sg13g2_xor2_1 _4189_ (.B(_1238_),
    .A(net1214),
    .X(_1239_));
 sg13g2_xnor2_1 _4190_ (.Y(_1240_),
    .A(_1194_),
    .B(_1236_));
 sg13g2_nand2_2 _4191_ (.Y(_1241_),
    .A(_1239_),
    .B(_1240_));
 sg13g2_nor2_1 _4192_ (.A(_1239_),
    .B(_1240_),
    .Y(_1242_));
 sg13g2_nand3b_1 _4193_ (.B(net1211),
    .C(_1241_),
    .Y(_1243_),
    .A_N(_1242_));
 sg13g2_nand4_1 _4194_ (.B(net1209),
    .C(_0801_),
    .A(_0625_),
    .Y(_1244_),
    .D(_0898_));
 sg13g2_a21oi_1 _4195_ (.A1(_1175_),
    .A2(_1187_),
    .Y(_1245_),
    .B1(_1244_));
 sg13g2_a21oi_2 _4196_ (.B1(net1220),
    .Y(_1246_),
    .A2(_1147_),
    .A1(net1221));
 sg13g2_nor2_1 _4197_ (.A(_1078_),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_a21oi_1 _4198_ (.A1(_0920_),
    .A2(_1246_),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_nand3_1 _4199_ (.B(_1245_),
    .C(_1248_),
    .A(_1243_),
    .Y(_1249_));
 sg13g2_a21oi_2 _4200_ (.B1(_1246_),
    .Y(_1250_),
    .A2(net1194),
    .A1(_0967_));
 sg13g2_nand2_2 _4201_ (.Y(_1251_),
    .A(_0629_),
    .B(_1250_));
 sg13g2_xnor2_1 _4202_ (.Y(_1252_),
    .A(_0629_),
    .B(_1246_));
 sg13g2_inv_2 _4203_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_nor2_2 _4204_ (.A(_1250_),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_o21ai_1 _4205_ (.B1(_1253_),
    .Y(_1255_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .A2(_1250_));
 sg13g2_and2_1 _4206_ (.A(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .B(_1250_),
    .X(_1256_));
 sg13g2_a22oi_1 _4207_ (.Y(_1257_),
    .B1(_1256_),
    .B2(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .A2(_1254_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[2] ));
 sg13g2_nand2_1 _4208_ (.Y(_1258_),
    .A(_1255_),
    .B(_1257_));
 sg13g2_o21ai_1 _4209_ (.B1(_1258_),
    .Y(_1259_),
    .A1(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .A2(_1251_));
 sg13g2_or2_1 _4210_ (.X(_1260_),
    .B(_1259_),
    .A(_1249_));
 sg13g2_inv_1 _4211_ (.Y(_1261_),
    .A(_1260_));
 sg13g2_o21ai_1 _4212_ (.B1(_1253_),
    .Y(_1262_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .A2(_1250_));
 sg13g2_a22oi_1 _4213_ (.Y(_1263_),
    .B1(_1256_),
    .B2(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .A2(_1254_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[3] ));
 sg13g2_nand2_1 _4214_ (.Y(_1264_),
    .A(_1262_),
    .B(_1263_));
 sg13g2_o21ai_1 _4215_ (.B1(_1264_),
    .Y(_1265_),
    .A1(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .A2(_1251_));
 sg13g2_nor2_2 _4216_ (.A(_1249_),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_inv_1 _4217_ (.Y(_1267_),
    .A(_1266_));
 sg13g2_nor2_1 _4218_ (.A(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .B(_1251_),
    .Y(_1268_));
 sg13g2_o21ai_1 _4219_ (.B1(_1253_),
    .Y(_1269_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .A2(_1250_));
 sg13g2_a22oi_1 _4220_ (.Y(_1270_),
    .B1(_1256_),
    .B2(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .A2(_1254_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[1] ));
 sg13g2_a21oi_2 _4221_ (.B1(_1268_),
    .Y(_1271_),
    .A2(_1270_),
    .A1(_1269_));
 sg13g2_inv_1 _4222_ (.Y(_1272_),
    .A(_1271_));
 sg13g2_nor2_1 _4223_ (.A(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .B(_1251_),
    .Y(_1273_));
 sg13g2_o21ai_1 _4224_ (.B1(_1253_),
    .Y(_1274_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .A2(_1250_));
 sg13g2_a22oi_1 _4225_ (.Y(_1275_),
    .B1(_1256_),
    .B2(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .A2(_1254_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[0] ));
 sg13g2_a21oi_1 _4226_ (.A1(_1274_),
    .A2(_1275_),
    .Y(_1276_),
    .B1(_1273_));
 sg13g2_nand2b_2 _4227_ (.Y(_1277_),
    .B(_1276_),
    .A_N(_1249_));
 sg13g2_nor2_1 _4228_ (.A(_1272_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_nand2b_1 _4229_ (.Y(_1279_),
    .B(_1271_),
    .A_N(_1249_));
 sg13g2_and2_1 _4230_ (.A(_1277_),
    .B(_1279_),
    .X(_1280_));
 sg13g2_nor2_1 _4231_ (.A(_1278_),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_nor3_1 _4232_ (.A(_1260_),
    .B(_1266_),
    .C(_1281_),
    .Y(_1282_));
 sg13g2_nor3_1 _4233_ (.A(_0627_),
    .B(_1241_),
    .C(_1282_),
    .Y(_1283_));
 sg13g2_and2_1 _4234_ (.A(_0627_),
    .B(_1240_),
    .X(_1284_));
 sg13g2_inv_1 _4235_ (.Y(_1285_),
    .A(_1284_));
 sg13g2_o21ai_1 _4236_ (.B1(_1243_),
    .Y(_1286_),
    .A1(net1211),
    .A2(_1241_));
 sg13g2_nor2_1 _4237_ (.A(_1239_),
    .B(_1285_),
    .Y(_1287_));
 sg13g2_nand2_1 _4238_ (.Y(_1288_),
    .A(_1260_),
    .B(_1279_));
 sg13g2_nor2_1 _4239_ (.A(_1271_),
    .B(_1277_),
    .Y(_1289_));
 sg13g2_inv_1 _4240_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_nand2_1 _4241_ (.Y(_1291_),
    .A(_1260_),
    .B(_1290_));
 sg13g2_or2_1 _4242_ (.X(_1292_),
    .B(_1278_),
    .A(_1260_));
 sg13g2_a21oi_1 _4243_ (.A1(_1291_),
    .A2(_1292_),
    .Y(_1293_),
    .B1(_1266_));
 sg13g2_xnor2_1 _4244_ (.Y(_1294_),
    .A(_1288_),
    .B(_1293_));
 sg13g2_nor3_1 _4245_ (.A(_1261_),
    .B(_1266_),
    .C(_1290_),
    .Y(_1295_));
 sg13g2_a21oi_1 _4246_ (.A1(net1211),
    .A2(_1239_),
    .Y(_1296_),
    .B1(_1240_));
 sg13g2_a221oi_1 _4247_ (.B2(_1296_),
    .C1(_1186_),
    .B1(_1295_),
    .A1(_1287_),
    .Y(_1297_),
    .A2(_1294_));
 sg13g2_nand3_1 _4248_ (.B(_1291_),
    .C(_1292_),
    .A(_1267_),
    .Y(_1298_));
 sg13g2_nand2_1 _4249_ (.Y(_1299_),
    .A(_1287_),
    .B(_1298_));
 sg13g2_o21ai_1 _4250_ (.B1(_1277_),
    .Y(_1300_),
    .A1(_1260_),
    .A2(_1271_));
 sg13g2_a22oi_1 _4251_ (.Y(_1301_),
    .B1(_1300_),
    .B2(_1267_),
    .A2(_1289_),
    .A1(_1260_));
 sg13g2_nand3b_1 _4252_ (.B(_1239_),
    .C(_0627_),
    .Y(_1302_),
    .A_N(_1240_));
 sg13g2_nor2_1 _4253_ (.A(_1266_),
    .B(_1280_),
    .Y(_1303_));
 sg13g2_a21oi_1 _4254_ (.A1(_1292_),
    .A2(_1303_),
    .Y(_1304_),
    .B1(_1302_));
 sg13g2_or2_1 _4255_ (.X(_1305_),
    .B(_1304_),
    .A(_1202_));
 sg13g2_a21oi_1 _4256_ (.A1(_1242_),
    .A2(_1301_),
    .Y(_1306_),
    .B1(_1305_));
 sg13g2_a21oi_1 _4257_ (.A1(_1299_),
    .A2(_1306_),
    .Y(_1307_),
    .B1(_1297_));
 sg13g2_nor3_1 _4258_ (.A(_1283_),
    .B(_1286_),
    .C(_1307_),
    .Y(_1308_));
 sg13g2_a221oi_1 _4259_ (.B2(_1281_),
    .C1(_1240_),
    .B1(_1267_),
    .A1(net1212),
    .Y(_1309_),
    .A2(_1239_));
 sg13g2_a21oi_1 _4260_ (.A1(_1243_),
    .A2(_1285_),
    .Y(_1310_),
    .B1(_1295_));
 sg13g2_o21ai_1 _4261_ (.B1(_1211_),
    .Y(_1311_),
    .A1(_0627_),
    .A2(_1241_));
 sg13g2_a21oi_1 _4262_ (.A1(_1242_),
    .A2(_1261_),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_o21ai_1 _4263_ (.B1(_1312_),
    .Y(_1313_),
    .A1(_1291_),
    .A2(_1302_));
 sg13g2_nor3_1 _4264_ (.A(_1309_),
    .B(_1310_),
    .C(_1313_),
    .Y(_1314_));
 sg13g2_nand3_1 _4265_ (.B(_1280_),
    .C(_1286_),
    .A(_1187_),
    .Y(_1315_));
 sg13g2_nor3_1 _4266_ (.A(_1260_),
    .B(_1266_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_or4_1 _4267_ (.A(_0902_),
    .B(_1135_),
    .C(_1160_),
    .D(_1249_),
    .X(_1317_));
 sg13g2_nor4_1 _4268_ (.A(_1308_),
    .B(_1314_),
    .C(_1316_),
    .D(_1317_),
    .Y(_1318_));
 sg13g2_or2_1 _4269_ (.X(_1319_),
    .B(_1318_),
    .A(_1232_));
 sg13g2_or2_1 _4270_ (.X(uo_out[4]),
    .B(_1319_),
    .A(_1138_));
 sg13g2_nand2_1 _4271_ (.Y(_1320_),
    .A(\vga_tetris.boardMem.board_12[3] ),
    .B(net1016));
 sg13g2_a22oi_1 _4272_ (.Y(_1321_),
    .B1(net998),
    .B2(\vga_tetris.boardMem.board_7[3] ),
    .A2(net1008),
    .A1(\vga_tetris.boardMem.board_9[3] ));
 sg13g2_a22oi_1 _4273_ (.Y(_1322_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_3[3] ),
    .A2(net1010),
    .A1(\vga_tetris.boardMem.board_14[3] ));
 sg13g2_nand2_1 _4274_ (.Y(_1323_),
    .A(_1320_),
    .B(_1322_));
 sg13g2_a22oi_1 _4275_ (.Y(_1324_),
    .B1(net996),
    .B2(\vga_tetris.boardMem.board_4[3] ),
    .A2(net1012),
    .A1(\vga_tetris.boardMem.board_6[3] ));
 sg13g2_a22oi_1 _4276_ (.Y(_1325_),
    .B1(net990),
    .B2(\vga_tetris.boardMem.board_2[3] ),
    .A2(net1018),
    .A1(\vga_tetris.boardMem.board_5[3] ));
 sg13g2_a22oi_1 _4277_ (.Y(_1326_),
    .B1(net1002),
    .B2(\vga_tetris.boardMem.board_10[3] ),
    .A2(net1024),
    .A1(\vga_tetris.boardMem.board_15[3] ));
 sg13g2_a22oi_1 _4278_ (.Y(_1327_),
    .B1(net994),
    .B2(\vga_tetris.boardMem.board_13[3] ),
    .A2(net1022),
    .A1(\vga_tetris.boardMem.board_17[3] ));
 sg13g2_a22oi_1 _4279_ (.Y(_1328_),
    .B1(net1014),
    .B2(\vga_tetris.boardMem.board_16[3] ),
    .A2(net1020),
    .A1(\vga_tetris.boardMem.board_1[3] ));
 sg13g2_nand4_1 _4280_ (.B(_1326_),
    .C(_1327_),
    .A(_1325_),
    .Y(_1329_),
    .D(_1328_));
 sg13g2_a22oi_1 _4281_ (.Y(_1330_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_18[3] ),
    .A2(net1006),
    .A1(\vga_tetris.boardMem.board_8[3] ));
 sg13g2_a22oi_1 _4282_ (.Y(_1331_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_19[3] ),
    .A2(net1004),
    .A1(\vga_tetris.boardMem.board_11[3] ));
 sg13g2_nand4_1 _4283_ (.B(_1324_),
    .C(_1330_),
    .A(_1321_),
    .Y(_1332_),
    .D(_1331_));
 sg13g2_or4_1 _4284_ (.A(net845),
    .B(_1323_),
    .C(_1329_),
    .D(_1332_),
    .X(_1333_));
 sg13g2_a21oi_1 _4285_ (.A1(_0676_),
    .A2(net847),
    .Y(_1334_),
    .B1(net1085));
 sg13g2_nand2_2 _4286_ (.Y(_1335_),
    .A(_1333_),
    .B(_1334_));
 sg13g2_nand3_1 _4287_ (.B(net1062),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_2[5] ),
    .Y(_1336_));
 sg13g2_nand3_1 _4288_ (.B(net1053),
    .C(net1045),
    .A(\vga_tetris.boardMem.board_5[5] ),
    .Y(_1337_));
 sg13g2_nand3_1 _4289_ (.B(net1051),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_9[5] ),
    .Y(_1338_));
 sg13g2_nand3_1 _4290_ (.B(net1069),
    .C(net1045),
    .A(\vga_tetris.boardMem.board_7[5] ),
    .Y(_1339_));
 sg13g2_nand3_1 _4291_ (.B(net1033),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_10[5] ),
    .Y(_1340_));
 sg13g2_nand3_1 _4292_ (.B(net1074),
    .C(net1069),
    .A(\vga_tetris.boardMem.board_15[5] ),
    .Y(_1341_));
 sg13g2_nand3_1 _4293_ (.B(net1057),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[5] ),
    .Y(_1342_));
 sg13g2_nand3_1 _4294_ (.B(net1074),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_12[5] ),
    .Y(_1343_));
 sg13g2_nand3_1 _4295_ (.B(net1059),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[5] ),
    .Y(_1344_));
 sg13g2_nand3_1 _4296_ (.B(net1045),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_6[5] ),
    .Y(_1345_));
 sg13g2_nand3_1 _4297_ (.B(_0839_),
    .C(net1057),
    .A(\vga_tetris.boardMem.board_17[5] ),
    .Y(_1346_));
 sg13g2_nand3_1 _4298_ (.B(net1074),
    .C(net1053),
    .A(\vga_tetris.boardMem.board_13[5] ),
    .Y(_1347_));
 sg13g2_nand3_1 _4299_ (.B(net1069),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_11[5] ),
    .Y(_1348_));
 sg13g2_nand3_1 _4300_ (.B(net1066),
    .C(net1062),
    .A(\vga_tetris.boardMem.board_3[5] ),
    .Y(_1349_));
 sg13g2_nand3_1 _4301_ (.B(net1040),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_8[5] ),
    .Y(_1350_));
 sg13g2_nand3_1 _4302_ (.B(net1045),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_4[5] ),
    .Y(_1351_));
 sg13g2_and3_1 _4303_ (.X(_1352_),
    .A(\vga_tetris.boardMem.board_14[5] ),
    .B(net1078),
    .C(net1037));
 sg13g2_nand4_1 _4304_ (.B(_1338_),
    .C(_1340_),
    .A(_1336_),
    .Y(_1353_),
    .D(_1343_));
 sg13g2_a21oi_1 _4305_ (.A1(net986),
    .A2(net985),
    .Y(_1354_),
    .B1(_1353_));
 sg13g2_and4_1 _4306_ (.A(_1341_),
    .B(_1344_),
    .C(_1346_),
    .D(_1349_),
    .X(_1355_));
 sg13g2_and4_1 _4307_ (.A(_1339_),
    .B(_1342_),
    .C(_1348_),
    .D(_1350_),
    .X(_1356_));
 sg13g2_a221oi_1 _4308_ (.B2(\vga_tetris.boardMem.board_19[5] ),
    .C1(_1352_),
    .B1(net987),
    .A1(\vga_tetris.boardMem.board_1[5] ),
    .Y(_1357_),
    .A2(net1019));
 sg13g2_and4_1 _4309_ (.A(_1337_),
    .B(_1345_),
    .C(_1347_),
    .D(_1351_),
    .X(_1358_));
 sg13g2_and4_1 _4310_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .D(_1358_),
    .X(_1359_));
 sg13g2_a221oi_1 _4311_ (.B2(_1359_),
    .C1(net1083),
    .B1(_1354_),
    .A1(_0678_),
    .Y(_1360_),
    .A2(net843));
 sg13g2_nand3_1 _4312_ (.B(_0920_),
    .C(_1360_),
    .A(_0918_),
    .Y(_1361_));
 sg13g2_o21ai_1 _4313_ (.B1(_1361_),
    .Y(_1362_),
    .A1(_0922_),
    .A2(_1335_));
 sg13g2_nand3_1 _4314_ (.B(net1057),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[7] ),
    .Y(_1363_));
 sg13g2_nand3_1 _4315_ (.B(net1053),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_9[7] ),
    .Y(_1364_));
 sg13g2_nand3_1 _4316_ (.B(net1046),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_6[7] ),
    .Y(_1365_));
 sg13g2_nand3_1 _4317_ (.B(net1039),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_8[7] ),
    .Y(_1366_));
 sg13g2_nand3_1 _4318_ (.B(net1067),
    .C(net1063),
    .A(\vga_tetris.boardMem.board_3[7] ),
    .Y(_1367_));
 sg13g2_nand3_1 _4319_ (.B(net1067),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_7[7] ),
    .Y(_1368_));
 sg13g2_nand3_1 _4320_ (.B(net1034),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_10[7] ),
    .Y(_1369_));
 sg13g2_nand3_1 _4321_ (.B(net1060),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[7] ),
    .Y(_1370_));
 sg13g2_nand3_1 _4322_ (.B(net1068),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_11[7] ),
    .Y(_1371_));
 sg13g2_nand3_1 _4323_ (.B(net1052),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_5[7] ),
    .Y(_1372_));
 sg13g2_nand3_1 _4324_ (.B(net1073),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_12[7] ),
    .Y(_1373_));
 sg13g2_nand3_1 _4325_ (.B(net1046),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_4[7] ),
    .Y(_1374_));
 sg13g2_nand3_1 _4326_ (.B(net1073),
    .C(net1051),
    .A(\vga_tetris.boardMem.board_13[7] ),
    .Y(_1375_));
 sg13g2_nand3_1 _4327_ (.B(net1062),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_2[7] ),
    .Y(_1376_));
 sg13g2_nand3_1 _4328_ (.B(net1075),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_14[7] ),
    .Y(_1377_));
 sg13g2_nand3_1 _4329_ (.B(_0836_),
    .C(net1060),
    .A(\vga_tetris.boardMem.board_19[7] ),
    .Y(_1378_));
 sg13g2_nand3_1 _4330_ (.B(net1075),
    .C(net1067),
    .A(\vga_tetris.boardMem.board_15[7] ),
    .Y(_1379_));
 sg13g2_nand3_1 _4331_ (.B(_0839_),
    .C(net1060),
    .A(\vga_tetris.boardMem.board_17[7] ),
    .Y(_1380_));
 sg13g2_nand3_1 _4332_ (.B(net1062),
    .C(net1052),
    .A(\vga_tetris.boardMem.board_1[7] ),
    .Y(_1381_));
 sg13g2_nand4_1 _4333_ (.B(_1370_),
    .C(_1371_),
    .A(_1364_),
    .Y(_1382_),
    .D(_1380_));
 sg13g2_a21oi_1 _4334_ (.A1(net986),
    .A2(net985),
    .Y(_1383_),
    .B1(_1382_));
 sg13g2_nand4_1 _4335_ (.B(_1368_),
    .C(_1369_),
    .A(_1367_),
    .Y(_1384_),
    .D(_1379_));
 sg13g2_nand4_1 _4336_ (.B(_1373_),
    .C(_1375_),
    .A(_1365_),
    .Y(_1385_),
    .D(_1376_));
 sg13g2_nand3_1 _4337_ (.B(_1372_),
    .C(_1378_),
    .A(_1366_),
    .Y(_1386_));
 sg13g2_nand4_1 _4338_ (.B(_1374_),
    .C(_1377_),
    .A(_1363_),
    .Y(_1387_),
    .D(_1381_));
 sg13g2_nor4_2 _4339_ (.A(_1384_),
    .B(_1385_),
    .C(_1386_),
    .Y(_1388_),
    .D(_1387_));
 sg13g2_a221oi_1 _4340_ (.B2(_1388_),
    .C1(net1083),
    .B1(_1383_),
    .A1(_0680_),
    .Y(_1389_),
    .A2(net843));
 sg13g2_nand3_1 _4341_ (.B(_0967_),
    .C(_1389_),
    .A(_0920_),
    .Y(_1390_));
 sg13g2_a22oi_1 _4342_ (.Y(_1391_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[13] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[13] ));
 sg13g2_nand2_1 _4343_ (.Y(_1392_),
    .A(\vga_tetris.boardMem.board_9[13] ),
    .B(net1007));
 sg13g2_a22oi_1 _4344_ (.Y(_1393_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[13] ),
    .A2(net1005),
    .A1(\vga_tetris.boardMem.board_8[13] ));
 sg13g2_a22oi_1 _4345_ (.Y(_1394_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[13] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[13] ));
 sg13g2_nand2_1 _4346_ (.Y(_1395_),
    .A(_1392_),
    .B(_1394_));
 sg13g2_a22oi_1 _4347_ (.Y(_1396_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[13] ),
    .A2(net1011),
    .A1(\vga_tetris.boardMem.board_6[13] ));
 sg13g2_a22oi_1 _4348_ (.Y(_1397_),
    .B1(net1003),
    .B2(\vga_tetris.boardMem.board_11[13] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[13] ));
 sg13g2_a22oi_1 _4349_ (.Y(_1398_),
    .B1(net1000),
    .B2(\vga_tetris.boardMem.board_18[13] ),
    .A2(net1015),
    .A1(\vga_tetris.boardMem.board_12[13] ));
 sg13g2_a22oi_1 _4350_ (.Y(_1399_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[13] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[13] ));
 sg13g2_a22oi_1 _4351_ (.Y(_1400_),
    .B1(net1021),
    .B2(\vga_tetris.boardMem.board_17[13] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[13] ));
 sg13g2_nand4_1 _4352_ (.B(_1398_),
    .C(_1399_),
    .A(_1397_),
    .Y(_1401_),
    .D(_1400_));
 sg13g2_a22oi_1 _4353_ (.Y(_1402_),
    .B1(net997),
    .B2(\vga_tetris.boardMem.board_7[13] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_10[13] ));
 sg13g2_nand4_1 _4354_ (.B(_1393_),
    .C(_1396_),
    .A(_1391_),
    .Y(_1403_),
    .D(_1402_));
 sg13g2_or4_1 _4355_ (.A(net844),
    .B(_1395_),
    .C(_1401_),
    .D(_1403_),
    .X(_1404_));
 sg13g2_a21oi_2 _4356_ (.B1(net1085),
    .Y(_1405_),
    .A2(net844),
    .A1(_0686_));
 sg13g2_nand2_1 _4357_ (.Y(_1406_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_and4_1 _4358_ (.A(_0917_),
    .B(_0918_),
    .C(_1404_),
    .D(_1405_),
    .X(_1407_));
 sg13g2_nand2_1 _4359_ (.Y(_1408_),
    .A(\vga_tetris.boardMem.board_6[1] ),
    .B(net1012));
 sg13g2_a22oi_1 _4360_ (.Y(_1409_),
    .B1(net994),
    .B2(\vga_tetris.boardMem.board_13[1] ),
    .A2(net996),
    .A1(\vga_tetris.boardMem.board_4[1] ));
 sg13g2_a22oi_1 _4361_ (.Y(_1410_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_19[1] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_7[1] ));
 sg13g2_nand2_1 _4362_ (.Y(_1411_),
    .A(_1408_),
    .B(_1410_));
 sg13g2_a22oi_1 _4363_ (.Y(_1412_),
    .B1(net1004),
    .B2(\vga_tetris.boardMem.board_11[1] ),
    .A2(net1016),
    .A1(\vga_tetris.boardMem.board_12[1] ));
 sg13g2_a22oi_1 _4364_ (.Y(_1413_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_3[1] ),
    .A2(net1014),
    .A1(\vga_tetris.boardMem.board_16[1] ));
 sg13g2_a22oi_1 _4365_ (.Y(_1414_),
    .B1(net1018),
    .B2(\vga_tetris.boardMem.board_5[1] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[1] ));
 sg13g2_a22oi_1 _4366_ (.Y(_1415_),
    .B1(net1010),
    .B2(\vga_tetris.boardMem.board_14[1] ),
    .A2(net1024),
    .A1(\vga_tetris.boardMem.board_15[1] ));
 sg13g2_a22oi_1 _4367_ (.Y(_1416_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_18[1] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_10[1] ));
 sg13g2_nand4_1 _4368_ (.B(_1414_),
    .C(_1415_),
    .A(_1413_),
    .Y(_1417_),
    .D(_1416_));
 sg13g2_a22oi_1 _4369_ (.Y(_1418_),
    .B1(net1005),
    .B2(\vga_tetris.boardMem.board_8[1] ),
    .A2(net1022),
    .A1(\vga_tetris.boardMem.board_17[1] ));
 sg13g2_a22oi_1 _4370_ (.Y(_1419_),
    .B1(net990),
    .B2(\vga_tetris.boardMem.board_2[1] ),
    .A2(net1008),
    .A1(\vga_tetris.boardMem.board_9[1] ));
 sg13g2_nand4_1 _4371_ (.B(_1412_),
    .C(_1418_),
    .A(_1409_),
    .Y(_1420_),
    .D(_1419_));
 sg13g2_or4_1 _4372_ (.A(net846),
    .B(_1411_),
    .C(_1417_),
    .D(_1420_),
    .X(_1421_));
 sg13g2_a21oi_1 _4373_ (.A1(_0674_),
    .A2(net846),
    .Y(_1422_),
    .B1(net1084));
 sg13g2_nand2_2 _4374_ (.Y(_1423_),
    .A(_1421_),
    .B(_1422_));
 sg13g2_inv_1 _4375_ (.Y(_1424_),
    .A(_1423_));
 sg13g2_nand3_1 _4376_ (.B(net1041),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_8[19] ),
    .Y(_1425_));
 sg13g2_nand3_1 _4377_ (.B(net1058),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[19] ),
    .Y(_1426_));
 sg13g2_nand3_1 _4378_ (.B(net1064),
    .C(net1036),
    .A(\vga_tetris.boardMem.board_2[19] ),
    .Y(_1427_));
 sg13g2_and3_1 _4379_ (.X(_1428_),
    .A(\vga_tetris.boardMem.board_12[19] ),
    .B(net1077),
    .C(net1041));
 sg13g2_nand3_1 _4380_ (.B(net1049),
    .C(net1036),
    .A(\vga_tetris.boardMem.board_6[19] ),
    .Y(_1429_));
 sg13g2_nand3_1 _4381_ (.B(net1065),
    .C(net1055),
    .A(\vga_tetris.boardMem.board_1[19] ),
    .Y(_1430_));
 sg13g2_nand3_1 _4382_ (.B(_0836_),
    .C(net1058),
    .A(\vga_tetris.boardMem.board_19[19] ),
    .Y(_1431_));
 sg13g2_nand3_1 _4383_ (.B(net1049),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_4[19] ),
    .Y(_1432_));
 sg13g2_nand3_1 _4384_ (.B(net1077),
    .C(net1036),
    .A(\vga_tetris.boardMem.board_14[19] ),
    .Y(_1433_));
 sg13g2_nand3_1 _4385_ (.B(net1054),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_9[19] ),
    .Y(_1434_));
 sg13g2_nand3_1 _4386_ (.B(net1077),
    .C(net1070),
    .A(\vga_tetris.boardMem.board_15[19] ),
    .Y(_1435_));
 sg13g2_nand3_1 _4387_ (.B(net1070),
    .C(net1064),
    .A(\vga_tetris.boardMem.board_3[19] ),
    .Y(_1436_));
 sg13g2_nand3_1 _4388_ (.B(net1070),
    .C(net1049),
    .A(\vga_tetris.boardMem.board_7[19] ),
    .Y(_1437_));
 sg13g2_nand3_1 _4389_ (.B(net1070),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_11[19] ),
    .Y(_1438_));
 sg13g2_nand3_1 _4390_ (.B(net1054),
    .C(net1049),
    .A(\vga_tetris.boardMem.board_5[19] ),
    .Y(_1439_));
 sg13g2_nand3_1 _4391_ (.B(net1077),
    .C(net1054),
    .A(\vga_tetris.boardMem.board_13[19] ),
    .Y(_1440_));
 sg13g2_nand3_1 _4392_ (.B(net1036),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_10[19] ),
    .Y(_1441_));
 sg13g2_nand4_1 _4393_ (.B(_1430_),
    .C(_1432_),
    .A(_1429_),
    .Y(_1442_),
    .D(_1439_));
 sg13g2_a21oi_1 _4394_ (.A1(_0871_),
    .A2(_0874_),
    .Y(_1443_),
    .B1(_1442_));
 sg13g2_and4_1 _4395_ (.A(_1425_),
    .B(_1431_),
    .C(_1433_),
    .D(_1440_),
    .X(_1444_));
 sg13g2_and4_1 _4396_ (.A(_1434_),
    .B(_1436_),
    .C(_1437_),
    .D(_1438_),
    .X(_1445_));
 sg13g2_a221oi_1 _4397_ (.B2(\vga_tetris.boardMem.board_18[19] ),
    .C1(_1428_),
    .B1(net1000),
    .A1(\vga_tetris.boardMem.board_17[19] ),
    .Y(_1446_),
    .A2(net1021));
 sg13g2_and4_1 _4398_ (.A(_1426_),
    .B(_1427_),
    .C(_1435_),
    .D(_1441_),
    .X(_1447_));
 sg13g2_and4_1 _4399_ (.A(_1444_),
    .B(_1445_),
    .C(_1446_),
    .D(_1447_),
    .X(_1448_));
 sg13g2_a221oi_1 _4400_ (.B2(_1448_),
    .C1(net1083),
    .B1(_1443_),
    .A1(_0692_),
    .Y(_1449_),
    .A2(net843));
 sg13g2_a22oi_1 _4401_ (.Y(_1450_),
    .B1(net1001),
    .B2(\vga_tetris.boardMem.board_10[9] ),
    .A2(net1019),
    .A1(\vga_tetris.boardMem.board_1[9] ));
 sg13g2_a22oi_1 _4402_ (.Y(_1451_),
    .B1(net987),
    .B2(\vga_tetris.boardMem.board_19[9] ),
    .A2(net1011),
    .A1(\vga_tetris.boardMem.board_6[9] ));
 sg13g2_nand2_1 _4403_ (.Y(_1452_),
    .A(\vga_tetris.boardMem.board_9[9] ),
    .B(net1007));
 sg13g2_a22oi_1 _4404_ (.Y(_1453_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[9] ),
    .A2(net1009),
    .A1(\vga_tetris.boardMem.board_14[9] ));
 sg13g2_a22oi_1 _4405_ (.Y(_1454_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_3[9] ),
    .A2(net1023),
    .A1(\vga_tetris.boardMem.board_15[9] ));
 sg13g2_a22oi_1 _4406_ (.Y(_1455_),
    .B1(net995),
    .B2(\vga_tetris.boardMem.board_4[9] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_7[9] ));
 sg13g2_a22oi_1 _4407_ (.Y(_1456_),
    .B1(net1000),
    .B2(\vga_tetris.boardMem.board_18[9] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[9] ));
 sg13g2_nand2_1 _4408_ (.Y(_1457_),
    .A(_1452_),
    .B(_1456_));
 sg13g2_a22oi_1 _4409_ (.Y(_1458_),
    .B1(net1003),
    .B2(\vga_tetris.boardMem.board_11[9] ),
    .A2(net1005),
    .A1(\vga_tetris.boardMem.board_8[9] ));
 sg13g2_a22oi_1 _4410_ (.Y(_1459_),
    .B1(net993),
    .B2(\vga_tetris.boardMem.board_13[9] ),
    .A2(net1013),
    .A1(\vga_tetris.boardMem.board_16[9] ));
 sg13g2_a22oi_1 _4411_ (.Y(_1460_),
    .B1(net1015),
    .B2(\vga_tetris.boardMem.board_12[9] ),
    .A2(net1021),
    .A1(\vga_tetris.boardMem.board_17[9] ));
 sg13g2_nand4_1 _4412_ (.B(_1458_),
    .C(_1459_),
    .A(_1450_),
    .Y(_1461_),
    .D(_1460_));
 sg13g2_nand4_1 _4413_ (.B(_1453_),
    .C(_1454_),
    .A(_1451_),
    .Y(_1462_),
    .D(_1455_));
 sg13g2_or4_1 _4414_ (.A(net846),
    .B(_1457_),
    .C(_1461_),
    .D(_1462_),
    .X(_1463_));
 sg13g2_a21oi_1 _4415_ (.A1(_0682_),
    .A2(net846),
    .Y(_1464_),
    .B1(net1084));
 sg13g2_and2_1 _4416_ (.A(_1463_),
    .B(_1464_),
    .X(_1465_));
 sg13g2_nand2_1 _4417_ (.Y(_1466_),
    .A(_1463_),
    .B(_1464_));
 sg13g2_nand2b_1 _4418_ (.Y(_1467_),
    .B(_1465_),
    .A_N(_1049_));
 sg13g2_a22oi_1 _4419_ (.Y(_1468_),
    .B1(net1010),
    .B2(\vga_tetris.boardMem.board_14[17] ),
    .A2(net1018),
    .A1(\vga_tetris.boardMem.board_5[17] ));
 sg13g2_a22oi_1 _4420_ (.Y(_1469_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_19[17] ),
    .A2(net1020),
    .A1(\vga_tetris.boardMem.board_1[17] ));
 sg13g2_a22oi_1 _4421_ (.Y(_1470_),
    .B1(net990),
    .B2(\vga_tetris.boardMem.board_2[17] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_7[17] ));
 sg13g2_a22oi_1 _4422_ (.Y(_1471_),
    .B1(net996),
    .B2(\vga_tetris.boardMem.board_4[17] ),
    .A2(net1022),
    .A1(\vga_tetris.boardMem.board_17[17] ));
 sg13g2_nand4_1 _4423_ (.B(_1469_),
    .C(_1470_),
    .A(_1468_),
    .Y(_1472_),
    .D(_1471_));
 sg13g2_a22oi_1 _4424_ (.Y(_1473_),
    .B1(net1008),
    .B2(\vga_tetris.boardMem.board_9[17] ),
    .A2(net1016),
    .A1(\vga_tetris.boardMem.board_12[17] ));
 sg13g2_a22oi_1 _4425_ (.Y(_1474_),
    .B1(net994),
    .B2(\vga_tetris.boardMem.board_13[17] ),
    .A2(net1014),
    .A1(\vga_tetris.boardMem.board_16[17] ));
 sg13g2_a22oi_1 _4426_ (.Y(_1475_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_3[17] ),
    .A2(net1012),
    .A1(\vga_tetris.boardMem.board_6[17] ));
 sg13g2_a22oi_1 _4427_ (.Y(_1476_),
    .B1(net1004),
    .B2(\vga_tetris.boardMem.board_11[17] ),
    .A2(net1024),
    .A1(\vga_tetris.boardMem.board_15[17] ));
 sg13g2_and4_1 _4428_ (.A(_1473_),
    .B(_1474_),
    .C(_1475_),
    .D(_1476_),
    .X(_1477_));
 sg13g2_nand2_1 _4429_ (.Y(_1478_),
    .A(\vga_tetris.boardMem.board_8[17] ),
    .B(net1006));
 sg13g2_a22oi_1 _4430_ (.Y(_1479_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_18[17] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_10[17] ));
 sg13g2_nand4_1 _4431_ (.B(_1477_),
    .C(_1478_),
    .A(_0876_),
    .Y(_1480_),
    .D(_1479_));
 sg13g2_a21oi_1 _4432_ (.A1(_0690_),
    .A2(net845),
    .Y(_1481_),
    .B1(net1085));
 sg13g2_o21ai_1 _4433_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_1472_),
    .A2(_1480_));
 sg13g2_nor2_1 _4434_ (.A(_1096_),
    .B(_1482_),
    .Y(_1483_));
 sg13g2_a22oi_1 _4435_ (.Y(_1484_),
    .B1(net994),
    .B2(\vga_tetris.boardMem.board_13[15] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_7[15] ));
 sg13g2_a22oi_1 _4436_ (.Y(_1485_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_3[15] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_10[15] ));
 sg13g2_nand2_1 _4437_ (.Y(_1486_),
    .A(\vga_tetris.boardMem.board_16[15] ),
    .B(net1013));
 sg13g2_a22oi_1 _4438_ (.Y(_1487_),
    .B1(net1004),
    .B2(\vga_tetris.boardMem.board_11[15] ),
    .A2(net1024),
    .A1(\vga_tetris.boardMem.board_15[15] ));
 sg13g2_a22oi_1 _4439_ (.Y(_1488_),
    .B1(net996),
    .B2(\vga_tetris.boardMem.board_4[15] ),
    .A2(net1010),
    .A1(\vga_tetris.boardMem.board_14[15] ));
 sg13g2_a22oi_1 _4440_ (.Y(_1489_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_2[15] ),
    .A2(net1022),
    .A1(\vga_tetris.boardMem.board_17[15] ));
 sg13g2_a22oi_1 _4441_ (.Y(_1490_),
    .B1(net1011),
    .B2(\vga_tetris.boardMem.board_6[15] ),
    .A2(net1016),
    .A1(\vga_tetris.boardMem.board_12[15] ));
 sg13g2_nand4_1 _4442_ (.B(_1488_),
    .C(_1489_),
    .A(_1487_),
    .Y(_1491_),
    .D(_1490_));
 sg13g2_nand2_1 _4443_ (.Y(_1492_),
    .A(_1484_),
    .B(_1486_));
 sg13g2_a22oi_1 _4444_ (.Y(_1493_),
    .B1(net1000),
    .B2(\vga_tetris.boardMem.board_18[15] ),
    .A2(net1020),
    .A1(\vga_tetris.boardMem.board_1[15] ));
 sg13g2_a22oi_1 _4445_ (.Y(_1494_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_19[15] ),
    .A2(net1006),
    .A1(\vga_tetris.boardMem.board_8[15] ));
 sg13g2_a22oi_1 _4446_ (.Y(_1495_),
    .B1(net1007),
    .B2(\vga_tetris.boardMem.board_9[15] ),
    .A2(net1017),
    .A1(\vga_tetris.boardMem.board_5[15] ));
 sg13g2_nand4_1 _4447_ (.B(_1493_),
    .C(_1494_),
    .A(_1485_),
    .Y(_1496_),
    .D(_1495_));
 sg13g2_or4_1 _4448_ (.A(net845),
    .B(_1491_),
    .C(_1492_),
    .D(_1496_),
    .X(_1497_));
 sg13g2_a21oi_1 _4449_ (.A1(_0688_),
    .A2(net847),
    .Y(_1498_),
    .B1(net1084));
 sg13g2_nand2_2 _4450_ (.Y(_1499_),
    .A(_1497_),
    .B(_1498_));
 sg13g2_nor2_1 _4451_ (.A(_0969_),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_nand3_1 _4452_ (.B(net1062),
    .C(net1051),
    .A(\vga_tetris.boardMem.board_1[11] ),
    .Y(_1501_));
 sg13g2_nand3_1 _4453_ (.B(net1059),
    .C(_0853_),
    .A(\vga_tetris.boardMem.board_18[11] ),
    .Y(_1502_));
 sg13g2_nand3_1 _4454_ (.B(net1073),
    .C(net1066),
    .A(\vga_tetris.boardMem.board_15[11] ),
    .Y(_1503_));
 sg13g2_nand3_1 _4455_ (.B(net1062),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_2[11] ),
    .Y(_1504_));
 sg13g2_nand3_1 _4456_ (.B(net1032),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_10[11] ),
    .Y(_1505_));
 sg13g2_nand3_1 _4457_ (.B(net1051),
    .C(net1044),
    .A(\vga_tetris.boardMem.board_5[11] ),
    .Y(_1506_));
 sg13g2_nand3_1 _4458_ (.B(net1074),
    .C(net1042),
    .A(\vga_tetris.boardMem.board_12[11] ),
    .Y(_1507_));
 sg13g2_nand3_1 _4459_ (.B(net1057),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_16[11] ),
    .Y(_1508_));
 sg13g2_nand3_1 _4460_ (.B(net1044),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_4[11] ),
    .Y(_1509_));
 sg13g2_nand3_1 _4461_ (.B(net1044),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_6[11] ),
    .Y(_1510_));
 sg13g2_nand3_1 _4462_ (.B(_0836_),
    .C(net1057),
    .A(\vga_tetris.boardMem.board_19[11] ),
    .Y(_1511_));
 sg13g2_nand3_1 _4463_ (.B(_0839_),
    .C(net1059),
    .A(\vga_tetris.boardMem.board_17[11] ),
    .Y(_1512_));
 sg13g2_nand3_1 _4464_ (.B(net1066),
    .C(net1062),
    .A(\vga_tetris.boardMem.board_3[11] ),
    .Y(_1513_));
 sg13g2_nand3_1 _4465_ (.B(net1051),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_9[11] ),
    .Y(_1514_));
 sg13g2_nand3_1 _4466_ (.B(net1073),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_14[11] ),
    .Y(_1515_));
 sg13g2_nand3_1 _4467_ (.B(net1073),
    .C(net1051),
    .A(\vga_tetris.boardMem.board_13[11] ),
    .Y(_1516_));
 sg13g2_nand3_1 _4468_ (.B(net1040),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_8[11] ),
    .Y(_1517_));
 sg13g2_nand3_1 _4469_ (.B(net1066),
    .C(net1044),
    .A(\vga_tetris.boardMem.board_7[11] ),
    .Y(_1518_));
 sg13g2_nand3_1 _4470_ (.B(net1066),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_11[11] ),
    .Y(_1519_));
 sg13g2_nand4_1 _4471_ (.B(_1506_),
    .C(_1507_),
    .A(_1502_),
    .Y(_1520_),
    .D(_1512_));
 sg13g2_a21oi_1 _4472_ (.A1(net986),
    .A2(net985),
    .Y(_1521_),
    .B1(_1520_));
 sg13g2_nand4_1 _4473_ (.B(_1505_),
    .C(_1511_),
    .A(_1501_),
    .Y(_1522_),
    .D(_1518_));
 sg13g2_nand4_1 _4474_ (.B(_1510_),
    .C(_1513_),
    .A(_1509_),
    .Y(_1523_),
    .D(_1514_));
 sg13g2_nand3_1 _4475_ (.B(_1508_),
    .C(_1517_),
    .A(_1504_),
    .Y(_1524_));
 sg13g2_nand4_1 _4476_ (.B(_1515_),
    .C(_1516_),
    .A(_1503_),
    .Y(_1525_),
    .D(_1519_));
 sg13g2_nor4_2 _4477_ (.A(_1522_),
    .B(_1523_),
    .C(_1524_),
    .Y(_1526_),
    .D(_1525_));
 sg13g2_a221oi_1 _4478_ (.B2(_1526_),
    .C1(net1083),
    .B1(_1521_),
    .A1(_0684_),
    .Y(_1527_),
    .A2(net843));
 sg13g2_nand2_1 _4479_ (.Y(_1528_),
    .A(_1032_),
    .B(_1527_));
 sg13g2_a221oi_1 _4480_ (.B2(_1079_),
    .C1(_1407_),
    .B1(_1449_),
    .A1(_0987_),
    .Y(_1529_),
    .A2(_1424_));
 sg13g2_nand4_1 _4481_ (.B(_1467_),
    .C(_1528_),
    .A(_1390_),
    .Y(_1530_),
    .D(_1529_));
 sg13g2_nor4_2 _4482_ (.A(_1362_),
    .B(_1483_),
    .C(_1500_),
    .Y(_1531_),
    .D(_1530_));
 sg13g2_a21o_2 _4483_ (.A2(_1531_),
    .A1(_1138_),
    .B1(_1319_),
    .X(uo_out[0]));
 sg13g2_nor4_2 _4484_ (.A(_1137_),
    .B(_1160_),
    .C(_1230_),
    .Y(uo_out[6]),
    .D(_1531_));
 sg13g2_a21o_2 _4485_ (.A2(uo_out[6]),
    .A1(_1130_),
    .B1(_1318_),
    .X(uo_out[1]));
 sg13g2_nand3_1 _4486_ (.B(_1231_),
    .C(_1531_),
    .A(_1138_),
    .Y(_1532_));
 sg13g2_nand2b_2 _4487_ (.Y(uo_out[5]),
    .B(_1532_),
    .A_N(uo_out[1]));
 sg13g2_nor2b_2 _4488_ (.A(_1130_),
    .B_N(uo_out[6]),
    .Y(uo_out[2]));
 sg13g2_nand3_1 _4489_ (.B(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .C(net1669),
    .A(net1682),
    .Y(_1533_));
 sg13g2_nor3_1 _4490_ (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .C(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .Y(_1534_));
 sg13g2_nor3_1 _4491_ (.A(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .B(_1133_),
    .C(_1534_),
    .Y(_1535_));
 sg13g2_nand2_1 _4492_ (.Y(vga_hs),
    .A(_1533_),
    .B(_1535_));
 sg13g2_nand3b_1 _4493_ (.B(net1622),
    .C(net1599),
    .Y(_1536_),
    .A_N(\vga_tetris.vgaController.verticalCounterQ[2] ));
 sg13g2_or4_1 _4494_ (.A(net1853),
    .B(net1667),
    .C(_1131_),
    .D(_1536_),
    .X(\vga_tetris._vgaController_io_vSync ));
 sg13g2_nor3_2 _4495_ (.A(net1233),
    .B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .C(net1789),
    .Y(_1537_));
 sg13g2_nand2_1 _4496_ (.Y(_1538_),
    .A(_0741_),
    .B(_1537_));
 sg13g2_o21ai_1 _4497_ (.B1(_1538_),
    .Y(_1539_),
    .A1(_0729_),
    .A2(_0737_));
 sg13g2_nor2b_1 _4498_ (.A(_0813_),
    .B_N(net1169),
    .Y(_1540_));
 sg13g2_nand4_1 _4499_ (.B(_0782_),
    .C(_0827_),
    .A(_0775_),
    .Y(_1541_),
    .D(_1540_));
 sg13g2_inv_1 _4500_ (.Y(_1542_),
    .A(_1541_));
 sg13g2_or2_1 _4501_ (.X(_1543_),
    .B(_0749_),
    .A(_0737_));
 sg13g2_nand2_1 _4502_ (.Y(_1544_),
    .A(_1541_),
    .B(_1543_));
 sg13g2_nor3_2 _4503_ (.A(_0699_),
    .B(_0740_),
    .C(_0749_),
    .Y(_1545_));
 sg13g2_nor2_2 _4504_ (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1546_));
 sg13g2_nand2b_2 _4505_ (.Y(_1547_),
    .B(_1546_),
    .A_N(net1237));
 sg13g2_nor2_2 _4506_ (.A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .B(_1547_),
    .Y(_1548_));
 sg13g2_nand2b_1 _4507_ (.Y(_1549_),
    .B(_0763_),
    .A_N(_0759_));
 sg13g2_inv_1 _4508_ (.Y(_1550_),
    .A(_1549_));
 sg13g2_nor4_1 _4509_ (.A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .B(net1235),
    .C(_1547_),
    .D(_1549_),
    .Y(_1551_));
 sg13g2_nor2_1 _4510_ (.A(_1031_),
    .B(_1527_),
    .Y(_1552_));
 sg13g2_inv_2 _4511_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_nor4_2 _4512_ (.A(net1239),
    .B(net1240),
    .C(_0701_),
    .Y(_1554_),
    .D(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ));
 sg13g2_nand2_2 _4513_ (.Y(_1555_),
    .A(_1095_),
    .B(_1482_));
 sg13g2_nand2_2 _4514_ (.Y(_1556_),
    .A(_0700_),
    .B(net1240));
 sg13g2_nand2_2 _4515_ (.Y(_1557_),
    .A(_0701_),
    .B(net1232));
 sg13g2_nor2_2 _4516_ (.A(_1556_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_nor2_2 _4517_ (.A(net1231),
    .B(net1232),
    .Y(_1559_));
 sg13g2_nor2b_2 _4518_ (.A(_1556_),
    .B_N(_1559_),
    .Y(_1560_));
 sg13g2_a22oi_1 _4519_ (.Y(_1561_),
    .B1(_1497_),
    .B2(_1498_),
    .A2(_0984_),
    .A1(_0983_));
 sg13g2_nand2_2 _4520_ (.Y(_1562_),
    .A(_0985_),
    .B(_1499_));
 sg13g2_nor2_2 _4521_ (.A(_0966_),
    .B(_1389_),
    .Y(_1563_));
 sg13g2_nand2_1 _4522_ (.Y(_1564_),
    .A(net1231),
    .B(net1232));
 sg13g2_a21oi_1 _4523_ (.A1(net1231),
    .A2(net1232),
    .Y(_1565_),
    .B1(net1240));
 sg13g2_inv_1 _4524_ (.Y(_1566_),
    .A(_1565_));
 sg13g2_nor2_1 _4525_ (.A(net1240),
    .B(net1231),
    .Y(_1567_));
 sg13g2_nor3_1 _4526_ (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .B(net1231),
    .C(net1232),
    .Y(_1568_));
 sg13g2_nand2b_2 _4527_ (.Y(_1569_),
    .B(_1559_),
    .A_N(net1240));
 sg13g2_nor2_2 _4528_ (.A(net1239),
    .B(_1569_),
    .Y(_1570_));
 sg13g2_nand2_1 _4529_ (.Y(_1571_),
    .A(_0700_),
    .B(_1568_));
 sg13g2_o21ai_1 _4530_ (.B1(_1571_),
    .Y(_1572_),
    .A1(_0700_),
    .A2(_1565_));
 sg13g2_nor2b_1 _4531_ (.A(_1563_),
    .B_N(_1572_),
    .Y(_1573_));
 sg13g2_a22oi_1 _4532_ (.Y(_1574_),
    .B1(_1404_),
    .B2(_1405_),
    .A2(_0915_),
    .A1(_0888_));
 sg13g2_nand2b_2 _4533_ (.Y(_1575_),
    .B(_1406_),
    .A_N(_0916_));
 sg13g2_nor3_2 _4534_ (.A(net1239),
    .B(net1240),
    .C(_1564_),
    .Y(_1576_));
 sg13g2_nor3_2 _4535_ (.A(net1239),
    .B(net1240),
    .C(_1557_),
    .Y(_1577_));
 sg13g2_a22oi_1 _4536_ (.Y(_1578_),
    .B1(_1463_),
    .B2(_1464_),
    .A2(_1047_),
    .A1(_1046_));
 sg13g2_nand2_2 _4537_ (.Y(_1579_),
    .A(_1048_),
    .B(_1466_));
 sg13g2_a22oi_1 _4538_ (.Y(_1580_),
    .B1(_1575_),
    .B2(_1576_),
    .A2(_1562_),
    .A1(_1560_));
 sg13g2_a21oi_1 _4539_ (.A1(_1553_),
    .A2(_1554_),
    .Y(_1581_),
    .B1(_1573_));
 sg13g2_a22oi_1 _4540_ (.Y(_1582_),
    .B1(_1577_),
    .B2(_1579_),
    .A2(_1558_),
    .A1(_1555_));
 sg13g2_nand3_1 _4541_ (.B(_1581_),
    .C(_1582_),
    .A(_1580_),
    .Y(_1583_));
 sg13g2_nor2_1 _4542_ (.A(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .B(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .Y(_1584_));
 sg13g2_nand2_1 _4543_ (.Y(_1585_),
    .A(_0662_),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ));
 sg13g2_nor2_2 _4544_ (.A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_nor2_1 _4545_ (.A(net1237),
    .B(_1546_),
    .Y(_1587_));
 sg13g2_a21oi_1 _4546_ (.A1(net1237),
    .A2(_1586_),
    .Y(_1588_),
    .B1(_1587_));
 sg13g2_nor3_1 _4547_ (.A(net1235),
    .B(_1549_),
    .C(_1588_),
    .Y(_1589_));
 sg13g2_nor2b_1 _4548_ (.A(_0763_),
    .B_N(_0759_),
    .Y(_1590_));
 sg13g2_inv_1 _4549_ (.Y(_1591_),
    .A(_1590_));
 sg13g2_and3_2 _4550_ (.X(_1592_),
    .A(_0660_),
    .B(net1237),
    .C(_1546_));
 sg13g2_nor2_1 _4551_ (.A(net1843),
    .B(net1236),
    .Y(_1593_));
 sg13g2_nor3_2 _4552_ (.A(net1237),
    .B(_0662_),
    .C(_0663_),
    .Y(_1594_));
 sg13g2_nor2_2 _4553_ (.A(_0660_),
    .B(net1236),
    .Y(_1595_));
 sg13g2_a22oi_1 _4554_ (.Y(_1596_),
    .B1(_1594_),
    .B2(_1595_),
    .A2(_1592_),
    .A1(_0661_));
 sg13g2_nor2_1 _4555_ (.A(_0759_),
    .B(_0763_),
    .Y(_1597_));
 sg13g2_nor3_2 _4556_ (.A(net1238),
    .B(_0662_),
    .C(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1598_));
 sg13g2_nand3_1 _4557_ (.B(_1597_),
    .C(_1598_),
    .A(_1595_),
    .Y(_1599_));
 sg13g2_o21ai_1 _4558_ (.B1(_1599_),
    .Y(_1600_),
    .A1(_1591_),
    .A2(_1596_));
 sg13g2_or3_1 _4559_ (.A(net1091),
    .B(_1589_),
    .C(_1600_),
    .X(_1601_));
 sg13g2_nor2_1 _4560_ (.A(_0700_),
    .B(_1566_),
    .Y(_1602_));
 sg13g2_o21ai_1 _4561_ (.B1(_1602_),
    .Y(_1603_),
    .A1(net1231),
    .A2(net1087));
 sg13g2_nor2b_1 _4562_ (.A(_1584_),
    .B_N(_1603_),
    .Y(_1604_));
 sg13g2_and2_1 _4563_ (.A(net1237),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .X(_1605_));
 sg13g2_nand2_2 _4564_ (.Y(_1606_),
    .A(net1238),
    .B(net1745));
 sg13g2_a21oi_1 _4565_ (.A1(_0663_),
    .A2(_1593_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_and2_1 _4566_ (.A(net1235),
    .B(_1598_),
    .X(_1608_));
 sg13g2_nand2_1 _4567_ (.Y(_1609_),
    .A(_0660_),
    .B(net1235));
 sg13g2_nor2_1 _4568_ (.A(_0660_),
    .B(_0661_),
    .Y(_1610_));
 sg13g2_nand2_1 _4569_ (.Y(_1611_),
    .A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .B(net1235));
 sg13g2_nor2_1 _4570_ (.A(net1238),
    .B(_1585_),
    .Y(_1612_));
 sg13g2_a22oi_1 _4571_ (.Y(_1613_),
    .B1(_1610_),
    .B2(_1612_),
    .A2(_1548_),
    .A1(net1236));
 sg13g2_nand3_1 _4572_ (.B(net1238),
    .C(_1586_),
    .A(net1235),
    .Y(_1614_));
 sg13g2_a21oi_1 _4573_ (.A1(_0660_),
    .A2(_1594_),
    .Y(_1615_),
    .B1(_1608_));
 sg13g2_nand3_1 _4574_ (.B(_1614_),
    .C(_1615_),
    .A(_1613_),
    .Y(_1616_));
 sg13g2_o21ai_1 _4575_ (.B1(_1597_),
    .Y(_1617_),
    .A1(_1605_),
    .A2(_1616_));
 sg13g2_o21ai_1 _4576_ (.B1(_1611_),
    .Y(_1618_),
    .A1(_1548_),
    .A2(_1594_));
 sg13g2_nor3_1 _4577_ (.A(_1592_),
    .B(_1605_),
    .C(_1612_),
    .Y(_1619_));
 sg13g2_nand2_1 _4578_ (.Y(_1620_),
    .A(_1598_),
    .B(_1609_));
 sg13g2_nand4_1 _4579_ (.B(_1618_),
    .C(_1619_),
    .A(_1614_),
    .Y(_1621_),
    .D(_1620_));
 sg13g2_nand2_1 _4580_ (.Y(_1622_),
    .A(_1550_),
    .B(_1621_));
 sg13g2_a21oi_1 _4581_ (.A1(_1617_),
    .A2(_1622_),
    .Y(_1623_),
    .B1(_1607_));
 sg13g2_nand2b_2 _4582_ (.Y(_1624_),
    .B(_1609_),
    .A_N(_1595_));
 sg13g2_a21oi_1 _4583_ (.A1(net1237),
    .A2(_1586_),
    .Y(_1625_),
    .B1(_1598_));
 sg13g2_or2_1 _4584_ (.X(_1626_),
    .B(_1625_),
    .A(_1624_));
 sg13g2_o21ai_1 _4585_ (.B1(net1235),
    .Y(_1627_),
    .A1(_1592_),
    .A2(_1594_));
 sg13g2_nand3_1 _4586_ (.B(_1626_),
    .C(_1627_),
    .A(_1613_),
    .Y(_1628_));
 sg13g2_a22oi_1 _4587_ (.Y(_1629_),
    .B1(_1590_),
    .B2(_1628_),
    .A2(_1548_),
    .A1(net1235));
 sg13g2_nand2b_2 _4588_ (.Y(_1630_),
    .B(_1629_),
    .A_N(_1623_));
 sg13g2_or2_1 _4589_ (.X(_1631_),
    .B(_1608_),
    .A(_1586_));
 sg13g2_a221oi_1 _4590_ (.B2(_1610_),
    .C1(_1631_),
    .B1(_1594_),
    .A1(_0661_),
    .Y(_1632_),
    .A2(_1592_));
 sg13g2_nand2b_1 _4591_ (.Y(_1633_),
    .B(_1590_),
    .A_N(_1632_));
 sg13g2_o21ai_1 _4592_ (.B1(_1624_),
    .Y(_1634_),
    .A1(_1608_),
    .A2(_1612_));
 sg13g2_nand3_1 _4593_ (.B(_1627_),
    .C(_1634_),
    .A(_1606_),
    .Y(_1635_));
 sg13g2_o21ai_1 _4594_ (.B1(_1609_),
    .Y(_1636_),
    .A1(_1548_),
    .A2(_1594_));
 sg13g2_o21ai_1 _4595_ (.B1(_1611_),
    .Y(_1637_),
    .A1(_1586_),
    .A2(_1598_));
 sg13g2_nand3_1 _4596_ (.B(_1636_),
    .C(_1637_),
    .A(_1619_),
    .Y(_1638_));
 sg13g2_a22oi_1 _4597_ (.Y(_1639_),
    .B1(_1638_),
    .B2(_1550_),
    .A2(_1635_),
    .A1(_1597_));
 sg13g2_o21ai_1 _4598_ (.B1(_1633_),
    .Y(_1640_),
    .A1(_1607_),
    .A2(_1639_));
 sg13g2_nor3_1 _4599_ (.A(net1087),
    .B(net1081),
    .C(net1086),
    .Y(_1641_));
 sg13g2_a21oi_1 _4600_ (.A1(_0784_),
    .A2(_1604_),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_nand3_1 _4601_ (.B(net1231),
    .C(net1232),
    .A(net1240),
    .Y(_1643_));
 sg13g2_nor2_2 _4602_ (.A(net1239),
    .B(_1643_),
    .Y(_1644_));
 sg13g2_a221oi_1 _4603_ (.B2(net1091),
    .C1(_1584_),
    .B1(_1644_),
    .A1(net1239),
    .Y(_1645_),
    .A2(_1566_));
 sg13g2_nand2b_1 _4604_ (.Y(_1646_),
    .B(_1645_),
    .A_N(_1642_));
 sg13g2_nor2_1 _4605_ (.A(_1123_),
    .B(_1360_),
    .Y(_1647_));
 sg13g2_inv_1 _4606_ (.Y(_1648_),
    .A(_1647_));
 sg13g2_nor2b_1 _4607_ (.A(_1563_),
    .B_N(_1577_),
    .Y(_1649_));
 sg13g2_a21oi_1 _4608_ (.A1(_1572_),
    .A2(_1648_),
    .Y(_1650_),
    .B1(_1649_));
 sg13g2_a22oi_1 _4609_ (.Y(_1651_),
    .B1(_1579_),
    .B2(_1554_),
    .A2(_1562_),
    .A1(_1558_));
 sg13g2_nor3_2 _4610_ (.A(_0701_),
    .B(net1232),
    .C(_1556_),
    .Y(_1652_));
 sg13g2_a22oi_1 _4611_ (.Y(_1653_),
    .B1(_1652_),
    .B2(_1555_),
    .A2(_1575_),
    .A1(_1560_));
 sg13g2_nor2_2 _4612_ (.A(_1076_),
    .B(_1449_),
    .Y(_1654_));
 sg13g2_a21oi_1 _4613_ (.A1(net1090),
    .A2(_1652_),
    .Y(_1655_),
    .B1(_1644_));
 sg13g2_nor2_1 _4614_ (.A(_1654_),
    .B(_1655_),
    .Y(_1656_));
 sg13g2_a21oi_1 _4615_ (.A1(_1553_),
    .A2(_1576_),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_nand4_1 _4616_ (.B(_1651_),
    .C(_1653_),
    .A(_1650_),
    .Y(_1658_),
    .D(_1657_));
 sg13g2_a22oi_1 _4617_ (.Y(_1659_),
    .B1(_1652_),
    .B2(net1090),
    .A2(_1644_),
    .A1(net1087));
 sg13g2_a221oi_1 _4618_ (.B2(_1658_),
    .C1(_1646_),
    .B1(_1601_),
    .A1(net1090),
    .Y(_1660_),
    .A2(_1583_));
 sg13g2_nor2_2 _4619_ (.A(_0700_),
    .B(_1569_),
    .Y(_1661_));
 sg13g2_nor2b_1 _4620_ (.A(_1654_),
    .B_N(_1661_),
    .Y(_1662_));
 sg13g2_a22oi_1 _4621_ (.Y(_1663_),
    .B1(_1333_),
    .B2(_1334_),
    .A2(_0937_),
    .A1(_0936_));
 sg13g2_nand2_1 _4622_ (.Y(_1664_),
    .A(_0938_),
    .B(_1335_));
 sg13g2_a21oi_1 _4623_ (.A1(_1572_),
    .A2(_1664_),
    .Y(_1665_),
    .B1(_1662_));
 sg13g2_a22oi_1 _4624_ (.Y(_1666_),
    .B1(_1652_),
    .B2(_1562_),
    .A2(_1644_),
    .A1(_1555_));
 sg13g2_nand2_1 _4625_ (.Y(_1667_),
    .A(_1665_),
    .B(_1666_));
 sg13g2_nand3_1 _4626_ (.B(net1232),
    .C(_1567_),
    .A(net1239),
    .Y(_1668_));
 sg13g2_nand2_1 _4627_ (.Y(_1669_),
    .A(_1577_),
    .B(_1648_));
 sg13g2_a22oi_1 _4628_ (.Y(_1670_),
    .B1(_1576_),
    .B2(_1579_),
    .A2(_1560_),
    .A1(_1553_));
 sg13g2_nor2b_1 _4629_ (.A(_1563_),
    .B_N(_1554_),
    .Y(_1671_));
 sg13g2_a21oi_1 _4630_ (.A1(_1558_),
    .A2(_1575_),
    .Y(_1672_),
    .B1(_1671_));
 sg13g2_nand4_1 _4631_ (.B(_1669_),
    .C(_1670_),
    .A(_1668_),
    .Y(_1673_),
    .D(_1672_));
 sg13g2_o21ai_1 _4632_ (.B1(net1086),
    .Y(_1674_),
    .A1(_1667_),
    .A2(_1673_));
 sg13g2_a22oi_1 _4633_ (.Y(_1675_),
    .B1(_1421_),
    .B2(_1422_),
    .A2(_1002_),
    .A1(_1001_));
 sg13g2_nand2_1 _4634_ (.Y(_1676_),
    .A(_1003_),
    .B(_1423_));
 sg13g2_nor2_1 _4635_ (.A(_1654_),
    .B(_1668_),
    .Y(_1677_));
 sg13g2_nor2b_1 _4636_ (.A(_1563_),
    .B_N(_1576_),
    .Y(_1678_));
 sg13g2_a22oi_1 _4637_ (.Y(_1679_),
    .B1(_1661_),
    .B2(_1555_),
    .A2(_1648_),
    .A1(_1554_));
 sg13g2_a22oi_1 _4638_ (.Y(_1680_),
    .B1(_1652_),
    .B2(_1575_),
    .A2(_1644_),
    .A1(_1562_));
 sg13g2_nand2_1 _4639_ (.Y(_1681_),
    .A(_1679_),
    .B(_1680_));
 sg13g2_a21oi_1 _4640_ (.A1(_1572_),
    .A2(_1676_),
    .Y(_1682_),
    .B1(_1678_));
 sg13g2_a21oi_1 _4641_ (.A1(_1560_),
    .A2(_1579_),
    .Y(_1683_),
    .B1(_1677_));
 sg13g2_a22oi_1 _4642_ (.Y(_1684_),
    .B1(_1577_),
    .B2(_1664_),
    .A2(_1558_),
    .A1(_1553_));
 sg13g2_nand3_1 _4643_ (.B(_1683_),
    .C(_1684_),
    .A(_1682_),
    .Y(_1685_));
 sg13g2_o21ai_1 _4644_ (.B1(net1081),
    .Y(_1686_),
    .A1(_1681_),
    .A2(_1685_));
 sg13g2_nand3_1 _4645_ (.B(_1674_),
    .C(_1686_),
    .A(_1660_),
    .Y(_1687_));
 sg13g2_inv_2 _4646_ (.Y(_1688_),
    .A(_1687_));
 sg13g2_nand4_1 _4647_ (.B(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .C(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .Y(_1689_),
    .D(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ));
 sg13g2_o21ai_1 _4648_ (.B1(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .Y(_1690_),
    .A1(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ));
 sg13g2_nor3_1 _4649_ (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .B(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .C(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .Y(_1691_));
 sg13g2_a22oi_1 _4650_ (.Y(_1692_),
    .B1(_1690_),
    .B2(_1691_),
    .A2(_1689_),
    .A1(_0702_));
 sg13g2_nand2_1 _4651_ (.Y(_1693_),
    .A(_0742_),
    .B(_1692_));
 sg13g2_a21oi_1 _4652_ (.A1(_0742_),
    .A2(_1692_),
    .Y(_1694_),
    .B1(_1545_));
 sg13g2_and2_1 _4653_ (.A(_0741_),
    .B(_0745_),
    .X(_1695_));
 sg13g2_nand2_2 _4654_ (.Y(_1696_),
    .A(_0741_),
    .B(_0745_));
 sg13g2_nand2_1 _4655_ (.Y(_1697_),
    .A(net1226),
    .B(_1537_));
 sg13g2_and2_1 _4656_ (.A(net1241),
    .B(_1537_),
    .X(_1698_));
 sg13g2_nand2_2 _4657_ (.Y(_1699_),
    .A(net1226),
    .B(net1187));
 sg13g2_inv_1 _4658_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_o21ai_1 _4659_ (.B1(_1696_),
    .Y(_1701_),
    .A1(net1227),
    .A2(_1699_));
 sg13g2_nand2_2 _4660_ (.Y(_1702_),
    .A(\vga_tetris._inputs_io_leftButtonActive ),
    .B(_1571_));
 sg13g2_inv_1 _4661_ (.Y(_1703_),
    .A(_1702_));
 sg13g2_nand3_1 _4662_ (.B(_1668_),
    .C(_1702_),
    .A(\vga_tetris._inputs_io_rightButtonActive ),
    .Y(_1704_));
 sg13g2_nor2_2 _4663_ (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .B(_1696_),
    .Y(_1705_));
 sg13g2_nand2_1 _4664_ (.Y(_1706_),
    .A(_1704_),
    .B(_1705_));
 sg13g2_nand2_1 _4665_ (.Y(_1707_),
    .A(_1701_),
    .B(_1706_));
 sg13g2_a22oi_1 _4666_ (.Y(_1708_),
    .B1(_1694_),
    .B2(_1707_),
    .A2(_1688_),
    .A1(_1545_));
 sg13g2_nor2_2 _4667_ (.A(_0728_),
    .B(_0749_),
    .Y(_1709_));
 sg13g2_or2_1 _4668_ (.X(_1710_),
    .B(_0749_),
    .A(_0728_));
 sg13g2_nand2_2 _4669_ (.Y(_1711_),
    .A(net1799),
    .B(_0754_));
 sg13g2_nor2_2 _4670_ (.A(\vga_tetris.tetrisLogic.stateQ[0] ),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_nor3_1 _4671_ (.A(_1708_),
    .B(_1709_),
    .C(_1712_),
    .Y(_1713_));
 sg13g2_a22oi_1 _4672_ (.Y(_1714_),
    .B1(_1713_),
    .B2(_1541_),
    .A2(_1544_),
    .A1(_1538_));
 sg13g2_or2_1 _4673_ (.X(_1715_),
    .B(_0738_),
    .A(_0699_));
 sg13g2_nand4_1 _4674_ (.B(_1699_),
    .C(_1711_),
    .A(_1696_),
    .Y(_1716_),
    .D(_1715_));
 sg13g2_nand4_1 _4675_ (.B(_0668_),
    .C(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .A(net1241),
    .Y(_1717_),
    .D(_0739_));
 sg13g2_inv_1 _4676_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_nand2_1 _4677_ (.Y(_1719_),
    .A(_1710_),
    .B(_1717_));
 sg13g2_nor2_1 _4678_ (.A(_0742_),
    .B(_1545_),
    .Y(_1720_));
 sg13g2_nor4_1 _4679_ (.A(_0742_),
    .B(_1545_),
    .C(_1716_),
    .D(_1719_),
    .Y(_1721_));
 sg13g2_nand2b_1 _4680_ (.Y(_1722_),
    .B(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .A_N(_0747_));
 sg13g2_nand2_2 _4681_ (.Y(_1723_),
    .A(net1878),
    .B(_0718_));
 sg13g2_nor2_1 _4682_ (.A(net1181),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_or2_1 _4683_ (.X(_1725_),
    .B(_0748_),
    .A(_0699_));
 sg13g2_nand3_1 _4684_ (.B(_0735_),
    .C(_1537_),
    .A(net1226),
    .Y(_1726_));
 sg13g2_and2_1 _4685_ (.A(_1725_),
    .B(_1726_),
    .X(_1727_));
 sg13g2_a21oi_1 _4686_ (.A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .A2(_0752_),
    .Y(_1728_),
    .B1(_1724_));
 sg13g2_and4_1 _4687_ (.A(_1721_),
    .B(_1722_),
    .C(_1727_),
    .D(_1728_),
    .X(_1729_));
 sg13g2_nand2_2 _4688_ (.Y(_1730_),
    .A(_1541_),
    .B(_1729_));
 sg13g2_o21ai_1 _4689_ (.B1(net1265),
    .Y(_1731_),
    .A1(net1880),
    .A2(_1730_));
 sg13g2_nand2_1 _4690_ (.Y(_1732_),
    .A(net1234),
    .B(_0743_));
 sg13g2_o21ai_1 _4691_ (.B1(_1543_),
    .Y(_1733_),
    .A1(net1241),
    .A2(_1732_));
 sg13g2_nor2_1 _4692_ (.A(_1714_),
    .B(_1731_),
    .Y(_0000_));
 sg13g2_or2_1 _4693_ (.X(_1734_),
    .B(_1715_),
    .A(_1687_));
 sg13g2_nand2_1 _4694_ (.Y(_1735_),
    .A(_1702_),
    .B(_1705_));
 sg13g2_nand2b_1 _4695_ (.Y(_1736_),
    .B(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .A_N(net1227));
 sg13g2_o21ai_1 _4696_ (.B1(_1696_),
    .Y(_1737_),
    .A1(_1699_),
    .A2(_1736_));
 sg13g2_nand2_1 _4697_ (.Y(_1738_),
    .A(_1735_),
    .B(_1737_));
 sg13g2_nor3_1 _4698_ (.A(_1712_),
    .B(_1718_),
    .C(_1724_),
    .Y(_1739_));
 sg13g2_nand4_1 _4699_ (.B(_1715_),
    .C(_1738_),
    .A(_1693_),
    .Y(_1740_),
    .D(_1739_));
 sg13g2_nand2_1 _4700_ (.Y(_1741_),
    .A(_1734_),
    .B(_1740_));
 sg13g2_nor2_1 _4701_ (.A(_1687_),
    .B(_1725_),
    .Y(_1742_));
 sg13g2_or2_1 _4702_ (.X(_1743_),
    .B(_1742_),
    .A(_1729_));
 sg13g2_a21oi_1 _4703_ (.A1(_1725_),
    .A2(_1741_),
    .Y(_1744_),
    .B1(_1743_));
 sg13g2_nor2_1 _4704_ (.A(_0667_),
    .B(_1730_),
    .Y(_1745_));
 sg13g2_nor3_1 _4705_ (.A(net1162),
    .B(_1744_),
    .C(_1745_),
    .Y(_1746_));
 sg13g2_nor2_1 _4706_ (.A(net1251),
    .B(_1746_),
    .Y(_0001_));
 sg13g2_nand2_1 _4707_ (.Y(_1747_),
    .A(net1265),
    .B(_1543_));
 sg13g2_or2_1 _4708_ (.X(_1748_),
    .B(net1162),
    .A(net1252));
 sg13g2_nand4_1 _4709_ (.B(_1722_),
    .C(_1735_),
    .A(_1720_),
    .Y(_1749_),
    .D(_1739_));
 sg13g2_a21oi_1 _4710_ (.A1(net1789),
    .A2(_1721_),
    .Y(_1750_),
    .B1(_1749_));
 sg13g2_nor2_1 _4711_ (.A(_1748_),
    .B(net1790),
    .Y(_0002_));
 sg13g2_a21o_1 _4712_ (.A2(_1725_),
    .A1(_1715_),
    .B1(_1688_),
    .X(_1751_));
 sg13g2_nand2_1 _4713_ (.Y(_1752_),
    .A(net1269),
    .B(_1710_));
 sg13g2_nand2_2 _4714_ (.Y(_1753_),
    .A(net1265),
    .B(_1751_));
 sg13g2_nor2_1 _4715_ (.A(_1709_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_nor2_1 _4716_ (.A(_0699_),
    .B(_1688_),
    .Y(_1755_));
 sg13g2_nand4_1 _4717_ (.B(\vga_tetris.tetrisLogic.stateQ[0] ),
    .C(_0745_),
    .A(net1242),
    .Y(_1756_),
    .D(_1755_));
 sg13g2_nand2_1 _4718_ (.Y(_1757_),
    .A(_1566_),
    .B(_1643_));
 sg13g2_nand3_1 _4719_ (.B(_0739_),
    .C(_1755_),
    .A(_0735_),
    .Y(_1758_));
 sg13g2_xnor2_1 _4720_ (.Y(_1759_),
    .A(net1910),
    .B(_1559_));
 sg13g2_or2_1 _4721_ (.X(_1760_),
    .B(_1759_),
    .A(_1702_));
 sg13g2_o21ai_1 _4722_ (.B1(_1760_),
    .Y(_1761_),
    .A1(_1704_),
    .A2(_1757_));
 sg13g2_nor4_2 _4723_ (.A(net1227),
    .B(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .C(_0729_),
    .Y(_1762_),
    .D(_1697_));
 sg13g2_a21o_1 _4724_ (.A2(_1668_),
    .A1(\vga_tetris._inputs_io_rightButtonActive ),
    .B1(_1703_),
    .X(_1763_));
 sg13g2_nand2_1 _4725_ (.Y(_1764_),
    .A(_1695_),
    .B(_1763_));
 sg13g2_nand2_1 _4726_ (.Y(_1765_),
    .A(_1705_),
    .B(_1763_));
 sg13g2_a21oi_1 _4727_ (.A1(_1705_),
    .A2(_1763_),
    .Y(_1766_),
    .B1(_1762_));
 sg13g2_a22oi_1 _4728_ (.Y(_1767_),
    .B1(_1766_),
    .B2(net1910),
    .A2(_1761_),
    .A1(_1705_));
 sg13g2_mux2_1 _4729_ (.A0(_1757_),
    .A1(_1767_),
    .S(_1756_),
    .X(_1768_));
 sg13g2_mux2_1 _4730_ (.A0(_1759_),
    .A1(_1768_),
    .S(_1758_),
    .X(_1769_));
 sg13g2_nor2b_1 _4731_ (.A(_1769_),
    .B_N(_1754_),
    .Y(_0003_));
 sg13g2_nand3_1 _4732_ (.B(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .C(_1569_),
    .A(\vga_tetris._inputs_io_leftButtonActive ),
    .Y(_1770_));
 sg13g2_xnor2_1 _4733_ (.Y(_1771_),
    .A(_0700_),
    .B(_1643_));
 sg13g2_o21ai_1 _4734_ (.B1(_1770_),
    .Y(_1772_),
    .A1(_1704_),
    .A2(_1771_));
 sg13g2_a22oi_1 _4735_ (.Y(_1773_),
    .B1(_1772_),
    .B2(_1705_),
    .A2(_1766_),
    .A1(net1908));
 sg13g2_xnor2_1 _4736_ (.Y(_1774_),
    .A(_0700_),
    .B(_1568_));
 sg13g2_mux2_1 _4737_ (.A0(_1771_),
    .A1(_1773_),
    .S(_1756_),
    .X(_1775_));
 sg13g2_o21ai_1 _4738_ (.B1(_1754_),
    .Y(_1776_),
    .A1(_1758_),
    .A2(_1774_));
 sg13g2_a21oi_1 _4739_ (.A1(_1758_),
    .A2(_1775_),
    .Y(_0004_),
    .B1(_1776_));
 sg13g2_and3_1 _4740_ (.X(_1777_),
    .A(net646),
    .B(net1351),
    .C(net738));
 sg13g2_and2_1 _4741_ (.A(net1522),
    .B(_1777_),
    .X(_1778_));
 sg13g2_and2_1 _4742_ (.A(net1787),
    .B(_1778_),
    .X(_1779_));
 sg13g2_nor3_1 _4743_ (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .C(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .Y(_1780_));
 sg13g2_nand4_1 _4744_ (.B(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .C(_1779_),
    .A(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .Y(_1781_),
    .D(_1780_));
 sg13g2_nand2_1 _4745_ (.Y(_1782_),
    .A(net1222),
    .B(_0906_));
 sg13g2_and2_1 _4746_ (.A(_0906_),
    .B(_0967_),
    .X(_1783_));
 sg13g2_inv_1 _4747_ (.Y(_1784_),
    .A(_1783_));
 sg13g2_nand2_1 _4748_ (.Y(_1785_),
    .A(net1219),
    .B(_1783_));
 sg13g2_nand2b_1 _4749_ (.Y(_1786_),
    .B(_1785_),
    .A_N(net1218));
 sg13g2_o21ai_1 _4750_ (.B1(net1809),
    .Y(_1787_),
    .A1(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .A2(_1786_));
 sg13g2_nor2_2 _4751_ (.A(_1781_),
    .B(net1089),
    .Y(_1788_));
 sg13g2_nor2_2 _4752_ (.A(net1245),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_o21ai_1 _4753_ (.B1(net1259),
    .Y(_1790_),
    .A1(_1781_),
    .A2(net1089));
 sg13g2_nor2_1 _4754_ (.A(net646),
    .B(net1088),
    .Y(_0005_));
 sg13g2_o21ai_1 _4755_ (.B1(_1789_),
    .Y(_1791_),
    .A1(net646),
    .A2(net1351));
 sg13g2_a21oi_1 _4756_ (.A1(net646),
    .A2(net1351),
    .Y(_0006_),
    .B1(_1791_));
 sg13g2_a21oi_1 _4757_ (.A1(net646),
    .A2(\vga_tetris.vgaController.horizontalCounterQ[1] ),
    .Y(_1792_),
    .B1(net738));
 sg13g2_nor3_1 _4758_ (.A(_1777_),
    .B(net1088),
    .C(net739),
    .Y(_0007_));
 sg13g2_nor2_1 _4759_ (.A(net1522),
    .B(_1777_),
    .Y(_1793_));
 sg13g2_nor3_1 _4760_ (.A(net1245),
    .B(_1778_),
    .C(_1793_),
    .Y(_0008_));
 sg13g2_o21ai_1 _4761_ (.B1(net1259),
    .Y(_1794_),
    .A1(net1787),
    .A2(_1778_));
 sg13g2_nor2_1 _4762_ (.A(_1779_),
    .B(_1794_),
    .Y(_0009_));
 sg13g2_and2_1 _4763_ (.A(net1682),
    .B(_1779_),
    .X(_1795_));
 sg13g2_nor2_1 _4764_ (.A(net1682),
    .B(_1779_),
    .Y(_1796_));
 sg13g2_nor3_1 _4765_ (.A(net1088),
    .B(_1795_),
    .C(net1683),
    .Y(_0010_));
 sg13g2_nor2_1 _4766_ (.A(net1669),
    .B(_1795_),
    .Y(_1797_));
 sg13g2_nor2b_1 _4767_ (.A(_1533_),
    .B_N(_1778_),
    .Y(_1798_));
 sg13g2_nor3_1 _4768_ (.A(net1088),
    .B(net1670),
    .C(_1798_),
    .Y(_0011_));
 sg13g2_and2_1 _4769_ (.A(net1695),
    .B(_1798_),
    .X(_1799_));
 sg13g2_nor2_1 _4770_ (.A(net1695),
    .B(_1798_),
    .Y(_1800_));
 sg13g2_nor3_1 _4771_ (.A(net1088),
    .B(_1799_),
    .C(net1696),
    .Y(_0012_));
 sg13g2_nand2_1 _4772_ (.Y(_1801_),
    .A(net1794),
    .B(_1799_));
 sg13g2_o21ai_1 _4773_ (.B1(_1789_),
    .Y(_1802_),
    .A1(net1794),
    .A2(_1799_));
 sg13g2_nor2b_1 _4774_ (.A(net1795),
    .B_N(_1801_),
    .Y(_0013_));
 sg13g2_xor2_1 _4775_ (.B(_1801_),
    .A(net1760),
    .X(_1803_));
 sg13g2_nor2_1 _4776_ (.A(_1790_),
    .B(net1761),
    .Y(_0014_));
 sg13g2_nor4_1 _4777_ (.A(\vga_tetris.msTimer.msTimerQ[9] ),
    .B(\vga_tetris.msTimer.msTimerQ[11] ),
    .C(\vga_tetris.msTimer.msTimerQ[10] ),
    .D(net1913),
    .Y(_1804_));
 sg13g2_o21ai_1 _4778_ (.B1(\vga_tetris.msTimer.msTimerQ[5] ),
    .Y(_1805_),
    .A1(\vga_tetris.msTimer.msTimerQ[3] ),
    .A2(\vga_tetris.msTimer.msTimerQ[4] ));
 sg13g2_nor2b_1 _4779_ (.A(\vga_tetris.msTimer.msTimerQ[6] ),
    .B_N(_1805_),
    .Y(_1806_));
 sg13g2_nand2_1 _4780_ (.Y(_1807_),
    .A(net1653),
    .B(net1743));
 sg13g2_o21ai_1 _4781_ (.B1(net1914),
    .Y(_1808_),
    .A1(_1806_),
    .A2(_1807_));
 sg13g2_nand3_1 _4782_ (.B(net1385),
    .C(_1808_),
    .A(net1346),
    .Y(_1809_));
 sg13g2_nand2_2 _4783_ (.Y(_1810_),
    .A(net1270),
    .B(_1809_));
 sg13g2_inv_2 _4784_ (.Y(_1811_),
    .A(net1158));
 sg13g2_nor2_1 _4785_ (.A(net647),
    .B(net1158),
    .Y(_0015_));
 sg13g2_xnor2_1 _4786_ (.Y(_1812_),
    .A(net1744),
    .B(net647));
 sg13g2_nor2_1 _4787_ (.A(net1158),
    .B(_1812_),
    .Y(_0016_));
 sg13g2_and3_1 _4788_ (.X(_1813_),
    .A(\vga_tetris.msTimer.msTimerQ[1] ),
    .B(net647),
    .C(net1355));
 sg13g2_a21oi_1 _4789_ (.A1(\vga_tetris.msTimer.msTimerQ[1] ),
    .A2(net647),
    .Y(_1814_),
    .B1(net1355));
 sg13g2_nor3_1 _4790_ (.A(net1158),
    .B(_1813_),
    .C(net1356),
    .Y(_0017_));
 sg13g2_and2_1 _4791_ (.A(net1658),
    .B(_1813_),
    .X(_1815_));
 sg13g2_nor2_1 _4792_ (.A(net1658),
    .B(_1813_),
    .Y(_1816_));
 sg13g2_nor3_1 _4793_ (.A(net1158),
    .B(_1815_),
    .C(net1659),
    .Y(_0018_));
 sg13g2_and2_1 _4794_ (.A(net1703),
    .B(_1815_),
    .X(_1817_));
 sg13g2_nor2_1 _4795_ (.A(net1703),
    .B(_1815_),
    .Y(_1818_));
 sg13g2_nor3_1 _4796_ (.A(_1810_),
    .B(_1817_),
    .C(net1704),
    .Y(_0019_));
 sg13g2_and2_1 _4797_ (.A(net1685),
    .B(_1817_),
    .X(_1819_));
 sg13g2_nor2_1 _4798_ (.A(net1685),
    .B(_1817_),
    .Y(_1820_));
 sg13g2_nor3_1 _4799_ (.A(_1810_),
    .B(_1819_),
    .C(net1686),
    .Y(_0020_));
 sg13g2_and2_1 _4800_ (.A(net1640),
    .B(_1819_),
    .X(_1821_));
 sg13g2_nor2_1 _4801_ (.A(net1640),
    .B(_1819_),
    .Y(_1822_));
 sg13g2_nor3_1 _4802_ (.A(net1158),
    .B(_1821_),
    .C(net1641),
    .Y(_0021_));
 sg13g2_nor2_1 _4803_ (.A(net1653),
    .B(_1821_),
    .Y(_1823_));
 sg13g2_and2_1 _4804_ (.A(net1653),
    .B(_1821_),
    .X(_1824_));
 sg13g2_nor3_1 _4805_ (.A(net1158),
    .B(net1654),
    .C(_1824_),
    .Y(_0022_));
 sg13g2_nor2b_1 _4806_ (.A(_1807_),
    .B_N(_1821_),
    .Y(_1825_));
 sg13g2_o21ai_1 _4807_ (.B1(_1811_),
    .Y(_1826_),
    .A1(net1743),
    .A2(_1824_));
 sg13g2_nor2_1 _4808_ (.A(_1825_),
    .B(_1826_),
    .Y(_0023_));
 sg13g2_and2_1 _4809_ (.A(net1759),
    .B(_1825_),
    .X(_1827_));
 sg13g2_o21ai_1 _4810_ (.B1(_1811_),
    .Y(_1828_),
    .A1(net1759),
    .A2(_1825_));
 sg13g2_nor2_1 _4811_ (.A(_1827_),
    .B(_1828_),
    .Y(_0024_));
 sg13g2_and2_1 _4812_ (.A(net1770),
    .B(_1827_),
    .X(_1829_));
 sg13g2_o21ai_1 _4813_ (.B1(_1811_),
    .Y(_1830_),
    .A1(net1770),
    .A2(_1827_));
 sg13g2_nor2_1 _4814_ (.A(_1829_),
    .B(_1830_),
    .Y(_0025_));
 sg13g2_and2_1 _4815_ (.A(net1780),
    .B(_1829_),
    .X(_1831_));
 sg13g2_o21ai_1 _4816_ (.B1(_1811_),
    .Y(_1832_),
    .A1(net1780),
    .A2(_1829_));
 sg13g2_nor2_1 _4817_ (.A(_1831_),
    .B(_1832_),
    .Y(_0026_));
 sg13g2_and2_1 _4818_ (.A(net1747),
    .B(_1831_),
    .X(_1833_));
 sg13g2_o21ai_1 _4819_ (.B1(_1811_),
    .Y(_1834_),
    .A1(net1747),
    .A2(_1831_));
 sg13g2_nor2_1 _4820_ (.A(_1833_),
    .B(net1748),
    .Y(_0027_));
 sg13g2_o21ai_1 _4821_ (.B1(_1811_),
    .Y(_1835_),
    .A1(net1346),
    .A2(_1833_));
 sg13g2_a21oi_1 _4822_ (.A1(net1346),
    .A2(_1833_),
    .Y(_0028_),
    .B1(_1835_));
 sg13g2_a21oi_1 _4823_ (.A1(net1346),
    .A2(_1833_),
    .Y(_1836_),
    .B1(net1385));
 sg13g2_nor2_1 _4824_ (.A(net1158),
    .B(net1386),
    .Y(_0029_));
 sg13g2_o21ai_1 _4825_ (.B1(_1694_),
    .Y(_1837_),
    .A1(_1687_),
    .A2(_1717_));
 sg13g2_nor3_1 _4826_ (.A(net1170),
    .B(_1742_),
    .C(_1837_),
    .Y(_1838_));
 sg13g2_a21oi_2 _4827_ (.B1(_1542_),
    .Y(_1839_),
    .A2(_1838_),
    .A1(_1734_));
 sg13g2_a21oi_1 _4828_ (.A1(_0668_),
    .A2(net1187),
    .Y(_1840_),
    .B1(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ));
 sg13g2_nor3_1 _4829_ (.A(net1227),
    .B(_1699_),
    .C(_1840_),
    .Y(_1841_));
 sg13g2_nand3_1 _4830_ (.B(_1715_),
    .C(_1725_),
    .A(_1710_),
    .Y(_1842_));
 sg13g2_nor4_2 _4831_ (.A(net1170),
    .B(_1837_),
    .C(_1841_),
    .Y(_1843_),
    .D(_1842_));
 sg13g2_inv_1 _4832_ (.Y(_1844_),
    .A(_1843_));
 sg13g2_o21ai_1 _4833_ (.B1(net1267),
    .Y(_1845_),
    .A1(net1376),
    .A2(_1839_));
 sg13g2_a21oi_1 _4834_ (.A1(net1376),
    .A2(_1844_),
    .Y(_0030_),
    .B1(_1845_));
 sg13g2_and2_1 _4835_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0750_),
    .X(_1846_));
 sg13g2_xor2_1 _4836_ (.B(_0750_),
    .A(net1812),
    .X(_1847_));
 sg13g2_xnor2_1 _4837_ (.Y(_1848_),
    .A(_0666_),
    .B(_1847_));
 sg13g2_a22oi_1 _4838_ (.Y(_1849_),
    .B1(_1848_),
    .B2(_1839_),
    .A2(_1843_),
    .A1(net1812));
 sg13g2_nor2_1 _4839_ (.A(net1251),
    .B(_1849_),
    .Y(_0031_));
 sg13g2_nand2_1 _4840_ (.Y(_1850_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .B(_0750_));
 sg13g2_nor2_1 _4841_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .B(_0750_),
    .Y(_1851_));
 sg13g2_xnor2_1 _4842_ (.Y(_1852_),
    .A(_0665_),
    .B(_0750_));
 sg13g2_a21oi_1 _4843_ (.A1(net1376),
    .A2(_1847_),
    .Y(_1853_),
    .B1(_1846_));
 sg13g2_xnor2_1 _4844_ (.Y(_1854_),
    .A(_1852_),
    .B(_1853_));
 sg13g2_a22oi_1 _4845_ (.Y(_1855_),
    .B1(_1854_),
    .B2(_1839_),
    .A2(_1843_),
    .A1(net1797));
 sg13g2_nor2_1 _4846_ (.A(net1247),
    .B(_1855_),
    .Y(_0032_));
 sg13g2_and2_1 _4847_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .B(_0750_),
    .X(_1856_));
 sg13g2_xnor2_1 _4848_ (.Y(_1857_),
    .A(_0664_),
    .B(_0750_));
 sg13g2_o21ai_1 _4849_ (.B1(_1850_),
    .Y(_1858_),
    .A1(_1851_),
    .A2(_1853_));
 sg13g2_xor2_1 _4850_ (.B(_1858_),
    .A(_1857_),
    .X(_1859_));
 sg13g2_a22oi_1 _4851_ (.Y(_1860_),
    .B1(_1859_),
    .B2(_1839_),
    .A2(_1843_),
    .A1(net1755));
 sg13g2_nor2_1 _4852_ (.A(net1247),
    .B(net1756),
    .Y(_0033_));
 sg13g2_a21oi_1 _4853_ (.A1(_1857_),
    .A2(_1858_),
    .Y(_1861_),
    .B1(_1856_));
 sg13g2_xor2_1 _4854_ (.B(_0750_),
    .A(net1823),
    .X(_1862_));
 sg13g2_xnor2_1 _4855_ (.Y(_1863_),
    .A(_1861_),
    .B(_1862_));
 sg13g2_a22oi_1 _4856_ (.Y(_1864_),
    .B1(_1863_),
    .B2(_1839_),
    .A2(_1843_),
    .A1(net1823));
 sg13g2_nor2_1 _4857_ (.A(net1247),
    .B(_1864_),
    .Y(_0034_));
 sg13g2_nor2_1 _4858_ (.A(_1709_),
    .B(_1762_),
    .Y(_1865_));
 sg13g2_a21oi_1 _4859_ (.A1(net1618),
    .A2(net1610),
    .Y(_1866_),
    .B1(_1710_));
 sg13g2_a22oi_1 _4860_ (.Y(_1867_),
    .B1(_1866_),
    .B2(net1624),
    .A2(_1865_),
    .A1(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ));
 sg13g2_nor2_1 _4861_ (.A(_1753_),
    .B(net1625),
    .Y(_0035_));
 sg13g2_a22oi_1 _4862_ (.Y(_1868_),
    .B1(_1865_),
    .B2(net1745),
    .A2(_1709_),
    .A1(net1610));
 sg13g2_nor2_1 _4863_ (.A(_1753_),
    .B(_1868_),
    .Y(_0036_));
 sg13g2_a22oi_1 _4864_ (.Y(_1869_),
    .B1(_1865_),
    .B2(net1655),
    .A2(_1709_),
    .A1(net1618));
 sg13g2_nor2_1 _4865_ (.A(_1753_),
    .B(net1656),
    .Y(_0037_));
 sg13g2_nand4_1 _4866_ (.B(_0668_),
    .C(_0745_),
    .A(net1242),
    .Y(_1870_),
    .D(_1755_));
 sg13g2_inv_1 _4867_ (.Y(_1871_),
    .A(_1870_));
 sg13g2_nor3_1 _4868_ (.A(net1236),
    .B(net1237),
    .C(_1546_),
    .Y(_1872_));
 sg13g2_nand2_2 _4869_ (.Y(_1873_),
    .A(net1650),
    .B(_1695_));
 sg13g2_and2_1 _4870_ (.A(_1870_),
    .B(_1873_),
    .X(_1874_));
 sg13g2_a22oi_1 _4871_ (.Y(_1875_),
    .B1(_1871_),
    .B2(_1595_),
    .A2(_1606_),
    .A1(_1593_));
 sg13g2_o21ai_1 _4872_ (.B1(_1870_),
    .Y(_1876_),
    .A1(_1872_),
    .A2(_1873_));
 sg13g2_a221oi_1 _4873_ (.B2(_1876_),
    .C1(_1752_),
    .B1(_1875_),
    .A1(_0661_),
    .Y(_0038_),
    .A2(_1874_));
 sg13g2_nor2_1 _4874_ (.A(net1843),
    .B(_1872_),
    .Y(_1877_));
 sg13g2_nor2_1 _4875_ (.A(_1595_),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_nand4_1 _4876_ (.B(_1587_),
    .C(_1624_),
    .A(net1650),
    .Y(_1879_),
    .D(_1695_));
 sg13g2_a22oi_1 _4877_ (.Y(_1880_),
    .B1(_1878_),
    .B2(_1871_),
    .A2(_1874_),
    .A1(net1843));
 sg13g2_a21oi_1 _4878_ (.A1(_1879_),
    .A2(_1880_),
    .Y(_0039_),
    .B1(_1752_));
 sg13g2_a221oi_1 _4879_ (.B2(_1736_),
    .C1(_1695_),
    .B1(_1700_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .Y(_1881_),
    .A2(_0752_));
 sg13g2_a221oi_1 _4880_ (.B2(_1705_),
    .C1(_1881_),
    .B1(_1702_),
    .A1(_0739_),
    .Y(_1882_),
    .A2(_0741_));
 sg13g2_nand2b_1 _4881_ (.Y(_1883_),
    .B(_0742_),
    .A_N(_1692_));
 sg13g2_nand2b_2 _4882_ (.Y(_1884_),
    .B(_1883_),
    .A_N(_1545_));
 sg13g2_o21ai_1 _4883_ (.B1(_1711_),
    .Y(_1885_),
    .A1(net1181),
    .A2(_1723_));
 sg13g2_nor4_1 _4884_ (.A(_1743_),
    .B(_1882_),
    .C(_1884_),
    .D(_1885_),
    .Y(_1886_));
 sg13g2_nor2_1 _4885_ (.A(net1796),
    .B(_1730_),
    .Y(_1887_));
 sg13g2_nor3_1 _4886_ (.A(_1748_),
    .B(_1886_),
    .C(_1887_),
    .Y(_0040_));
 sg13g2_nor2_1 _4887_ (.A(net1234),
    .B(_1730_),
    .Y(_1888_));
 sg13g2_o21ai_1 _4888_ (.B1(_1700_),
    .Y(_1889_),
    .A1(net1227),
    .A2(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ));
 sg13g2_a21oi_1 _4889_ (.A1(_1711_),
    .A2(_1889_),
    .Y(_1890_),
    .B1(_1712_));
 sg13g2_nor3_1 _4890_ (.A(_1729_),
    .B(_1842_),
    .C(_1890_),
    .Y(_1891_));
 sg13g2_nor3_1 _4891_ (.A(_1748_),
    .B(_1888_),
    .C(_1891_),
    .Y(_0041_));
 sg13g2_nand3_1 _4892_ (.B(_1758_),
    .C(_1765_),
    .A(_1756_),
    .Y(_1892_));
 sg13g2_nor2_1 _4893_ (.A(net1905),
    .B(_1762_),
    .Y(_1893_));
 sg13g2_nand2_1 _4894_ (.Y(_1894_),
    .A(_1710_),
    .B(_1751_));
 sg13g2_xnor2_1 _4895_ (.Y(_1895_),
    .A(_1892_),
    .B(_1893_));
 sg13g2_o21ai_1 _4896_ (.B1(net1267),
    .Y(_1896_),
    .A1(_1894_),
    .A2(_1895_));
 sg13g2_inv_1 _4897_ (.Y(_0042_),
    .A(_1896_));
 sg13g2_nor2b_2 _4898_ (.A(_1559_),
    .B_N(_1564_),
    .Y(_1897_));
 sg13g2_or2_1 _4899_ (.X(_1898_),
    .B(_1762_),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ));
 sg13g2_o21ai_1 _4900_ (.B1(_1705_),
    .Y(_1899_),
    .A1(_1703_),
    .A2(_1897_));
 sg13g2_a21oi_1 _4901_ (.A1(_1704_),
    .A2(_1897_),
    .Y(_1900_),
    .B1(_1899_));
 sg13g2_a21oi_1 _4902_ (.A1(_1765_),
    .A2(_1898_),
    .Y(_1901_),
    .B1(_1900_));
 sg13g2_o21ai_1 _4903_ (.B1(_1758_),
    .Y(_1902_),
    .A1(_1756_),
    .A2(_1897_));
 sg13g2_a21oi_1 _4904_ (.A1(_1756_),
    .A2(_1901_),
    .Y(_1903_),
    .B1(_1902_));
 sg13g2_nor2_1 _4905_ (.A(_1758_),
    .B(_1897_),
    .Y(_1904_));
 sg13g2_nor3_1 _4906_ (.A(_1894_),
    .B(_1903_),
    .C(_1904_),
    .Y(_1905_));
 sg13g2_nor2_1 _4907_ (.A(net1251),
    .B(_1905_),
    .Y(_0043_));
 sg13g2_a21o_2 _4908_ (.A2(net1162),
    .A1(_1692_),
    .B1(net1252),
    .X(_1906_));
 sg13g2_xnor2_1 _4909_ (.Y(_1907_),
    .A(net1728),
    .B(net1226));
 sg13g2_nor2_1 _4910_ (.A(_1906_),
    .B(_1907_),
    .Y(_0044_));
 sg13g2_a21oi_1 _4911_ (.A1(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .A2(net1226),
    .Y(_1908_),
    .B1(net1548));
 sg13g2_and3_1 _4912_ (.X(_1909_),
    .A(net1548),
    .B(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .C(net1226));
 sg13g2_nor3_1 _4913_ (.A(_1906_),
    .B(net1549),
    .C(_1909_),
    .Y(_0045_));
 sg13g2_nor2_1 _4914_ (.A(net1678),
    .B(_1909_),
    .Y(_1910_));
 sg13g2_and2_1 _4915_ (.A(net1678),
    .B(_1909_),
    .X(_1911_));
 sg13g2_nor3_1 _4916_ (.A(_1906_),
    .B(net1679),
    .C(_1911_),
    .Y(_0046_));
 sg13g2_nor2_1 _4917_ (.A(net1712),
    .B(_1911_),
    .Y(_1912_));
 sg13g2_and2_1 _4918_ (.A(net1712),
    .B(_1911_),
    .X(_1913_));
 sg13g2_nor3_1 _4919_ (.A(_1906_),
    .B(net1713),
    .C(_1913_),
    .Y(_0047_));
 sg13g2_nor2_1 _4920_ (.A(net1741),
    .B(_1913_),
    .Y(_1914_));
 sg13g2_and2_1 _4921_ (.A(net1741),
    .B(_1913_),
    .X(_1915_));
 sg13g2_nor3_1 _4922_ (.A(_1906_),
    .B(_1914_),
    .C(_1915_),
    .Y(_0048_));
 sg13g2_xnor2_1 _4923_ (.Y(_1916_),
    .A(net1735),
    .B(_1915_));
 sg13g2_nor2_1 _4924_ (.A(_1906_),
    .B(net1736),
    .Y(_0049_));
 sg13g2_xnor2_1 _4925_ (.Y(_1917_),
    .A(net1601),
    .B(net1666));
 sg13g2_xnor2_1 _4926_ (.Y(_1918_),
    .A(net1631),
    .B(net1524));
 sg13g2_xnor2_1 _4927_ (.Y(_1919_),
    .A(_1917_),
    .B(_1918_));
 sg13g2_a21oi_1 _4928_ (.A1(net1624),
    .A2(net1182),
    .Y(_1920_),
    .B1(net1254));
 sg13g2_o21ai_1 _4929_ (.B1(_1920_),
    .Y(_0050_),
    .A1(net1183),
    .A2(_1919_));
 sg13g2_o21ai_1 _4930_ (.B1(net1270),
    .Y(_1921_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .A2(net1183));
 sg13g2_a21oi_1 _4931_ (.A1(_0658_),
    .A2(net1185),
    .Y(_0051_),
    .B1(_1921_));
 sg13g2_o21ai_1 _4932_ (.B1(net1270),
    .Y(_1922_),
    .A1(net1610),
    .A2(net1186));
 sg13g2_a21oi_1 _4933_ (.A1(_0657_),
    .A2(net1186),
    .Y(_0052_),
    .B1(_1922_));
 sg13g2_o21ai_1 _4934_ (.B1(net1270),
    .Y(_1923_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .A2(net1186));
 sg13g2_a21oi_1 _4935_ (.A1(_0656_),
    .A2(net1186),
    .Y(_0053_),
    .B1(_1923_));
 sg13g2_o21ai_1 _4936_ (.B1(net1269),
    .Y(_1924_),
    .A1(net1331),
    .A2(net1186));
 sg13g2_a21oi_1 _4937_ (.A1(_0655_),
    .A2(net1186),
    .Y(_0054_),
    .B1(_1924_));
 sg13g2_a21oi_1 _4938_ (.A1(net1399),
    .A2(net1185),
    .Y(_1925_),
    .B1(net1255));
 sg13g2_o21ai_1 _4939_ (.B1(_1925_),
    .Y(_0055_),
    .A1(_0655_),
    .A2(net1186));
 sg13g2_a21oi_1 _4940_ (.A1(net1410),
    .A2(net1185),
    .Y(_1926_),
    .B1(net1256));
 sg13g2_o21ai_1 _4941_ (.B1(_1926_),
    .Y(_0056_),
    .A1(_0654_),
    .A2(net1185));
 sg13g2_a21oi_1 _4942_ (.A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .A2(net1185),
    .Y(_1927_),
    .B1(net1256));
 sg13g2_o21ai_1 _4943_ (.B1(_1927_),
    .Y(_0057_),
    .A1(_0653_),
    .A2(net1184));
 sg13g2_o21ai_1 _4944_ (.B1(net1270),
    .Y(_1928_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .A2(net1185));
 sg13g2_a21oi_1 _4945_ (.A1(_0652_),
    .A2(net1184),
    .Y(_0058_),
    .B1(_1928_));
 sg13g2_o21ai_1 _4946_ (.B1(net1270),
    .Y(_1929_),
    .A1(net1367),
    .A2(net1184));
 sg13g2_a21oi_1 _4947_ (.A1(_0651_),
    .A2(net1184),
    .Y(_0059_),
    .B1(_1929_));
 sg13g2_a21oi_1 _4948_ (.A1(net1524),
    .A2(net1184),
    .Y(_1930_),
    .B1(net1256));
 sg13g2_o21ai_1 _4949_ (.B1(_1930_),
    .Y(_0060_),
    .A1(_0651_),
    .A2(net1184));
 sg13g2_a21oi_1 _4950_ (.A1(net1676),
    .A2(net1184),
    .Y(_1931_),
    .B1(net1256));
 sg13g2_o21ai_1 _4951_ (.B1(_1931_),
    .Y(_0061_),
    .A1(_0650_),
    .A2(net1184));
 sg13g2_o21ai_1 _4952_ (.B1(net1270),
    .Y(_1932_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .A2(net1182));
 sg13g2_a21oi_1 _4953_ (.A1(_0649_),
    .A2(net1183),
    .Y(_0062_),
    .B1(_1932_));
 sg13g2_a21oi_1 _4954_ (.A1(net1666),
    .A2(net1182),
    .Y(_1933_),
    .B1(net1254));
 sg13g2_o21ai_1 _4955_ (.B1(_1933_),
    .Y(_0063_),
    .A1(_0649_),
    .A2(net1182));
 sg13g2_o21ai_1 _4956_ (.B1(net1268),
    .Y(_1934_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .A2(net1182));
 sg13g2_a21oi_1 _4957_ (.A1(_0648_),
    .A2(net1182),
    .Y(_0064_),
    .B1(_1934_));
 sg13g2_a21oi_1 _4958_ (.A1(net1601),
    .A2(net1182),
    .Y(_1935_),
    .B1(net1254));
 sg13g2_o21ai_1 _4959_ (.B1(_1935_),
    .Y(_0065_),
    .A1(_0648_),
    .A2(net1182));
 sg13g2_nand2b_2 _4960_ (.Y(_1936_),
    .B(net744),
    .A_N(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ));
 sg13g2_nand2_1 _4961_ (.Y(_1937_),
    .A(net1700),
    .B(net1850));
 sg13g2_nor3_1 _4962_ (.A(net1253),
    .B(_1936_),
    .C(net1701),
    .Y(_0066_));
 sg13g2_or2_1 _4963_ (.X(_1938_),
    .B(_1884_),
    .A(net1723));
 sg13g2_nor2_1 _4964_ (.A(net744),
    .B(_1938_),
    .Y(_1939_));
 sg13g2_o21ai_1 _4965_ (.B1(net1198),
    .Y(_1940_),
    .A1(_1936_),
    .A2(net1701));
 sg13g2_nor3_1 _4966_ (.A(net1253),
    .B(_1939_),
    .C(_1940_),
    .Y(_0067_));
 sg13g2_nand2_1 _4967_ (.Y(_1941_),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .B(net1268));
 sg13g2_a21oi_1 _4968_ (.A1(net744),
    .A2(_1938_),
    .Y(_0068_),
    .B1(_1941_));
 sg13g2_nor2b_1 _4969_ (.A(_1936_),
    .B_N(_1937_),
    .Y(_1942_));
 sg13g2_o21ai_1 _4970_ (.B1(net1806),
    .Y(_1943_),
    .A1(_1938_),
    .A2(_1942_));
 sg13g2_nand2b_1 _4971_ (.Y(_1944_),
    .B(_1936_),
    .A_N(net1806));
 sg13g2_and3_1 _4972_ (.X(_0069_),
    .A(net1267),
    .B(net1807),
    .C(_1944_));
 sg13g2_o21ai_1 _4973_ (.B1(_1942_),
    .Y(_1945_),
    .A1(net1700),
    .A2(net1806));
 sg13g2_o21ai_1 _4974_ (.B1(_1945_),
    .Y(_1946_),
    .A1(_0647_),
    .A2(_1938_));
 sg13g2_and2_1 _4975_ (.A(net1268),
    .B(_1946_),
    .X(_0070_));
 sg13g2_nand2_1 _4976_ (.Y(_1947_),
    .A(_1570_),
    .B(net1082));
 sg13g2_a21oi_1 _4977_ (.A1(net1238),
    .A2(_1546_),
    .Y(_1948_),
    .B1(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ));
 sg13g2_o21ai_1 _4978_ (.B1(_1948_),
    .Y(_1949_),
    .A1(net1238),
    .A2(_1585_));
 sg13g2_mux2_1 _4979_ (.A0(net1167),
    .A1(_1003_),
    .S(_1947_),
    .X(_1950_));
 sg13g2_nor2_1 _4980_ (.A(net1200),
    .B(_1950_),
    .Y(_1951_));
 sg13g2_a21oi_1 _4981_ (.A1(net1596),
    .A2(net1200),
    .Y(_1952_),
    .B1(_1951_));
 sg13g2_nor2_1 _4982_ (.A(net1251),
    .B(net1597),
    .Y(_0071_));
 sg13g2_a21oi_1 _4983_ (.A1(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .A2(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1953_),
    .B1(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ));
 sg13g2_nand3_1 _4984_ (.B(_1606_),
    .C(_1953_),
    .A(_1547_),
    .Y(_1954_));
 sg13g2_mux2_1 _4985_ (.A0(net1166),
    .A1(_1423_),
    .S(_1947_),
    .X(_1955_));
 sg13g2_nor2_1 _4986_ (.A(net1198),
    .B(_1955_),
    .Y(_1956_));
 sg13g2_a21oi_1 _4987_ (.A1(net1509),
    .A2(net1198),
    .Y(_1957_),
    .B1(_1956_));
 sg13g2_nor2_1 _4988_ (.A(net1253),
    .B(_1957_),
    .Y(_0072_));
 sg13g2_and2_1 _4989_ (.A(_1570_),
    .B(_1640_),
    .X(_1958_));
 sg13g2_a21o_2 _4990_ (.A2(net1082),
    .A1(_1577_),
    .B1(_1958_),
    .X(_1959_));
 sg13g2_nand2b_1 _4991_ (.Y(_1960_),
    .B(_0938_),
    .A_N(_1959_));
 sg13g2_a21oi_1 _4992_ (.A1(net1167),
    .A2(_1959_),
    .Y(_1961_),
    .B1(net1199));
 sg13g2_a22oi_1 _4993_ (.Y(_1962_),
    .B1(_1960_),
    .B2(_1961_),
    .A2(net1199),
    .A1(net1746));
 sg13g2_nor2_1 _4994_ (.A(net1254),
    .B(_1962_),
    .Y(_0073_));
 sg13g2_nand2b_1 _4995_ (.Y(_1963_),
    .B(_1335_),
    .A_N(_1959_));
 sg13g2_a21oi_1 _4996_ (.A1(net1166),
    .A2(_1959_),
    .Y(_1964_),
    .B1(net1199));
 sg13g2_a22oi_1 _4997_ (.Y(_1965_),
    .B1(_1963_),
    .B2(_1964_),
    .A2(net1199),
    .A1(net1672));
 sg13g2_nor2_1 _4998_ (.A(net1253),
    .B(_1965_),
    .Y(_0074_));
 sg13g2_nand2_1 _4999_ (.Y(_1966_),
    .A(net1391),
    .B(net1197));
 sg13g2_nand2_1 _5000_ (.Y(_1967_),
    .A(_1570_),
    .B(net1087));
 sg13g2_a22oi_1 _5001_ (.Y(_1968_),
    .B1(net1086),
    .B2(_1577_),
    .A2(net1081),
    .A1(_1554_));
 sg13g2_nand2_2 _5002_ (.Y(_1969_),
    .A(_1967_),
    .B(_1968_));
 sg13g2_a21oi_1 _5003_ (.A1(net1167),
    .A2(_1969_),
    .Y(_1970_),
    .B1(net1197));
 sg13g2_o21ai_1 _5004_ (.B1(_1970_),
    .Y(_1971_),
    .A1(_1123_),
    .A2(_1969_));
 sg13g2_a21oi_1 _5005_ (.A1(_1966_),
    .A2(_1971_),
    .Y(_0075_),
    .B1(net1247));
 sg13g2_nand2_1 _5006_ (.Y(_1972_),
    .A(net1466),
    .B(net1197));
 sg13g2_a21oi_1 _5007_ (.A1(net1166),
    .A2(_1969_),
    .Y(_1973_),
    .B1(_0889_));
 sg13g2_o21ai_1 _5008_ (.B1(_1973_),
    .Y(_1974_),
    .A1(_1360_),
    .A2(_1969_));
 sg13g2_a21oi_1 _5009_ (.A1(_1972_),
    .A2(_1974_),
    .Y(_0076_),
    .B1(net1247));
 sg13g2_nand2_1 _5010_ (.Y(_1975_),
    .A(net1398),
    .B(net1195));
 sg13g2_a22oi_1 _5011_ (.Y(_1976_),
    .B1(_1576_),
    .B2(net1081),
    .A2(_1570_),
    .A1(net1090));
 sg13g2_a22oi_1 _5012_ (.Y(_1977_),
    .B1(net1086),
    .B2(_1554_),
    .A2(net1087),
    .A1(_1577_));
 sg13g2_nand2_2 _5013_ (.Y(_1978_),
    .A(_1976_),
    .B(_1977_));
 sg13g2_a21oi_1 _5014_ (.A1(net1167),
    .A2(_1978_),
    .Y(_1979_),
    .B1(net1195));
 sg13g2_o21ai_1 _5015_ (.B1(_1979_),
    .Y(_1980_),
    .A1(_0966_),
    .A2(_1978_));
 sg13g2_a21oi_1 _5016_ (.A1(_1975_),
    .A2(_1980_),
    .Y(_0077_),
    .B1(net1246));
 sg13g2_nand2_1 _5017_ (.Y(_1981_),
    .A(net1393),
    .B(net1195));
 sg13g2_a21oi_1 _5018_ (.A1(net1166),
    .A2(_1978_),
    .Y(_1982_),
    .B1(net1195));
 sg13g2_o21ai_1 _5019_ (.B1(_1982_),
    .Y(_1983_),
    .A1(_1389_),
    .A2(_1978_));
 sg13g2_a21oi_1 _5020_ (.A1(_1981_),
    .A2(_1983_),
    .Y(_0078_),
    .B1(net1246));
 sg13g2_a22oi_1 _5021_ (.Y(_1984_),
    .B1(net1081),
    .B2(_1560_),
    .A2(_1577_),
    .A1(net1090));
 sg13g2_a22oi_1 _5022_ (.Y(_1985_),
    .B1(net1086),
    .B2(_1576_),
    .A2(net1087),
    .A1(_1554_));
 sg13g2_nand2_2 _5023_ (.Y(_1986_),
    .A(_1984_),
    .B(_1985_));
 sg13g2_nand2b_1 _5024_ (.Y(_1987_),
    .B(_1048_),
    .A_N(_1986_));
 sg13g2_a21oi_1 _5025_ (.A1(net1167),
    .A2(_1986_),
    .Y(_1988_),
    .B1(net1200));
 sg13g2_a22oi_1 _5026_ (.Y(_1989_),
    .B1(_1987_),
    .B2(_1988_),
    .A2(net1200),
    .A1(net1633));
 sg13g2_nor2_1 _5027_ (.A(net1251),
    .B(net1634),
    .Y(_0079_));
 sg13g2_nand2_1 _5028_ (.Y(_1990_),
    .A(net1381),
    .B(net1200));
 sg13g2_a21oi_1 _5029_ (.A1(_1954_),
    .A2(_1986_),
    .Y(_1991_),
    .B1(net1200));
 sg13g2_o21ai_1 _5030_ (.B1(_1991_),
    .Y(_1992_),
    .A1(_1465_),
    .A2(_1986_));
 sg13g2_a21oi_1 _5031_ (.A1(_1990_),
    .A2(_1992_),
    .Y(_0080_),
    .B1(net1251));
 sg13g2_nand2_1 _5032_ (.Y(_1993_),
    .A(net1515),
    .B(net1195));
 sg13g2_a21oi_2 _5033_ (.B1(_1567_),
    .Y(_1994_),
    .A2(_1557_),
    .A1(_0700_));
 sg13g2_a22oi_1 _5034_ (.Y(_1995_),
    .B1(net1081),
    .B2(_1994_),
    .A2(_1554_),
    .A1(net1090));
 sg13g2_a22oi_1 _5035_ (.Y(_1996_),
    .B1(net1086),
    .B2(_1560_),
    .A2(net1087),
    .A1(_1576_));
 sg13g2_nand2_2 _5036_ (.Y(_1997_),
    .A(_1995_),
    .B(_1996_));
 sg13g2_a21oi_1 _5037_ (.A1(net1167),
    .A2(_1997_),
    .Y(_1998_),
    .B1(net1195));
 sg13g2_o21ai_1 _5038_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_1031_),
    .A2(_1997_));
 sg13g2_a21oi_1 _5039_ (.A1(_1993_),
    .A2(_1999_),
    .Y(_0081_),
    .B1(net1246));
 sg13g2_nand2_1 _5040_ (.Y(_2000_),
    .A(net1423),
    .B(net1195));
 sg13g2_a21oi_1 _5041_ (.A1(net1166),
    .A2(_1997_),
    .Y(_2001_),
    .B1(net1196));
 sg13g2_o21ai_1 _5042_ (.B1(_2001_),
    .Y(_2002_),
    .A1(_1527_),
    .A2(_1997_));
 sg13g2_a21oi_1 _5043_ (.A1(_2000_),
    .A2(_2002_),
    .Y(_0082_),
    .B1(net1246));
 sg13g2_nand2_1 _5044_ (.Y(_2003_),
    .A(net1430),
    .B(net1197));
 sg13g2_a22oi_1 _5045_ (.Y(_2004_),
    .B1(net1081),
    .B2(_1652_),
    .A2(_1576_),
    .A1(net1090));
 sg13g2_a22oi_1 _5046_ (.Y(_2005_),
    .B1(net1086),
    .B2(_1994_),
    .A2(net1087),
    .A1(_1560_));
 sg13g2_nand2_2 _5047_ (.Y(_2006_),
    .A(_2004_),
    .B(_2005_));
 sg13g2_a21oi_1 _5048_ (.A1(net1167),
    .A2(_2006_),
    .Y(_2007_),
    .B1(net1197));
 sg13g2_o21ai_1 _5049_ (.B1(_2007_),
    .Y(_2008_),
    .A1(_0916_),
    .A2(_2006_));
 sg13g2_a21oi_1 _5050_ (.A1(_2003_),
    .A2(_2008_),
    .Y(_0083_),
    .B1(net1251));
 sg13g2_nand2b_1 _5051_ (.Y(_2009_),
    .B(_1406_),
    .A_N(_2006_));
 sg13g2_a21oi_1 _5052_ (.A1(net1166),
    .A2(_2006_),
    .Y(_2010_),
    .B1(net1197));
 sg13g2_a22oi_1 _5053_ (.Y(_2011_),
    .B1(_2009_),
    .B2(_2010_),
    .A2(net1197),
    .A1(net1643));
 sg13g2_nor2_1 _5054_ (.A(net1251),
    .B(net1644),
    .Y(_0084_));
 sg13g2_a22oi_1 _5055_ (.Y(_2012_),
    .B1(net1082),
    .B2(_1644_),
    .A2(_1560_),
    .A1(net1091));
 sg13g2_a22oi_1 _5056_ (.Y(_2013_),
    .B1(_1994_),
    .B2(_1601_),
    .A2(_1652_),
    .A1(_1640_));
 sg13g2_nand2_2 _5057_ (.Y(_2014_),
    .A(_2012_),
    .B(_2013_));
 sg13g2_nand2b_1 _5058_ (.Y(_2015_),
    .B(_0985_),
    .A_N(_2014_));
 sg13g2_a21oi_1 _5059_ (.A1(_1949_),
    .A2(_2014_),
    .Y(_2016_),
    .B1(net1199));
 sg13g2_a22oi_1 _5060_ (.Y(_2017_),
    .B1(_2015_),
    .B2(_2016_),
    .A2(net1199),
    .A1(net1651));
 sg13g2_nor2_1 _5061_ (.A(net1253),
    .B(net1652),
    .Y(_0085_));
 sg13g2_nand2b_1 _5062_ (.Y(_2018_),
    .B(_1499_),
    .A_N(_2014_));
 sg13g2_a21oi_1 _5063_ (.A1(_1954_),
    .A2(_2014_),
    .Y(_2019_),
    .B1(net1199));
 sg13g2_a22oi_1 _5064_ (.Y(_2020_),
    .B1(_2018_),
    .B2(_2019_),
    .A2(net1198),
    .A1(net1648));
 sg13g2_nor2_1 _5065_ (.A(net1253),
    .B(net1649),
    .Y(_0086_));
 sg13g2_a22oi_1 _5066_ (.Y(_2021_),
    .B1(_1994_),
    .B2(net1090),
    .A2(_1661_),
    .A1(net1082));
 sg13g2_a22oi_1 _5067_ (.Y(_2022_),
    .B1(_1652_),
    .B2(_1601_),
    .A2(_1644_),
    .A1(_1640_));
 sg13g2_nand2_2 _5068_ (.Y(_2023_),
    .A(_2021_),
    .B(_2022_));
 sg13g2_nand2b_1 _5069_ (.Y(_2024_),
    .B(_1095_),
    .A_N(_2023_));
 sg13g2_a21oi_1 _5070_ (.A1(_1949_),
    .A2(_2023_),
    .Y(_2025_),
    .B1(net1198));
 sg13g2_a22oi_1 _5071_ (.Y(_2026_),
    .B1(_2024_),
    .B2(_2025_),
    .A2(net1198),
    .A1(net1638));
 sg13g2_nor2_1 _5072_ (.A(net1253),
    .B(net1639),
    .Y(_0087_));
 sg13g2_nand2b_1 _5073_ (.Y(_2027_),
    .B(_1482_),
    .A_N(_2023_));
 sg13g2_a21oi_1 _5074_ (.A1(net1166),
    .A2(_2023_),
    .Y(_2028_),
    .B1(net1198));
 sg13g2_a22oi_1 _5075_ (.Y(_2029_),
    .B1(_2027_),
    .B2(_2028_),
    .A2(net1198),
    .A1(net1630));
 sg13g2_nor2_1 _5076_ (.A(net1253),
    .B(_2029_),
    .Y(_0088_));
 sg13g2_nand2_1 _5077_ (.Y(_2030_),
    .A(net1484),
    .B(net1196));
 sg13g2_nand2b_1 _5078_ (.Y(_2031_),
    .B(net1081),
    .A_N(_1668_));
 sg13g2_nand2_1 _5079_ (.Y(_2032_),
    .A(net1086),
    .B(_1661_));
 sg13g2_nand3_1 _5080_ (.B(_2031_),
    .C(_2032_),
    .A(_1659_),
    .Y(_2033_));
 sg13g2_a21oi_1 _5081_ (.A1(net1167),
    .A2(_2033_),
    .Y(_2034_),
    .B1(net1196));
 sg13g2_o21ai_1 _5082_ (.B1(_2034_),
    .Y(_2035_),
    .A1(_1076_),
    .A2(_2033_));
 sg13g2_a21oi_1 _5083_ (.A1(_2030_),
    .A2(_2035_),
    .Y(_0089_),
    .B1(net1246));
 sg13g2_nand2_1 _5084_ (.Y(_2036_),
    .A(net1414),
    .B(net1195));
 sg13g2_a21oi_1 _5085_ (.A1(net1166),
    .A2(_2033_),
    .Y(_2037_),
    .B1(net1196));
 sg13g2_o21ai_1 _5086_ (.B1(_2037_),
    .Y(_2038_),
    .A1(_1449_),
    .A2(_2033_));
 sg13g2_a21oi_1 _5087_ (.A1(_2036_),
    .A2(_2038_),
    .Y(_0090_),
    .B1(net1246));
 sg13g2_nand2_1 _5088_ (.Y(_2039_),
    .A(net1714),
    .B(net1388));
 sg13g2_o21ai_1 _5089_ (.B1(net1227),
    .Y(_2040_),
    .A1(net1732),
    .A2(_2039_));
 sg13g2_nand3_1 _5090_ (.B(_1543_),
    .C(_2040_),
    .A(net1227),
    .Y(_2041_));
 sg13g2_o21ai_1 _5091_ (.B1(net1750),
    .Y(_2042_),
    .A1(net1227),
    .A2(_1699_));
 sg13g2_a21oi_1 _5092_ (.A1(_2041_),
    .A2(net1751),
    .Y(_0091_),
    .B1(net1252));
 sg13g2_nor2b_1 _5093_ (.A(_1719_),
    .B_N(_1873_),
    .Y(_2043_));
 sg13g2_nand4_1 _5094_ (.B(_1734_),
    .C(_1764_),
    .A(_1693_),
    .Y(_2044_),
    .D(_2043_));
 sg13g2_a21oi_1 _5095_ (.A1(net1437),
    .A2(net1285),
    .Y(_2045_),
    .B1(_1687_));
 sg13g2_nand2_1 _5096_ (.Y(_2046_),
    .A(net1602),
    .B(net1265));
 sg13g2_a21oi_1 _5097_ (.A1(net1602),
    .A2(_2045_),
    .Y(_2047_),
    .B1(_2044_));
 sg13g2_nor2_1 _5098_ (.A(net1252),
    .B(_2047_),
    .Y(_0092_));
 sg13g2_nor3_1 _5099_ (.A(net1799),
    .B(_0706_),
    .C(_1884_),
    .Y(_2048_));
 sg13g2_o21ai_1 _5100_ (.B1(net1269),
    .Y(_2049_),
    .A1(net1723),
    .A2(net1800));
 sg13g2_inv_1 _5101_ (.Y(_0093_),
    .A(_2049_));
 sg13g2_a21o_1 _5102_ (.A2(_1687_),
    .A1(_0646_),
    .B1(_2046_),
    .X(_2050_));
 sg13g2_a21oi_1 _5103_ (.A1(net1285),
    .A2(_2045_),
    .Y(_0094_),
    .B1(_2050_));
 sg13g2_a21oi_1 _5104_ (.A1(net1285),
    .A2(_1688_),
    .Y(_2051_),
    .B1(net1437));
 sg13g2_nor2_1 _5105_ (.A(_2046_),
    .B(_2051_),
    .Y(_0095_));
 sg13g2_a21oi_1 _5106_ (.A1(net1230),
    .A2(_1723_),
    .Y(_2052_),
    .B1(_1712_));
 sg13g2_nor2_1 _5107_ (.A(net1247),
    .B(net1879),
    .Y(_0096_));
 sg13g2_or4_1 _5108_ (.A(_1563_),
    .B(_1654_),
    .C(_1663_),
    .D(_1675_),
    .X(_2053_));
 sg13g2_or4_1 _5109_ (.A(_1561_),
    .B(_1574_),
    .C(_1578_),
    .D(_1647_),
    .X(_2054_));
 sg13g2_a21o_2 _5110_ (.A2(_1482_),
    .A1(_1095_),
    .B1(_1552_),
    .X(_2055_));
 sg13g2_or3_1 _5111_ (.A(_2053_),
    .B(_2054_),
    .C(_2055_),
    .X(_2056_));
 sg13g2_and2_1 _5112_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .X(_2057_));
 sg13g2_nand4_1 _5113_ (.B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .C(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .Y(_2058_),
    .D(_2057_));
 sg13g2_or2_1 _5114_ (.X(_2059_),
    .B(_2058_),
    .A(_0894_));
 sg13g2_or2_1 _5115_ (.X(_2060_),
    .B(_2059_),
    .A(_2056_));
 sg13g2_inv_1 _5116_ (.Y(_2061_),
    .A(_2060_));
 sg13g2_nor3_1 _5117_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B(net1229),
    .C(net1873),
    .Y(_2062_));
 sg13g2_nand2_1 _5118_ (.Y(_2063_),
    .A(_0670_),
    .B(_2062_));
 sg13g2_nor2_2 _5119_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_inv_1 _5120_ (.Y(_2065_),
    .A(_2064_));
 sg13g2_nor2_2 _5121_ (.A(_0724_),
    .B(_2064_),
    .Y(_2066_));
 sg13g2_nor2_2 _5122_ (.A(net1903),
    .B(_1712_),
    .Y(_2067_));
 sg13g2_or2_1 _5123_ (.X(_2068_),
    .B(_1712_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ));
 sg13g2_nor2_1 _5124_ (.A(net1896),
    .B(net1156),
    .Y(_2069_));
 sg13g2_nor2_1 _5125_ (.A(net1161),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_o21ai_1 _5126_ (.B1(_2070_),
    .Y(_2071_),
    .A1(net1229),
    .A2(_2060_));
 sg13g2_a21oi_1 _5127_ (.A1(_0671_),
    .A2(_2066_),
    .Y(_2072_),
    .B1(net1203));
 sg13g2_a221oi_1 _5128_ (.B2(_2072_),
    .C1(net1249),
    .B1(_2071_),
    .A1(net1203),
    .Y(_0097_),
    .A2(_2069_));
 sg13g2_o21ai_1 _5129_ (.B1(net1204),
    .Y(_2073_),
    .A1(net1882),
    .A2(net1157));
 sg13g2_o21ai_1 _5130_ (.B1(_2060_),
    .Y(_2074_),
    .A1(net1882),
    .A2(net1156));
 sg13g2_a21oi_1 _5131_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .A2(_2061_),
    .Y(_2075_),
    .B1(net1161));
 sg13g2_nor2_1 _5132_ (.A(net1896),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2076_));
 sg13g2_nor2_1 _5133_ (.A(_2057_),
    .B(_2076_),
    .Y(_2077_));
 sg13g2_a22oi_1 _5134_ (.Y(_2078_),
    .B1(_2077_),
    .B2(net1161),
    .A2(_2075_),
    .A1(_2074_));
 sg13g2_nand2_1 _5135_ (.Y(_2079_),
    .A(net1230),
    .B(_2078_));
 sg13g2_a21oi_1 _5136_ (.A1(_2073_),
    .A2(_2079_),
    .Y(_0098_),
    .B1(net1248));
 sg13g2_nand2b_1 _5137_ (.Y(_2080_),
    .B(_2067_),
    .A_N(net1906));
 sg13g2_nand2_1 _5138_ (.Y(_2081_),
    .A(net1204),
    .B(_2080_));
 sg13g2_mux2_1 _5139_ (.A0(net1873),
    .A1(_2080_),
    .S(_2060_),
    .X(_2082_));
 sg13g2_nor3_1 _5140_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .C(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2083_));
 sg13g2_xnor2_1 _5141_ (.Y(_2084_),
    .A(net1906),
    .B(_2076_));
 sg13g2_a21oi_1 _5142_ (.A1(net1161),
    .A2(_2084_),
    .Y(_2085_),
    .B1(net1204));
 sg13g2_o21ai_1 _5143_ (.B1(_2085_),
    .Y(_2086_),
    .A1(net1161),
    .A2(_2082_));
 sg13g2_a21oi_1 _5144_ (.A1(_2081_),
    .A2(_2086_),
    .Y(_0099_),
    .B1(net1249));
 sg13g2_o21ai_1 _5145_ (.B1(net1203),
    .Y(_2087_),
    .A1(net1886),
    .A2(net1157));
 sg13g2_o21ai_1 _5146_ (.B1(_2060_),
    .Y(_2088_),
    .A1(net1886),
    .A2(net1156));
 sg13g2_a21oi_1 _5147_ (.A1(net1827),
    .A2(_2061_),
    .Y(_2089_),
    .B1(_2066_));
 sg13g2_nor2b_1 _5148_ (.A(net1886),
    .B_N(_2083_),
    .Y(_2090_));
 sg13g2_xnor2_1 _5149_ (.Y(_2091_),
    .A(net1886),
    .B(_2083_));
 sg13g2_a22oi_1 _5150_ (.Y(_2092_),
    .B1(_2091_),
    .B2(net1161),
    .A2(_2089_),
    .A1(_2088_));
 sg13g2_nand2_1 _5151_ (.Y(_2093_),
    .A(net1230),
    .B(_2092_));
 sg13g2_a21oi_1 _5152_ (.A1(_2087_),
    .A2(_2093_),
    .Y(_0100_),
    .B1(net1248));
 sg13g2_nor2_1 _5153_ (.A(net1889),
    .B(net1156),
    .Y(_2094_));
 sg13g2_nor2_1 _5154_ (.A(net1161),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_o21ai_1 _5155_ (.B1(_2095_),
    .Y(_2096_),
    .A1(net1851),
    .A2(_2060_));
 sg13g2_xor2_1 _5156_ (.B(_2090_),
    .A(net1889),
    .X(_2097_));
 sg13g2_a21oi_1 _5157_ (.A1(net1161),
    .A2(_2097_),
    .Y(_2098_),
    .B1(net1203));
 sg13g2_a221oi_1 _5158_ (.B2(_2098_),
    .C1(net1248),
    .B1(_2096_),
    .A1(net1203),
    .Y(_0101_),
    .A2(_2094_));
 sg13g2_nor2_1 _5159_ (.A(net1904),
    .B(net1156),
    .Y(_2099_));
 sg13g2_o21ai_1 _5160_ (.B1(net1204),
    .Y(_2100_),
    .A1(net1904),
    .A2(net1156));
 sg13g2_nand2_1 _5161_ (.Y(_2101_),
    .A(net1709),
    .B(_0892_));
 sg13g2_and3_2 _5162_ (.X(_2102_),
    .A(net1230),
    .B(_1723_),
    .C(_2101_));
 sg13g2_a21oi_1 _5163_ (.A1(_2056_),
    .A2(_2058_),
    .Y(_2103_),
    .B1(_2064_));
 sg13g2_nor2_1 _5164_ (.A(_0894_),
    .B(_2103_),
    .Y(_2104_));
 sg13g2_o21ai_1 _5165_ (.B1(_0722_),
    .Y(_2105_),
    .A1(_0894_),
    .A2(_2103_));
 sg13g2_nor3_1 _5166_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .C(net1918),
    .Y(_2106_));
 sg13g2_and2_1 _5167_ (.A(_0643_),
    .B(_2106_),
    .X(_2107_));
 sg13g2_and2_1 _5168_ (.A(_0642_),
    .B(_2107_),
    .X(_2108_));
 sg13g2_a21oi_1 _5169_ (.A1(net1193),
    .A2(_2108_),
    .Y(_2109_),
    .B1(_0891_));
 sg13g2_o21ai_1 _5170_ (.B1(_2109_),
    .Y(_2110_),
    .A1(_2099_),
    .A2(_2105_));
 sg13g2_nand2_1 _5171_ (.Y(_2111_),
    .A(_2102_),
    .B(_2110_));
 sg13g2_a22oi_1 _5172_ (.Y(_2112_),
    .B1(_2108_),
    .B2(net1193),
    .A2(_2064_),
    .A1(net1188));
 sg13g2_o21ai_1 _5173_ (.B1(_2112_),
    .Y(_2113_),
    .A1(_2059_),
    .A2(_2065_));
 sg13g2_nor2_1 _5174_ (.A(net1204),
    .B(_2102_),
    .Y(_2114_));
 sg13g2_nor2_1 _5175_ (.A(net1156),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_a22oi_1 _5176_ (.Y(_2116_),
    .B1(_2115_),
    .B2(net1709),
    .A2(_2113_),
    .A1(_2102_));
 sg13g2_and2_1 _5177_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B(_2067_),
    .X(_2117_));
 sg13g2_nand2_1 _5178_ (.Y(_2118_),
    .A(net1878),
    .B(_2067_));
 sg13g2_and2_1 _5179_ (.A(_2102_),
    .B(_2112_),
    .X(_2119_));
 sg13g2_o21ai_1 _5180_ (.B1(_2119_),
    .Y(_2120_),
    .A1(_2105_),
    .A2(_2117_));
 sg13g2_o21ai_1 _5181_ (.B1(_2120_),
    .Y(_2121_),
    .A1(net1230),
    .A2(_2118_));
 sg13g2_nand4_1 _5182_ (.B(_2111_),
    .C(_2116_),
    .A(_2100_),
    .Y(_2122_),
    .D(_2121_));
 sg13g2_a21oi_1 _5183_ (.A1(_0893_),
    .A2(_2122_),
    .Y(_2123_),
    .B1(net1188));
 sg13g2_nor2_1 _5184_ (.A(_2064_),
    .B(_2123_),
    .Y(_2124_));
 sg13g2_nor3_2 _5185_ (.A(net1203),
    .B(_2064_),
    .C(_2123_),
    .Y(_2125_));
 sg13g2_nor3_1 _5186_ (.A(net1229),
    .B(net1157),
    .C(_2125_),
    .Y(_2126_));
 sg13g2_a21oi_1 _5187_ (.A1(net1229),
    .A2(_2125_),
    .Y(_2127_),
    .B1(net1249));
 sg13g2_nor2b_1 _5188_ (.A(_2126_),
    .B_N(_2127_),
    .Y(_0102_));
 sg13g2_xor2_1 _5189_ (.B(net1229),
    .A(net1891),
    .X(_2128_));
 sg13g2_nand2b_1 _5190_ (.Y(_2129_),
    .B(_2067_),
    .A_N(net1891));
 sg13g2_o21ai_1 _5191_ (.B1(net1263),
    .Y(_2130_),
    .A1(_2125_),
    .A2(_2129_));
 sg13g2_a21oi_1 _5192_ (.A1(_2125_),
    .A2(net1892),
    .Y(_0103_),
    .B1(_2130_));
 sg13g2_o21ai_1 _5193_ (.B1(net1873),
    .Y(_2131_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ));
 sg13g2_nor2b_1 _5194_ (.A(_2062_),
    .B_N(_2131_),
    .Y(_2132_));
 sg13g2_nand2_1 _5195_ (.Y(_2133_),
    .A(net1873),
    .B(_2067_));
 sg13g2_mux2_1 _5196_ (.A0(net1874),
    .A1(_2132_),
    .S(_2125_),
    .X(_2134_));
 sg13g2_nor2_1 _5197_ (.A(net1249),
    .B(net1875),
    .Y(_0104_));
 sg13g2_xnor2_1 _5198_ (.Y(_2135_),
    .A(net1827),
    .B(_2062_));
 sg13g2_nor2_1 _5199_ (.A(_0670_),
    .B(net1157),
    .Y(_2136_));
 sg13g2_o21ai_1 _5200_ (.B1(net1263),
    .Y(_2137_),
    .A1(_2125_),
    .A2(_2136_));
 sg13g2_a21oi_1 _5201_ (.A1(_2125_),
    .A2(net1828),
    .Y(_0105_),
    .B1(_2137_));
 sg13g2_nor2_1 _5202_ (.A(net1851),
    .B(net1156),
    .Y(_2138_));
 sg13g2_or2_1 _5203_ (.X(_2139_),
    .B(_2138_),
    .A(_2124_));
 sg13g2_a21oi_1 _5204_ (.A1(net1851),
    .A2(_2063_),
    .Y(_2140_),
    .B1(net1203));
 sg13g2_a221oi_1 _5205_ (.B2(_2140_),
    .C1(net1248),
    .B1(_2139_),
    .A1(net1203),
    .Y(_0106_),
    .A2(_2138_));
 sg13g2_nor2_1 _5206_ (.A(net1190),
    .B(_2108_),
    .Y(_2141_));
 sg13g2_a21oi_2 _5207_ (.B1(_2141_),
    .Y(_2142_),
    .A2(_2064_),
    .A1(net1188));
 sg13g2_inv_1 _5208_ (.Y(_2143_),
    .A(net1155));
 sg13g2_o21ai_1 _5209_ (.B1(net1230),
    .Y(_2144_),
    .A1(_2104_),
    .A2(_2143_));
 sg13g2_nand2_1 _5210_ (.Y(_2145_),
    .A(net1229),
    .B(_0671_));
 sg13g2_nand2b_1 _5211_ (.Y(_2146_),
    .B(net1917),
    .A_N(net1229));
 sg13g2_a21o_1 _5212_ (.A2(_2146_),
    .A1(_2145_),
    .B1(_2143_),
    .X(_2147_));
 sg13g2_o21ai_1 _5213_ (.B1(_2147_),
    .Y(_2148_),
    .A1(net1688),
    .A2(net1155));
 sg13g2_o21ai_1 _5214_ (.B1(net1262),
    .Y(_2149_),
    .A1(net842),
    .A2(_2148_));
 sg13g2_a21oi_1 _5215_ (.A1(_0645_),
    .A2(net842),
    .Y(_0107_),
    .B1(_2149_));
 sg13g2_nand2b_1 _5216_ (.Y(_2150_),
    .B(_2144_),
    .A_N(net1855));
 sg13g2_xnor2_1 _5217_ (.Y(_2151_),
    .A(net1855),
    .B(net1688));
 sg13g2_nor2b_1 _5218_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2152_));
 sg13g2_xnor2_1 _5219_ (.Y(_2153_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ));
 sg13g2_xnor2_1 _5220_ (.Y(_2154_),
    .A(_2145_),
    .B(_2153_));
 sg13g2_nand2_1 _5221_ (.Y(_2155_),
    .A(net1155),
    .B(_2154_));
 sg13g2_o21ai_1 _5222_ (.B1(_2155_),
    .Y(_2156_),
    .A1(net1155),
    .A2(_2151_));
 sg13g2_nand2b_1 _5223_ (.Y(_2157_),
    .B(_2156_),
    .A_N(_2144_));
 sg13g2_and3_1 _5224_ (.X(_0108_),
    .A(net1262),
    .B(_2150_),
    .C(_2157_));
 sg13g2_o21ai_1 _5225_ (.B1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .Y(_2158_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ));
 sg13g2_nor2b_1 _5226_ (.A(net1919),
    .B_N(_2158_),
    .Y(_2159_));
 sg13g2_nand2b_1 _5227_ (.Y(_2160_),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ));
 sg13g2_xnor2_1 _5228_ (.Y(_2161_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ));
 sg13g2_a21oi_1 _5229_ (.A1(_2145_),
    .A2(_2153_),
    .Y(_2162_),
    .B1(_2152_));
 sg13g2_nand2b_1 _5230_ (.Y(_2163_),
    .B(_2161_),
    .A_N(_2162_));
 sg13g2_nand2b_1 _5231_ (.Y(_2164_),
    .B(_2162_),
    .A_N(_2161_));
 sg13g2_nand3_1 _5232_ (.B(_2163_),
    .C(_2164_),
    .A(net1155),
    .Y(_2165_));
 sg13g2_o21ai_1 _5233_ (.B1(_2165_),
    .Y(_2166_),
    .A1(_2142_),
    .A2(_2159_));
 sg13g2_o21ai_1 _5234_ (.B1(net1262),
    .Y(_2167_),
    .A1(net842),
    .A2(_2166_));
 sg13g2_a21oi_1 _5235_ (.A1(_0644_),
    .A2(net842),
    .Y(_0109_),
    .B1(_2167_));
 sg13g2_xnor2_1 _5236_ (.Y(_2168_),
    .A(net1729),
    .B(_2106_));
 sg13g2_xor2_1 _5237_ (.B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .X(_2169_));
 sg13g2_nand3_1 _5238_ (.B(_2163_),
    .C(_2169_),
    .A(_2160_),
    .Y(_2170_));
 sg13g2_a21oi_1 _5239_ (.A1(_2160_),
    .A2(_2163_),
    .Y(_2171_),
    .B1(_2169_));
 sg13g2_nand3b_1 _5240_ (.B(net1155),
    .C(_2170_),
    .Y(_2172_),
    .A_N(_2171_));
 sg13g2_o21ai_1 _5241_ (.B1(_2172_),
    .Y(_2173_),
    .A1(_2142_),
    .A2(_2168_));
 sg13g2_o21ai_1 _5242_ (.B1(net1262),
    .Y(_2174_),
    .A1(net842),
    .A2(_2173_));
 sg13g2_a21oi_1 _5243_ (.A1(_0643_),
    .A2(net842),
    .Y(_0110_),
    .B1(_2174_));
 sg13g2_a21oi_1 _5244_ (.A1(_0670_),
    .A2(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .Y(_2175_),
    .B1(_2171_));
 sg13g2_xor2_1 _5245_ (.B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .X(_2176_));
 sg13g2_xnor2_1 _5246_ (.Y(_2177_),
    .A(_2175_),
    .B(_2176_));
 sg13g2_nor2_1 _5247_ (.A(_0642_),
    .B(_2107_),
    .Y(_2178_));
 sg13g2_nor3_1 _5248_ (.A(_2108_),
    .B(net1155),
    .C(_2178_),
    .Y(_2179_));
 sg13g2_a21oi_1 _5249_ (.A1(net1155),
    .A2(_2177_),
    .Y(_2180_),
    .B1(_2179_));
 sg13g2_o21ai_1 _5250_ (.B1(net1262),
    .Y(_2181_),
    .A1(net842),
    .A2(_2180_));
 sg13g2_a21oi_1 _5251_ (.A1(_0642_),
    .A2(net842),
    .Y(_0111_),
    .B1(_2181_));
 sg13g2_a21oi_1 _5252_ (.A1(_2100_),
    .A2(_2111_),
    .Y(_0112_),
    .B1(net1248));
 sg13g2_and2_1 _5253_ (.A(net1263),
    .B(_2121_),
    .X(_0113_));
 sg13g2_nor2_1 _5254_ (.A(net1248),
    .B(_2116_),
    .Y(_0114_));
 sg13g2_nor3_2 _5255_ (.A(net1204),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .C(_0722_),
    .Y(_2182_));
 sg13g2_nand2_2 _5256_ (.Y(_2183_),
    .A(net1230),
    .B(_0891_));
 sg13g2_o21ai_1 _5257_ (.B1(net1267),
    .Y(_2184_),
    .A1(net1719),
    .A2(net1165));
 sg13g2_a21oi_1 _5258_ (.A1(_1003_),
    .A2(net1165),
    .Y(_0115_),
    .B1(_2184_));
 sg13g2_o21ai_1 _5259_ (.B1(net1268),
    .Y(_2185_),
    .A1(net1742),
    .A2(net1164));
 sg13g2_a21oi_1 _5260_ (.A1(_1423_),
    .A2(net1164),
    .Y(_0116_),
    .B1(_2185_));
 sg13g2_o21ai_1 _5261_ (.B1(net1268),
    .Y(_2186_),
    .A1(net1689),
    .A2(net1164));
 sg13g2_a21oi_1 _5262_ (.A1(_0938_),
    .A2(net1163),
    .Y(_0117_),
    .B1(_2186_));
 sg13g2_o21ai_1 _5263_ (.B1(net1271),
    .Y(_2187_),
    .A1(net1699),
    .A2(net1164));
 sg13g2_a21oi_1 _5264_ (.A1(_1335_),
    .A2(net1163),
    .Y(_0118_),
    .B1(_2187_));
 sg13g2_o21ai_1 _5265_ (.B1(net1261),
    .Y(_2188_),
    .A1(_1123_),
    .A2(_2183_));
 sg13g2_a21oi_1 _5266_ (.A1(_0641_),
    .A2(net1160),
    .Y(_0119_),
    .B1(_2188_));
 sg13g2_o21ai_1 _5267_ (.B1(net1264),
    .Y(_2189_),
    .A1(_1360_),
    .A2(net1160));
 sg13g2_a21oi_1 _5268_ (.A1(_0640_),
    .A2(net1160),
    .Y(_0120_),
    .B1(_2189_));
 sg13g2_o21ai_1 _5269_ (.B1(net1261),
    .Y(_2190_),
    .A1(_0966_),
    .A2(net1159));
 sg13g2_a21oi_1 _5270_ (.A1(_0639_),
    .A2(net1159),
    .Y(_0121_),
    .B1(_2190_));
 sg13g2_o21ai_1 _5271_ (.B1(net1261),
    .Y(_2191_),
    .A1(_1389_),
    .A2(net1159));
 sg13g2_a21oi_1 _5272_ (.A1(_0638_),
    .A2(net1159),
    .Y(_0122_),
    .B1(_2191_));
 sg13g2_o21ai_1 _5273_ (.B1(net1267),
    .Y(_2192_),
    .A1(net1694),
    .A2(net1165));
 sg13g2_a21oi_1 _5274_ (.A1(_1048_),
    .A2(net1165),
    .Y(_0123_),
    .B1(_2192_));
 sg13g2_o21ai_1 _5275_ (.B1(net1267),
    .Y(_2193_),
    .A1(net1681),
    .A2(net1165));
 sg13g2_a21oi_1 _5276_ (.A1(_1466_),
    .A2(net1165),
    .Y(_0124_),
    .B1(_2193_));
 sg13g2_o21ai_1 _5277_ (.B1(net1261),
    .Y(_2194_),
    .A1(_1031_),
    .A2(net1160));
 sg13g2_a21oi_1 _5278_ (.A1(_0637_),
    .A2(net1159),
    .Y(_0125_),
    .B1(_2194_));
 sg13g2_o21ai_1 _5279_ (.B1(net1261),
    .Y(_2195_),
    .A1(_1527_),
    .A2(net1159));
 sg13g2_a21oi_1 _5280_ (.A1(_0636_),
    .A2(net1159),
    .Y(_0126_),
    .B1(_2195_));
 sg13g2_o21ai_1 _5281_ (.B1(net1261),
    .Y(_2196_),
    .A1(_0916_),
    .A2(net1160));
 sg13g2_a21oi_1 _5282_ (.A1(_0635_),
    .A2(net1160),
    .Y(_0127_),
    .B1(_2196_));
 sg13g2_o21ai_1 _5283_ (.B1(net1267),
    .Y(_2197_),
    .A1(net1705),
    .A2(net1165));
 sg13g2_a21oi_1 _5284_ (.A1(_1406_),
    .A2(net1165),
    .Y(_0128_),
    .B1(_2197_));
 sg13g2_o21ai_1 _5285_ (.B1(net1271),
    .Y(_2198_),
    .A1(net1740),
    .A2(net1163));
 sg13g2_a21oi_1 _5286_ (.A1(_0985_),
    .A2(net1163),
    .Y(_0129_),
    .B1(_2198_));
 sg13g2_o21ai_1 _5287_ (.B1(net1268),
    .Y(_2199_),
    .A1(net1675),
    .A2(net1164));
 sg13g2_a21oi_1 _5288_ (.A1(_1499_),
    .A2(net1164),
    .Y(_0130_),
    .B1(_2199_));
 sg13g2_o21ai_1 _5289_ (.B1(net1268),
    .Y(_2200_),
    .A1(net1716),
    .A2(net1163));
 sg13g2_a21oi_1 _5290_ (.A1(_1095_),
    .A2(net1163),
    .Y(_0131_),
    .B1(_2200_));
 sg13g2_o21ai_1 _5291_ (.B1(net1268),
    .Y(_2201_),
    .A1(net1697),
    .A2(net1163));
 sg13g2_a21oi_1 _5292_ (.A1(_1482_),
    .A2(net1163),
    .Y(_0132_),
    .B1(_2201_));
 sg13g2_o21ai_1 _5293_ (.B1(net1261),
    .Y(_2202_),
    .A1(_1076_),
    .A2(net1160));
 sg13g2_a21oi_1 _5294_ (.A1(_0634_),
    .A2(net1159),
    .Y(_0133_),
    .B1(_2202_));
 sg13g2_o21ai_1 _5295_ (.B1(net1261),
    .Y(_2203_),
    .A1(_1449_),
    .A2(_2183_));
 sg13g2_a21oi_1 _5296_ (.A1(_0633_),
    .A2(_2183_),
    .Y(_0134_),
    .B1(_2203_));
 sg13g2_nand4_1 _5297_ (.B(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .C(_0714_),
    .A(_0707_),
    .Y(_2204_),
    .D(\vga_tetris._tetrisLogic_io_score_3[3] ));
 sg13g2_nand3_1 _5298_ (.B(_0893_),
    .C(_2204_),
    .A(net1230),
    .Y(_2205_));
 sg13g2_nor4_2 _5299_ (.A(_2053_),
    .B(_2054_),
    .C(_2055_),
    .Y(_2206_),
    .D(_2205_));
 sg13g2_and2_1 _5300_ (.A(net1661),
    .B(_2206_),
    .X(_2207_));
 sg13g2_a21oi_1 _5301_ (.A1(net1661),
    .A2(_2206_),
    .Y(_2208_),
    .B1(net1898));
 sg13g2_a21oi_1 _5302_ (.A1(_0713_),
    .A2(_2208_),
    .Y(_2209_),
    .B1(_0712_));
 sg13g2_a21o_1 _5303_ (.A2(_2208_),
    .A1(_0713_),
    .B1(_0712_),
    .X(_2210_));
 sg13g2_a21oi_1 _5304_ (.A1(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .A2(_2209_),
    .Y(_2211_),
    .B1(net1830));
 sg13g2_a21oi_2 _5305_ (.B1(_0710_),
    .Y(_2212_),
    .A2(_2211_),
    .A1(_0711_));
 sg13g2_a21oi_1 _5306_ (.A1(net1753),
    .A2(_2212_),
    .Y(_2213_),
    .B1(net1839));
 sg13g2_a21oi_2 _5307_ (.B1(_0708_),
    .Y(_2214_),
    .A2(_2213_),
    .A1(_0709_));
 sg13g2_nor2_1 _5308_ (.A(net1720),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_nand2_2 _5309_ (.Y(_2216_),
    .A(net1265),
    .B(_2041_));
 sg13g2_and2_1 _5310_ (.A(net1720),
    .B(_2214_),
    .X(_2217_));
 sg13g2_nor3_1 _5311_ (.A(net1721),
    .B(net1153),
    .C(_2217_),
    .Y(_0135_));
 sg13g2_nand3_1 _5312_ (.B(net1720),
    .C(_2214_),
    .A(net1829),
    .Y(_2218_));
 sg13g2_nand2_1 _5313_ (.Y(_2219_),
    .A(_0714_),
    .B(_2218_));
 sg13g2_xnor2_1 _5314_ (.Y(_2220_),
    .A(net1829),
    .B(_2217_));
 sg13g2_inv_1 _5315_ (.Y(_2221_),
    .A(_2220_));
 sg13g2_nand3_1 _5316_ (.B(net1763),
    .C(_2220_),
    .A(net1737),
    .Y(_2222_));
 sg13g2_or2_1 _5317_ (.X(_2223_),
    .B(_2220_),
    .A(net1737));
 sg13g2_a21oi_1 _5318_ (.A1(net1764),
    .A2(_2223_),
    .Y(_0136_),
    .B1(net1153));
 sg13g2_nor2_1 _5319_ (.A(_0714_),
    .B(_2218_),
    .Y(_2224_));
 sg13g2_and2_1 _5320_ (.A(net1737),
    .B(_2224_),
    .X(_2225_));
 sg13g2_nand2_1 _5321_ (.Y(_2226_),
    .A(net1737),
    .B(_2224_));
 sg13g2_xnor2_1 _5322_ (.Y(_2227_),
    .A(_0714_),
    .B(_2218_));
 sg13g2_a21o_1 _5323_ (.A2(_2220_),
    .A1(net1737),
    .B1(_2227_),
    .X(_2228_));
 sg13g2_a21oi_1 _5324_ (.A1(net1738),
    .A2(_2228_),
    .Y(_0137_),
    .B1(net1153));
 sg13g2_o21ai_1 _5325_ (.B1(_2227_),
    .Y(_2229_),
    .A1(net1737),
    .A2(_2224_));
 sg13g2_nor4_1 _5326_ (.A(net1153),
    .B(_2221_),
    .C(_2225_),
    .D(_2229_),
    .Y(_0138_));
 sg13g2_and3_2 _5327_ (.X(_2230_),
    .A(net1228),
    .B(net1388),
    .C(net1692));
 sg13g2_a21oi_1 _5328_ (.A1(net1228),
    .A2(\vga_tetris._inputs_io_downButtonActive ),
    .Y(_2231_),
    .B1(net1388));
 sg13g2_nor3_1 _5329_ (.A(_1747_),
    .B(_2230_),
    .C(net1389),
    .Y(_0139_));
 sg13g2_nand2_1 _5330_ (.Y(_2232_),
    .A(net1714),
    .B(_2230_));
 sg13g2_xnor2_1 _5331_ (.Y(_2233_),
    .A(net1714),
    .B(_2230_));
 sg13g2_nor2_1 _5332_ (.A(_1747_),
    .B(net1715),
    .Y(_0140_));
 sg13g2_xor2_1 _5333_ (.B(_2232_),
    .A(net1732),
    .X(_2234_));
 sg13g2_nor2_1 _5334_ (.A(_1747_),
    .B(_2234_),
    .Y(_0141_));
 sg13g2_nor2_1 _5335_ (.A(_2045_),
    .B(_2046_),
    .Y(_0142_));
 sg13g2_xnor2_1 _5336_ (.Y(_2235_),
    .A(net1753),
    .B(_2212_));
 sg13g2_nor2_1 _5337_ (.A(net1153),
    .B(net1754),
    .Y(_0143_));
 sg13g2_and3_2 _5338_ (.X(_2236_),
    .A(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .B(net1753),
    .C(_2212_));
 sg13g2_or2_1 _5339_ (.X(_2237_),
    .B(_2236_),
    .A(_2213_));
 sg13g2_nand2_1 _5340_ (.Y(_2238_),
    .A(_2214_),
    .B(_2237_));
 sg13g2_nand2b_1 _5341_ (.Y(_2239_),
    .B(_0708_),
    .A_N(_2237_));
 sg13g2_a21oi_1 _5342_ (.A1(net1840),
    .A2(_2239_),
    .Y(_0144_),
    .B1(net1153));
 sg13g2_a21oi_1 _5343_ (.A1(net1784),
    .A2(_2236_),
    .Y(_2240_),
    .B1(_2238_));
 sg13g2_nand3_1 _5344_ (.B(net1784),
    .C(_2236_),
    .A(_0708_),
    .Y(_2241_));
 sg13g2_o21ai_1 _5345_ (.B1(_2241_),
    .Y(_2242_),
    .A1(net1784),
    .A2(_2236_));
 sg13g2_nor3_1 _5346_ (.A(net1153),
    .B(net1785),
    .C(_2242_),
    .Y(_0145_));
 sg13g2_a21oi_1 _5347_ (.A1(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .A2(_2236_),
    .Y(_2243_),
    .B1(net1453));
 sg13g2_nor3_1 _5348_ (.A(_2214_),
    .B(net1153),
    .C(net1454),
    .Y(_0146_));
 sg13g2_xnor2_1 _5349_ (.Y(_2244_),
    .A(net1733),
    .B(_2209_));
 sg13g2_nor2_1 _5350_ (.A(net1154),
    .B(net1734),
    .Y(_0147_));
 sg13g2_and3_2 _5351_ (.X(_2245_),
    .A(net1733),
    .B(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .C(_2209_));
 sg13g2_or2_1 _5352_ (.X(_2246_),
    .B(_2245_),
    .A(net1831));
 sg13g2_nand2_1 _5353_ (.Y(_2247_),
    .A(_2212_),
    .B(_2246_));
 sg13g2_nand2b_1 _5354_ (.Y(_2248_),
    .B(_0710_),
    .A_N(_2246_));
 sg13g2_a21oi_1 _5355_ (.A1(net1832),
    .A2(_2248_),
    .Y(_0148_),
    .B1(net1154));
 sg13g2_a21oi_1 _5356_ (.A1(net1773),
    .A2(_2245_),
    .Y(_2249_),
    .B1(_2247_));
 sg13g2_nand3_1 _5357_ (.B(net1773),
    .C(_2245_),
    .A(_0710_),
    .Y(_2250_));
 sg13g2_o21ai_1 _5358_ (.B1(_2250_),
    .Y(_2251_),
    .A1(net1773),
    .A2(_2245_));
 sg13g2_nor3_1 _5359_ (.A(net1154),
    .B(net1774),
    .C(_2251_),
    .Y(_0149_));
 sg13g2_a21oi_1 _5360_ (.A1(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .A2(_2245_),
    .Y(_2252_),
    .B1(net1404));
 sg13g2_nor3_1 _5361_ (.A(_2212_),
    .B(net1154),
    .C(net1405),
    .Y(_0150_));
 sg13g2_nor2_1 _5362_ (.A(net1661),
    .B(_2206_),
    .Y(_2253_));
 sg13g2_nor3_1 _5363_ (.A(_2207_),
    .B(net1154),
    .C(net1662),
    .Y(_0151_));
 sg13g2_xor2_1 _5364_ (.B(_2207_),
    .A(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .X(_2254_));
 sg13g2_nor2_1 _5365_ (.A(_2210_),
    .B(_2254_),
    .Y(_2255_));
 sg13g2_a21oi_1 _5366_ (.A1(_0712_),
    .A2(_2254_),
    .Y(_2256_),
    .B1(_2255_));
 sg13g2_nor2_1 _5367_ (.A(net1154),
    .B(net1859),
    .Y(_0152_));
 sg13g2_nand3_1 _5368_ (.B(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .C(_2207_),
    .A(net1791),
    .Y(_2257_));
 sg13g2_a21oi_1 _5369_ (.A1(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .A2(_2207_),
    .Y(_2258_),
    .B1(net1791));
 sg13g2_nor2_1 _5370_ (.A(net1154),
    .B(_2258_),
    .Y(_2259_));
 sg13g2_o21ai_1 _5371_ (.B1(_2259_),
    .Y(_2260_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .A2(net1792));
 sg13g2_a21oi_1 _5372_ (.A1(_2255_),
    .A2(net1792),
    .Y(_0153_),
    .B1(_2260_));
 sg13g2_a21oi_1 _5373_ (.A1(_0712_),
    .A2(net1792),
    .Y(_2261_),
    .B1(net1154));
 sg13g2_and2_1 _5374_ (.A(_2210_),
    .B(_2261_),
    .X(_0154_));
 sg13g2_a21oi_1 _5375_ (.A1(_1543_),
    .A2(_2040_),
    .Y(_0155_),
    .B1(net1252));
 sg13g2_nand2_1 _5376_ (.Y(_2262_),
    .A(_0816_),
    .B(_0830_));
 sg13g2_o21ai_1 _5377_ (.B1(net1179),
    .Y(_2263_),
    .A1(_0719_),
    .A2(net1188));
 sg13g2_o21ai_1 _5378_ (.B1(_2263_),
    .Y(_2264_),
    .A1(net1175),
    .A2(_1936_));
 sg13g2_a21o_2 _5379_ (.A2(_2264_),
    .A1(_0784_),
    .B1(net1168),
    .X(_2265_));
 sg13g2_nor3_1 _5380_ (.A(_0787_),
    .B(_0793_),
    .C(_0799_),
    .Y(_2266_));
 sg13g2_nand2_2 _5381_ (.Y(_2267_),
    .A(_2265_),
    .B(_2266_));
 sg13g2_nor2_1 _5382_ (.A(_2262_),
    .B(_2267_),
    .Y(_2268_));
 sg13g2_nor2_1 _5383_ (.A(net1523),
    .B(net981),
    .Y(_2269_));
 sg13g2_nand2_1 _5384_ (.Y(_2270_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .B(net1191));
 sg13g2_a21oi_1 _5385_ (.A1(net1178),
    .A2(_2270_),
    .Y(_2271_),
    .B1(net1170));
 sg13g2_o21ai_1 _5386_ (.B1(_2271_),
    .Y(_2272_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ),
    .A2(net1178));
 sg13g2_a21oi_1 _5387_ (.A1(net981),
    .A2(net1151),
    .Y(_0156_),
    .B1(_2269_));
 sg13g2_nor2_1 _5388_ (.A(net1576),
    .B(net983),
    .Y(_2273_));
 sg13g2_nand2_1 _5389_ (.Y(_2274_),
    .A(net1915),
    .B(net1191));
 sg13g2_a21oi_1 _5390_ (.A1(net1176),
    .A2(_2274_),
    .Y(_2275_),
    .B1(net1170));
 sg13g2_o21ai_1 _5391_ (.B1(_2275_),
    .Y(_2276_),
    .A1(net1509),
    .A2(net1176));
 sg13g2_a21oi_1 _5392_ (.A1(net983),
    .A2(net1148),
    .Y(_0157_),
    .B1(_2273_));
 sg13g2_nor2_1 _5393_ (.A(net1568),
    .B(net982),
    .Y(_2277_));
 sg13g2_nand2_1 _5394_ (.Y(_2278_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .B(net1191));
 sg13g2_a21oi_1 _5395_ (.A1(net1177),
    .A2(_2278_),
    .Y(_2279_),
    .B1(net1171));
 sg13g2_o21ai_1 _5396_ (.B1(_2279_),
    .Y(_2280_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .A2(net1177));
 sg13g2_a21oi_1 _5397_ (.A1(net982),
    .A2(net1145),
    .Y(_0158_),
    .B1(_2277_));
 sg13g2_nor2_1 _5398_ (.A(net1562),
    .B(net982),
    .Y(_2281_));
 sg13g2_nand2_1 _5399_ (.Y(_2282_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ),
    .B(net1191));
 sg13g2_a21oi_1 _5400_ (.A1(net1177),
    .A2(_2282_),
    .Y(_2283_),
    .B1(net1171));
 sg13g2_o21ai_1 _5401_ (.B1(_2283_),
    .Y(_2284_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ),
    .A2(net1177));
 sg13g2_a21oi_1 _5402_ (.A1(net982),
    .A2(net1142),
    .Y(_0159_),
    .B1(_2281_));
 sg13g2_nor2_1 _5403_ (.A(net1588),
    .B(net984),
    .Y(_2285_));
 sg13g2_nand2_1 _5404_ (.Y(_2286_),
    .A(net818),
    .B(net1190));
 sg13g2_a21oi_1 _5405_ (.A1(net1175),
    .A2(_2286_),
    .Y(_2287_),
    .B1(net1169));
 sg13g2_o21ai_1 _5406_ (.B1(_2287_),
    .Y(_2288_),
    .A1(net1391),
    .A2(net1175));
 sg13g2_a21oi_1 _5407_ (.A1(net984),
    .A2(net1138),
    .Y(_0160_),
    .B1(_2285_));
 sg13g2_nor2_1 _5408_ (.A(net1518),
    .B(net980),
    .Y(_2289_));
 sg13g2_nand2_1 _5409_ (.Y(_2290_),
    .A(net821),
    .B(net1189));
 sg13g2_a21oi_1 _5410_ (.A1(net1173),
    .A2(_2290_),
    .Y(_2291_),
    .B1(net1168));
 sg13g2_o21ai_1 _5411_ (.B1(_2291_),
    .Y(_2292_),
    .A1(net1916),
    .A2(net1175));
 sg13g2_a21oi_1 _5412_ (.A1(net980),
    .A2(net1137),
    .Y(_0161_),
    .B1(_2289_));
 sg13g2_nor2_1 _5413_ (.A(net1578),
    .B(net978),
    .Y(_2293_));
 sg13g2_nand2_1 _5414_ (.Y(_2294_),
    .A(net1302),
    .B(net1189));
 sg13g2_a21oi_1 _5415_ (.A1(net1172),
    .A2(_2294_),
    .Y(_2295_),
    .B1(net1168));
 sg13g2_o21ai_1 _5416_ (.B1(_2295_),
    .Y(_2296_),
    .A1(net1398),
    .A2(net1172));
 sg13g2_a21oi_1 _5417_ (.A1(net978),
    .A2(net1132),
    .Y(_0162_),
    .B1(_2293_));
 sg13g2_nor2_1 _5418_ (.A(net1543),
    .B(net978),
    .Y(_2297_));
 sg13g2_nand2_1 _5419_ (.Y(_2298_),
    .A(net756),
    .B(net1189));
 sg13g2_a21oi_1 _5420_ (.A1(net1172),
    .A2(_2298_),
    .Y(_2299_),
    .B1(net1168));
 sg13g2_o21ai_1 _5421_ (.B1(_2299_),
    .Y(_2300_),
    .A1(net1393),
    .A2(net1172));
 sg13g2_a21oi_1 _5422_ (.A1(net978),
    .A2(net1130),
    .Y(_0163_),
    .B1(_2297_));
 sg13g2_nor2_1 _5423_ (.A(net1615),
    .B(net981),
    .Y(_2301_));
 sg13g2_nand2_1 _5424_ (.Y(_2302_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .B(net1191));
 sg13g2_a21oi_1 _5425_ (.A1(net1178),
    .A2(_2302_),
    .Y(_2303_),
    .B1(net1170));
 sg13g2_o21ai_1 _5426_ (.B1(_2303_),
    .Y(_2304_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ),
    .A2(net1178));
 sg13g2_a21oi_1 _5427_ (.A1(net981),
    .A2(net1128),
    .Y(_0164_),
    .B1(_2301_));
 sg13g2_nor2_1 _5428_ (.A(net1536),
    .B(net981),
    .Y(_2305_));
 sg13g2_nand2_1 _5429_ (.Y(_2306_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .B(net1190));
 sg13g2_a21oi_1 _5430_ (.A1(net1178),
    .A2(_2306_),
    .Y(_2307_),
    .B1(net1169));
 sg13g2_o21ai_1 _5431_ (.B1(_2307_),
    .Y(_2308_),
    .A1(net1381),
    .A2(net1178));
 sg13g2_a21oi_1 _5432_ (.A1(net981),
    .A2(net1123),
    .Y(_0165_),
    .B1(_2305_));
 sg13g2_nor2_1 _5433_ (.A(net1486),
    .B(net979),
    .Y(_2309_));
 sg13g2_nand2_1 _5434_ (.Y(_2310_),
    .A(net1383),
    .B(net1189));
 sg13g2_a21oi_1 _5435_ (.A1(net1172),
    .A2(_2310_),
    .Y(_2311_),
    .B1(net1168));
 sg13g2_o21ai_1 _5436_ (.B1(_2311_),
    .Y(_2312_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .A2(net1172));
 sg13g2_a21oi_1 _5437_ (.A1(net979),
    .A2(net1121),
    .Y(_0166_),
    .B1(_2309_));
 sg13g2_nor2_1 _5438_ (.A(net1458),
    .B(net978),
    .Y(_2313_));
 sg13g2_nand2_1 _5439_ (.Y(_2314_),
    .A(net1369),
    .B(net1189));
 sg13g2_a21oi_1 _5440_ (.A1(net1172),
    .A2(_2314_),
    .Y(_2315_),
    .B1(net1168));
 sg13g2_o21ai_1 _5441_ (.B1(_2315_),
    .Y(_2316_),
    .A1(net1423),
    .A2(net1172));
 sg13g2_a21oi_1 _5442_ (.A1(net978),
    .A2(net1118),
    .Y(_0167_),
    .B1(_2313_));
 sg13g2_nor2_1 _5443_ (.A(net1428),
    .B(net980),
    .Y(_2317_));
 sg13g2_nand2_1 _5444_ (.Y(_2318_),
    .A(net1287),
    .B(net1192));
 sg13g2_a21oi_1 _5445_ (.A1(net1175),
    .A2(_2318_),
    .Y(_2319_),
    .B1(net1169));
 sg13g2_o21ai_1 _5446_ (.B1(_2319_),
    .Y(_2320_),
    .A1(net1430),
    .A2(net1175));
 sg13g2_a21oi_1 _5447_ (.A1(net980),
    .A2(net1115),
    .Y(_0168_),
    .B1(_2317_));
 sg13g2_nor2_1 _5448_ (.A(net1614),
    .B(net980),
    .Y(_2321_));
 sg13g2_nand2_1 _5449_ (.Y(_2322_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .B(net1190));
 sg13g2_a21oi_1 _5450_ (.A1(net1175),
    .A2(_2322_),
    .Y(_2323_),
    .B1(net1169));
 sg13g2_o21ai_1 _5451_ (.B1(_2323_),
    .Y(_2324_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ),
    .A2(net1175));
 sg13g2_a21oi_1 _5452_ (.A1(net980),
    .A2(net1113),
    .Y(_0169_),
    .B1(_2321_));
 sg13g2_nor2_1 _5453_ (.A(net1503),
    .B(net982),
    .Y(_2325_));
 sg13g2_nand2_1 _5454_ (.Y(_2326_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .B(net1191));
 sg13g2_a21oi_1 _5455_ (.A1(net1177),
    .A2(_2326_),
    .Y(_2327_),
    .B1(net1170));
 sg13g2_o21ai_1 _5456_ (.B1(_2327_),
    .Y(_2328_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .A2(net1177));
 sg13g2_a21oi_1 _5457_ (.A1(net982),
    .A2(net1110),
    .Y(_0170_),
    .B1(_2325_));
 sg13g2_nor2_1 _5458_ (.A(net1584),
    .B(net981),
    .Y(_2329_));
 sg13g2_nand2_1 _5459_ (.Y(_2330_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .B(net1191));
 sg13g2_a21oi_1 _5460_ (.A1(net1176),
    .A2(_2330_),
    .Y(_2331_),
    .B1(net1170));
 sg13g2_o21ai_1 _5461_ (.B1(_2331_),
    .Y(_2332_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .A2(net1176));
 sg13g2_a21oi_1 _5462_ (.A1(net981),
    .A2(net1107),
    .Y(_0171_),
    .B1(_2329_));
 sg13g2_nor2_1 _5463_ (.A(net1436),
    .B(net983),
    .Y(_2333_));
 sg13g2_nand2_1 _5464_ (.Y(_2334_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .B(net1191));
 sg13g2_a21oi_1 _5465_ (.A1(net1176),
    .A2(_2334_),
    .Y(_2335_),
    .B1(net1170));
 sg13g2_o21ai_1 _5466_ (.B1(_2335_),
    .Y(_2336_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .A2(net1176));
 sg13g2_a21oi_1 _5467_ (.A1(net983),
    .A2(net1102),
    .Y(_0172_),
    .B1(_2333_));
 sg13g2_nor2_1 _5468_ (.A(net1590),
    .B(net982),
    .Y(_2337_));
 sg13g2_nand2_1 _5469_ (.Y(_2338_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .B(net1192));
 sg13g2_a21oi_1 _5470_ (.A1(net1176),
    .A2(_2338_),
    .Y(_2339_),
    .B1(net1171));
 sg13g2_o21ai_1 _5471_ (.B1(_2339_),
    .Y(_2340_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .A2(net1176));
 sg13g2_a21oi_1 _5472_ (.A1(net982),
    .A2(net1100),
    .Y(_0173_),
    .B1(_2337_));
 sg13g2_nor2_1 _5473_ (.A(net1577),
    .B(net979),
    .Y(_2341_));
 sg13g2_nand2_1 _5474_ (.Y(_2342_),
    .A(net1384),
    .B(net1189));
 sg13g2_a21oi_1 _5475_ (.A1(net1174),
    .A2(_2342_),
    .Y(_2343_),
    .B1(net1168));
 sg13g2_o21ai_1 _5476_ (.B1(_2343_),
    .Y(_2344_),
    .A1(net1484),
    .A2(net1173));
 sg13g2_a21oi_1 _5477_ (.A1(net979),
    .A2(net1096),
    .Y(_0174_),
    .B1(_2341_));
 sg13g2_nor2_1 _5478_ (.A(net1589),
    .B(net978),
    .Y(_2345_));
 sg13g2_nand2_1 _5479_ (.Y(_2346_),
    .A(net1279),
    .B(net1189));
 sg13g2_a21oi_1 _5480_ (.A1(net1173),
    .A2(_2346_),
    .Y(_2347_),
    .B1(net1168));
 sg13g2_o21ai_1 _5481_ (.B1(_2347_),
    .Y(_2348_),
    .A1(net1414),
    .A2(net1173));
 sg13g2_a21oi_1 _5482_ (.A1(net978),
    .A2(net1093),
    .Y(_0175_),
    .B1(_2345_));
 sg13g2_a21oi_1 _5483_ (.A1(net1650),
    .A2(net1162),
    .Y(_2349_),
    .B1(net1255));
 sg13g2_a21oi_2 _5484_ (.B1(net3),
    .Y(_2350_),
    .A2(net1162),
    .A1(net1650));
 sg13g2_nand2_2 _5485_ (.Y(_2351_),
    .A(net1269),
    .B(_2350_));
 sg13g2_nand4_1 _5486_ (.B(\vga_tetris.msTimer.msTimerQ[3] ),
    .C(\vga_tetris.msTimer.msTimerQ[13] ),
    .A(_0693_),
    .Y(_2352_),
    .D(\vga_tetris.msTimer.msTimerQ[14] ));
 sg13g2_nor4_1 _5487_ (.A(\vga_tetris.msTimer.msTimerQ[1] ),
    .B(\vga_tetris.msTimer.msTimerQ[0] ),
    .C(_1807_),
    .D(_2352_),
    .Y(_2353_));
 sg13g2_nor4_1 _5488_ (.A(\vga_tetris.msTimer.msTimerQ[4] ),
    .B(_0694_),
    .C(\vga_tetris.msTimer.msTimerQ[6] ),
    .D(\vga_tetris.msTimer.msTimerQ[11] ),
    .Y(_2354_));
 sg13g2_nand3_1 _5489_ (.B(_2353_),
    .C(_2354_),
    .A(_1804_),
    .Y(_2355_));
 sg13g2_nor2_1 _5490_ (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .B(_2355_),
    .Y(_2356_));
 sg13g2_and3_2 _5491_ (.X(_2357_),
    .A(_1804_),
    .B(_2353_),
    .C(_2354_));
 sg13g2_nor2b_1 _5492_ (.A(net1650),
    .B_N(_2357_),
    .Y(_2358_));
 sg13g2_xnor2_1 _5493_ (.Y(_2359_),
    .A(net1725),
    .B(_2358_));
 sg13g2_nor2_1 _5494_ (.A(_2351_),
    .B(_2359_),
    .Y(_0176_));
 sg13g2_a21oi_1 _5495_ (.A1(\vga_tetris.inputs.buttonTimerQ_0[0] ),
    .A2(_2358_),
    .Y(_2360_),
    .B1(net1361));
 sg13g2_and3_2 _5496_ (.X(_2361_),
    .A(net1361),
    .B(net1725),
    .C(_2356_));
 sg13g2_nor3_1 _5497_ (.A(_2351_),
    .B(net1362),
    .C(_2361_),
    .Y(_0177_));
 sg13g2_nand2_1 _5498_ (.Y(_2362_),
    .A(net1847),
    .B(_2361_));
 sg13g2_o21ai_1 _5499_ (.B1(_2350_),
    .Y(_2363_),
    .A1(net1847),
    .A2(_2361_));
 sg13g2_nand2b_1 _5500_ (.Y(_2364_),
    .B(_2362_),
    .A_N(_2363_));
 sg13g2_nor2_1 _5501_ (.A(net1255),
    .B(_2364_),
    .Y(_0178_));
 sg13g2_and3_1 _5502_ (.X(_2365_),
    .A(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .B(\vga_tetris.inputs.buttonTimerQ_0[2] ),
    .C(_2361_));
 sg13g2_xnor2_1 _5503_ (.Y(_2366_),
    .A(net1845),
    .B(_2362_));
 sg13g2_and3_1 _5504_ (.X(_0179_),
    .A(net1269),
    .B(_2350_),
    .C(net1846));
 sg13g2_and2_1 _5505_ (.A(net1813),
    .B(_2365_),
    .X(_2367_));
 sg13g2_o21ai_1 _5506_ (.B1(_2350_),
    .Y(_2368_),
    .A1(net1813),
    .A2(_2365_));
 sg13g2_nor3_1 _5507_ (.A(net1255),
    .B(_2367_),
    .C(net1814),
    .Y(_0180_));
 sg13g2_and2_1 _5508_ (.A(net1822),
    .B(_2367_),
    .X(_2369_));
 sg13g2_o21ai_1 _5509_ (.B1(_2350_),
    .Y(_2370_),
    .A1(net1822),
    .A2(_2367_));
 sg13g2_nor3_1 _5510_ (.A(net1255),
    .B(_2369_),
    .C(_2370_),
    .Y(_0181_));
 sg13g2_nor2_1 _5511_ (.A(net1635),
    .B(_2369_),
    .Y(_2371_));
 sg13g2_and2_1 _5512_ (.A(net1635),
    .B(_2369_),
    .X(_2372_));
 sg13g2_nor3_1 _5513_ (.A(_2351_),
    .B(net1636),
    .C(_2372_),
    .Y(_0182_));
 sg13g2_xnor2_1 _5514_ (.Y(_2373_),
    .A(net1626),
    .B(_2372_));
 sg13g2_nor2_1 _5515_ (.A(_2351_),
    .B(net1627),
    .Y(_0183_));
 sg13g2_nand2_1 _5516_ (.Y(_2374_),
    .A(net1866),
    .B(net1162));
 sg13g2_nand2b_2 _5517_ (.Y(_2375_),
    .B(_2374_),
    .A_N(net1));
 sg13g2_or2_1 _5518_ (.X(_2376_),
    .B(_2375_),
    .A(net1255));
 sg13g2_nor2_1 _5519_ (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .B(_2355_),
    .Y(_2377_));
 sg13g2_nor2b_1 _5520_ (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .B_N(_2357_),
    .Y(_2378_));
 sg13g2_nor2_1 _5521_ (.A(net1663),
    .B(_2378_),
    .Y(_2379_));
 sg13g2_and2_1 _5522_ (.A(net1663),
    .B(_2378_),
    .X(_2380_));
 sg13g2_nor3_1 _5523_ (.A(_2376_),
    .B(net1664),
    .C(_2380_),
    .Y(_0184_));
 sg13g2_xnor2_1 _5524_ (.Y(_2381_),
    .A(net1726),
    .B(_2380_));
 sg13g2_nor2_1 _5525_ (.A(_2376_),
    .B(net1727),
    .Y(_0185_));
 sg13g2_a21oi_1 _5526_ (.A1(net1726),
    .A2(_2380_),
    .Y(_2382_),
    .B1(net1838));
 sg13g2_and4_1 _5527_ (.A(net1838),
    .B(net1726),
    .C(net1663),
    .D(_2377_),
    .X(_2383_));
 sg13g2_nor3_1 _5528_ (.A(_2375_),
    .B(_2382_),
    .C(_2383_),
    .Y(_2384_));
 sg13g2_and2_1 _5529_ (.A(net1269),
    .B(_2384_),
    .X(_0186_));
 sg13g2_nand4_1 _5530_ (.B(net1838),
    .C(net1726),
    .A(net1856),
    .Y(_2385_),
    .D(_2380_));
 sg13g2_o21ai_1 _5531_ (.B1(_2385_),
    .Y(_2386_),
    .A1(net1856),
    .A2(_2383_));
 sg13g2_nor2_1 _5532_ (.A(_2375_),
    .B(_2386_),
    .Y(_2387_));
 sg13g2_nor3_1 _5533_ (.A(net1255),
    .B(_2375_),
    .C(_2386_),
    .Y(_0187_));
 sg13g2_a21oi_1 _5534_ (.A1(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .A2(_2383_),
    .Y(_2388_),
    .B1(net1824));
 sg13g2_and3_1 _5535_ (.X(_2389_),
    .A(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .B(net1824),
    .C(_2383_));
 sg13g2_nor3_1 _5536_ (.A(_2375_),
    .B(net1825),
    .C(_2389_),
    .Y(_2390_));
 sg13g2_and2_1 _5537_ (.A(net1269),
    .B(net1826),
    .X(_0188_));
 sg13g2_nor2_1 _5538_ (.A(net1767),
    .B(_2389_),
    .Y(_2391_));
 sg13g2_and2_1 _5539_ (.A(net1767),
    .B(_2389_),
    .X(_2392_));
 sg13g2_nor4_1 _5540_ (.A(net1255),
    .B(_2375_),
    .C(net1768),
    .D(_2392_),
    .Y(_0189_));
 sg13g2_nand2_1 _5541_ (.Y(_2393_),
    .A(\vga_tetris.inputs.buttonTimerQ_1[6] ),
    .B(_2392_));
 sg13g2_xnor2_1 _5542_ (.Y(_2394_),
    .A(net1730),
    .B(_2392_));
 sg13g2_nor2_1 _5543_ (.A(_2376_),
    .B(net1731),
    .Y(_0190_));
 sg13g2_xor2_1 _5544_ (.B(_2393_),
    .A(net1673),
    .X(_2395_));
 sg13g2_nor2_1 _5545_ (.A(_2376_),
    .B(net1674),
    .Y(_0191_));
 sg13g2_nand2_1 _5546_ (.Y(_2396_),
    .A(net1871),
    .B(_1733_));
 sg13g2_a21oi_2 _5547_ (.B1(net2),
    .Y(_2397_),
    .A2(_1733_),
    .A1(\vga_tetris._inputs_io_rightButtonActive ));
 sg13g2_nand2b_1 _5548_ (.Y(_2398_),
    .B(_2396_),
    .A_N(net2));
 sg13g2_nand2_2 _5549_ (.Y(_2399_),
    .A(net1266),
    .B(_2397_));
 sg13g2_nor2_1 _5550_ (.A(\vga_tetris._inputs_io_rightButtonActive ),
    .B(_2355_),
    .Y(_2400_));
 sg13g2_and2_1 _5551_ (.A(_0695_),
    .B(_2357_),
    .X(_2401_));
 sg13g2_nor2_1 _5552_ (.A(net1645),
    .B(_2401_),
    .Y(_2402_));
 sg13g2_and2_1 _5553_ (.A(net1645),
    .B(_2401_),
    .X(_2403_));
 sg13g2_nor3_1 _5554_ (.A(_2399_),
    .B(net1646),
    .C(_2403_),
    .Y(_0192_));
 sg13g2_nand2_1 _5555_ (.Y(_2404_),
    .A(net1717),
    .B(_2403_));
 sg13g2_xnor2_1 _5556_ (.Y(_2405_),
    .A(net1717),
    .B(_2403_));
 sg13g2_nor2_1 _5557_ (.A(_2399_),
    .B(_2405_),
    .Y(_0193_));
 sg13g2_a21oi_1 _5558_ (.A1(net1717),
    .A2(_2403_),
    .Y(_2406_),
    .B1(net1836));
 sg13g2_and4_1 _5559_ (.A(net1836),
    .B(net1717),
    .C(net1645),
    .D(_2400_),
    .X(_2407_));
 sg13g2_nor3_1 _5560_ (.A(_2398_),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_));
 sg13g2_and2_1 _5561_ (.A(net1266),
    .B(net1837),
    .X(_0194_));
 sg13g2_nor2_1 _5562_ (.A(net1876),
    .B(_2407_),
    .Y(_2409_));
 sg13g2_nor3_1 _5563_ (.A(_0696_),
    .B(_0697_),
    .C(_2404_),
    .Y(_2410_));
 sg13g2_nor3_1 _5564_ (.A(_2398_),
    .B(_2409_),
    .C(_2410_),
    .Y(_2411_));
 sg13g2_and2_1 _5565_ (.A(net1266),
    .B(net1877),
    .X(_0195_));
 sg13g2_and3_2 _5566_ (.X(_2412_),
    .A(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .B(net1816),
    .C(_2407_));
 sg13g2_o21ai_1 _5567_ (.B1(_2397_),
    .Y(_2413_),
    .A1(net1816),
    .A2(_2410_));
 sg13g2_nor2_1 _5568_ (.A(_2412_),
    .B(_2413_),
    .Y(_2414_));
 sg13g2_nor3_1 _5569_ (.A(net1252),
    .B(_2412_),
    .C(net1817),
    .Y(_0196_));
 sg13g2_o21ai_1 _5570_ (.B1(_2397_),
    .Y(_2415_),
    .A1(net1841),
    .A2(_2412_));
 sg13g2_a21oi_1 _5571_ (.A1(net1841),
    .A2(_2412_),
    .Y(_2416_),
    .B1(_2415_));
 sg13g2_and2_1 _5572_ (.A(net1265),
    .B(net1842),
    .X(_0197_));
 sg13g2_a21oi_1 _5573_ (.A1(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .A2(_2412_),
    .Y(_2417_),
    .B1(net1424));
 sg13g2_nand3_1 _5574_ (.B(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .C(_2412_),
    .A(net1424),
    .Y(_2418_));
 sg13g2_nand2b_1 _5575_ (.Y(_2419_),
    .B(_2418_),
    .A_N(_2399_));
 sg13g2_nor2_1 _5576_ (.A(net1425),
    .B(_2419_),
    .Y(_0198_));
 sg13g2_xor2_1 _5577_ (.B(_2418_),
    .A(net1706),
    .X(_2420_));
 sg13g2_nor2_1 _5578_ (.A(_2399_),
    .B(net1707),
    .Y(_0199_));
 sg13g2_a21o_2 _5579_ (.A2(net1162),
    .A1(net1692),
    .B1(net4),
    .X(_2421_));
 sg13g2_and2_1 _5580_ (.A(_0702_),
    .B(_2357_),
    .X(_2422_));
 sg13g2_nor3_1 _5581_ (.A(net1692),
    .B(_0704_),
    .C(_2355_),
    .Y(_2423_));
 sg13g2_xnor2_1 _5582_ (.Y(_2424_),
    .A(net1798),
    .B(_2422_));
 sg13g2_nor2_1 _5583_ (.A(net1092),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_nor3_1 _5584_ (.A(net1252),
    .B(net1092),
    .C(_2424_),
    .Y(_0200_));
 sg13g2_nor2_1 _5585_ (.A(net1865),
    .B(_2423_),
    .Y(_2426_));
 sg13g2_and2_1 _5586_ (.A(net1865),
    .B(_2423_),
    .X(_2427_));
 sg13g2_nor3_1 _5587_ (.A(_2421_),
    .B(_2426_),
    .C(_2427_),
    .Y(_2428_));
 sg13g2_and2_1 _5588_ (.A(net1265),
    .B(_2428_),
    .X(_0201_));
 sg13g2_nor2_1 _5589_ (.A(net1870),
    .B(_2427_),
    .Y(_2429_));
 sg13g2_and2_1 _5590_ (.A(net1870),
    .B(_2427_),
    .X(_2430_));
 sg13g2_and4_1 _5591_ (.A(net1798),
    .B(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .C(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .D(_2422_),
    .X(_2431_));
 sg13g2_nor3_1 _5592_ (.A(_2421_),
    .B(_2429_),
    .C(_2430_),
    .Y(_2432_));
 sg13g2_and2_1 _5593_ (.A(net1265),
    .B(_2432_),
    .X(_0202_));
 sg13g2_xnor2_1 _5594_ (.Y(_2433_),
    .A(net1801),
    .B(_2431_));
 sg13g2_nor2_1 _5595_ (.A(net1092),
    .B(_2433_),
    .Y(_2434_));
 sg13g2_nor3_1 _5596_ (.A(net1248),
    .B(net1092),
    .C(net1802),
    .Y(_0203_));
 sg13g2_a21oi_1 _5597_ (.A1(net1801),
    .A2(_2431_),
    .Y(_2435_),
    .B1(net1834));
 sg13g2_and3_1 _5598_ (.X(_2436_),
    .A(net1801),
    .B(net1834),
    .C(_2430_));
 sg13g2_nor3_1 _5599_ (.A(net1092),
    .B(net1835),
    .C(_2436_),
    .Y(_2437_));
 sg13g2_and2_1 _5600_ (.A(net1262),
    .B(_2437_),
    .X(_0204_));
 sg13g2_nor2_1 _5601_ (.A(net1888),
    .B(_2436_),
    .Y(_2438_));
 sg13g2_and2_1 _5602_ (.A(net1888),
    .B(_2436_),
    .X(_2439_));
 sg13g2_nand4_1 _5603_ (.B(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .C(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .A(net1801),
    .Y(_2440_),
    .D(_2431_));
 sg13g2_nor3_1 _5604_ (.A(net1092),
    .B(_2438_),
    .C(_2439_),
    .Y(_2441_));
 sg13g2_and2_1 _5605_ (.A(net1262),
    .B(_2441_),
    .X(_0205_));
 sg13g2_nor2_1 _5606_ (.A(net1867),
    .B(_2439_),
    .Y(_2442_));
 sg13g2_nor2_1 _5607_ (.A(_0705_),
    .B(_2440_),
    .Y(_2443_));
 sg13g2_nor3_1 _5608_ (.A(net1092),
    .B(net1868),
    .C(_2443_),
    .Y(_2444_));
 sg13g2_and2_1 _5609_ (.A(net1262),
    .B(_2444_),
    .X(_0206_));
 sg13g2_a21oi_1 _5610_ (.A1(net1803),
    .A2(_2443_),
    .Y(_2445_),
    .B1(net1092));
 sg13g2_o21ai_1 _5611_ (.B1(net1804),
    .Y(_2446_),
    .A1(net1803),
    .A2(_2443_));
 sg13g2_nor2_1 _5612_ (.A(net1249),
    .B(net1805),
    .Y(_0207_));
 sg13g2_o21ai_1 _5613_ (.B1(_2364_),
    .Y(_2447_),
    .A1(_2367_),
    .A2(_2368_));
 sg13g2_a21oi_1 _5614_ (.A1(_2350_),
    .A2(_2366_),
    .Y(_2448_),
    .B1(_2447_));
 sg13g2_nor4_1 _5615_ (.A(_0698_),
    .B(_2369_),
    .C(_2370_),
    .D(_2448_),
    .Y(_2449_));
 sg13g2_o21ai_1 _5616_ (.B1(_2349_),
    .Y(_2450_),
    .A1(net1650),
    .A2(_2449_));
 sg13g2_nand2b_1 _5617_ (.Y(_0208_),
    .B(_2450_),
    .A_N(_0183_));
 sg13g2_nor3_1 _5618_ (.A(_2384_),
    .B(_2387_),
    .C(_2390_),
    .Y(_2451_));
 sg13g2_nor4_1 _5619_ (.A(_2375_),
    .B(_2391_),
    .C(_2392_),
    .D(_2451_),
    .Y(_2452_));
 sg13g2_a21o_1 _5620_ (.A2(_2452_),
    .A1(net1730),
    .B1(net1866),
    .X(_2453_));
 sg13g2_nand3_1 _5621_ (.B(_2374_),
    .C(_2453_),
    .A(net1269),
    .Y(_2454_));
 sg13g2_nand2b_1 _5622_ (.Y(_0209_),
    .B(_2454_),
    .A_N(_0191_));
 sg13g2_nor3_1 _5623_ (.A(_2408_),
    .B(_2411_),
    .C(_2414_),
    .Y(_2455_));
 sg13g2_nand2_1 _5624_ (.Y(_2456_),
    .A(net1424),
    .B(_2416_));
 sg13g2_o21ai_1 _5625_ (.B1(_0695_),
    .Y(_2457_),
    .A1(_2455_),
    .A2(_2456_));
 sg13g2_nand3_1 _5626_ (.B(_2396_),
    .C(_2457_),
    .A(net1266),
    .Y(_2458_));
 sg13g2_nand2b_1 _5627_ (.Y(_0210_),
    .B(_2458_),
    .A_N(net1708));
 sg13g2_nor4_1 _5628_ (.A(net1692),
    .B(_2425_),
    .C(_2428_),
    .D(_2432_),
    .Y(_2459_));
 sg13g2_nand2b_1 _5629_ (.Y(_2460_),
    .B(_2459_),
    .A_N(_2434_));
 sg13g2_nor4_1 _5630_ (.A(_2437_),
    .B(_2441_),
    .C(_2444_),
    .D(_2460_),
    .Y(_2461_));
 sg13g2_a221oi_1 _5631_ (.B2(_2461_),
    .C1(net1249),
    .B1(_2446_),
    .A1(net1692),
    .Y(_0211_),
    .A2(net1162));
 sg13g2_or2_1 _5632_ (.X(_2462_),
    .B(net1854),
    .A(net1246));
 sg13g2_nor3_1 _5633_ (.A(net1206),
    .B(net1226),
    .C(_2462_),
    .Y(_0212_));
 sg13g2_nand2_1 _5634_ (.Y(_2463_),
    .A(_0799_),
    .B(_2265_));
 sg13g2_or3_1 _5635_ (.A(_0816_),
    .B(_0830_),
    .C(_2463_),
    .X(_2464_));
 sg13g2_nor3_2 _5636_ (.A(_0787_),
    .B(_0793_),
    .C(_2464_),
    .Y(_2465_));
 sg13g2_nor2_1 _5637_ (.A(net1501),
    .B(net977),
    .Y(_2466_));
 sg13g2_a21oi_1 _5638_ (.A1(net1151),
    .A2(net977),
    .Y(_0213_),
    .B1(_2466_));
 sg13g2_nor2_1 _5639_ (.A(net1537),
    .B(net977),
    .Y(_2467_));
 sg13g2_a21oi_1 _5640_ (.A1(net1149),
    .A2(net977),
    .Y(_0214_),
    .B1(_2467_));
 sg13g2_nor2_1 _5641_ (.A(net1594),
    .B(net975),
    .Y(_2468_));
 sg13g2_a21oi_1 _5642_ (.A1(_2280_),
    .A2(net975),
    .Y(_0215_),
    .B1(_2468_));
 sg13g2_nor2_1 _5643_ (.A(net1407),
    .B(net975),
    .Y(_2469_));
 sg13g2_a21oi_1 _5644_ (.A1(_2284_),
    .A2(net975),
    .Y(_0216_),
    .B1(_2469_));
 sg13g2_nor2_1 _5645_ (.A(net1517),
    .B(net973),
    .Y(_2470_));
 sg13g2_a21oi_1 _5646_ (.A1(net1140),
    .A2(net973),
    .Y(_0217_),
    .B1(_2470_));
 sg13g2_nor2_1 _5647_ (.A(net1395),
    .B(net971),
    .Y(_2471_));
 sg13g2_a21oi_1 _5648_ (.A1(_2292_),
    .A2(net971),
    .Y(_0218_),
    .B1(_2471_));
 sg13g2_nor2_1 _5649_ (.A(net1485),
    .B(net971),
    .Y(_2472_));
 sg13g2_a21oi_1 _5650_ (.A1(net1134),
    .A2(net971),
    .Y(_0219_),
    .B1(_2472_));
 sg13g2_nor2_1 _5651_ (.A(net1440),
    .B(net971),
    .Y(_2473_));
 sg13g2_a21oi_1 _5652_ (.A1(net1131),
    .A2(net971),
    .Y(_0220_),
    .B1(_2473_));
 sg13g2_nor2_1 _5653_ (.A(net1527),
    .B(net977),
    .Y(_2474_));
 sg13g2_a21oi_1 _5654_ (.A1(net1128),
    .A2(net977),
    .Y(_0221_),
    .B1(_2474_));
 sg13g2_nor2_1 _5655_ (.A(net1489),
    .B(net977),
    .Y(_2475_));
 sg13g2_a21oi_1 _5656_ (.A1(_2308_),
    .A2(net974),
    .Y(_0222_),
    .B1(_2475_));
 sg13g2_nor2_1 _5657_ (.A(net1511),
    .B(net972),
    .Y(_2476_));
 sg13g2_a21oi_1 _5658_ (.A1(net1122),
    .A2(net972),
    .Y(_0223_),
    .B1(_2476_));
 sg13g2_nor2_1 _5659_ (.A(net1447),
    .B(net971),
    .Y(_2477_));
 sg13g2_a21oi_1 _5660_ (.A1(net1119),
    .A2(net971),
    .Y(_0224_),
    .B1(_2477_));
 sg13g2_nor2_1 _5661_ (.A(net1439),
    .B(net974),
    .Y(_2478_));
 sg13g2_a21oi_1 _5662_ (.A1(net1116),
    .A2(net974),
    .Y(_0225_),
    .B1(_2478_));
 sg13g2_nor2_1 _5663_ (.A(net1546),
    .B(net974),
    .Y(_2479_));
 sg13g2_a21oi_1 _5664_ (.A1(_2324_),
    .A2(net974),
    .Y(_0226_),
    .B1(_2479_));
 sg13g2_nor2_1 _5665_ (.A(net1539),
    .B(net975),
    .Y(_2480_));
 sg13g2_a21oi_1 _5666_ (.A1(_2328_),
    .A2(net975),
    .Y(_0227_),
    .B1(_2480_));
 sg13g2_nor2_1 _5667_ (.A(net1421),
    .B(net976),
    .Y(_2481_));
 sg13g2_a21oi_1 _5668_ (.A1(_2332_),
    .A2(net976),
    .Y(_0228_),
    .B1(_2481_));
 sg13g2_nor2_1 _5669_ (.A(net1416),
    .B(net975),
    .Y(_2482_));
 sg13g2_a21oi_1 _5670_ (.A1(net1102),
    .A2(net975),
    .Y(_0229_),
    .B1(_2482_));
 sg13g2_nor2_1 _5671_ (.A(net1417),
    .B(net976),
    .Y(_2483_));
 sg13g2_a21oi_1 _5672_ (.A1(net1099),
    .A2(net976),
    .Y(_0230_),
    .B1(_2483_));
 sg13g2_nor2_1 _5673_ (.A(net1469),
    .B(net972),
    .Y(_2484_));
 sg13g2_a21oi_1 _5674_ (.A1(net1098),
    .A2(net972),
    .Y(_0231_),
    .B1(_2484_));
 sg13g2_nor2_1 _5675_ (.A(net1526),
    .B(net973),
    .Y(_2485_));
 sg13g2_a21oi_1 _5676_ (.A1(net1095),
    .A2(net973),
    .Y(_0232_),
    .B1(_2485_));
 sg13g2_o21ai_1 _5677_ (.B1(_0816_),
    .Y(_2486_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_or2_1 _5678_ (.X(_2487_),
    .B(_2486_),
    .A(_2463_));
 sg13g2_nor3_1 _5679_ (.A(_0787_),
    .B(_0793_),
    .C(_2487_),
    .Y(_2488_));
 sg13g2_nor2_1 _5680_ (.A(net1612),
    .B(net969),
    .Y(_2489_));
 sg13g2_a21oi_1 _5681_ (.A1(net1151),
    .A2(net969),
    .Y(_0233_),
    .B1(_2489_));
 sg13g2_nor2_1 _5682_ (.A(net1448),
    .B(net969),
    .Y(_2490_));
 sg13g2_a21oi_1 _5683_ (.A1(net1149),
    .A2(net969),
    .Y(_0234_),
    .B1(_2490_));
 sg13g2_nor2_1 _5684_ (.A(net1500),
    .B(net967),
    .Y(_2491_));
 sg13g2_a21oi_1 _5685_ (.A1(net1146),
    .A2(net967),
    .Y(_0235_),
    .B1(_2491_));
 sg13g2_nor2_1 _5686_ (.A(net1471),
    .B(net967),
    .Y(_2492_));
 sg13g2_a21oi_1 _5687_ (.A1(net1143),
    .A2(net967),
    .Y(_0236_),
    .B1(_2492_));
 sg13g2_nor2_1 _5688_ (.A(net1462),
    .B(net965),
    .Y(_2493_));
 sg13g2_a21oi_1 _5689_ (.A1(net1139),
    .A2(net965),
    .Y(_0237_),
    .B1(_2493_));
 sg13g2_nor2_1 _5690_ (.A(net1504),
    .B(net965),
    .Y(_2494_));
 sg13g2_a21oi_1 _5691_ (.A1(net1137),
    .A2(net965),
    .Y(_0238_),
    .B1(_2494_));
 sg13g2_nor2_1 _5692_ (.A(net1609),
    .B(net964),
    .Y(_2495_));
 sg13g2_a21oi_1 _5693_ (.A1(net1134),
    .A2(net964),
    .Y(_0239_),
    .B1(_2495_));
 sg13g2_nor2_1 _5694_ (.A(net1569),
    .B(net964),
    .Y(_2496_));
 sg13g2_a21oi_1 _5695_ (.A1(net1130),
    .A2(net964),
    .Y(_0240_),
    .B1(_2496_));
 sg13g2_nor2_1 _5696_ (.A(net1585),
    .B(net969),
    .Y(_2497_));
 sg13g2_a21oi_1 _5697_ (.A1(net1126),
    .A2(net969),
    .Y(_0241_),
    .B1(_2497_));
 sg13g2_nor2_1 _5698_ (.A(net1559),
    .B(net969),
    .Y(_2498_));
 sg13g2_a21oi_1 _5699_ (.A1(net1125),
    .A2(net969),
    .Y(_0242_),
    .B1(_2498_));
 sg13g2_nor2_1 _5700_ (.A(net1487),
    .B(net966),
    .Y(_2499_));
 sg13g2_a21oi_1 _5701_ (.A1(net1120),
    .A2(net966),
    .Y(_0243_),
    .B1(_2499_));
 sg13g2_nor2_1 _5702_ (.A(net1497),
    .B(net964),
    .Y(_2500_));
 sg13g2_a21oi_1 _5703_ (.A1(net1118),
    .A2(net964),
    .Y(_0244_),
    .B1(_2500_));
 sg13g2_nor2_1 _5704_ (.A(net1525),
    .B(net966),
    .Y(_2501_));
 sg13g2_a21oi_1 _5705_ (.A1(net1114),
    .A2(net966),
    .Y(_0245_),
    .B1(_2501_));
 sg13g2_nor2_1 _5706_ (.A(net1456),
    .B(net965),
    .Y(_2502_));
 sg13g2_a21oi_1 _5707_ (.A1(net1112),
    .A2(net965),
    .Y(_0246_),
    .B1(_2502_));
 sg13g2_nor2_1 _5708_ (.A(net1556),
    .B(net967),
    .Y(_2503_));
 sg13g2_a21oi_1 _5709_ (.A1(net1108),
    .A2(net967),
    .Y(_0247_),
    .B1(_2503_));
 sg13g2_nor2_1 _5710_ (.A(net1581),
    .B(net967),
    .Y(_2504_));
 sg13g2_a21oi_1 _5711_ (.A1(net1106),
    .A2(net967),
    .Y(_0248_),
    .B1(_2504_));
 sg13g2_nor2_1 _5712_ (.A(net1606),
    .B(net968),
    .Y(_2505_));
 sg13g2_a21oi_1 _5713_ (.A1(net1104),
    .A2(net968),
    .Y(_0249_),
    .B1(_2505_));
 sg13g2_nor2_1 _5714_ (.A(net1542),
    .B(net968),
    .Y(_2506_));
 sg13g2_a21oi_1 _5715_ (.A1(net1100),
    .A2(net968),
    .Y(_0250_),
    .B1(_2506_));
 sg13g2_nor2_1 _5716_ (.A(net1402),
    .B(net964),
    .Y(_2507_));
 sg13g2_a21oi_1 _5717_ (.A1(net1096),
    .A2(net964),
    .Y(_0251_),
    .B1(_2507_));
 sg13g2_nor2_1 _5718_ (.A(net1553),
    .B(net965),
    .Y(_2508_));
 sg13g2_a21oi_1 _5719_ (.A1(net1094),
    .A2(net965),
    .Y(_0252_),
    .B1(_2508_));
 sg13g2_nand2b_1 _5720_ (.Y(_2509_),
    .B(_0830_),
    .A_N(_0816_));
 sg13g2_or2_1 _5721_ (.X(_2510_),
    .B(_2509_),
    .A(_2463_));
 sg13g2_nor3_1 _5722_ (.A(_0787_),
    .B(_0793_),
    .C(_2510_),
    .Y(_2511_));
 sg13g2_nor2_1 _5723_ (.A(net1478),
    .B(net962),
    .Y(_2512_));
 sg13g2_a21oi_1 _5724_ (.A1(net1150),
    .A2(net962),
    .Y(_0253_),
    .B1(_2512_));
 sg13g2_nor2_1 _5725_ (.A(net1505),
    .B(net962),
    .Y(_2513_));
 sg13g2_a21oi_1 _5726_ (.A1(net1147),
    .A2(net962),
    .Y(_0254_),
    .B1(_2513_));
 sg13g2_nor2_1 _5727_ (.A(net1510),
    .B(net960),
    .Y(_2514_));
 sg13g2_a21oi_1 _5728_ (.A1(net1145),
    .A2(net960),
    .Y(_0255_),
    .B1(_2514_));
 sg13g2_nor2_1 _5729_ (.A(net1613),
    .B(net961),
    .Y(_2515_));
 sg13g2_a21oi_1 _5730_ (.A1(net1142),
    .A2(net961),
    .Y(_0256_),
    .B1(_2515_));
 sg13g2_nor2_1 _5731_ (.A(net1473),
    .B(net963),
    .Y(_2516_));
 sg13g2_a21oi_1 _5732_ (.A1(net1139),
    .A2(net963),
    .Y(_0257_),
    .B1(_2516_));
 sg13g2_nor2_1 _5733_ (.A(net1593),
    .B(net957),
    .Y(_2517_));
 sg13g2_a21oi_1 _5734_ (.A1(net1135),
    .A2(net957),
    .Y(_0258_),
    .B1(_2517_));
 sg13g2_nor2_1 _5735_ (.A(net1493),
    .B(net957),
    .Y(_2518_));
 sg13g2_a21oi_1 _5736_ (.A1(net1132),
    .A2(net957),
    .Y(_0259_),
    .B1(_2518_));
 sg13g2_nor2_1 _5737_ (.A(net1555),
    .B(net957),
    .Y(_2519_));
 sg13g2_a21oi_1 _5738_ (.A1(net1129),
    .A2(net957),
    .Y(_0260_),
    .B1(_2519_));
 sg13g2_nor2_1 _5739_ (.A(net1397),
    .B(net962),
    .Y(_2520_));
 sg13g2_a21oi_1 _5740_ (.A1(net1126),
    .A2(net962),
    .Y(_0261_),
    .B1(_2520_));
 sg13g2_nor2_1 _5741_ (.A(net1506),
    .B(net962),
    .Y(_2521_));
 sg13g2_a21oi_1 _5742_ (.A1(net1123),
    .A2(net962),
    .Y(_0262_),
    .B1(_2521_));
 sg13g2_nor2_1 _5743_ (.A(net1533),
    .B(net958),
    .Y(_2522_));
 sg13g2_a21oi_1 _5744_ (.A1(net1121),
    .A2(net958),
    .Y(_0263_),
    .B1(_2522_));
 sg13g2_nor2_1 _5745_ (.A(net1394),
    .B(net957),
    .Y(_2523_));
 sg13g2_a21oi_1 _5746_ (.A1(net1118),
    .A2(net957),
    .Y(_0264_),
    .B1(_2523_));
 sg13g2_nor2_1 _5747_ (.A(net1620),
    .B(net959),
    .Y(_2524_));
 sg13g2_a21oi_1 _5748_ (.A1(net1116),
    .A2(net959),
    .Y(_0265_),
    .B1(_2524_));
 sg13g2_nor2_1 _5749_ (.A(net1529),
    .B(net959),
    .Y(_2525_));
 sg13g2_a21oi_1 _5750_ (.A1(net1111),
    .A2(net959),
    .Y(_0266_),
    .B1(_2525_));
 sg13g2_nor2_1 _5751_ (.A(net1598),
    .B(net960),
    .Y(_2526_));
 sg13g2_a21oi_1 _5752_ (.A1(net1110),
    .A2(net960),
    .Y(_0267_),
    .B1(_2526_));
 sg13g2_nor2_1 _5753_ (.A(net1561),
    .B(net960),
    .Y(_2527_));
 sg13g2_a21oi_1 _5754_ (.A1(net1106),
    .A2(net960),
    .Y(_0268_),
    .B1(_2527_));
 sg13g2_nor2_1 _5755_ (.A(net1461),
    .B(net960),
    .Y(_2528_));
 sg13g2_a21oi_1 _5756_ (.A1(net1103),
    .A2(net960),
    .Y(_0269_),
    .B1(_2528_));
 sg13g2_nor2_1 _5757_ (.A(net1587),
    .B(net961),
    .Y(_2529_));
 sg13g2_a21oi_1 _5758_ (.A1(net1100),
    .A2(net961),
    .Y(_0270_),
    .B1(_2529_));
 sg13g2_nor2_1 _5759_ (.A(net1541),
    .B(net958),
    .Y(_2530_));
 sg13g2_a21oi_1 _5760_ (.A1(net1097),
    .A2(net958),
    .Y(_0271_),
    .B1(_2530_));
 sg13g2_nor2_1 _5761_ (.A(net1560),
    .B(net959),
    .Y(_2531_));
 sg13g2_a21oi_1 _5762_ (.A1(net1094),
    .A2(net959),
    .Y(_0272_),
    .B1(_2531_));
 sg13g2_or2_1 _5763_ (.X(_2532_),
    .B(_2463_),
    .A(_2262_));
 sg13g2_nor3_1 _5764_ (.A(_0787_),
    .B(_0793_),
    .C(_2532_),
    .Y(_2533_));
 sg13g2_nor2_1 _5765_ (.A(net1608),
    .B(net955),
    .Y(_2534_));
 sg13g2_a21oi_1 _5766_ (.A1(net1151),
    .A2(net955),
    .Y(_0273_),
    .B1(_2534_));
 sg13g2_nor2_1 _5767_ (.A(net1575),
    .B(net954),
    .Y(_2535_));
 sg13g2_a21oi_1 _5768_ (.A1(net1148),
    .A2(net954),
    .Y(_0274_),
    .B1(_2535_));
 sg13g2_nor2_1 _5769_ (.A(net1534),
    .B(net953),
    .Y(_2536_));
 sg13g2_a21oi_1 _5770_ (.A1(net1146),
    .A2(net953),
    .Y(_0275_),
    .B1(_2536_));
 sg13g2_nor2_1 _5771_ (.A(net1535),
    .B(net953),
    .Y(_2537_));
 sg13g2_a21oi_1 _5772_ (.A1(net1143),
    .A2(net953),
    .Y(_0276_),
    .B1(_2537_));
 sg13g2_nor2_1 _5773_ (.A(net1502),
    .B(net956),
    .Y(_2538_));
 sg13g2_a21oi_1 _5774_ (.A1(net1138),
    .A2(net956),
    .Y(_0277_),
    .B1(_2538_));
 sg13g2_nor2_1 _5775_ (.A(net1520),
    .B(net951),
    .Y(_2539_));
 sg13g2_a21oi_1 _5776_ (.A1(net1136),
    .A2(net951),
    .Y(_0278_),
    .B1(_2539_));
 sg13g2_nor2_1 _5777_ (.A(net1442),
    .B(net951),
    .Y(_2540_));
 sg13g2_a21oi_1 _5778_ (.A1(net1134),
    .A2(net951),
    .Y(_0279_),
    .B1(_2540_));
 sg13g2_nor2_1 _5779_ (.A(net1563),
    .B(net952),
    .Y(_2541_));
 sg13g2_a21oi_1 _5780_ (.A1(net1129),
    .A2(net952),
    .Y(_0280_),
    .B1(_2541_));
 sg13g2_nor2_1 _5781_ (.A(net1564),
    .B(net955),
    .Y(_2542_));
 sg13g2_a21oi_1 _5782_ (.A1(net1128),
    .A2(net955),
    .Y(_0281_),
    .B1(_2542_));
 sg13g2_nor2_1 _5783_ (.A(net1554),
    .B(net955),
    .Y(_2543_));
 sg13g2_a21oi_1 _5784_ (.A1(net1125),
    .A2(net955),
    .Y(_0282_),
    .B1(_2543_));
 sg13g2_nor2_1 _5785_ (.A(net1572),
    .B(net952),
    .Y(_2544_));
 sg13g2_a21oi_1 _5786_ (.A1(net1120),
    .A2(net952),
    .Y(_0283_),
    .B1(_2544_));
 sg13g2_nor2_1 _5787_ (.A(net1629),
    .B(net952),
    .Y(_2545_));
 sg13g2_a21oi_1 _5788_ (.A1(net1117),
    .A2(net952),
    .Y(_0284_),
    .B1(_2545_));
 sg13g2_nor2_1 _5789_ (.A(net1477),
    .B(net951),
    .Y(_2546_));
 sg13g2_a21oi_1 _5790_ (.A1(net1114),
    .A2(net951),
    .Y(_0285_),
    .B1(_2546_));
 sg13g2_nor2_1 _5791_ (.A(net1498),
    .B(net955),
    .Y(_2547_));
 sg13g2_a21oi_1 _5792_ (.A1(net1112),
    .A2(net955),
    .Y(_0286_),
    .B1(_2547_));
 sg13g2_nor2_1 _5793_ (.A(net1507),
    .B(net953),
    .Y(_2548_));
 sg13g2_a21oi_1 _5794_ (.A1(net1109),
    .A2(net953),
    .Y(_0287_),
    .B1(_2548_));
 sg13g2_nor2_1 _5795_ (.A(net1532),
    .B(net953),
    .Y(_2549_));
 sg13g2_a21oi_1 _5796_ (.A1(net1107),
    .A2(net953),
    .Y(_0288_),
    .B1(_2549_));
 sg13g2_nor2_1 _5797_ (.A(net1573),
    .B(net954),
    .Y(_2550_));
 sg13g2_a21oi_1 _5798_ (.A1(net1102),
    .A2(net954),
    .Y(_0289_),
    .B1(_2550_));
 sg13g2_nor2_1 _5799_ (.A(net1460),
    .B(net954),
    .Y(_2551_));
 sg13g2_a21oi_1 _5800_ (.A1(net1099),
    .A2(net954),
    .Y(_0290_),
    .B1(_2551_));
 sg13g2_nor2_1 _5801_ (.A(net1521),
    .B(net952),
    .Y(_2552_));
 sg13g2_a21oi_1 _5802_ (.A1(net1096),
    .A2(net952),
    .Y(_0291_),
    .B1(_2552_));
 sg13g2_nor2_1 _5803_ (.A(net1492),
    .B(net951),
    .Y(_2553_));
 sg13g2_a21oi_1 _5804_ (.A1(net1095),
    .A2(net951),
    .Y(_0292_),
    .B1(_2553_));
 sg13g2_nand2b_1 _5805_ (.Y(_2554_),
    .B(_0793_),
    .A_N(_0787_));
 sg13g2_or2_1 _5806_ (.X(_2555_),
    .B(_2554_),
    .A(_2464_));
 sg13g2_nand2_1 _5807_ (.Y(_2556_),
    .A(net795),
    .B(net949));
 sg13g2_o21ai_1 _5808_ (.B1(_2556_),
    .Y(_0293_),
    .A1(net1150),
    .A2(net949));
 sg13g2_nand2_1 _5809_ (.Y(_2557_),
    .A(net834),
    .B(net949));
 sg13g2_o21ai_1 _5810_ (.B1(_2557_),
    .Y(_0294_),
    .A1(net1147),
    .A2(net949));
 sg13g2_nand2_1 _5811_ (.Y(_2558_),
    .A(net835),
    .B(net947));
 sg13g2_o21ai_1 _5812_ (.B1(_2558_),
    .Y(_0295_),
    .A1(net1144),
    .A2(net947));
 sg13g2_nand2_1 _5813_ (.Y(_2559_),
    .A(net1293),
    .B(net948));
 sg13g2_o21ai_1 _5814_ (.B1(_2559_),
    .Y(_0296_),
    .A1(net1141),
    .A2(net948));
 sg13g2_nand2_1 _5815_ (.Y(_2560_),
    .A(net668),
    .B(net950));
 sg13g2_o21ai_1 _5816_ (.B1(_2560_),
    .Y(_0297_),
    .A1(net1138),
    .A2(net950));
 sg13g2_nand2_1 _5817_ (.Y(_2561_),
    .A(net1348),
    .B(net944));
 sg13g2_o21ai_1 _5818_ (.B1(_2561_),
    .Y(_0298_),
    .A1(net1135),
    .A2(net944));
 sg13g2_nand2_1 _5819_ (.Y(_2562_),
    .A(net759),
    .B(net944));
 sg13g2_o21ai_1 _5820_ (.B1(_2562_),
    .Y(_0299_),
    .A1(net1133),
    .A2(net944));
 sg13g2_nand2_1 _5821_ (.Y(_2563_),
    .A(net1324),
    .B(net944));
 sg13g2_o21ai_1 _5822_ (.B1(_2563_),
    .Y(_0300_),
    .A1(net1131),
    .A2(net944));
 sg13g2_nand2_1 _5823_ (.Y(_2564_),
    .A(net1306),
    .B(net949));
 sg13g2_o21ai_1 _5824_ (.B1(_2564_),
    .Y(_0301_),
    .A1(net1126),
    .A2(net949));
 sg13g2_nand2_1 _5825_ (.Y(_2565_),
    .A(net736),
    .B(net949));
 sg13g2_o21ai_1 _5826_ (.B1(_2565_),
    .Y(_0302_),
    .A1(net1123),
    .A2(net949));
 sg13g2_nand2_1 _5827_ (.Y(_2566_),
    .A(net696),
    .B(net945));
 sg13g2_o21ai_1 _5828_ (.B1(_2566_),
    .Y(_0303_),
    .A1(net1122),
    .A2(net945));
 sg13g2_nand2_1 _5829_ (.Y(_2567_),
    .A(net686),
    .B(net944));
 sg13g2_o21ai_1 _5830_ (.B1(_2567_),
    .Y(_0304_),
    .A1(net1119),
    .A2(net944));
 sg13g2_nand2_1 _5831_ (.Y(_2568_),
    .A(net663),
    .B(net946));
 sg13g2_o21ai_1 _5832_ (.B1(_2568_),
    .Y(_0305_),
    .A1(net1115),
    .A2(net946));
 sg13g2_nand2_1 _5833_ (.Y(_2569_),
    .A(net1341),
    .B(net946));
 sg13g2_o21ai_1 _5834_ (.B1(_2569_),
    .Y(_0306_),
    .A1(net1111),
    .A2(net946));
 sg13g2_nand2_1 _5835_ (.Y(_2570_),
    .A(net667),
    .B(net947));
 sg13g2_o21ai_1 _5836_ (.B1(_2570_),
    .Y(_0307_),
    .A1(net1108),
    .A2(net947));
 sg13g2_nand2_1 _5837_ (.Y(_2571_),
    .A(net1379),
    .B(net947));
 sg13g2_o21ai_1 _5838_ (.B1(_2571_),
    .Y(_0308_),
    .A1(net1105),
    .A2(net947));
 sg13g2_nand2_1 _5839_ (.Y(_2572_),
    .A(net699),
    .B(net948));
 sg13g2_o21ai_1 _5840_ (.B1(_2572_),
    .Y(_0309_),
    .A1(net1102),
    .A2(net948));
 sg13g2_nand2_1 _5841_ (.Y(_2573_),
    .A(net727),
    .B(net947));
 sg13g2_o21ai_1 _5842_ (.B1(_2573_),
    .Y(_0310_),
    .A1(net1101),
    .A2(net947));
 sg13g2_nand2_1 _5843_ (.Y(_2574_),
    .A(net839),
    .B(net945));
 sg13g2_o21ai_1 _5844_ (.B1(_2574_),
    .Y(_0311_),
    .A1(net1096),
    .A2(net945));
 sg13g2_nand2_1 _5845_ (.Y(_2575_),
    .A(net1360),
    .B(net946));
 sg13g2_o21ai_1 _5846_ (.B1(_2575_),
    .Y(_0312_),
    .A1(net1093),
    .A2(net946));
 sg13g2_or2_1 _5847_ (.X(_2576_),
    .B(_2554_),
    .A(_2487_));
 sg13g2_nand2_1 _5848_ (.Y(_2577_),
    .A(net1345),
    .B(net942));
 sg13g2_o21ai_1 _5849_ (.B1(_2577_),
    .Y(_0313_),
    .A1(net1151),
    .A2(net942));
 sg13g2_nand2_1 _5850_ (.Y(_2578_),
    .A(net765),
    .B(net940));
 sg13g2_o21ai_1 _5851_ (.B1(_2578_),
    .Y(_0314_),
    .A1(net1149),
    .A2(net940));
 sg13g2_nand2_1 _5852_ (.Y(_2579_),
    .A(net716),
    .B(net941));
 sg13g2_o21ai_1 _5853_ (.B1(_2579_),
    .Y(_0315_),
    .A1(net1146),
    .A2(net941));
 sg13g2_nand2_1 _5854_ (.Y(_2580_),
    .A(net838),
    .B(net941));
 sg13g2_o21ai_1 _5855_ (.B1(_2580_),
    .Y(_0316_),
    .A1(net1141),
    .A2(net941));
 sg13g2_nand2_1 _5856_ (.Y(_2581_),
    .A(net1327),
    .B(net943));
 sg13g2_o21ai_1 _5857_ (.B1(_2581_),
    .Y(_0317_),
    .A1(net1139),
    .A2(net943));
 sg13g2_nand2_1 _5858_ (.Y(_2582_),
    .A(net656),
    .B(net937));
 sg13g2_o21ai_1 _5859_ (.B1(_2582_),
    .Y(_0318_),
    .A1(net1136),
    .A2(net937));
 sg13g2_nand2_1 _5860_ (.Y(_2583_),
    .A(net801),
    .B(net937));
 sg13g2_o21ai_1 _5861_ (.B1(_2583_),
    .Y(_0319_),
    .A1(net1133),
    .A2(net937));
 sg13g2_nand2_1 _5862_ (.Y(_2584_),
    .A(net1291),
    .B(net937));
 sg13g2_o21ai_1 _5863_ (.B1(_2584_),
    .Y(_0320_),
    .A1(net1130),
    .A2(net937));
 sg13g2_nand2_1 _5864_ (.Y(_2585_),
    .A(net675),
    .B(net940));
 sg13g2_o21ai_1 _5865_ (.B1(_2585_),
    .Y(_0321_),
    .A1(net1127),
    .A2(net940));
 sg13g2_nand2_1 _5866_ (.Y(_2586_),
    .A(net833),
    .B(net940));
 sg13g2_o21ai_1 _5867_ (.B1(_2586_),
    .Y(_0322_),
    .A1(net1125),
    .A2(net940));
 sg13g2_nand2_1 _5868_ (.Y(_2587_),
    .A(net825),
    .B(net938));
 sg13g2_o21ai_1 _5869_ (.B1(_2587_),
    .Y(_0323_),
    .A1(net1121),
    .A2(net938));
 sg13g2_nand2_1 _5870_ (.Y(_2588_),
    .A(net793),
    .B(net937));
 sg13g2_o21ai_1 _5871_ (.B1(_2588_),
    .Y(_0324_),
    .A1(net1119),
    .A2(net937));
 sg13g2_nand2_1 _5872_ (.Y(_2589_),
    .A(net1337),
    .B(net939));
 sg13g2_o21ai_1 _5873_ (.B1(_2589_),
    .Y(_0325_),
    .A1(net1114),
    .A2(net939));
 sg13g2_nand2_1 _5874_ (.Y(_2590_),
    .A(net812),
    .B(net939));
 sg13g2_o21ai_1 _5875_ (.B1(_2590_),
    .Y(_0326_),
    .A1(net1112),
    .A2(net939));
 sg13g2_nand2_1 _5876_ (.Y(_2591_),
    .A(net1377),
    .B(net941));
 sg13g2_o21ai_1 _5877_ (.B1(_2591_),
    .Y(_0327_),
    .A1(net1110),
    .A2(net941));
 sg13g2_nand2_1 _5878_ (.Y(_2592_),
    .A(net1281),
    .B(net940));
 sg13g2_o21ai_1 _5879_ (.B1(_2592_),
    .Y(_0328_),
    .A1(net1106),
    .A2(net940));
 sg13g2_nand2_1 _5880_ (.Y(_2593_),
    .A(net1326),
    .B(net941));
 sg13g2_o21ai_1 _5881_ (.B1(_2593_),
    .Y(_0329_),
    .A1(net1102),
    .A2(net941));
 sg13g2_nand2_1 _5882_ (.Y(_2594_),
    .A(net703),
    .B(net942));
 sg13g2_o21ai_1 _5883_ (.B1(_2594_),
    .Y(_0330_),
    .A1(net1100),
    .A2(net942));
 sg13g2_nand2_1 _5884_ (.Y(_2595_),
    .A(net694),
    .B(net938));
 sg13g2_o21ai_1 _5885_ (.B1(_2595_),
    .Y(_0331_),
    .A1(net1096),
    .A2(net938));
 sg13g2_nand2_1 _5886_ (.Y(_2596_),
    .A(net809),
    .B(net939));
 sg13g2_o21ai_1 _5887_ (.B1(_2596_),
    .Y(_0332_),
    .A1(net1094),
    .A2(net939));
 sg13g2_or2_1 _5888_ (.X(_2597_),
    .B(_2554_),
    .A(_2510_));
 sg13g2_nand2_1 _5889_ (.Y(_2598_),
    .A(net767),
    .B(net935));
 sg13g2_o21ai_1 _5890_ (.B1(_2598_),
    .Y(_0333_),
    .A1(net1150),
    .A2(net935));
 sg13g2_nand2_1 _5891_ (.Y(_2599_),
    .A(net761),
    .B(net933));
 sg13g2_o21ai_1 _5892_ (.B1(_2599_),
    .Y(_0334_),
    .A1(net1148),
    .A2(net933));
 sg13g2_nand2_1 _5893_ (.Y(_2600_),
    .A(net1284),
    .B(net933));
 sg13g2_o21ai_1 _5894_ (.B1(_2600_),
    .Y(_0335_),
    .A1(net1144),
    .A2(net933));
 sg13g2_nand2_1 _5895_ (.Y(_2601_),
    .A(net785),
    .B(net934));
 sg13g2_o21ai_1 _5896_ (.B1(_2601_),
    .Y(_0336_),
    .A1(net1141),
    .A2(net934));
 sg13g2_nand2_1 _5897_ (.Y(_2602_),
    .A(net734),
    .B(net932));
 sg13g2_o21ai_1 _5898_ (.B1(_2602_),
    .Y(_0337_),
    .A1(net1138),
    .A2(net932));
 sg13g2_nand2_1 _5899_ (.Y(_2603_),
    .A(net1320),
    .B(net930));
 sg13g2_o21ai_1 _5900_ (.B1(_2603_),
    .Y(_0338_),
    .A1(net1135),
    .A2(net930));
 sg13g2_nand2_1 _5901_ (.Y(_2604_),
    .A(net1315),
    .B(net930));
 sg13g2_o21ai_1 _5902_ (.B1(_2604_),
    .Y(_0339_),
    .A1(net1133),
    .A2(net930));
 sg13g2_nand2_1 _5903_ (.Y(_2605_),
    .A(net1365),
    .B(net931));
 sg13g2_o21ai_1 _5904_ (.B1(_2605_),
    .Y(_0340_),
    .A1(net1129),
    .A2(net931));
 sg13g2_nand2_1 _5905_ (.Y(_2606_),
    .A(net721),
    .B(net935));
 sg13g2_o21ai_1 _5906_ (.B1(_2606_),
    .Y(_0341_),
    .A1(net1126),
    .A2(net935));
 sg13g2_nand2_1 _5907_ (.Y(_2607_),
    .A(net1342),
    .B(net935));
 sg13g2_o21ai_1 _5908_ (.B1(_2607_),
    .Y(_0342_),
    .A1(net1123),
    .A2(net935));
 sg13g2_nand2_1 _5909_ (.Y(_2608_),
    .A(net710),
    .B(net931));
 sg13g2_o21ai_1 _5910_ (.B1(_2608_),
    .Y(_0343_),
    .A1(net1122),
    .A2(net931));
 sg13g2_nand2_1 _5911_ (.Y(_2609_),
    .A(net1319),
    .B(net930));
 sg13g2_o21ai_1 _5912_ (.B1(_2609_),
    .Y(_0344_),
    .A1(net1118),
    .A2(net930));
 sg13g2_nand2_1 _5913_ (.Y(_2610_),
    .A(net1323),
    .B(net935));
 sg13g2_o21ai_1 _5914_ (.B1(_2610_),
    .Y(_0345_),
    .A1(net1115),
    .A2(net935));
 sg13g2_nand2_1 _5915_ (.Y(_2611_),
    .A(net1328),
    .B(net932));
 sg13g2_o21ai_1 _5916_ (.B1(_2611_),
    .Y(_0346_),
    .A1(net1111),
    .A2(net932));
 sg13g2_nand2_1 _5917_ (.Y(_2612_),
    .A(net779),
    .B(net933));
 sg13g2_o21ai_1 _5918_ (.B1(_2612_),
    .Y(_0347_),
    .A1(net1108),
    .A2(net933));
 sg13g2_nand2_1 _5919_ (.Y(_2613_),
    .A(net707),
    .B(net933));
 sg13g2_o21ai_1 _5920_ (.B1(_2613_),
    .Y(_0348_),
    .A1(net1105),
    .A2(net933));
 sg13g2_nand2_1 _5921_ (.Y(_2614_),
    .A(net755),
    .B(net934));
 sg13g2_o21ai_1 _5922_ (.B1(_2614_),
    .Y(_0349_),
    .A1(net1102),
    .A2(net934));
 sg13g2_nand2_1 _5923_ (.Y(_2615_),
    .A(net683),
    .B(net934));
 sg13g2_o21ai_1 _5924_ (.B1(_2615_),
    .Y(_0350_),
    .A1(net1099),
    .A2(net934));
 sg13g2_nand2_1 _5925_ (.Y(_2616_),
    .A(net685),
    .B(net930));
 sg13g2_o21ai_1 _5926_ (.B1(_2616_),
    .Y(_0351_),
    .A1(net1096),
    .A2(net930));
 sg13g2_nand2_1 _5927_ (.Y(_2617_),
    .A(net1387),
    .B(net932));
 sg13g2_o21ai_1 _5928_ (.B1(_2617_),
    .Y(_0352_),
    .A1(net1093),
    .A2(net932));
 sg13g2_or2_1 _5929_ (.X(_2618_),
    .B(_2554_),
    .A(_2532_));
 sg13g2_nand2_1 _5930_ (.Y(_2619_),
    .A(net760),
    .B(net929));
 sg13g2_o21ai_1 _5931_ (.B1(_2619_),
    .Y(_0353_),
    .A1(net1151),
    .A2(net929));
 sg13g2_nand2_1 _5932_ (.Y(_2620_),
    .A(net773),
    .B(net928));
 sg13g2_o21ai_1 _5933_ (.B1(_2620_),
    .Y(_0354_),
    .A1(net1148),
    .A2(net929));
 sg13g2_nand2_1 _5934_ (.Y(_2621_),
    .A(net1318),
    .B(net928));
 sg13g2_o21ai_1 _5935_ (.B1(_2621_),
    .Y(_0355_),
    .A1(net1144),
    .A2(net928));
 sg13g2_nand2_1 _5936_ (.Y(_2622_),
    .A(net671),
    .B(net929));
 sg13g2_o21ai_1 _5937_ (.B1(_2622_),
    .Y(_0356_),
    .A1(net1141),
    .A2(net928));
 sg13g2_nand2_1 _5938_ (.Y(_2623_),
    .A(net692),
    .B(net926));
 sg13g2_o21ai_1 _5939_ (.B1(_2623_),
    .Y(_0357_),
    .A1(net1138),
    .A2(net926));
 sg13g2_nand2_1 _5940_ (.Y(_2624_),
    .A(net650),
    .B(net924));
 sg13g2_o21ai_1 _5941_ (.B1(_2624_),
    .Y(_0358_),
    .A1(net1135),
    .A2(net924));
 sg13g2_nand2_1 _5942_ (.Y(_2625_),
    .A(net1282),
    .B(net924));
 sg13g2_o21ai_1 _5943_ (.B1(_2625_),
    .Y(_0359_),
    .A1(net1132),
    .A2(net924));
 sg13g2_nand2_1 _5944_ (.Y(_2626_),
    .A(net1298),
    .B(net925));
 sg13g2_o21ai_1 _5945_ (.B1(_2626_),
    .Y(_0360_),
    .A1(net1129),
    .A2(net925));
 sg13g2_nand2_1 _5946_ (.Y(_2627_),
    .A(net670),
    .B(net927));
 sg13g2_o21ai_1 _5947_ (.B1(_2627_),
    .Y(_0361_),
    .A1(net1127),
    .A2(net927));
 sg13g2_nand2_1 _5948_ (.Y(_2628_),
    .A(net742),
    .B(net927));
 sg13g2_o21ai_1 _5949_ (.B1(_2628_),
    .Y(_0362_),
    .A1(net1123),
    .A2(net927));
 sg13g2_nand2_1 _5950_ (.Y(_2629_),
    .A(net1344),
    .B(net925));
 sg13g2_o21ai_1 _5951_ (.B1(_2629_),
    .Y(_0363_),
    .A1(net1120),
    .A2(net925));
 sg13g2_nand2_1 _5952_ (.Y(_2630_),
    .A(net824),
    .B(net924));
 sg13g2_o21ai_1 _5953_ (.B1(_2630_),
    .Y(_0364_),
    .A1(net1117),
    .A2(net924));
 sg13g2_nand2_1 _5954_ (.Y(_2631_),
    .A(net1333),
    .B(net926));
 sg13g2_o21ai_1 _5955_ (.B1(_2631_),
    .Y(_0365_),
    .A1(net1116),
    .A2(net926));
 sg13g2_nand2_1 _5956_ (.Y(_2632_),
    .A(net698),
    .B(net927));
 sg13g2_o21ai_1 _5957_ (.B1(_2632_),
    .Y(_0366_),
    .A1(net1111),
    .A2(net927));
 sg13g2_nand2_1 _5958_ (.Y(_2633_),
    .A(net1366),
    .B(net928));
 sg13g2_o21ai_1 _5959_ (.B1(_2633_),
    .Y(_0367_),
    .A1(net1110),
    .A2(net928));
 sg13g2_nand2_1 _5960_ (.Y(_2634_),
    .A(net840),
    .B(net927));
 sg13g2_o21ai_1 _5961_ (.B1(_2634_),
    .Y(_0368_),
    .A1(net1105),
    .A2(net927));
 sg13g2_nand2_1 _5962_ (.Y(_2635_),
    .A(net830),
    .B(net928));
 sg13g2_o21ai_1 _5963_ (.B1(_2635_),
    .Y(_0369_),
    .A1(net1103),
    .A2(net928));
 sg13g2_nand2_1 _5964_ (.Y(_2636_),
    .A(net804),
    .B(net929));
 sg13g2_o21ai_1 _5965_ (.B1(_2636_),
    .Y(_0370_),
    .A1(net1100),
    .A2(net929));
 sg13g2_nand2_1 _5966_ (.Y(_2637_),
    .A(net700),
    .B(net924));
 sg13g2_o21ai_1 _5967_ (.B1(_2637_),
    .Y(_0371_),
    .A1(net1098),
    .A2(net924));
 sg13g2_nand2_1 _5968_ (.Y(_2638_),
    .A(net714),
    .B(net926));
 sg13g2_o21ai_1 _5969_ (.B1(_2638_),
    .Y(_0372_),
    .A1(net1093),
    .A2(net926));
 sg13g2_nand2b_1 _5970_ (.Y(_2639_),
    .B(_0787_),
    .A_N(_0793_));
 sg13g2_or2_1 _5971_ (.X(_2640_),
    .B(_2639_),
    .A(_2464_));
 sg13g2_nand2_1 _5972_ (.Y(_2641_),
    .A(net1317),
    .B(net923));
 sg13g2_o21ai_1 _5973_ (.B1(_2641_),
    .Y(_0373_),
    .A1(net1151),
    .A2(net923));
 sg13g2_nand2_1 _5974_ (.Y(_2642_),
    .A(net688),
    .B(net920));
 sg13g2_o21ai_1 _5975_ (.B1(_2642_),
    .Y(_0374_),
    .A1(net1147),
    .A2(net920));
 sg13g2_nand2_1 _5976_ (.Y(_2643_),
    .A(net672),
    .B(net921));
 sg13g2_o21ai_1 _5977_ (.B1(_2643_),
    .Y(_0375_),
    .A1(_2280_),
    .A2(net921));
 sg13g2_nand2_1 _5978_ (.Y(_2644_),
    .A(net802),
    .B(net922));
 sg13g2_o21ai_1 _5979_ (.B1(_2644_),
    .Y(_0376_),
    .A1(net1143),
    .A2(net922));
 sg13g2_nand2_1 _5980_ (.Y(_2645_),
    .A(net788),
    .B(net919));
 sg13g2_o21ai_1 _5981_ (.B1(_2645_),
    .Y(_0377_),
    .A1(net1140),
    .A2(net919));
 sg13g2_nand2_1 _5982_ (.Y(_2646_),
    .A(net792),
    .B(net917));
 sg13g2_o21ai_1 _5983_ (.B1(_2646_),
    .Y(_0378_),
    .A1(net1135),
    .A2(net917));
 sg13g2_nand2_1 _5984_ (.Y(_2647_),
    .A(net787),
    .B(net917));
 sg13g2_o21ai_1 _5985_ (.B1(_2647_),
    .Y(_0379_),
    .A1(net1133),
    .A2(net917));
 sg13g2_nand2_1 _5986_ (.Y(_2648_),
    .A(net649),
    .B(net918));
 sg13g2_o21ai_1 _5987_ (.B1(_2648_),
    .Y(_0380_),
    .A1(net1129),
    .A2(net918));
 sg13g2_nand2_1 _5988_ (.Y(_2649_),
    .A(net1294),
    .B(net920));
 sg13g2_o21ai_1 _5989_ (.B1(_2649_),
    .Y(_0381_),
    .A1(net1126),
    .A2(net920));
 sg13g2_nand2_1 _5990_ (.Y(_2650_),
    .A(net766),
    .B(net920));
 sg13g2_o21ai_1 _5991_ (.B1(_2650_),
    .Y(_0382_),
    .A1(net1124),
    .A2(net920));
 sg13g2_nand2_1 _5992_ (.Y(_2651_),
    .A(net723),
    .B(net918));
 sg13g2_o21ai_1 _5993_ (.B1(_2651_),
    .Y(_0383_),
    .A1(net1120),
    .A2(net918));
 sg13g2_nand2_1 _5994_ (.Y(_2652_),
    .A(net717),
    .B(net917));
 sg13g2_o21ai_1 _5995_ (.B1(_2652_),
    .Y(_0384_),
    .A1(net1117),
    .A2(net917));
 sg13g2_nand2_1 _5996_ (.Y(_2653_),
    .A(net719),
    .B(net920));
 sg13g2_o21ai_1 _5997_ (.B1(_2653_),
    .Y(_0385_),
    .A1(net1116),
    .A2(net923));
 sg13g2_nand2_1 _5998_ (.Y(_2654_),
    .A(net690),
    .B(net920));
 sg13g2_o21ai_1 _5999_ (.B1(_2654_),
    .Y(_0386_),
    .A1(net1113),
    .A2(net919));
 sg13g2_nand2_1 _6000_ (.Y(_2655_),
    .A(net1343),
    .B(net921));
 sg13g2_o21ai_1 _6001_ (.B1(_2655_),
    .Y(_0387_),
    .A1(net1109),
    .A2(net921));
 sg13g2_nand2_1 _6002_ (.Y(_2656_),
    .A(net808),
    .B(net921));
 sg13g2_o21ai_1 _6003_ (.B1(_2656_),
    .Y(_0388_),
    .A1(net1106),
    .A2(net921));
 sg13g2_nand2_1 _6004_ (.Y(_2657_),
    .A(net718),
    .B(net921));
 sg13g2_o21ai_1 _6005_ (.B1(_2657_),
    .Y(_0389_),
    .A1(net1103),
    .A2(net921));
 sg13g2_nand2_1 _6006_ (.Y(_2658_),
    .A(net778),
    .B(net922));
 sg13g2_o21ai_1 _6007_ (.B1(_2658_),
    .Y(_0390_),
    .A1(net1099),
    .A2(net922));
 sg13g2_nand2_1 _6008_ (.Y(_2659_),
    .A(net1289),
    .B(net917));
 sg13g2_o21ai_1 _6009_ (.B1(_2659_),
    .Y(_0391_),
    .A1(net1098),
    .A2(net917));
 sg13g2_nand2_1 _6010_ (.Y(_2660_),
    .A(net1322),
    .B(net919));
 sg13g2_o21ai_1 _6011_ (.B1(_2660_),
    .Y(_0392_),
    .A1(net1093),
    .A2(net919));
 sg13g2_or2_1 _6012_ (.X(_2661_),
    .B(_2639_),
    .A(_2487_));
 sg13g2_nand2_1 _6013_ (.Y(_2662_),
    .A(net1290),
    .B(net916));
 sg13g2_o21ai_1 _6014_ (.B1(_2662_),
    .Y(_0393_),
    .A1(net1150),
    .A2(net916));
 sg13g2_nand2_1 _6015_ (.Y(_2663_),
    .A(net666),
    .B(net914));
 sg13g2_o21ai_1 _6016_ (.B1(_2663_),
    .Y(_0394_),
    .A1(net1147),
    .A2(net915));
 sg13g2_nand2_1 _6017_ (.Y(_2664_),
    .A(net1380),
    .B(net914));
 sg13g2_o21ai_1 _6018_ (.B1(_2664_),
    .Y(_0395_),
    .A1(net1146),
    .A2(net914));
 sg13g2_nand2_1 _6019_ (.Y(_2665_),
    .A(net816),
    .B(net915));
 sg13g2_o21ai_1 _6020_ (.B1(_2665_),
    .Y(_0396_),
    .A1(net1141),
    .A2(net915));
 sg13g2_nand2_1 _6021_ (.Y(_2666_),
    .A(net733),
    .B(net913));
 sg13g2_o21ai_1 _6022_ (.B1(_2666_),
    .Y(_0397_),
    .A1(net1139),
    .A2(net913));
 sg13g2_nand2_1 _6023_ (.Y(_2667_),
    .A(net1305),
    .B(net911));
 sg13g2_o21ai_1 _6024_ (.B1(_2667_),
    .Y(_0398_),
    .A1(net1136),
    .A2(net911));
 sg13g2_nand2_1 _6025_ (.Y(_2668_),
    .A(net775),
    .B(net911));
 sg13g2_o21ai_1 _6026_ (.B1(_2668_),
    .Y(_0399_),
    .A1(net1133),
    .A2(net911));
 sg13g2_nand2_1 _6027_ (.Y(_2669_),
    .A(net776),
    .B(net912));
 sg13g2_o21ai_1 _6028_ (.B1(_2669_),
    .Y(_0400_),
    .A1(net1131),
    .A2(net912));
 sg13g2_nand2_1 _6029_ (.Y(_2670_),
    .A(net684),
    .B(net916));
 sg13g2_o21ai_1 _6030_ (.B1(_2670_),
    .Y(_0401_),
    .A1(net1127),
    .A2(net916));
 sg13g2_nand2_1 _6031_ (.Y(_2671_),
    .A(net655),
    .B(net916));
 sg13g2_o21ai_1 _6032_ (.B1(_2671_),
    .Y(_0402_),
    .A1(net1125),
    .A2(net916));
 sg13g2_nand2_1 _6033_ (.Y(_2672_),
    .A(net677),
    .B(net912));
 sg13g2_o21ai_1 _6034_ (.B1(_2672_),
    .Y(_0403_),
    .A1(net1122),
    .A2(net912));
 sg13g2_nand2_1 _6035_ (.Y(_2673_),
    .A(net841),
    .B(net911));
 sg13g2_o21ai_1 _6036_ (.B1(_2673_),
    .Y(_0404_),
    .A1(net1118),
    .A2(net911));
 sg13g2_nand2_1 _6037_ (.Y(_2674_),
    .A(net661),
    .B(net913));
 sg13g2_o21ai_1 _6038_ (.B1(_2674_),
    .Y(_0405_),
    .A1(net1114),
    .A2(net913));
 sg13g2_nand2_1 _6039_ (.Y(_2675_),
    .A(net652),
    .B(net913));
 sg13g2_o21ai_1 _6040_ (.B1(_2675_),
    .Y(_0406_),
    .A1(net1112),
    .A2(net913));
 sg13g2_nand2_1 _6041_ (.Y(_2676_),
    .A(net799),
    .B(net914));
 sg13g2_o21ai_1 _6042_ (.B1(_2676_),
    .Y(_0407_),
    .A1(net1108),
    .A2(net914));
 sg13g2_nand2_1 _6043_ (.Y(_2677_),
    .A(net709),
    .B(net914));
 sg13g2_o21ai_1 _6044_ (.B1(_2677_),
    .Y(_0408_),
    .A1(net1106),
    .A2(net914));
 sg13g2_nand2_1 _6045_ (.Y(_2678_),
    .A(net725),
    .B(net914));
 sg13g2_o21ai_1 _6046_ (.B1(_2678_),
    .Y(_0409_),
    .A1(net1103),
    .A2(net915));
 sg13g2_nand2_1 _6047_ (.Y(_2679_),
    .A(net659),
    .B(net915));
 sg13g2_o21ai_1 _6048_ (.B1(_2679_),
    .Y(_0410_),
    .A1(net1099),
    .A2(net915));
 sg13g2_nand2_1 _6049_ (.Y(_2680_),
    .A(net713),
    .B(net912));
 sg13g2_o21ai_1 _6050_ (.B1(_2680_),
    .Y(_0411_),
    .A1(net1098),
    .A2(net912));
 sg13g2_nand2_1 _6051_ (.Y(_2681_),
    .A(net815),
    .B(net911));
 sg13g2_o21ai_1 _6052_ (.B1(_2681_),
    .Y(_0412_),
    .A1(net1094),
    .A2(net911));
 sg13g2_or2_1 _6053_ (.X(_2682_),
    .B(_2639_),
    .A(_2510_));
 sg13g2_nand2_1 _6054_ (.Y(_2683_),
    .A(net1275),
    .B(net907));
 sg13g2_o21ai_1 _6055_ (.B1(_2683_),
    .Y(_0413_),
    .A1(net1150),
    .A2(net907));
 sg13g2_nand2_1 _6056_ (.Y(_2684_),
    .A(net1338),
    .B(net909));
 sg13g2_o21ai_1 _6057_ (.B1(_2684_),
    .Y(_0414_),
    .A1(net1149),
    .A2(net909));
 sg13g2_nand2_1 _6058_ (.Y(_2685_),
    .A(net660),
    .B(net908));
 sg13g2_o21ai_1 _6059_ (.B1(_2685_),
    .Y(_0415_),
    .A1(net1144),
    .A2(net908));
 sg13g2_nand2_1 _6060_ (.Y(_2686_),
    .A(net651),
    .B(net909));
 sg13g2_o21ai_1 _6061_ (.B1(_2686_),
    .Y(_0416_),
    .A1(net1143),
    .A2(net909));
 sg13g2_nand2_1 _6062_ (.Y(_2687_),
    .A(net708),
    .B(net906));
 sg13g2_o21ai_1 _6063_ (.B1(_2687_),
    .Y(_0417_),
    .A1(net1138),
    .A2(net906));
 sg13g2_nand2_1 _6064_ (.Y(_2688_),
    .A(net706),
    .B(net906));
 sg13g2_o21ai_1 _6065_ (.B1(_2688_),
    .Y(_0418_),
    .A1(net1136),
    .A2(_2682_));
 sg13g2_nand2_1 _6066_ (.Y(_2689_),
    .A(net774),
    .B(net905));
 sg13g2_o21ai_1 _6067_ (.B1(_2689_),
    .Y(_0419_),
    .A1(net1132),
    .A2(net905));
 sg13g2_nand2_1 _6068_ (.Y(_2690_),
    .A(net1316),
    .B(net905));
 sg13g2_o21ai_1 _6069_ (.B1(_2690_),
    .Y(_0420_),
    .A1(net1129),
    .A2(net905));
 sg13g2_nand2_1 _6070_ (.Y(_2691_),
    .A(net771),
    .B(net907));
 sg13g2_o21ai_1 _6071_ (.B1(_2691_),
    .Y(_0421_),
    .A1(net1126),
    .A2(net907));
 sg13g2_nand2_1 _6072_ (.Y(_2692_),
    .A(net811),
    .B(net907));
 sg13g2_o21ai_1 _6073_ (.B1(_2692_),
    .Y(_0422_),
    .A1(net1125),
    .A2(net907));
 sg13g2_nand2_1 _6074_ (.Y(_2693_),
    .A(net722),
    .B(net906));
 sg13g2_o21ai_1 _6075_ (.B1(_2693_),
    .Y(_0423_),
    .A1(net1120),
    .A2(net906));
 sg13g2_nand2_1 _6076_ (.Y(_2694_),
    .A(net1313),
    .B(net905));
 sg13g2_o21ai_1 _6077_ (.B1(_2694_),
    .Y(_0424_),
    .A1(net1117),
    .A2(net905));
 sg13g2_nand2_1 _6078_ (.Y(_2695_),
    .A(net1308),
    .B(net910));
 sg13g2_o21ai_1 _6079_ (.B1(_2695_),
    .Y(_0425_),
    .A1(net1115),
    .A2(net910));
 sg13g2_nand2_1 _6080_ (.Y(_2696_),
    .A(net828),
    .B(net907));
 sg13g2_o21ai_1 _6081_ (.B1(_2696_),
    .Y(_0426_),
    .A1(net1111),
    .A2(net907));
 sg13g2_nand2_1 _6082_ (.Y(_2697_),
    .A(net741),
    .B(net908));
 sg13g2_o21ai_1 _6083_ (.B1(_2697_),
    .Y(_0427_),
    .A1(net1108),
    .A2(net908));
 sg13g2_nand2_1 _6084_ (.Y(_2698_),
    .A(net743),
    .B(net908));
 sg13g2_o21ai_1 _6085_ (.B1(_2698_),
    .Y(_0428_),
    .A1(net1107),
    .A2(net908));
 sg13g2_nand2_1 _6086_ (.Y(_2699_),
    .A(net751),
    .B(net909));
 sg13g2_o21ai_1 _6087_ (.B1(_2699_),
    .Y(_0429_),
    .A1(net1102),
    .A2(net909));
 sg13g2_nand2_1 _6088_ (.Y(_2700_),
    .A(net746),
    .B(net908));
 sg13g2_o21ai_1 _6089_ (.B1(_2700_),
    .Y(_0430_),
    .A1(net1101),
    .A2(net908));
 sg13g2_nand2_1 _6090_ (.Y(_2701_),
    .A(net826),
    .B(net905));
 sg13g2_o21ai_1 _6091_ (.B1(_2701_),
    .Y(_0431_),
    .A1(net1098),
    .A2(net905));
 sg13g2_nand2_1 _6092_ (.Y(_2702_),
    .A(net1283),
    .B(net906));
 sg13g2_o21ai_1 _6093_ (.B1(_2702_),
    .Y(_0432_),
    .A1(net1093),
    .A2(net906));
 sg13g2_or2_1 _6094_ (.X(_2703_),
    .B(_2639_),
    .A(_2532_));
 sg13g2_nand2_1 _6095_ (.Y(_2704_),
    .A(net783),
    .B(net901));
 sg13g2_o21ai_1 _6096_ (.B1(_2704_),
    .Y(_0433_),
    .A1(net1150),
    .A2(net901));
 sg13g2_nand2_1 _6097_ (.Y(_2705_),
    .A(net831),
    .B(net901));
 sg13g2_o21ai_1 _6098_ (.B1(_2705_),
    .Y(_0434_),
    .A1(net1147),
    .A2(net901));
 sg13g2_nand2_1 _6099_ (.Y(_2706_),
    .A(net1310),
    .B(net902));
 sg13g2_o21ai_1 _6100_ (.B1(_2706_),
    .Y(_0435_),
    .A1(net1146),
    .A2(net902));
 sg13g2_nand2_1 _6101_ (.Y(_2707_),
    .A(net1292),
    .B(net902));
 sg13g2_o21ai_1 _6102_ (.B1(_2707_),
    .Y(_0436_),
    .A1(net1141),
    .A2(net902));
 sg13g2_nand2_1 _6103_ (.Y(_2708_),
    .A(net731),
    .B(net904));
 sg13g2_o21ai_1 _6104_ (.B1(_2708_),
    .Y(_0437_),
    .A1(net1138),
    .A2(net904));
 sg13g2_nand2_1 _6105_ (.Y(_2709_),
    .A(net763),
    .B(net899));
 sg13g2_o21ai_1 _6106_ (.B1(_2709_),
    .Y(_0438_),
    .A1(net1135),
    .A2(net899));
 sg13g2_nand2_1 _6107_ (.Y(_2710_),
    .A(net676),
    .B(net898));
 sg13g2_o21ai_1 _6108_ (.B1(_2710_),
    .Y(_0439_),
    .A1(net1132),
    .A2(net898));
 sg13g2_nand2_1 _6109_ (.Y(_2711_),
    .A(net836),
    .B(net899));
 sg13g2_o21ai_1 _6110_ (.B1(_2711_),
    .Y(_0440_),
    .A1(net1131),
    .A2(net899));
 sg13g2_nand2_1 _6111_ (.Y(_2712_),
    .A(net832),
    .B(net901));
 sg13g2_o21ai_1 _6112_ (.B1(_2712_),
    .Y(_0441_),
    .A1(net1127),
    .A2(net901));
 sg13g2_nand2_1 _6113_ (.Y(_2713_),
    .A(net729),
    .B(net901));
 sg13g2_o21ai_1 _6114_ (.B1(_2713_),
    .Y(_0442_),
    .A1(net1124),
    .A2(net901));
 sg13g2_nand2_1 _6115_ (.Y(_2714_),
    .A(net823),
    .B(net898));
 sg13g2_o21ai_1 _6116_ (.B1(_2714_),
    .Y(_0443_),
    .A1(net1120),
    .A2(net898));
 sg13g2_nand2_1 _6117_ (.Y(_2715_),
    .A(net681),
    .B(net898));
 sg13g2_o21ai_1 _6118_ (.B1(_2715_),
    .Y(_0444_),
    .A1(net1117),
    .A2(net898));
 sg13g2_nand2_1 _6119_ (.Y(_2716_),
    .A(net695),
    .B(net900));
 sg13g2_o21ai_1 _6120_ (.B1(_2716_),
    .Y(_0445_),
    .A1(net1114),
    .A2(net900));
 sg13g2_nand2_1 _6121_ (.Y(_2717_),
    .A(net691),
    .B(net900));
 sg13g2_o21ai_1 _6122_ (.B1(_2717_),
    .Y(_0446_),
    .A1(net1112),
    .A2(net900));
 sg13g2_nand2_1 _6123_ (.Y(_2718_),
    .A(net1321),
    .B(net902));
 sg13g2_o21ai_1 _6124_ (.B1(_2718_),
    .Y(_0447_),
    .A1(net1110),
    .A2(net902));
 sg13g2_nand2_1 _6125_ (.Y(_2719_),
    .A(net772),
    .B(net903));
 sg13g2_o21ai_1 _6126_ (.B1(_2719_),
    .Y(_0448_),
    .A1(net1105),
    .A2(net903));
 sg13g2_nand2_1 _6127_ (.Y(_2720_),
    .A(net1371),
    .B(net902));
 sg13g2_o21ai_1 _6128_ (.B1(_2720_),
    .Y(_0449_),
    .A1(net1103),
    .A2(net902));
 sg13g2_nand2_1 _6129_ (.Y(_2721_),
    .A(net1278),
    .B(net903));
 sg13g2_o21ai_1 _6130_ (.B1(_2721_),
    .Y(_0450_),
    .A1(net1100),
    .A2(net903));
 sg13g2_nand2_1 _6131_ (.Y(_2722_),
    .A(net682),
    .B(net898));
 sg13g2_o21ai_1 _6132_ (.B1(_2722_),
    .Y(_0451_),
    .A1(net1098),
    .A2(net898));
 sg13g2_nand2_1 _6133_ (.Y(_2723_),
    .A(net701),
    .B(net900));
 sg13g2_o21ai_1 _6134_ (.B1(_2723_),
    .Y(_0452_),
    .A1(net1095),
    .A2(net900));
 sg13g2_nand2_1 _6135_ (.Y(_2724_),
    .A(_0787_),
    .B(_0793_));
 sg13g2_or2_1 _6136_ (.X(_2725_),
    .B(_2724_),
    .A(_2464_));
 sg13g2_nand2_1 _6137_ (.Y(_2726_),
    .A(net664),
    .B(net896));
 sg13g2_o21ai_1 _6138_ (.B1(_2726_),
    .Y(_0453_),
    .A1(net1152),
    .A2(net896));
 sg13g2_nand2_1 _6139_ (.Y(_2727_),
    .A(net712),
    .B(net895));
 sg13g2_o21ai_1 _6140_ (.B1(_2727_),
    .Y(_0454_),
    .A1(net1147),
    .A2(net895));
 sg13g2_nand2_1 _6141_ (.Y(_2728_),
    .A(net724),
    .B(net894));
 sg13g2_o21ai_1 _6142_ (.B1(_2728_),
    .Y(_0455_),
    .A1(net1144),
    .A2(net894));
 sg13g2_nand2_1 _6143_ (.Y(_2729_),
    .A(net693),
    .B(net895));
 sg13g2_o21ai_1 _6144_ (.B1(_2729_),
    .Y(_0456_),
    .A1(net1143),
    .A2(net895));
 sg13g2_nand2_1 _6145_ (.Y(_2730_),
    .A(net657),
    .B(net893));
 sg13g2_o21ai_1 _6146_ (.B1(_2730_),
    .Y(_0457_),
    .A1(net1139),
    .A2(net893));
 sg13g2_nand2_1 _6147_ (.Y(_2731_),
    .A(net800),
    .B(net891));
 sg13g2_o21ai_1 _6148_ (.B1(_2731_),
    .Y(_0458_),
    .A1(net1135),
    .A2(net891));
 sg13g2_nand2_1 _6149_ (.Y(_2732_),
    .A(net732),
    .B(net891));
 sg13g2_o21ai_1 _6150_ (.B1(_2732_),
    .Y(_0459_),
    .A1(net1132),
    .A2(net891));
 sg13g2_nand2_1 _6151_ (.Y(_2733_),
    .A(net1309),
    .B(net891));
 sg13g2_o21ai_1 _6152_ (.B1(_2733_),
    .Y(_0460_),
    .A1(net1130),
    .A2(net891));
 sg13g2_nand2_1 _6153_ (.Y(_2734_),
    .A(net796),
    .B(net894));
 sg13g2_o21ai_1 _6154_ (.B1(_2734_),
    .Y(_0461_),
    .A1(net1126),
    .A2(net894));
 sg13g2_nand2_1 _6155_ (.Y(_2735_),
    .A(net827),
    .B(net896));
 sg13g2_o21ai_1 _6156_ (.B1(_2735_),
    .Y(_0462_),
    .A1(net1124),
    .A2(net896));
 sg13g2_nand2_1 _6157_ (.Y(_2736_),
    .A(net726),
    .B(net892));
 sg13g2_o21ai_1 _6158_ (.B1(_2736_),
    .Y(_0463_),
    .A1(net1121),
    .A2(net892));
 sg13g2_nand2_1 _6159_ (.Y(_2737_),
    .A(net679),
    .B(net892));
 sg13g2_o21ai_1 _6160_ (.B1(_2737_),
    .Y(_0464_),
    .A1(net1119),
    .A2(net892));
 sg13g2_nand2_1 _6161_ (.Y(_2738_),
    .A(net820),
    .B(net896));
 sg13g2_o21ai_1 _6162_ (.B1(_2738_),
    .Y(_0465_),
    .A1(net1115),
    .A2(net896));
 sg13g2_nand2_1 _6163_ (.Y(_2739_),
    .A(net705),
    .B(net896));
 sg13g2_o21ai_1 _6164_ (.B1(_2739_),
    .Y(_0466_),
    .A1(net1113),
    .A2(net896));
 sg13g2_nand2_1 _6165_ (.Y(_2740_),
    .A(net768),
    .B(net894));
 sg13g2_o21ai_1 _6166_ (.B1(_2740_),
    .Y(_0467_),
    .A1(net1108),
    .A2(net894));
 sg13g2_nand2_1 _6167_ (.Y(_2741_),
    .A(net1301),
    .B(net894));
 sg13g2_o21ai_1 _6168_ (.B1(_2741_),
    .Y(_0468_),
    .A1(net1105),
    .A2(net894));
 sg13g2_nand2_1 _6169_ (.Y(_2742_),
    .A(net762),
    .B(net895));
 sg13g2_o21ai_1 _6170_ (.B1(_2742_),
    .Y(_0469_),
    .A1(net1102),
    .A2(net895));
 sg13g2_nand2_1 _6171_ (.Y(_2743_),
    .A(net829),
    .B(net895));
 sg13g2_o21ai_1 _6172_ (.B1(_2743_),
    .Y(_0470_),
    .A1(net1099),
    .A2(net895));
 sg13g2_nand2_1 _6173_ (.Y(_2744_),
    .A(net805),
    .B(net891));
 sg13g2_o21ai_1 _6174_ (.B1(_2744_),
    .Y(_0471_),
    .A1(net1096),
    .A2(net891));
 sg13g2_nand2_1 _6175_ (.Y(_2745_),
    .A(net1273),
    .B(net893));
 sg13g2_o21ai_1 _6176_ (.B1(_2745_),
    .Y(_0472_),
    .A1(net1095),
    .A2(net893));
 sg13g2_or2_1 _6177_ (.X(_2746_),
    .B(_2724_),
    .A(_2487_));
 sg13g2_nand2_1 _6178_ (.Y(_2747_),
    .A(net752),
    .B(net889));
 sg13g2_o21ai_1 _6179_ (.B1(_2747_),
    .Y(_0473_),
    .A1(net1152),
    .A2(net889));
 sg13g2_nand2_1 _6180_ (.Y(_2748_),
    .A(net662),
    .B(net886));
 sg13g2_o21ai_1 _6181_ (.B1(_2748_),
    .Y(_0474_),
    .A1(net1147),
    .A2(net886));
 sg13g2_nand2_1 _6182_ (.Y(_2749_),
    .A(net764),
    .B(net887));
 sg13g2_o21ai_1 _6183_ (.B1(_2749_),
    .Y(_0475_),
    .A1(net1144),
    .A2(net887));
 sg13g2_nand2_1 _6184_ (.Y(_2750_),
    .A(net1330),
    .B(net888));
 sg13g2_o21ai_1 _6185_ (.B1(_2750_),
    .Y(_0476_),
    .A1(net1141),
    .A2(net888));
 sg13g2_nand2_1 _6186_ (.Y(_2751_),
    .A(net653),
    .B(net890));
 sg13g2_o21ai_1 _6187_ (.B1(_2751_),
    .Y(_0477_),
    .A1(net1140),
    .A2(net890));
 sg13g2_nand2_1 _6188_ (.Y(_2752_),
    .A(net754),
    .B(net884));
 sg13g2_o21ai_1 _6189_ (.B1(_2752_),
    .Y(_0478_),
    .A1(net1135),
    .A2(net884));
 sg13g2_nand2_1 _6190_ (.Y(_2753_),
    .A(net806),
    .B(net885));
 sg13g2_o21ai_1 _6191_ (.B1(_2753_),
    .Y(_0479_),
    .A1(net1134),
    .A2(net890));
 sg13g2_nand2_1 _6192_ (.Y(_2754_),
    .A(net1329),
    .B(net884));
 sg13g2_o21ai_1 _6193_ (.B1(_2754_),
    .Y(_0480_),
    .A1(net1129),
    .A2(net884));
 sg13g2_nand2_1 _6194_ (.Y(_2755_),
    .A(net814),
    .B(net886));
 sg13g2_o21ai_1 _6195_ (.B1(_2755_),
    .Y(_0481_),
    .A1(net1126),
    .A2(net886));
 sg13g2_nand2_1 _6196_ (.Y(_2756_),
    .A(net1276),
    .B(net886));
 sg13g2_o21ai_1 _6197_ (.B1(_2756_),
    .Y(_0482_),
    .A1(net1123),
    .A2(net886));
 sg13g2_nand2_1 _6198_ (.Y(_2757_),
    .A(net817),
    .B(net885));
 sg13g2_o21ai_1 _6199_ (.B1(_2757_),
    .Y(_0483_),
    .A1(net1120),
    .A2(net885));
 sg13g2_nand2_1 _6200_ (.Y(_2758_),
    .A(net1354),
    .B(net884));
 sg13g2_o21ai_1 _6201_ (.B1(_2758_),
    .Y(_0484_),
    .A1(net1117),
    .A2(net884));
 sg13g2_nand2_1 _6202_ (.Y(_2759_),
    .A(net704),
    .B(net886));
 sg13g2_o21ai_1 _6203_ (.B1(_2759_),
    .Y(_0485_),
    .A1(net1114),
    .A2(net885));
 sg13g2_nand2_1 _6204_ (.Y(_2760_),
    .A(net780),
    .B(net886));
 sg13g2_o21ai_1 _6205_ (.B1(_2760_),
    .Y(_0486_),
    .A1(net1111),
    .A2(net885));
 sg13g2_nand2_1 _6206_ (.Y(_2761_),
    .A(net1277),
    .B(net887));
 sg13g2_o21ai_1 _6207_ (.B1(_2761_),
    .Y(_0487_),
    .A1(net1109),
    .A2(net887));
 sg13g2_nand2_1 _6208_ (.Y(_2762_),
    .A(net689),
    .B(net887));
 sg13g2_o21ai_1 _6209_ (.B1(_2762_),
    .Y(_0488_),
    .A1(net1105),
    .A2(net887));
 sg13g2_nand2_1 _6210_ (.Y(_2763_),
    .A(net669),
    .B(net887));
 sg13g2_o21ai_1 _6211_ (.B1(_2763_),
    .Y(_0489_),
    .A1(net1103),
    .A2(net887));
 sg13g2_nand2_1 _6212_ (.Y(_2764_),
    .A(net750),
    .B(net888));
 sg13g2_o21ai_1 _6213_ (.B1(_2764_),
    .Y(_0490_),
    .A1(net1099),
    .A2(net888));
 sg13g2_nand2_1 _6214_ (.Y(_2765_),
    .A(net784),
    .B(net884));
 sg13g2_o21ai_1 _6215_ (.B1(_2765_),
    .Y(_0491_),
    .A1(net1096),
    .A2(net884));
 sg13g2_nand2_1 _6216_ (.Y(_2766_),
    .A(net1358),
    .B(net885));
 sg13g2_o21ai_1 _6217_ (.B1(_2766_),
    .Y(_0492_),
    .A1(net1093),
    .A2(net885));
 sg13g2_or2_1 _6218_ (.X(_2767_),
    .B(_2724_),
    .A(_2510_));
 sg13g2_nand2_1 _6219_ (.Y(_2768_),
    .A(net1296),
    .B(net879));
 sg13g2_o21ai_1 _6220_ (.B1(_2768_),
    .Y(_0493_),
    .A1(net1150),
    .A2(net882));
 sg13g2_nand2_1 _6221_ (.Y(_2769_),
    .A(net1299),
    .B(net881));
 sg13g2_o21ai_1 _6222_ (.B1(_2769_),
    .Y(_0494_),
    .A1(net1149),
    .A2(net879));
 sg13g2_nand2_1 _6223_ (.Y(_2770_),
    .A(net1304),
    .B(net880));
 sg13g2_o21ai_1 _6224_ (.B1(_2770_),
    .Y(_0495_),
    .A1(net1145),
    .A2(net880));
 sg13g2_nand2_1 _6225_ (.Y(_2771_),
    .A(net1300),
    .B(net880));
 sg13g2_o21ai_1 _6226_ (.B1(_2771_),
    .Y(_0496_),
    .A1(net1143),
    .A2(net880));
 sg13g2_nand2_1 _6227_ (.Y(_2772_),
    .A(net749),
    .B(net883));
 sg13g2_o21ai_1 _6228_ (.B1(_2772_),
    .Y(_0497_),
    .A1(net1138),
    .A2(net883));
 sg13g2_nand2_1 _6229_ (.Y(_2773_),
    .A(net797),
    .B(net878));
 sg13g2_o21ai_1 _6230_ (.B1(_2773_),
    .Y(_0498_),
    .A1(net1137),
    .A2(net878));
 sg13g2_nand2_1 _6231_ (.Y(_2774_),
    .A(net1359),
    .B(net877));
 sg13g2_o21ai_1 _6232_ (.B1(_2774_),
    .Y(_0499_),
    .A1(net1132),
    .A2(net877));
 sg13g2_nand2_1 _6233_ (.Y(_2775_),
    .A(net1352),
    .B(net877));
 sg13g2_o21ai_1 _6234_ (.B1(_2775_),
    .Y(_0500_),
    .A1(net1129),
    .A2(net877));
 sg13g2_nand2_1 _6235_ (.Y(_2776_),
    .A(net781),
    .B(net879));
 sg13g2_o21ai_1 _6236_ (.B1(_2776_),
    .Y(_0501_),
    .A1(net1127),
    .A2(net879));
 sg13g2_nand2_1 _6237_ (.Y(_2777_),
    .A(net798),
    .B(net879));
 sg13g2_o21ai_1 _6238_ (.B1(_2777_),
    .Y(_0502_),
    .A1(net1123),
    .A2(net879));
 sg13g2_nand2_1 _6239_ (.Y(_2778_),
    .A(net786),
    .B(net878));
 sg13g2_o21ai_1 _6240_ (.B1(_2778_),
    .Y(_0503_),
    .A1(net1121),
    .A2(net878));
 sg13g2_nand2_1 _6241_ (.Y(_2779_),
    .A(net1312),
    .B(net877));
 sg13g2_o21ai_1 _6242_ (.B1(_2779_),
    .Y(_0504_),
    .A1(net1117),
    .A2(net877));
 sg13g2_nand2_1 _6243_ (.Y(_2780_),
    .A(net1372),
    .B(net878));
 sg13g2_o21ai_1 _6244_ (.B1(_2780_),
    .Y(_0505_),
    .A1(net1116),
    .A2(net878));
 sg13g2_nand2_1 _6245_ (.Y(_2781_),
    .A(net1295),
    .B(net879));
 sg13g2_o21ai_1 _6246_ (.B1(_2781_),
    .Y(_0506_),
    .A1(net1111),
    .A2(net879));
 sg13g2_nand2_1 _6247_ (.Y(_2782_),
    .A(net791),
    .B(net880));
 sg13g2_o21ai_1 _6248_ (.B1(_2782_),
    .Y(_0507_),
    .A1(net1110),
    .A2(net880));
 sg13g2_nand2_1 _6249_ (.Y(_2783_),
    .A(net1307),
    .B(net880));
 sg13g2_o21ai_1 _6250_ (.B1(_2783_),
    .Y(_0508_),
    .A1(net1105),
    .A2(net880));
 sg13g2_nand2_1 _6251_ (.Y(_2784_),
    .A(net1339),
    .B(net881));
 sg13g2_o21ai_1 _6252_ (.B1(_2784_),
    .Y(_0509_),
    .A1(net1104),
    .A2(net881));
 sg13g2_nand2_1 _6253_ (.Y(_2785_),
    .A(net813),
    .B(net881));
 sg13g2_o21ai_1 _6254_ (.B1(_2785_),
    .Y(_0510_),
    .A1(net1100),
    .A2(net881));
 sg13g2_nand2_1 _6255_ (.Y(_2786_),
    .A(net1350),
    .B(net877));
 sg13g2_o21ai_1 _6256_ (.B1(_2786_),
    .Y(_0511_),
    .A1(net1097),
    .A2(net877));
 sg13g2_nand2_1 _6257_ (.Y(_2787_),
    .A(net1297),
    .B(net878));
 sg13g2_o21ai_1 _6258_ (.B1(_2787_),
    .Y(_0512_),
    .A1(net1093),
    .A2(net883));
 sg13g2_or2_1 _6259_ (.X(_2788_),
    .B(_2724_),
    .A(_2532_));
 sg13g2_nand2_1 _6260_ (.Y(_2789_),
    .A(net758),
    .B(net873));
 sg13g2_o21ai_1 _6261_ (.B1(_2789_),
    .Y(_0513_),
    .A1(net1151),
    .A2(net873));
 sg13g2_nand2_1 _6262_ (.Y(_2790_),
    .A(net1335),
    .B(net876));
 sg13g2_o21ai_1 _6263_ (.B1(_2790_),
    .Y(_0514_),
    .A1(_2276_),
    .A2(net876));
 sg13g2_nand2_1 _6264_ (.Y(_2791_),
    .A(net1375),
    .B(net874));
 sg13g2_o21ai_1 _6265_ (.B1(_2791_),
    .Y(_0515_),
    .A1(net1145),
    .A2(net874));
 sg13g2_nand2_1 _6266_ (.Y(_2792_),
    .A(net735),
    .B(net874));
 sg13g2_o21ai_1 _6267_ (.B1(_2792_),
    .Y(_0516_),
    .A1(net1143),
    .A2(net874));
 sg13g2_nand2_1 _6268_ (.Y(_2793_),
    .A(net1364),
    .B(net872));
 sg13g2_o21ai_1 _6269_ (.B1(_2793_),
    .Y(_0517_),
    .A1(net1139),
    .A2(net872));
 sg13g2_nand2_1 _6270_ (.Y(_2794_),
    .A(net1349),
    .B(net870));
 sg13g2_o21ai_1 _6271_ (.B1(_2794_),
    .Y(_0518_),
    .A1(net1136),
    .A2(net870));
 sg13g2_nand2_1 _6272_ (.Y(_2795_),
    .A(net737),
    .B(net870));
 sg13g2_o21ai_1 _6273_ (.B1(_2795_),
    .Y(_0519_),
    .A1(net1132),
    .A2(net870));
 sg13g2_nand2_1 _6274_ (.Y(_2796_),
    .A(net1314),
    .B(net871));
 sg13g2_o21ai_1 _6275_ (.B1(_2796_),
    .Y(_0520_),
    .A1(net1130),
    .A2(net871));
 sg13g2_nand2_1 _6276_ (.Y(_2797_),
    .A(net715),
    .B(net873));
 sg13g2_o21ai_1 _6277_ (.B1(_2797_),
    .Y(_0521_),
    .A1(net1127),
    .A2(net873));
 sg13g2_nand2_1 _6278_ (.Y(_2798_),
    .A(net810),
    .B(net873));
 sg13g2_o21ai_1 _6279_ (.B1(_2798_),
    .Y(_0522_),
    .A1(net1124),
    .A2(net873));
 sg13g2_nand2_1 _6280_ (.Y(_2799_),
    .A(net674),
    .B(net871));
 sg13g2_o21ai_1 _6281_ (.B1(_2799_),
    .Y(_0523_),
    .A1(net1120),
    .A2(net871));
 sg13g2_nand2_1 _6282_ (.Y(_2800_),
    .A(net658),
    .B(net870));
 sg13g2_o21ai_1 _6283_ (.B1(_2800_),
    .Y(_0524_),
    .A1(net1117),
    .A2(net870));
 sg13g2_nand2_1 _6284_ (.Y(_2801_),
    .A(net1374),
    .B(net872));
 sg13g2_o21ai_1 _6285_ (.B1(_2801_),
    .Y(_0525_),
    .A1(net1114),
    .A2(net872));
 sg13g2_nand2_1 _6286_ (.Y(_2802_),
    .A(net803),
    .B(net873));
 sg13g2_o21ai_1 _6287_ (.B1(_2802_),
    .Y(_0526_),
    .A1(net1112),
    .A2(net873));
 sg13g2_nand2_1 _6288_ (.Y(_2803_),
    .A(net730),
    .B(net874));
 sg13g2_o21ai_1 _6289_ (.B1(_2803_),
    .Y(_0527_),
    .A1(net1110),
    .A2(net874));
 sg13g2_nand2_1 _6290_ (.Y(_2804_),
    .A(net1311),
    .B(net874));
 sg13g2_o21ai_1 _6291_ (.B1(_2804_),
    .Y(_0528_),
    .A1(net1106),
    .A2(net874));
 sg13g2_nand2_1 _6292_ (.Y(_2805_),
    .A(net769),
    .B(net875));
 sg13g2_o21ai_1 _6293_ (.B1(_2805_),
    .Y(_0529_),
    .A1(net1104),
    .A2(net875));
 sg13g2_nand2_1 _6294_ (.Y(_2806_),
    .A(net748),
    .B(net875));
 sg13g2_o21ai_1 _6295_ (.B1(_2806_),
    .Y(_0530_),
    .A1(net1100),
    .A2(net875));
 sg13g2_nand2_1 _6296_ (.Y(_2807_),
    .A(net782),
    .B(net870));
 sg13g2_o21ai_1 _6297_ (.B1(_2807_),
    .Y(_0531_),
    .A1(net1097),
    .A2(net870));
 sg13g2_nand2_1 _6298_ (.Y(_2808_),
    .A(net790),
    .B(net872));
 sg13g2_o21ai_1 _6299_ (.B1(_2808_),
    .Y(_0532_),
    .A1(net1094),
    .A2(net872));
 sg13g2_nor3_1 _6300_ (.A(_0816_),
    .B(_0830_),
    .C(_2267_),
    .Y(_2809_));
 sg13g2_nor2_1 _6301_ (.A(net1591),
    .B(net868),
    .Y(_2810_));
 sg13g2_a21oi_1 _6302_ (.A1(net1152),
    .A2(net868),
    .Y(_0533_),
    .B1(_2810_));
 sg13g2_nor2_1 _6303_ (.A(net1538),
    .B(net867),
    .Y(_2811_));
 sg13g2_a21oi_1 _6304_ (.A1(net1148),
    .A2(net867),
    .Y(_0534_),
    .B1(_2811_));
 sg13g2_nor2_1 _6305_ (.A(net1480),
    .B(net866),
    .Y(_2812_));
 sg13g2_a21oi_1 _6306_ (.A1(net1144),
    .A2(net866),
    .Y(_0535_),
    .B1(_2812_));
 sg13g2_nor2_1 _6307_ (.A(net1468),
    .B(net866),
    .Y(_2813_));
 sg13g2_a21oi_1 _6308_ (.A1(net1143),
    .A2(net866),
    .Y(_0536_),
    .B1(_2813_));
 sg13g2_nor2_1 _6309_ (.A(net1412),
    .B(net865),
    .Y(_2814_));
 sg13g2_a21oi_1 _6310_ (.A1(net1139),
    .A2(net865),
    .Y(_0537_),
    .B1(_2814_));
 sg13g2_nor2_1 _6311_ (.A(net1483),
    .B(net863),
    .Y(_2815_));
 sg13g2_a21oi_1 _6312_ (.A1(net1136),
    .A2(net863),
    .Y(_0538_),
    .B1(_2815_));
 sg13g2_nor2_1 _6313_ (.A(net1429),
    .B(net863),
    .Y(_2816_));
 sg13g2_a21oi_1 _6314_ (.A1(net1133),
    .A2(net863),
    .Y(_0539_),
    .B1(_2816_));
 sg13g2_nor2_1 _6315_ (.A(net1427),
    .B(net863),
    .Y(_2817_));
 sg13g2_a21oi_1 _6316_ (.A1(net1130),
    .A2(net863),
    .Y(_0540_),
    .B1(_2817_));
 sg13g2_nor2_1 _6317_ (.A(net1472),
    .B(net868),
    .Y(_2818_));
 sg13g2_a21oi_1 _6318_ (.A1(net1127),
    .A2(net868),
    .Y(_0541_),
    .B1(_2818_));
 sg13g2_nor2_1 _6319_ (.A(net1551),
    .B(net868),
    .Y(_2819_));
 sg13g2_a21oi_1 _6320_ (.A1(net1123),
    .A2(net868),
    .Y(_0542_),
    .B1(_2819_));
 sg13g2_nor2_1 _6321_ (.A(net1514),
    .B(net864),
    .Y(_2820_));
 sg13g2_a21oi_1 _6322_ (.A1(net1121),
    .A2(net864),
    .Y(_0543_),
    .B1(_2820_));
 sg13g2_nor2_1 _6323_ (.A(net1435),
    .B(net863),
    .Y(_2821_));
 sg13g2_a21oi_1 _6324_ (.A1(net1118),
    .A2(net863),
    .Y(_0544_),
    .B1(_2821_));
 sg13g2_nor2_1 _6325_ (.A(net1516),
    .B(net868),
    .Y(_2822_));
 sg13g2_a21oi_1 _6326_ (.A1(net1115),
    .A2(net868),
    .Y(_0545_),
    .B1(_2822_));
 sg13g2_nor2_1 _6327_ (.A(net1621),
    .B(net865),
    .Y(_2823_));
 sg13g2_a21oi_1 _6328_ (.A1(net1111),
    .A2(net865),
    .Y(_0546_),
    .B1(_2823_));
 sg13g2_nor2_1 _6329_ (.A(net1413),
    .B(net866),
    .Y(_2824_));
 sg13g2_a21oi_1 _6330_ (.A1(net1108),
    .A2(net866),
    .Y(_0547_),
    .B1(_2824_));
 sg13g2_nor2_1 _6331_ (.A(net1441),
    .B(net866),
    .Y(_2825_));
 sg13g2_a21oi_1 _6332_ (.A1(net1105),
    .A2(net866),
    .Y(_0548_),
    .B1(_2825_));
 sg13g2_nor2_1 _6333_ (.A(net1481),
    .B(net867),
    .Y(_2826_));
 sg13g2_a21oi_1 _6334_ (.A1(net1104),
    .A2(net867),
    .Y(_0549_),
    .B1(_2826_));
 sg13g2_nor2_1 _6335_ (.A(net1586),
    .B(net867),
    .Y(_2827_));
 sg13g2_a21oi_1 _6336_ (.A1(net1099),
    .A2(net867),
    .Y(_0550_),
    .B1(_2827_));
 sg13g2_nor2_1 _6337_ (.A(net1513),
    .B(net864),
    .Y(_2828_));
 sg13g2_a21oi_1 _6338_ (.A1(net1097),
    .A2(net864),
    .Y(_0551_),
    .B1(_2828_));
 sg13g2_nor2_1 _6339_ (.A(net1495),
    .B(net865),
    .Y(_2829_));
 sg13g2_a21oi_1 _6340_ (.A1(net1094),
    .A2(net865),
    .Y(_0552_),
    .B1(_2829_));
 sg13g2_nor2_2 _6341_ (.A(_2267_),
    .B(_2486_),
    .Y(_2830_));
 sg13g2_nor2_1 _6342_ (.A(net1450),
    .B(net862),
    .Y(_2831_));
 sg13g2_a21oi_1 _6343_ (.A1(net1150),
    .A2(net862),
    .Y(_0553_),
    .B1(_2831_));
 sg13g2_nor2_1 _6344_ (.A(net1470),
    .B(net862),
    .Y(_2832_));
 sg13g2_a21oi_1 _6345_ (.A1(net1147),
    .A2(net862),
    .Y(_0554_),
    .B1(_2832_));
 sg13g2_nor2_1 _6346_ (.A(net1415),
    .B(net860),
    .Y(_2833_));
 sg13g2_a21oi_1 _6347_ (.A1(net1144),
    .A2(net860),
    .Y(_0555_),
    .B1(_2833_));
 sg13g2_nor2_1 _6348_ (.A(net1574),
    .B(net860),
    .Y(_2834_));
 sg13g2_a21oi_1 _6349_ (.A1(net1141),
    .A2(net860),
    .Y(_0556_),
    .B1(_2834_));
 sg13g2_nor2_1 _6350_ (.A(net1400),
    .B(net857),
    .Y(_2835_));
 sg13g2_a21oi_1 _6351_ (.A1(net1139),
    .A2(net857),
    .Y(_0557_),
    .B1(_2835_));
 sg13g2_nor2_1 _6352_ (.A(net1409),
    .B(net856),
    .Y(_2836_));
 sg13g2_a21oi_1 _6353_ (.A1(net1136),
    .A2(net856),
    .Y(_0558_),
    .B1(_2836_));
 sg13g2_nor2_1 _6354_ (.A(net1617),
    .B(net856),
    .Y(_2837_));
 sg13g2_a21oi_1 _6355_ (.A1(net1134),
    .A2(net856),
    .Y(_0559_),
    .B1(_2837_));
 sg13g2_nor2_1 _6356_ (.A(net1401),
    .B(net856),
    .Y(_2838_));
 sg13g2_a21oi_1 _6357_ (.A1(net1131),
    .A2(net856),
    .Y(_0560_),
    .B1(_2838_));
 sg13g2_nor2_1 _6358_ (.A(net1474),
    .B(net862),
    .Y(_2839_));
 sg13g2_a21oi_1 _6359_ (.A1(net1127),
    .A2(net862),
    .Y(_0561_),
    .B1(_2839_));
 sg13g2_nor2_1 _6360_ (.A(net1557),
    .B(net859),
    .Y(_2840_));
 sg13g2_a21oi_1 _6361_ (.A1(_2308_),
    .A2(net859),
    .Y(_0562_),
    .B1(_2840_));
 sg13g2_nor2_1 _6362_ (.A(net1418),
    .B(net858),
    .Y(_2841_));
 sg13g2_a21oi_1 _6363_ (.A1(net1122),
    .A2(net858),
    .Y(_0563_),
    .B1(_2841_));
 sg13g2_nor2_1 _6364_ (.A(net1494),
    .B(net856),
    .Y(_2842_));
 sg13g2_a21oi_1 _6365_ (.A1(net1119),
    .A2(net856),
    .Y(_0564_),
    .B1(_2842_));
 sg13g2_nor2_1 _6366_ (.A(net1403),
    .B(net859),
    .Y(_2843_));
 sg13g2_a21oi_1 _6367_ (.A1(net1114),
    .A2(net859),
    .Y(_0565_),
    .B1(_2843_));
 sg13g2_nor2_1 _6368_ (.A(net1582),
    .B(net859),
    .Y(_2844_));
 sg13g2_a21oi_1 _6369_ (.A1(net1112),
    .A2(net859),
    .Y(_0566_),
    .B1(_2844_));
 sg13g2_nor2_1 _6370_ (.A(net1420),
    .B(net860),
    .Y(_2845_));
 sg13g2_a21oi_1 _6371_ (.A1(net1108),
    .A2(net860),
    .Y(_0567_),
    .B1(_2845_));
 sg13g2_nor2_1 _6372_ (.A(net1479),
    .B(net860),
    .Y(_2846_));
 sg13g2_a21oi_1 _6373_ (.A1(net1106),
    .A2(net860),
    .Y(_0568_),
    .B1(_2846_));
 sg13g2_nor2_1 _6374_ (.A(net1488),
    .B(net861),
    .Y(_2847_));
 sg13g2_a21oi_1 _6375_ (.A1(net1103),
    .A2(net861),
    .Y(_0569_),
    .B1(_2847_));
 sg13g2_nor2_1 _6376_ (.A(net1579),
    .B(net861),
    .Y(_2848_));
 sg13g2_a21oi_1 _6377_ (.A1(net1101),
    .A2(net861),
    .Y(_0570_),
    .B1(_2848_));
 sg13g2_nor2_1 _6378_ (.A(net1443),
    .B(net858),
    .Y(_2849_));
 sg13g2_a21oi_1 _6379_ (.A1(_2344_),
    .A2(net858),
    .Y(_0571_),
    .B1(_2849_));
 sg13g2_nor2_1 _6380_ (.A(net1476),
    .B(net857),
    .Y(_2850_));
 sg13g2_a21oi_1 _6381_ (.A1(net1094),
    .A2(net857),
    .Y(_0572_),
    .B1(_2850_));
 sg13g2_nor2_1 _6382_ (.A(_2267_),
    .B(_2509_),
    .Y(_2851_));
 sg13g2_nor2_1 _6383_ (.A(net1544),
    .B(net854),
    .Y(_2852_));
 sg13g2_a21oi_1 _6384_ (.A1(net1152),
    .A2(net854),
    .Y(_0573_),
    .B1(_2852_));
 sg13g2_nor2_1 _6385_ (.A(net1433),
    .B(net854),
    .Y(_2853_));
 sg13g2_a21oi_1 _6386_ (.A1(net1149),
    .A2(net854),
    .Y(_0574_),
    .B1(_2853_));
 sg13g2_nor2_1 _6387_ (.A(net1570),
    .B(net852),
    .Y(_2854_));
 sg13g2_a21oi_1 _6388_ (.A1(net1146),
    .A2(net852),
    .Y(_0575_),
    .B1(_2854_));
 sg13g2_nor2_1 _6389_ (.A(net1508),
    .B(net852),
    .Y(_2855_));
 sg13g2_a21oi_1 _6390_ (.A1(net1142),
    .A2(net852),
    .Y(_0576_),
    .B1(_2855_));
 sg13g2_nor2_1 _6391_ (.A(net1459),
    .B(net849),
    .Y(_2856_));
 sg13g2_a21oi_1 _6392_ (.A1(net1140),
    .A2(net849),
    .Y(_0577_),
    .B1(_2856_));
 sg13g2_nor2_1 _6393_ (.A(net1451),
    .B(net848),
    .Y(_2857_));
 sg13g2_a21oi_1 _6394_ (.A1(_2292_),
    .A2(net848),
    .Y(_0578_),
    .B1(_2857_));
 sg13g2_nor2_1 _6395_ (.A(net1475),
    .B(net848),
    .Y(_2858_));
 sg13g2_a21oi_1 _6396_ (.A1(net1134),
    .A2(net848),
    .Y(_0579_),
    .B1(_2858_));
 sg13g2_nor2_1 _6397_ (.A(net1496),
    .B(net848),
    .Y(_2859_));
 sg13g2_a21oi_1 _6398_ (.A1(net1131),
    .A2(net848),
    .Y(_0580_),
    .B1(_2859_));
 sg13g2_nor2_1 _6399_ (.A(net1566),
    .B(net854),
    .Y(_2860_));
 sg13g2_a21oi_1 _6400_ (.A1(net1128),
    .A2(net854),
    .Y(_0581_),
    .B1(_2860_));
 sg13g2_nor2_1 _6401_ (.A(net1491),
    .B(net854),
    .Y(_2861_));
 sg13g2_a21oi_1 _6402_ (.A1(net1125),
    .A2(net854),
    .Y(_0582_),
    .B1(_2861_));
 sg13g2_nor2_1 _6403_ (.A(net1464),
    .B(net850),
    .Y(_2862_));
 sg13g2_a21oi_1 _6404_ (.A1(net1122),
    .A2(net850),
    .Y(_0583_),
    .B1(_2862_));
 sg13g2_nor2_1 _6405_ (.A(net1432),
    .B(net848),
    .Y(_2863_));
 sg13g2_a21oi_1 _6406_ (.A1(net1119),
    .A2(net848),
    .Y(_0584_),
    .B1(_2863_));
 sg13g2_nor2_1 _6407_ (.A(net1499),
    .B(net851),
    .Y(_2864_));
 sg13g2_a21oi_1 _6408_ (.A1(net1116),
    .A2(net851),
    .Y(_0585_),
    .B1(_2864_));
 sg13g2_nor2_1 _6409_ (.A(net1457),
    .B(net851),
    .Y(_2865_));
 sg13g2_a21oi_1 _6410_ (.A1(net1112),
    .A2(net851),
    .Y(_0586_),
    .B1(_2865_));
 sg13g2_nor2_1 _6411_ (.A(net1552),
    .B(net852),
    .Y(_2866_));
 sg13g2_a21oi_1 _6412_ (.A1(net1109),
    .A2(net852),
    .Y(_0587_),
    .B1(_2866_));
 sg13g2_nor2_1 _6413_ (.A(net1519),
    .B(net852),
    .Y(_2867_));
 sg13g2_a21oi_1 _6414_ (.A1(net1107),
    .A2(net852),
    .Y(_0588_),
    .B1(_2867_));
 sg13g2_nor2_1 _6415_ (.A(net1452),
    .B(net853),
    .Y(_2868_));
 sg13g2_a21oi_1 _6416_ (.A1(net1103),
    .A2(net853),
    .Y(_0589_),
    .B1(_2868_));
 sg13g2_nor2_1 _6417_ (.A(net1530),
    .B(net853),
    .Y(_2869_));
 sg13g2_a21oi_1 _6418_ (.A1(net1101),
    .A2(net853),
    .Y(_0590_),
    .B1(_2869_));
 sg13g2_nor2_1 _6419_ (.A(net1571),
    .B(net850),
    .Y(_2870_));
 sg13g2_a21oi_1 _6420_ (.A1(_2344_),
    .A2(net850),
    .Y(_0591_),
    .B1(_2870_));
 sg13g2_nor2_1 _6421_ (.A(net1463),
    .B(net849),
    .Y(_2871_));
 sg13g2_a21oi_1 _6422_ (.A1(net1095),
    .A2(net849),
    .Y(_0592_),
    .B1(_2871_));
 sg13g2_nor3_1 _6423_ (.A(net1204),
    .B(net1248),
    .C(net1710),
    .Y(_0593_));
 sg13g2_nor4_1 _6424_ (.A(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .B(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .C(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .D(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .Y(_2872_));
 sg13g2_nor4_1 _6425_ (.A(_0630_),
    .B(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .C(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .D(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .Y(_2873_));
 sg13g2_nand4_1 _6426_ (.B(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .C(_2872_),
    .A(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .Y(_2874_),
    .D(_2873_));
 sg13g2_and2_1 _6427_ (.A(_1788_),
    .B(_2874_),
    .X(_2875_));
 sg13g2_or4_1 _6428_ (.A(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .B(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .C(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .D(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .X(_2876_));
 sg13g2_nand4_1 _6429_ (.B(_0631_),
    .C(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .A(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .Y(_2877_),
    .D(\vga_tetris.vgaController.verticalCounterQ[2] ));
 sg13g2_nor4_1 _6430_ (.A(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .B(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .C(_2876_),
    .D(_2877_),
    .Y(_2878_));
 sg13g2_o21ai_1 _6431_ (.B1(net1259),
    .Y(_2879_),
    .A1(net1603),
    .A2(_2875_));
 sg13g2_a21oi_1 _6432_ (.A1(net1603),
    .A2(_1788_),
    .Y(_0594_),
    .B1(_2879_));
 sg13g2_a21oi_1 _6433_ (.A1(net1603),
    .A2(_1788_),
    .Y(_2880_),
    .B1(net1622));
 sg13g2_nand2_1 _6434_ (.Y(_2881_),
    .A(net1622),
    .B(net1603));
 sg13g2_nand2_1 _6435_ (.Y(_2882_),
    .A(net1259),
    .B(_2881_));
 sg13g2_a21oi_1 _6436_ (.A1(net1088),
    .A2(_2882_),
    .Y(_0595_),
    .B1(net1623));
 sg13g2_nand2_1 _6437_ (.Y(_2883_),
    .A(net1677),
    .B(_1789_));
 sg13g2_nand3_1 _6438_ (.B(net1622),
    .C(net1603),
    .A(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .Y(_2884_));
 sg13g2_xor2_1 _6439_ (.B(_2881_),
    .A(net1677),
    .X(_2885_));
 sg13g2_nand2_2 _6440_ (.Y(_2886_),
    .A(net1259),
    .B(_2875_));
 sg13g2_o21ai_1 _6441_ (.B1(_2883_),
    .Y(_0596_),
    .A1(_2885_),
    .A2(_2886_));
 sg13g2_nand2_1 _6442_ (.Y(_2887_),
    .A(net1599),
    .B(_1789_));
 sg13g2_nor2_1 _6443_ (.A(_0632_),
    .B(_2884_),
    .Y(_2888_));
 sg13g2_xnor2_1 _6444_ (.Y(_2889_),
    .A(_0632_),
    .B(_2884_));
 sg13g2_o21ai_1 _6445_ (.B1(_2887_),
    .Y(_0597_),
    .A1(_2886_),
    .A2(_2889_));
 sg13g2_a21oi_1 _6446_ (.A1(_1788_),
    .A2(_2888_),
    .Y(_2890_),
    .B1(net1667));
 sg13g2_and3_2 _6447_ (.X(_2891_),
    .A(net1667),
    .B(_1788_),
    .C(_2888_));
 sg13g2_nor3_1 _6448_ (.A(net1245),
    .B(net1668),
    .C(_2891_),
    .Y(_0598_));
 sg13g2_and2_1 _6449_ (.A(net1766),
    .B(_2891_),
    .X(_2892_));
 sg13g2_xnor2_1 _6450_ (.Y(_2893_),
    .A(net1766),
    .B(_2891_));
 sg13g2_nor2_1 _6451_ (.A(net1245),
    .B(_2893_),
    .Y(_0599_));
 sg13g2_xnor2_1 _6452_ (.Y(_2894_),
    .A(net1779),
    .B(_2892_));
 sg13g2_nor2_1 _6453_ (.A(net1245),
    .B(_2894_),
    .Y(_0600_));
 sg13g2_a21o_1 _6454_ (.A2(_2892_),
    .A1(net1779),
    .B1(net1833),
    .X(_2895_));
 sg13g2_nand3_1 _6455_ (.B(net1779),
    .C(_2892_),
    .A(net1833),
    .Y(_2896_));
 sg13g2_and3_1 _6456_ (.X(_0601_),
    .A(net1259),
    .B(_2895_),
    .C(_2896_));
 sg13g2_nand3_1 _6457_ (.B(_1132_),
    .C(_2888_),
    .A(net1667),
    .Y(_2897_));
 sg13g2_nand2_1 _6458_ (.Y(_2898_),
    .A(net1259),
    .B(_2897_));
 sg13g2_a22oi_1 _6459_ (.Y(_0602_),
    .B1(_2898_),
    .B2(_1790_),
    .A2(_2896_),
    .A1(_0631_));
 sg13g2_o21ai_1 _6460_ (.B1(_0630_),
    .Y(_2899_),
    .A1(_2886_),
    .A2(_2897_));
 sg13g2_nor2_1 _6461_ (.A(_0630_),
    .B(_2897_),
    .Y(_2900_));
 sg13g2_o21ai_1 _6462_ (.B1(net1088),
    .Y(_2901_),
    .A1(_2886_),
    .A2(_2900_));
 sg13g2_and2_1 _6463_ (.A(_2899_),
    .B(_2901_),
    .X(_0603_));
 sg13g2_xnor2_1 _6464_ (.Y(_2902_),
    .A(net1782),
    .B(net1089));
 sg13g2_nor2_1 _6465_ (.A(net1088),
    .B(net1783),
    .Y(_0604_));
 sg13g2_nor2b_2 _6466_ (.A(net1089),
    .B_N(_1781_),
    .Y(_2903_));
 sg13g2_xor2_1 _6467_ (.B(net1782),
    .A(net1788),
    .X(_2904_));
 sg13g2_a22oi_1 _6468_ (.Y(_2905_),
    .B1(_2904_),
    .B2(net1089),
    .A2(_2903_),
    .A1(net1788));
 sg13g2_nor2_1 _6469_ (.A(net1243),
    .B(_2905_),
    .Y(_0605_));
 sg13g2_a21oi_1 _6470_ (.A1(net1788),
    .A2(net1782),
    .Y(_2906_),
    .B1(net1225));
 sg13g2_nor2_1 _6471_ (.A(_0905_),
    .B(_2906_),
    .Y(_2907_));
 sg13g2_a22oi_1 _6472_ (.Y(_2908_),
    .B1(_2907_),
    .B2(net1089),
    .A2(_2903_),
    .A1(net1225));
 sg13g2_nor2_1 _6473_ (.A(net1243),
    .B(_2908_),
    .Y(_0606_));
 sg13g2_a22oi_1 _6474_ (.Y(_2909_),
    .B1(_2903_),
    .B2(net1819),
    .A2(net1089),
    .A1(_0907_));
 sg13g2_o21ai_1 _6475_ (.B1(net1260),
    .Y(_2910_),
    .A1(net1819),
    .A2(_0905_));
 sg13g2_nor2_1 _6476_ (.A(_2909_),
    .B(_2910_),
    .Y(_0607_));
 sg13g2_a22oi_1 _6477_ (.Y(_2911_),
    .B1(_2903_),
    .B2(net1221),
    .A2(net1089),
    .A1(_1782_));
 sg13g2_o21ai_1 _6478_ (.B1(net1260),
    .Y(_2912_),
    .A1(net1222),
    .A2(_0906_));
 sg13g2_nor2_1 _6479_ (.A(_2911_),
    .B(_2912_),
    .Y(_0608_));
 sg13g2_a22oi_1 _6480_ (.Y(_2913_),
    .B1(_2903_),
    .B2(net1220),
    .A2(_1787_),
    .A1(_1784_));
 sg13g2_a21oi_1 _6481_ (.A1(net1222),
    .A2(_0906_),
    .Y(_2914_),
    .B1(net1220));
 sg13g2_nor3_1 _6482_ (.A(net1246),
    .B(_2913_),
    .C(net1861),
    .Y(_0609_));
 sg13g2_a22oi_1 _6483_ (.Y(_2915_),
    .B1(_2903_),
    .B2(net1219),
    .A2(_1787_),
    .A1(_1785_));
 sg13g2_o21ai_1 _6484_ (.B1(net1260),
    .Y(_2916_),
    .A1(net1219),
    .A2(_1783_));
 sg13g2_nor2_1 _6485_ (.A(net1902),
    .B(_2916_),
    .Y(_0610_));
 sg13g2_nand3_1 _6486_ (.B(net1219),
    .C(_1783_),
    .A(net1218),
    .Y(_2917_));
 sg13g2_and2_1 _6487_ (.A(_1786_),
    .B(_2917_),
    .X(_2918_));
 sg13g2_a22oi_1 _6488_ (.Y(_2919_),
    .B1(_2918_),
    .B2(_0628_),
    .A2(_2903_),
    .A1(net1218));
 sg13g2_nor2_1 _6489_ (.A(net1244),
    .B(net1810),
    .Y(_0611_));
 sg13g2_nand2b_2 _6490_ (.Y(_2920_),
    .B(_0628_),
    .A_N(_2917_));
 sg13g2_nand3b_1 _6491_ (.B(_2920_),
    .C(net1776),
    .Y(_2921_),
    .A_N(_1788_));
 sg13g2_or2_1 _6492_ (.X(_2922_),
    .B(_2920_),
    .A(net1776));
 sg13g2_a21oi_1 _6493_ (.A1(net1777),
    .A2(_2922_),
    .Y(_0612_),
    .B1(net1243));
 sg13g2_o21ai_1 _6494_ (.B1(_2920_),
    .Y(_2923_),
    .A1(net1776),
    .A2(_1786_));
 sg13g2_nor2b_1 _6495_ (.A(_1139_),
    .B_N(_2923_),
    .Y(_2924_));
 sg13g2_nor2_1 _6496_ (.A(_2903_),
    .B(_2924_),
    .Y(_2925_));
 sg13g2_nor2_1 _6497_ (.A(net1244),
    .B(_2925_),
    .Y(_0613_));
 sg13g2_nand2b_1 _6498_ (.Y(_2926_),
    .B(_1156_),
    .A_N(net1210));
 sg13g2_a21oi_1 _6499_ (.A1(_1143_),
    .A2(_2926_),
    .Y(_2927_),
    .B1(net1657));
 sg13g2_and2_1 _6500_ (.A(_2875_),
    .B(_2927_),
    .X(_2928_));
 sg13g2_o21ai_1 _6501_ (.B1(_1788_),
    .Y(_2929_),
    .A1(_2878_),
    .A2(_2927_));
 sg13g2_inv_1 _6502_ (.Y(_2930_),
    .A(_2929_));
 sg13g2_o21ai_1 _6503_ (.B1(net1260),
    .Y(_2931_),
    .A1(net1619),
    .A2(net1080));
 sg13g2_a21oi_1 _6504_ (.A1(net1619),
    .A2(_2930_),
    .Y(_0614_),
    .B1(_2931_));
 sg13g2_xor2_1 _6505_ (.B(net1619),
    .A(net1821),
    .X(_2932_));
 sg13g2_a22oi_1 _6506_ (.Y(_2933_),
    .B1(_2932_),
    .B2(net1080),
    .A2(_2929_),
    .A1(net1821));
 sg13g2_nor2_1 _6507_ (.A(net1243),
    .B(_2933_),
    .Y(_0615_));
 sg13g2_xnor2_1 _6508_ (.Y(_2934_),
    .A(net1217),
    .B(_0908_));
 sg13g2_a22oi_1 _6509_ (.Y(_2935_),
    .B1(_2934_),
    .B2(net1080),
    .A2(_2929_),
    .A1(net1217));
 sg13g2_nor2_1 _6510_ (.A(net1243),
    .B(_2935_),
    .Y(_0616_));
 sg13g2_xnor2_1 _6511_ (.Y(_2936_),
    .A(net1215),
    .B(_0910_));
 sg13g2_a22oi_1 _6512_ (.Y(_2937_),
    .B1(_2936_),
    .B2(net1080),
    .A2(_2929_),
    .A1(net1215));
 sg13g2_nor2_1 _6513_ (.A(net1243),
    .B(_2937_),
    .Y(_0617_));
 sg13g2_xnor2_1 _6514_ (.Y(_2938_),
    .A(_0627_),
    .B(_0911_));
 sg13g2_a22oi_1 _6515_ (.Y(_2939_),
    .B1(_2938_),
    .B2(_2928_),
    .A2(_2929_),
    .A1(net1212));
 sg13g2_nor2_1 _6516_ (.A(net1243),
    .B(_2939_),
    .Y(_0618_));
 sg13g2_nand2_1 _6517_ (.Y(_2940_),
    .A(_0911_),
    .B(_1179_));
 sg13g2_a21oi_1 _6518_ (.A1(net1080),
    .A2(_2940_),
    .Y(_2941_),
    .B1(_2929_));
 sg13g2_o21ai_1 _6519_ (.B1(_2926_),
    .Y(_2942_),
    .A1(net1209),
    .A2(net1080));
 sg13g2_nor3_1 _6520_ (.A(net1244),
    .B(_2941_),
    .C(_2942_),
    .Y(_0619_));
 sg13g2_xnor2_1 _6521_ (.Y(_2943_),
    .A(net1208),
    .B(_2940_));
 sg13g2_a22oi_1 _6522_ (.Y(_2944_),
    .B1(_2943_),
    .B2(net1080),
    .A2(_2929_),
    .A1(net1208));
 sg13g2_nor2_1 _6523_ (.A(net1243),
    .B(_2944_),
    .Y(_0620_));
 sg13g2_nand4_1 _6524_ (.B(_0911_),
    .C(_1179_),
    .A(net1208),
    .Y(_2945_),
    .D(_2928_));
 sg13g2_nand2_1 _6525_ (.Y(_2946_),
    .A(_0716_),
    .B(net1080));
 sg13g2_a21o_1 _6526_ (.A2(_2946_),
    .A1(_2941_),
    .B1(net1244),
    .X(_2947_));
 sg13g2_a21oi_1 _6527_ (.A1(_0626_),
    .A2(_2945_),
    .Y(_0621_),
    .B1(_2947_));
 sg13g2_nand2b_1 _6528_ (.Y(_2948_),
    .B(net1207),
    .A_N(_2947_));
 sg13g2_nand2_1 _6529_ (.Y(_2949_),
    .A(net1260),
    .B(_1152_));
 sg13g2_o21ai_1 _6530_ (.B1(_2948_),
    .Y(_0622_),
    .A1(_2945_),
    .A2(_2949_));
 sg13g2_nor3_1 _6531_ (.A(_0625_),
    .B(net1244),
    .C(_2930_),
    .Y(_0623_));
 sg13g2_a21oi_1 _6532_ (.A1(net1202),
    .A2(net1226),
    .Y(_0624_),
    .B1(_2462_));
 sg13g2_dfrbpq_2 _6533_ (.RESET_B(net329),
    .D(net1881),
    .Q(\vga_tetris.tetrisLogic.stateQ[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6534_ (.RESET_B(net551),
    .D(_0001_),
    .Q(\vga_tetris.tetrisLogic.stateQ[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6535_ (.RESET_B(net549),
    .D(_0002_),
    .Q(\vga_tetris.tetrisLogic.stateQ[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6536_ (.RESET_B(net547),
    .D(_0003_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6537_ (.RESET_B(net546),
    .D(net1909),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6538_ (.RESET_B(net545),
    .D(_0005_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6539_ (.RESET_B(net544),
    .D(_0006_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6540_ (.RESET_B(net543),
    .D(net740),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6541_ (.RESET_B(net542),
    .D(_0008_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6542_ (.RESET_B(net541),
    .D(_0009_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6543_ (.RESET_B(net540),
    .D(net1684),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6544_ (.RESET_B(net539),
    .D(net1671),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6545_ (.RESET_B(net538),
    .D(_0012_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6546_ (.RESET_B(net537),
    .D(_0013_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6547_ (.RESET_B(net536),
    .D(_0014_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6548_ (.RESET_B(net535),
    .D(net648),
    .Q(\vga_tetris.msTimer.msTimerQ[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _6549_ (.RESET_B(net534),
    .D(_0016_),
    .Q(\vga_tetris.msTimer.msTimerQ[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6550_ (.RESET_B(net533),
    .D(net1357),
    .Q(\vga_tetris.msTimer.msTimerQ[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _6551_ (.RESET_B(net532),
    .D(net1660),
    .Q(\vga_tetris.msTimer.msTimerQ[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6552_ (.RESET_B(net531),
    .D(_0019_),
    .Q(\vga_tetris.msTimer.msTimerQ[4] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6553_ (.RESET_B(net530),
    .D(net1687),
    .Q(\vga_tetris.msTimer.msTimerQ[5] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6554_ (.RESET_B(net529),
    .D(net1642),
    .Q(\vga_tetris.msTimer.msTimerQ[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6555_ (.RESET_B(net528),
    .D(_0022_),
    .Q(\vga_tetris.msTimer.msTimerQ[7] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6556_ (.RESET_B(net527),
    .D(_0023_),
    .Q(\vga_tetris.msTimer.msTimerQ[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6557_ (.RESET_B(net526),
    .D(_0024_),
    .Q(\vga_tetris.msTimer.msTimerQ[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6558_ (.RESET_B(net525),
    .D(_0025_),
    .Q(\vga_tetris.msTimer.msTimerQ[10] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6559_ (.RESET_B(net524),
    .D(_0026_),
    .Q(\vga_tetris.msTimer.msTimerQ[11] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6560_ (.RESET_B(net523),
    .D(net1749),
    .Q(\vga_tetris.msTimer.msTimerQ[12] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6561_ (.RESET_B(net522),
    .D(net1347),
    .Q(\vga_tetris.msTimer.msTimerQ[13] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6562_ (.RESET_B(net521),
    .D(_0029_),
    .Q(\vga_tetris.msTimer.msTimerQ[14] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _6563_ (.RESET_B(net520),
    .D(_0030_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6564_ (.RESET_B(net518),
    .D(_0031_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6565_ (.RESET_B(net516),
    .D(_0032_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6566_ (.RESET_B(net514),
    .D(_0033_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6567_ (.RESET_B(net512),
    .D(_0034_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6568_ (.RESET_B(net510),
    .D(_0035_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6569_ (.RESET_B(net508),
    .D(_0036_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6570_ (.RESET_B(net506),
    .D(_0037_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6571_ (.RESET_B(net504),
    .D(_0038_),
    .Q(\vga_tetris.tetrisLogic.rotationQ[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6572_ (.RESET_B(net502),
    .D(net1844),
    .Q(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6573_ (.RESET_B(net500),
    .D(_0040_),
    .Q(\vga_tetris.tetrisLogic.stateQ[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6574_ (.RESET_B(net498),
    .D(net1895),
    .Q(\vga_tetris.tetrisLogic.stateQ[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6575_ (.RESET_B(net496),
    .D(_0042_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6576_ (.RESET_B(net495),
    .D(_0043_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6577_ (.RESET_B(net494),
    .D(_0044_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6578_ (.RESET_B(net493),
    .D(net1550),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6579_ (.RESET_B(net492),
    .D(net1680),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6580_ (.RESET_B(net491),
    .D(_0047_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6581_ (.RESET_B(net490),
    .D(_0048_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6582_ (.RESET_B(net489),
    .D(_0049_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6583_ (.RESET_B(net488),
    .D(_0050_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6584_ (.RESET_B(net486),
    .D(net1611),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6585_ (.RESET_B(net484),
    .D(_0052_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6586_ (.RESET_B(net482),
    .D(net1332),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6587_ (.RESET_B(net480),
    .D(_0054_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6588_ (.RESET_B(net478),
    .D(_0055_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6589_ (.RESET_B(net476),
    .D(_0056_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6590_ (.RESET_B(net474),
    .D(net1411),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6591_ (.RESET_B(net472),
    .D(net1368),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6592_ (.RESET_B(net470),
    .D(_0059_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6593_ (.RESET_B(net468),
    .D(_0060_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6594_ (.RESET_B(net466),
    .D(_0061_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6595_ (.RESET_B(net464),
    .D(net1632),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6596_ (.RESET_B(net462),
    .D(_0063_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6597_ (.RESET_B(net460),
    .D(net1446),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6598_ (.RESET_B(net458),
    .D(_0065_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6599_ (.RESET_B(net456),
    .D(net1702),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6600_ (.RESET_B(net455),
    .D(net1724),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6601_ (.RESET_B(net454),
    .D(net745),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6602_ (.RESET_B(net453),
    .D(net1808),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6603_ (.RESET_B(net451),
    .D(_0070_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6604_ (.RESET_B(net449),
    .D(_0071_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6605_ (.RESET_B(net447),
    .D(_0072_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6606_ (.RESET_B(net445),
    .D(_0073_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6607_ (.RESET_B(net443),
    .D(_0074_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6608_ (.RESET_B(net441),
    .D(net1392),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6609_ (.RESET_B(net439),
    .D(net1467),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6610_ (.RESET_B(net437),
    .D(_0077_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6611_ (.RESET_B(net435),
    .D(_0078_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6612_ (.RESET_B(net433),
    .D(_0079_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6613_ (.RESET_B(net431),
    .D(net1382),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6614_ (.RESET_B(net429),
    .D(_0081_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6615_ (.RESET_B(net427),
    .D(_0082_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6616_ (.RESET_B(net425),
    .D(net1431),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6617_ (.RESET_B(net423),
    .D(_0084_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6618_ (.RESET_B(net421),
    .D(_0085_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6619_ (.RESET_B(net419),
    .D(_0086_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6620_ (.RESET_B(net417),
    .D(_0087_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6621_ (.RESET_B(net415),
    .D(_0088_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6622_ (.RESET_B(net413),
    .D(_0089_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6623_ (.RESET_B(net411),
    .D(_0090_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6624_ (.RESET_B(net409),
    .D(net1752),
    .Q(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6625_ (.RESET_B(net408),
    .D(_0092_),
    .Q(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6626_ (.RESET_B(net407),
    .D(_0093_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6627_ (.RESET_B(net406),
    .D(net1286),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6628_ (.RESET_B(net404),
    .D(net1438),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6629_ (.RESET_B(net402),
    .D(_0096_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6630_ (.RESET_B(net401),
    .D(net1897),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6631_ (.RESET_B(net400),
    .D(net1883),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6632_ (.RESET_B(net399),
    .D(_0099_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6633_ (.RESET_B(net398),
    .D(net1887),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6634_ (.RESET_B(net397),
    .D(_0101_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6635_ (.RESET_B(net396),
    .D(_0102_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6636_ (.RESET_B(net395),
    .D(net1893),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6637_ (.RESET_B(net394),
    .D(_0104_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6638_ (.RESET_B(net393),
    .D(_0105_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6639_ (.RESET_B(net392),
    .D(net1852),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6640_ (.RESET_B(net391),
    .D(_0107_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6641_ (.RESET_B(net389),
    .D(_0108_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6642_ (.RESET_B(net387),
    .D(_0109_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6643_ (.RESET_B(net385),
    .D(_0110_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6644_ (.RESET_B(net383),
    .D(_0111_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6645_ (.RESET_B(net381),
    .D(_0112_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6646_ (.RESET_B(net380),
    .D(_0113_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6647_ (.RESET_B(net379),
    .D(_0114_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6648_ (.RESET_B(net378),
    .D(_0115_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6649_ (.RESET_B(net376),
    .D(_0116_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6650_ (.RESET_B(net374),
    .D(_0117_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6651_ (.RESET_B(net372),
    .D(_0118_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6652_ (.RESET_B(net370),
    .D(net819),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6653_ (.RESET_B(net368),
    .D(net822),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6654_ (.RESET_B(net366),
    .D(net1303),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6655_ (.RESET_B(net364),
    .D(net757),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6656_ (.RESET_B(net362),
    .D(_0123_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6657_ (.RESET_B(net360),
    .D(_0124_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6658_ (.RESET_B(net358),
    .D(_0125_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6659_ (.RESET_B(net356),
    .D(net1370),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6660_ (.RESET_B(net354),
    .D(net1288),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6661_ (.RESET_B(net352),
    .D(_0128_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6662_ (.RESET_B(net350),
    .D(_0129_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6663_ (.RESET_B(net348),
    .D(_0130_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6664_ (.RESET_B(net346),
    .D(_0131_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6665_ (.RESET_B(net344),
    .D(net1698),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6666_ (.RESET_B(net342),
    .D(_0133_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6667_ (.RESET_B(net340),
    .D(net1280),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6668_ (.RESET_B(net338),
    .D(net1722),
    .Q(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6669_ (.RESET_B(net337),
    .D(net1765),
    .Q(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6670_ (.RESET_B(net336),
    .D(net1739),
    .Q(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6671_ (.RESET_B(net335),
    .D(_0138_),
    .Q(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6672_ (.RESET_B(net334),
    .D(net1390),
    .Q(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6673_ (.RESET_B(net332),
    .D(_0140_),
    .Q(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6674_ (.RESET_B(net330),
    .D(_0141_),
    .Q(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6675_ (.RESET_B(net328),
    .D(_0142_),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6676_ (.RESET_B(net327),
    .D(_0143_),
    .Q(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6677_ (.RESET_B(net326),
    .D(_0144_),
    .Q(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6678_ (.RESET_B(net325),
    .D(net1786),
    .Q(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6679_ (.RESET_B(net324),
    .D(net1455),
    .Q(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6680_ (.RESET_B(net323),
    .D(_0147_),
    .Q(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6681_ (.RESET_B(net322),
    .D(_0148_),
    .Q(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6682_ (.RESET_B(net321),
    .D(net1775),
    .Q(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6683_ (.RESET_B(net320),
    .D(net1406),
    .Q(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6684_ (.RESET_B(net319),
    .D(_0151_),
    .Q(\vga_tetris._tetrisLogic_io_score_0[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6685_ (.RESET_B(net318),
    .D(_0152_),
    .Q(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6686_ (.RESET_B(net317),
    .D(net1793),
    .Q(\vga_tetris._tetrisLogic_io_score_0[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6687_ (.RESET_B(net316),
    .D(_0154_),
    .Q(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6688_ (.RESET_B(net315),
    .D(_0155_),
    .Q(\vga_tetris._tetrisLogic_io_gameOver ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6689_ (.RESET_B(net314),
    .D(_0156_),
    .Q(\vga_tetris.boardMem.board_19[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6690_ (.RESET_B(net313),
    .D(_0157_),
    .Q(\vga_tetris.boardMem.board_19[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6691_ (.RESET_B(net312),
    .D(_0158_),
    .Q(\vga_tetris.boardMem.board_19[2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6692_ (.RESET_B(net311),
    .D(_0159_),
    .Q(\vga_tetris.boardMem.board_19[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6693_ (.RESET_B(net310),
    .D(_0160_),
    .Q(\vga_tetris.boardMem.board_19[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _6694_ (.RESET_B(net309),
    .D(_0161_),
    .Q(\vga_tetris.boardMem.board_19[5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6695_ (.RESET_B(net308),
    .D(_0162_),
    .Q(\vga_tetris.boardMem.board_19[6] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6696_ (.RESET_B(net307),
    .D(_0163_),
    .Q(\vga_tetris.boardMem.board_19[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6697_ (.RESET_B(net306),
    .D(net1616),
    .Q(\vga_tetris.boardMem.board_19[8] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6698_ (.RESET_B(net305),
    .D(_0165_),
    .Q(\vga_tetris.boardMem.board_19[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6699_ (.RESET_B(net304),
    .D(_0166_),
    .Q(\vga_tetris.boardMem.board_19[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6700_ (.RESET_B(net303),
    .D(_0167_),
    .Q(\vga_tetris.boardMem.board_19[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6701_ (.RESET_B(net302),
    .D(_0168_),
    .Q(\vga_tetris.boardMem.board_19[12] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6702_ (.RESET_B(net301),
    .D(_0169_),
    .Q(\vga_tetris.boardMem.board_19[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6703_ (.RESET_B(net300),
    .D(_0170_),
    .Q(\vga_tetris.boardMem.board_19[14] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6704_ (.RESET_B(net299),
    .D(_0171_),
    .Q(\vga_tetris.boardMem.board_19[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6705_ (.RESET_B(net298),
    .D(_0172_),
    .Q(\vga_tetris.boardMem.board_19[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6706_ (.RESET_B(net297),
    .D(_0173_),
    .Q(\vga_tetris.boardMem.board_19[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6707_ (.RESET_B(net296),
    .D(_0174_),
    .Q(\vga_tetris.boardMem.board_19[18] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6708_ (.RESET_B(net295),
    .D(_0175_),
    .Q(\vga_tetris.boardMem.board_19[19] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6709_ (.RESET_B(net294),
    .D(_0176_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6710_ (.RESET_B(net293),
    .D(net1363),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6711_ (.RESET_B(net292),
    .D(_0178_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6712_ (.RESET_B(net291),
    .D(_0179_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6713_ (.RESET_B(net290),
    .D(net1815),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[4] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6714_ (.RESET_B(net289),
    .D(_0181_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6715_ (.RESET_B(net288),
    .D(net1637),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6716_ (.RESET_B(net287),
    .D(net1628),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[7] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6717_ (.RESET_B(net286),
    .D(net1665),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6718_ (.RESET_B(net285),
    .D(_0185_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6719_ (.RESET_B(net284),
    .D(_0186_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6720_ (.RESET_B(net283),
    .D(net1857),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6721_ (.RESET_B(net282),
    .D(_0188_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6722_ (.RESET_B(net281),
    .D(net1769),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6723_ (.RESET_B(net280),
    .D(_0190_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6724_ (.RESET_B(net279),
    .D(_0191_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6725_ (.RESET_B(net278),
    .D(net1647),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6726_ (.RESET_B(net277),
    .D(net1718),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6727_ (.RESET_B(net276),
    .D(_0194_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6728_ (.RESET_B(net275),
    .D(_0195_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6729_ (.RESET_B(net274),
    .D(net1818),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6730_ (.RESET_B(net273),
    .D(_0197_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6731_ (.RESET_B(net272),
    .D(net1426),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6732_ (.RESET_B(net271),
    .D(net1708),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6733_ (.RESET_B(net270),
    .D(_0200_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6734_ (.RESET_B(net269),
    .D(_0201_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6735_ (.RESET_B(net268),
    .D(_0202_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6736_ (.RESET_B(net267),
    .D(_0203_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6737_ (.RESET_B(net266),
    .D(_0204_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6738_ (.RESET_B(net265),
    .D(_0205_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6739_ (.RESET_B(net264),
    .D(_0206_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6740_ (.RESET_B(net263),
    .D(_0207_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6741_ (.RESET_B(net262),
    .D(_0208_),
    .Q(\vga_tetris._inputs_io_rotateButtonActive ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6742_ (.RESET_B(net261),
    .D(_0209_),
    .Q(\vga_tetris._inputs_io_leftButtonActive ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6743_ (.RESET_B(net260),
    .D(_0210_),
    .Q(\vga_tetris._inputs_io_rightButtonActive ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6744_ (.RESET_B(net259),
    .D(net1693),
    .Q(\vga_tetris._inputs_io_downButtonActive ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6745_ (.RESET_B(net258),
    .D(net1772),
    .Q(\vga_tetris.startTetrisLogicQ ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6746_ (.RESET_B(net257),
    .D(_0213_),
    .Q(\vga_tetris.boardMem.board_0[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6747_ (.RESET_B(net256),
    .D(_0214_),
    .Q(\vga_tetris.boardMem.board_0[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6748_ (.RESET_B(net255),
    .D(net1595),
    .Q(\vga_tetris.boardMem.board_0[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6749_ (.RESET_B(net254),
    .D(net1408),
    .Q(\vga_tetris.boardMem.board_0[3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6750_ (.RESET_B(net253),
    .D(_0217_),
    .Q(\vga_tetris.boardMem.board_0[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6751_ (.RESET_B(net252),
    .D(net1396),
    .Q(\vga_tetris.boardMem.board_0[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6752_ (.RESET_B(net251),
    .D(_0219_),
    .Q(\vga_tetris.boardMem.board_0[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6753_ (.RESET_B(net250),
    .D(_0220_),
    .Q(\vga_tetris.boardMem.board_0[7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6754_ (.RESET_B(net249),
    .D(net1528),
    .Q(\vga_tetris.boardMem.board_0[8] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6755_ (.RESET_B(net248),
    .D(net1490),
    .Q(\vga_tetris.boardMem.board_0[9] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6756_ (.RESET_B(net247),
    .D(net1512),
    .Q(\vga_tetris.boardMem.board_0[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6757_ (.RESET_B(net246),
    .D(_0224_),
    .Q(\vga_tetris.boardMem.board_0[11] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6758_ (.RESET_B(net245),
    .D(_0225_),
    .Q(\vga_tetris.boardMem.board_0[12] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6759_ (.RESET_B(net244),
    .D(net1547),
    .Q(\vga_tetris.boardMem.board_0[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6760_ (.RESET_B(net243),
    .D(net1540),
    .Q(\vga_tetris.boardMem.board_0[14] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6761_ (.RESET_B(net242),
    .D(net1422),
    .Q(\vga_tetris.boardMem.board_0[15] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6762_ (.RESET_B(net241),
    .D(_0229_),
    .Q(\vga_tetris.boardMem.board_0[16] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6763_ (.RESET_B(net240),
    .D(_0230_),
    .Q(\vga_tetris.boardMem.board_0[17] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6764_ (.RESET_B(net239),
    .D(_0231_),
    .Q(\vga_tetris.boardMem.board_0[18] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6765_ (.RESET_B(net238),
    .D(_0232_),
    .Q(\vga_tetris.boardMem.board_0[19] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6766_ (.RESET_B(net237),
    .D(_0233_),
    .Q(\vga_tetris.boardMem.board_1[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6767_ (.RESET_B(net236),
    .D(net1449),
    .Q(\vga_tetris.boardMem.board_1[1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6768_ (.RESET_B(net235),
    .D(_0235_),
    .Q(\vga_tetris.boardMem.board_1[2] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6769_ (.RESET_B(net234),
    .D(_0236_),
    .Q(\vga_tetris.boardMem.board_1[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6770_ (.RESET_B(net233),
    .D(_0237_),
    .Q(\vga_tetris.boardMem.board_1[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _6771_ (.RESET_B(net232),
    .D(_0238_),
    .Q(\vga_tetris.boardMem.board_1[5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6772_ (.RESET_B(net231),
    .D(_0239_),
    .Q(\vga_tetris.boardMem.board_1[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6773_ (.RESET_B(net230),
    .D(_0240_),
    .Q(\vga_tetris.boardMem.board_1[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6774_ (.RESET_B(net229),
    .D(_0241_),
    .Q(\vga_tetris.boardMem.board_1[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6775_ (.RESET_B(net228),
    .D(_0242_),
    .Q(\vga_tetris.boardMem.board_1[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6776_ (.RESET_B(net227),
    .D(_0243_),
    .Q(\vga_tetris.boardMem.board_1[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6777_ (.RESET_B(net226),
    .D(_0244_),
    .Q(\vga_tetris.boardMem.board_1[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6778_ (.RESET_B(net225),
    .D(_0245_),
    .Q(\vga_tetris.boardMem.board_1[12] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _6779_ (.RESET_B(net224),
    .D(_0246_),
    .Q(\vga_tetris.boardMem.board_1[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6780_ (.RESET_B(net223),
    .D(_0247_),
    .Q(\vga_tetris.boardMem.board_1[14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6781_ (.RESET_B(net222),
    .D(_0248_),
    .Q(\vga_tetris.boardMem.board_1[15] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6782_ (.RESET_B(net221),
    .D(net1607),
    .Q(\vga_tetris.boardMem.board_1[16] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6783_ (.RESET_B(net220),
    .D(_0250_),
    .Q(\vga_tetris.boardMem.board_1[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6784_ (.RESET_B(net219),
    .D(_0251_),
    .Q(\vga_tetris.boardMem.board_1[18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6785_ (.RESET_B(net218),
    .D(_0252_),
    .Q(\vga_tetris.boardMem.board_1[19] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _6786_ (.RESET_B(net217),
    .D(_0253_),
    .Q(\vga_tetris.boardMem.board_2[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _6787_ (.RESET_B(net216),
    .D(_0254_),
    .Q(\vga_tetris.boardMem.board_2[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6788_ (.RESET_B(net215),
    .D(_0255_),
    .Q(\vga_tetris.boardMem.board_2[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6789_ (.RESET_B(net214),
    .D(_0256_),
    .Q(\vga_tetris.boardMem.board_2[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6790_ (.RESET_B(net213),
    .D(_0257_),
    .Q(\vga_tetris.boardMem.board_2[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _6791_ (.RESET_B(net212),
    .D(_0258_),
    .Q(\vga_tetris.boardMem.board_2[5] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6792_ (.RESET_B(net211),
    .D(_0259_),
    .Q(\vga_tetris.boardMem.board_2[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6793_ (.RESET_B(net210),
    .D(_0260_),
    .Q(\vga_tetris.boardMem.board_2[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6794_ (.RESET_B(net209),
    .D(_0261_),
    .Q(\vga_tetris.boardMem.board_2[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6795_ (.RESET_B(net208),
    .D(_0262_),
    .Q(\vga_tetris.boardMem.board_2[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6796_ (.RESET_B(net207),
    .D(_0263_),
    .Q(\vga_tetris.boardMem.board_2[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6797_ (.RESET_B(net206),
    .D(_0264_),
    .Q(\vga_tetris.boardMem.board_2[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6798_ (.RESET_B(net205),
    .D(_0265_),
    .Q(\vga_tetris.boardMem.board_2[12] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6799_ (.RESET_B(net204),
    .D(_0266_),
    .Q(\vga_tetris.boardMem.board_2[13] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6800_ (.RESET_B(net203),
    .D(_0267_),
    .Q(\vga_tetris.boardMem.board_2[14] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6801_ (.RESET_B(net202),
    .D(_0268_),
    .Q(\vga_tetris.boardMem.board_2[15] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6802_ (.RESET_B(net201),
    .D(_0269_),
    .Q(\vga_tetris.boardMem.board_2[16] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6803_ (.RESET_B(net200),
    .D(_0270_),
    .Q(\vga_tetris.boardMem.board_2[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6804_ (.RESET_B(net199),
    .D(_0271_),
    .Q(\vga_tetris.boardMem.board_2[18] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6805_ (.RESET_B(net198),
    .D(_0272_),
    .Q(\vga_tetris.boardMem.board_2[19] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6806_ (.RESET_B(net197),
    .D(_0273_),
    .Q(\vga_tetris.boardMem.board_3[0] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _6807_ (.RESET_B(net196),
    .D(_0274_),
    .Q(\vga_tetris.boardMem.board_3[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6808_ (.RESET_B(net195),
    .D(_0275_),
    .Q(\vga_tetris.boardMem.board_3[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6809_ (.RESET_B(net194),
    .D(_0276_),
    .Q(\vga_tetris.boardMem.board_3[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6810_ (.RESET_B(net193),
    .D(_0277_),
    .Q(\vga_tetris.boardMem.board_3[4] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _6811_ (.RESET_B(net192),
    .D(_0278_),
    .Q(\vga_tetris.boardMem.board_3[5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6812_ (.RESET_B(net191),
    .D(_0279_),
    .Q(\vga_tetris.boardMem.board_3[6] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _6813_ (.RESET_B(net190),
    .D(_0280_),
    .Q(\vga_tetris.boardMem.board_3[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6814_ (.RESET_B(net189),
    .D(net1565),
    .Q(\vga_tetris.boardMem.board_3[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6815_ (.RESET_B(net188),
    .D(_0282_),
    .Q(\vga_tetris.boardMem.board_3[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6816_ (.RESET_B(net187),
    .D(_0283_),
    .Q(\vga_tetris.boardMem.board_3[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6817_ (.RESET_B(net186),
    .D(_0284_),
    .Q(\vga_tetris.boardMem.board_3[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6818_ (.RESET_B(net185),
    .D(_0285_),
    .Q(\vga_tetris.boardMem.board_3[12] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _6819_ (.RESET_B(net184),
    .D(_0286_),
    .Q(\vga_tetris.boardMem.board_3[13] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6820_ (.RESET_B(net183),
    .D(_0287_),
    .Q(\vga_tetris.boardMem.board_3[14] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6821_ (.RESET_B(net182),
    .D(_0288_),
    .Q(\vga_tetris.boardMem.board_3[15] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6822_ (.RESET_B(net181),
    .D(_0289_),
    .Q(\vga_tetris.boardMem.board_3[16] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6823_ (.RESET_B(net180),
    .D(_0290_),
    .Q(\vga_tetris.boardMem.board_3[17] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6824_ (.RESET_B(net179),
    .D(_0291_),
    .Q(\vga_tetris.boardMem.board_3[18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6825_ (.RESET_B(net178),
    .D(_0292_),
    .Q(\vga_tetris.boardMem.board_3[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _6826_ (.RESET_B(net177),
    .D(_0293_),
    .Q(\vga_tetris.boardMem.board_4[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _6827_ (.RESET_B(net176),
    .D(_0294_),
    .Q(\vga_tetris.boardMem.board_4[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6828_ (.RESET_B(net175),
    .D(_0295_),
    .Q(\vga_tetris.boardMem.board_4[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6829_ (.RESET_B(net174),
    .D(_0296_),
    .Q(\vga_tetris.boardMem.board_4[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6830_ (.RESET_B(net173),
    .D(_0297_),
    .Q(\vga_tetris.boardMem.board_4[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6831_ (.RESET_B(net172),
    .D(_0298_),
    .Q(\vga_tetris.boardMem.board_4[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6832_ (.RESET_B(net171),
    .D(_0299_),
    .Q(\vga_tetris.boardMem.board_4[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6833_ (.RESET_B(net170),
    .D(net1325),
    .Q(\vga_tetris.boardMem.board_4[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6834_ (.RESET_B(net169),
    .D(_0301_),
    .Q(\vga_tetris.boardMem.board_4[8] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6835_ (.RESET_B(net168),
    .D(_0302_),
    .Q(\vga_tetris.boardMem.board_4[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6836_ (.RESET_B(net167),
    .D(net697),
    .Q(\vga_tetris.boardMem.board_4[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6837_ (.RESET_B(net166),
    .D(net687),
    .Q(\vga_tetris.boardMem.board_4[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6838_ (.RESET_B(net165),
    .D(_0305_),
    .Q(\vga_tetris.boardMem.board_4[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _6839_ (.RESET_B(net164),
    .D(_0306_),
    .Q(\vga_tetris.boardMem.board_4[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6840_ (.RESET_B(net163),
    .D(_0307_),
    .Q(\vga_tetris.boardMem.board_4[14] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6841_ (.RESET_B(net162),
    .D(_0308_),
    .Q(\vga_tetris.boardMem.board_4[15] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6842_ (.RESET_B(net161),
    .D(_0309_),
    .Q(\vga_tetris.boardMem.board_4[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6843_ (.RESET_B(net160),
    .D(net728),
    .Q(\vga_tetris.boardMem.board_4[17] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6844_ (.RESET_B(net159),
    .D(_0311_),
    .Q(\vga_tetris.boardMem.board_4[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6845_ (.RESET_B(net158),
    .D(_0312_),
    .Q(\vga_tetris.boardMem.board_4[19] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6846_ (.RESET_B(net157),
    .D(_0313_),
    .Q(\vga_tetris.boardMem.board_5[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6847_ (.RESET_B(net156),
    .D(_0314_),
    .Q(\vga_tetris.boardMem.board_5[1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6848_ (.RESET_B(net155),
    .D(_0315_),
    .Q(\vga_tetris.boardMem.board_5[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6849_ (.RESET_B(net154),
    .D(_0316_),
    .Q(\vga_tetris.boardMem.board_5[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6850_ (.RESET_B(net153),
    .D(_0317_),
    .Q(\vga_tetris.boardMem.board_5[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _6851_ (.RESET_B(net152),
    .D(_0318_),
    .Q(\vga_tetris.boardMem.board_5[5] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _6852_ (.RESET_B(net151),
    .D(_0319_),
    .Q(\vga_tetris.boardMem.board_5[6] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _6853_ (.RESET_B(net150),
    .D(_0320_),
    .Q(\vga_tetris.boardMem.board_5[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6854_ (.RESET_B(net149),
    .D(_0321_),
    .Q(\vga_tetris.boardMem.board_5[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6855_ (.RESET_B(net148),
    .D(_0322_),
    .Q(\vga_tetris.boardMem.board_5[9] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6856_ (.RESET_B(net147),
    .D(_0323_),
    .Q(\vga_tetris.boardMem.board_5[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6857_ (.RESET_B(net146),
    .D(net794),
    .Q(\vga_tetris.boardMem.board_5[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6858_ (.RESET_B(net145),
    .D(_0325_),
    .Q(\vga_tetris.boardMem.board_5[12] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _6859_ (.RESET_B(net144),
    .D(_0326_),
    .Q(\vga_tetris.boardMem.board_5[13] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6860_ (.RESET_B(net143),
    .D(_0327_),
    .Q(\vga_tetris.boardMem.board_5[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6861_ (.RESET_B(net142),
    .D(_0328_),
    .Q(\vga_tetris.boardMem.board_5[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6862_ (.RESET_B(net141),
    .D(_0329_),
    .Q(\vga_tetris.boardMem.board_5[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6863_ (.RESET_B(net140),
    .D(_0330_),
    .Q(\vga_tetris.boardMem.board_5[17] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6864_ (.RESET_B(net139),
    .D(_0331_),
    .Q(\vga_tetris.boardMem.board_5[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6865_ (.RESET_B(net138),
    .D(_0332_),
    .Q(\vga_tetris.boardMem.board_5[19] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _6866_ (.RESET_B(net137),
    .D(_0333_),
    .Q(\vga_tetris.boardMem.board_6[0] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6867_ (.RESET_B(net136),
    .D(_0334_),
    .Q(\vga_tetris.boardMem.board_6[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6868_ (.RESET_B(net135),
    .D(_0335_),
    .Q(\vga_tetris.boardMem.board_6[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6869_ (.RESET_B(net134),
    .D(_0336_),
    .Q(\vga_tetris.boardMem.board_6[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6870_ (.RESET_B(net133),
    .D(_0337_),
    .Q(\vga_tetris.boardMem.board_6[4] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _6871_ (.RESET_B(net132),
    .D(_0338_),
    .Q(\vga_tetris.boardMem.board_6[5] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6872_ (.RESET_B(net131),
    .D(_0339_),
    .Q(\vga_tetris.boardMem.board_6[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6873_ (.RESET_B(net130),
    .D(_0340_),
    .Q(\vga_tetris.boardMem.board_6[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6874_ (.RESET_B(net129),
    .D(_0341_),
    .Q(\vga_tetris.boardMem.board_6[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6875_ (.RESET_B(net128),
    .D(_0342_),
    .Q(\vga_tetris.boardMem.board_6[9] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6876_ (.RESET_B(net127),
    .D(net711),
    .Q(\vga_tetris.boardMem.board_6[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6877_ (.RESET_B(net126),
    .D(_0344_),
    .Q(\vga_tetris.boardMem.board_6[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6878_ (.RESET_B(net125),
    .D(_0345_),
    .Q(\vga_tetris.boardMem.board_6[12] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6879_ (.RESET_B(net124),
    .D(_0346_),
    .Q(\vga_tetris.boardMem.board_6[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _6880_ (.RESET_B(net123),
    .D(_0347_),
    .Q(\vga_tetris.boardMem.board_6[14] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6881_ (.RESET_B(net122),
    .D(_0348_),
    .Q(\vga_tetris.boardMem.board_6[15] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6882_ (.RESET_B(net121),
    .D(_0349_),
    .Q(\vga_tetris.boardMem.board_6[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6883_ (.RESET_B(net120),
    .D(_0350_),
    .Q(\vga_tetris.boardMem.board_6[17] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6884_ (.RESET_B(net119),
    .D(_0351_),
    .Q(\vga_tetris.boardMem.board_6[18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6885_ (.RESET_B(net118),
    .D(_0352_),
    .Q(\vga_tetris.boardMem.board_6[19] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6886_ (.RESET_B(net117),
    .D(_0353_),
    .Q(\vga_tetris.boardMem.board_7[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6887_ (.RESET_B(net116),
    .D(_0354_),
    .Q(\vga_tetris.boardMem.board_7[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6888_ (.RESET_B(net115),
    .D(_0355_),
    .Q(\vga_tetris.boardMem.board_7[2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6889_ (.RESET_B(net114),
    .D(_0356_),
    .Q(\vga_tetris.boardMem.board_7[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6890_ (.RESET_B(net113),
    .D(_0357_),
    .Q(\vga_tetris.boardMem.board_7[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6891_ (.RESET_B(net112),
    .D(_0358_),
    .Q(\vga_tetris.boardMem.board_7[5] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6892_ (.RESET_B(net111),
    .D(_0359_),
    .Q(\vga_tetris.boardMem.board_7[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6893_ (.RESET_B(net110),
    .D(_0360_),
    .Q(\vga_tetris.boardMem.board_7[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6894_ (.RESET_B(net109),
    .D(_0361_),
    .Q(\vga_tetris.boardMem.board_7[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6895_ (.RESET_B(net108),
    .D(_0362_),
    .Q(\vga_tetris.boardMem.board_7[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6896_ (.RESET_B(net107),
    .D(_0363_),
    .Q(\vga_tetris.boardMem.board_7[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6897_ (.RESET_B(net106),
    .D(_0364_),
    .Q(\vga_tetris.boardMem.board_7[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6898_ (.RESET_B(net105),
    .D(net1334),
    .Q(\vga_tetris.boardMem.board_7[12] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _6899_ (.RESET_B(net104),
    .D(_0366_),
    .Q(\vga_tetris.boardMem.board_7[13] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6900_ (.RESET_B(net103),
    .D(_0367_),
    .Q(\vga_tetris.boardMem.board_7[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6901_ (.RESET_B(net102),
    .D(_0368_),
    .Q(\vga_tetris.boardMem.board_7[15] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6902_ (.RESET_B(net101),
    .D(_0369_),
    .Q(\vga_tetris.boardMem.board_7[16] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6903_ (.RESET_B(net100),
    .D(_0370_),
    .Q(\vga_tetris.boardMem.board_7[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6904_ (.RESET_B(net99),
    .D(_0371_),
    .Q(\vga_tetris.boardMem.board_7[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6905_ (.RESET_B(net98),
    .D(_0372_),
    .Q(\vga_tetris.boardMem.board_7[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _6906_ (.RESET_B(net97),
    .D(_0373_),
    .Q(\vga_tetris.boardMem.board_8[0] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _6907_ (.RESET_B(net96),
    .D(_0374_),
    .Q(\vga_tetris.boardMem.board_8[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6908_ (.RESET_B(net95),
    .D(net673),
    .Q(\vga_tetris.boardMem.board_8[2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6909_ (.RESET_B(net94),
    .D(_0376_),
    .Q(\vga_tetris.boardMem.board_8[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6910_ (.RESET_B(net93),
    .D(net789),
    .Q(\vga_tetris.boardMem.board_8[4] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _6911_ (.RESET_B(net92),
    .D(_0378_),
    .Q(\vga_tetris.boardMem.board_8[5] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6912_ (.RESET_B(net91),
    .D(_0379_),
    .Q(\vga_tetris.boardMem.board_8[6] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6913_ (.RESET_B(net90),
    .D(_0380_),
    .Q(\vga_tetris.boardMem.board_8[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6914_ (.RESET_B(net89),
    .D(_0381_),
    .Q(\vga_tetris.boardMem.board_8[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6915_ (.RESET_B(net88),
    .D(_0382_),
    .Q(\vga_tetris.boardMem.board_8[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6916_ (.RESET_B(net87),
    .D(_0383_),
    .Q(\vga_tetris.boardMem.board_8[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6917_ (.RESET_B(net86),
    .D(_0384_),
    .Q(\vga_tetris.boardMem.board_8[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6918_ (.RESET_B(net85),
    .D(net720),
    .Q(\vga_tetris.boardMem.board_8[12] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _6919_ (.RESET_B(net84),
    .D(_0386_),
    .Q(\vga_tetris.boardMem.board_8[13] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6920_ (.RESET_B(net83),
    .D(_0387_),
    .Q(\vga_tetris.boardMem.board_8[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6921_ (.RESET_B(net82),
    .D(_0388_),
    .Q(\vga_tetris.boardMem.board_8[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6922_ (.RESET_B(net81),
    .D(_0389_),
    .Q(\vga_tetris.boardMem.board_8[16] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6923_ (.RESET_B(net80),
    .D(_0390_),
    .Q(\vga_tetris.boardMem.board_8[17] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6924_ (.RESET_B(net79),
    .D(_0391_),
    .Q(\vga_tetris.boardMem.board_8[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6925_ (.RESET_B(net78),
    .D(_0392_),
    .Q(\vga_tetris.boardMem.board_8[19] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6926_ (.RESET_B(net77),
    .D(_0393_),
    .Q(\vga_tetris.boardMem.board_9[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _6927_ (.RESET_B(net76),
    .D(_0394_),
    .Q(\vga_tetris.boardMem.board_9[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6928_ (.RESET_B(net75),
    .D(_0395_),
    .Q(\vga_tetris.boardMem.board_9[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6929_ (.RESET_B(net74),
    .D(_0396_),
    .Q(\vga_tetris.boardMem.board_9[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6930_ (.RESET_B(net73),
    .D(_0397_),
    .Q(\vga_tetris.boardMem.board_9[4] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _6931_ (.RESET_B(net72),
    .D(_0398_),
    .Q(\vga_tetris.boardMem.board_9[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6932_ (.RESET_B(net71),
    .D(_0399_),
    .Q(\vga_tetris.boardMem.board_9[6] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _6933_ (.RESET_B(net70),
    .D(net777),
    .Q(\vga_tetris.boardMem.board_9[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6934_ (.RESET_B(net69),
    .D(_0401_),
    .Q(\vga_tetris.boardMem.board_9[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6935_ (.RESET_B(net68),
    .D(_0402_),
    .Q(\vga_tetris.boardMem.board_9[9] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6936_ (.RESET_B(net67),
    .D(net678),
    .Q(\vga_tetris.boardMem.board_9[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6937_ (.RESET_B(net66),
    .D(_0404_),
    .Q(\vga_tetris.boardMem.board_9[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6938_ (.RESET_B(net65),
    .D(_0405_),
    .Q(\vga_tetris.boardMem.board_9[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _6939_ (.RESET_B(net64),
    .D(_0406_),
    .Q(\vga_tetris.boardMem.board_9[13] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6940_ (.RESET_B(net63),
    .D(_0407_),
    .Q(\vga_tetris.boardMem.board_9[14] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6941_ (.RESET_B(net62),
    .D(_0408_),
    .Q(\vga_tetris.boardMem.board_9[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6942_ (.RESET_B(net61),
    .D(_0409_),
    .Q(\vga_tetris.boardMem.board_9[16] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6943_ (.RESET_B(net60),
    .D(_0410_),
    .Q(\vga_tetris.boardMem.board_9[17] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6944_ (.RESET_B(net59),
    .D(_0411_),
    .Q(\vga_tetris.boardMem.board_9[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6945_ (.RESET_B(net58),
    .D(_0412_),
    .Q(\vga_tetris.boardMem.board_9[19] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6946_ (.RESET_B(net57),
    .D(_0413_),
    .Q(\vga_tetris.boardMem.board_10[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _6947_ (.RESET_B(net56),
    .D(_0414_),
    .Q(\vga_tetris.boardMem.board_10[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6948_ (.RESET_B(net55),
    .D(_0415_),
    .Q(\vga_tetris.boardMem.board_10[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6949_ (.RESET_B(net54),
    .D(_0416_),
    .Q(\vga_tetris.boardMem.board_10[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6950_ (.RESET_B(net53),
    .D(_0417_),
    .Q(\vga_tetris.boardMem.board_10[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6951_ (.RESET_B(net52),
    .D(_0418_),
    .Q(\vga_tetris.boardMem.board_10[5] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6952_ (.RESET_B(net51),
    .D(_0419_),
    .Q(\vga_tetris.boardMem.board_10[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6953_ (.RESET_B(net50),
    .D(_0420_),
    .Q(\vga_tetris.boardMem.board_10[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6954_ (.RESET_B(net49),
    .D(_0421_),
    .Q(\vga_tetris.boardMem.board_10[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6955_ (.RESET_B(net48),
    .D(_0422_),
    .Q(\vga_tetris.boardMem.board_10[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6956_ (.RESET_B(net47),
    .D(_0423_),
    .Q(\vga_tetris.boardMem.board_10[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6957_ (.RESET_B(net46),
    .D(_0424_),
    .Q(\vga_tetris.boardMem.board_10[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6958_ (.RESET_B(net45),
    .D(_0425_),
    .Q(\vga_tetris.boardMem.board_10[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _6959_ (.RESET_B(net44),
    .D(_0426_),
    .Q(\vga_tetris.boardMem.board_10[13] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6960_ (.RESET_B(net43),
    .D(_0427_),
    .Q(\vga_tetris.boardMem.board_10[14] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6961_ (.RESET_B(net42),
    .D(_0428_),
    .Q(\vga_tetris.boardMem.board_10[15] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6962_ (.RESET_B(net41),
    .D(_0429_),
    .Q(\vga_tetris.boardMem.board_10[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6963_ (.RESET_B(net40),
    .D(net747),
    .Q(\vga_tetris.boardMem.board_10[17] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6964_ (.RESET_B(net39),
    .D(_0431_),
    .Q(\vga_tetris.boardMem.board_10[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6965_ (.RESET_B(net38),
    .D(_0432_),
    .Q(\vga_tetris.boardMem.board_10[19] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _6966_ (.RESET_B(net37),
    .D(_0433_),
    .Q(\vga_tetris.boardMem.board_11[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _6967_ (.RESET_B(net36),
    .D(_0434_),
    .Q(\vga_tetris.boardMem.board_11[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6968_ (.RESET_B(net35),
    .D(_0435_),
    .Q(\vga_tetris.boardMem.board_11[2] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6969_ (.RESET_B(net34),
    .D(_0436_),
    .Q(\vga_tetris.boardMem.board_11[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6970_ (.RESET_B(net33),
    .D(_0437_),
    .Q(\vga_tetris.boardMem.board_11[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6971_ (.RESET_B(net32),
    .D(_0438_),
    .Q(\vga_tetris.boardMem.board_11[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6972_ (.RESET_B(net31),
    .D(_0439_),
    .Q(\vga_tetris.boardMem.board_11[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6973_ (.RESET_B(net30),
    .D(net837),
    .Q(\vga_tetris.boardMem.board_11[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6974_ (.RESET_B(net29),
    .D(_0441_),
    .Q(\vga_tetris.boardMem.board_11[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6975_ (.RESET_B(net28),
    .D(_0442_),
    .Q(\vga_tetris.boardMem.board_11[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6976_ (.RESET_B(net27),
    .D(_0443_),
    .Q(\vga_tetris.boardMem.board_11[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6977_ (.RESET_B(net26),
    .D(_0444_),
    .Q(\vga_tetris.boardMem.board_11[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6978_ (.RESET_B(net25),
    .D(_0445_),
    .Q(\vga_tetris.boardMem.board_11[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _6979_ (.RESET_B(net24),
    .D(_0446_),
    .Q(\vga_tetris.boardMem.board_11[13] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _6980_ (.RESET_B(net23),
    .D(_0447_),
    .Q(\vga_tetris.boardMem.board_11[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6981_ (.RESET_B(net22),
    .D(_0448_),
    .Q(\vga_tetris.boardMem.board_11[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6982_ (.RESET_B(net21),
    .D(_0449_),
    .Q(\vga_tetris.boardMem.board_11[16] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6983_ (.RESET_B(net645),
    .D(_0450_),
    .Q(\vga_tetris.boardMem.board_11[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6984_ (.RESET_B(net644),
    .D(_0451_),
    .Q(\vga_tetris.boardMem.board_11[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6985_ (.RESET_B(net643),
    .D(net702),
    .Q(\vga_tetris.boardMem.board_11[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _6986_ (.RESET_B(net642),
    .D(net665),
    .Q(\vga_tetris.boardMem.board_12[0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6987_ (.RESET_B(net641),
    .D(_0454_),
    .Q(\vga_tetris.boardMem.board_12[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6988_ (.RESET_B(net640),
    .D(_0455_),
    .Q(\vga_tetris.boardMem.board_12[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6989_ (.RESET_B(net639),
    .D(_0456_),
    .Q(\vga_tetris.boardMem.board_12[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6990_ (.RESET_B(net638),
    .D(_0457_),
    .Q(\vga_tetris.boardMem.board_12[4] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _6991_ (.RESET_B(net637),
    .D(_0458_),
    .Q(\vga_tetris.boardMem.board_12[5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _6992_ (.RESET_B(net636),
    .D(_0459_),
    .Q(\vga_tetris.boardMem.board_12[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _6993_ (.RESET_B(net635),
    .D(_0460_),
    .Q(\vga_tetris.boardMem.board_12[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6994_ (.RESET_B(net634),
    .D(_0461_),
    .Q(\vga_tetris.boardMem.board_12[8] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6995_ (.RESET_B(net633),
    .D(_0462_),
    .Q(\vga_tetris.boardMem.board_12[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6996_ (.RESET_B(net632),
    .D(_0463_),
    .Q(\vga_tetris.boardMem.board_12[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6997_ (.RESET_B(net631),
    .D(net680),
    .Q(\vga_tetris.boardMem.board_12[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6998_ (.RESET_B(net630),
    .D(_0465_),
    .Q(\vga_tetris.boardMem.board_12[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _6999_ (.RESET_B(net629),
    .D(_0466_),
    .Q(\vga_tetris.boardMem.board_12[13] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _7000_ (.RESET_B(net628),
    .D(_0467_),
    .Q(\vga_tetris.boardMem.board_12[14] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _7001_ (.RESET_B(net627),
    .D(_0468_),
    .Q(\vga_tetris.boardMem.board_12[15] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _7002_ (.RESET_B(net626),
    .D(_0469_),
    .Q(\vga_tetris.boardMem.board_12[16] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _7003_ (.RESET_B(net625),
    .D(_0470_),
    .Q(\vga_tetris.boardMem.board_12[17] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _7004_ (.RESET_B(net624),
    .D(_0471_),
    .Q(\vga_tetris.boardMem.board_12[18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7005_ (.RESET_B(net623),
    .D(net1274),
    .Q(\vga_tetris.boardMem.board_12[19] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _7006_ (.RESET_B(net622),
    .D(net753),
    .Q(\vga_tetris.boardMem.board_13[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7007_ (.RESET_B(net621),
    .D(_0474_),
    .Q(\vga_tetris.boardMem.board_13[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _7008_ (.RESET_B(net620),
    .D(_0475_),
    .Q(\vga_tetris.boardMem.board_13[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _7009_ (.RESET_B(net619),
    .D(_0476_),
    .Q(\vga_tetris.boardMem.board_13[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7010_ (.RESET_B(net618),
    .D(net654),
    .Q(\vga_tetris.boardMem.board_13[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _7011_ (.RESET_B(net617),
    .D(_0478_),
    .Q(\vga_tetris.boardMem.board_13[5] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _7012_ (.RESET_B(net616),
    .D(net807),
    .Q(\vga_tetris.boardMem.board_13[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7013_ (.RESET_B(net615),
    .D(_0480_),
    .Q(\vga_tetris.boardMem.board_13[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7014_ (.RESET_B(net614),
    .D(_0481_),
    .Q(\vga_tetris.boardMem.board_13[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _7015_ (.RESET_B(net613),
    .D(_0482_),
    .Q(\vga_tetris.boardMem.board_13[9] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7016_ (.RESET_B(net612),
    .D(_0483_),
    .Q(\vga_tetris.boardMem.board_13[10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _7017_ (.RESET_B(net611),
    .D(_0484_),
    .Q(\vga_tetris.boardMem.board_13[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7018_ (.RESET_B(net610),
    .D(_0485_),
    .Q(\vga_tetris.boardMem.board_13[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7019_ (.RESET_B(net609),
    .D(_0486_),
    .Q(\vga_tetris.boardMem.board_13[13] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7020_ (.RESET_B(net608),
    .D(_0487_),
    .Q(\vga_tetris.boardMem.board_13[14] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _7021_ (.RESET_B(net607),
    .D(_0488_),
    .Q(\vga_tetris.boardMem.board_13[15] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _7022_ (.RESET_B(net606),
    .D(_0489_),
    .Q(\vga_tetris.boardMem.board_13[16] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _7023_ (.RESET_B(net605),
    .D(_0490_),
    .Q(\vga_tetris.boardMem.board_13[17] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _7024_ (.RESET_B(net604),
    .D(_0491_),
    .Q(\vga_tetris.boardMem.board_13[18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7025_ (.RESET_B(net603),
    .D(_0492_),
    .Q(\vga_tetris.boardMem.board_13[19] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _7026_ (.RESET_B(net602),
    .D(_0493_),
    .Q(\vga_tetris.boardMem.board_14[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7027_ (.RESET_B(net601),
    .D(_0494_),
    .Q(\vga_tetris.boardMem.board_14[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _7028_ (.RESET_B(net600),
    .D(_0495_),
    .Q(\vga_tetris.boardMem.board_14[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _7029_ (.RESET_B(net599),
    .D(_0496_),
    .Q(\vga_tetris.boardMem.board_14[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7030_ (.RESET_B(net598),
    .D(_0497_),
    .Q(\vga_tetris.boardMem.board_14[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _7031_ (.RESET_B(net597),
    .D(_0498_),
    .Q(\vga_tetris.boardMem.board_14[5] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _7032_ (.RESET_B(net596),
    .D(_0499_),
    .Q(\vga_tetris.boardMem.board_14[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7033_ (.RESET_B(net595),
    .D(_0500_),
    .Q(\vga_tetris.boardMem.board_14[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7034_ (.RESET_B(net594),
    .D(_0501_),
    .Q(\vga_tetris.boardMem.board_14[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _7035_ (.RESET_B(net593),
    .D(_0502_),
    .Q(\vga_tetris.boardMem.board_14[9] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7036_ (.RESET_B(net592),
    .D(_0503_),
    .Q(\vga_tetris.boardMem.board_14[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7037_ (.RESET_B(net591),
    .D(_0504_),
    .Q(\vga_tetris.boardMem.board_14[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7038_ (.RESET_B(net590),
    .D(net1373),
    .Q(\vga_tetris.boardMem.board_14[12] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _7039_ (.RESET_B(net589),
    .D(_0506_),
    .Q(\vga_tetris.boardMem.board_14[13] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7040_ (.RESET_B(net588),
    .D(_0507_),
    .Q(\vga_tetris.boardMem.board_14[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7041_ (.RESET_B(net587),
    .D(_0508_),
    .Q(\vga_tetris.boardMem.board_14[15] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _7042_ (.RESET_B(net586),
    .D(net1340),
    .Q(\vga_tetris.boardMem.board_14[16] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7043_ (.RESET_B(net585),
    .D(_0510_),
    .Q(\vga_tetris.boardMem.board_14[17] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7044_ (.RESET_B(net584),
    .D(_0511_),
    .Q(\vga_tetris.boardMem.board_14[18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7045_ (.RESET_B(net583),
    .D(_0512_),
    .Q(\vga_tetris.boardMem.board_14[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _7046_ (.RESET_B(net582),
    .D(_0513_),
    .Q(\vga_tetris.boardMem.board_15[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _7047_ (.RESET_B(net581),
    .D(net1336),
    .Q(\vga_tetris.boardMem.board_15[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _7048_ (.RESET_B(net580),
    .D(_0515_),
    .Q(\vga_tetris.boardMem.board_15[2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _7049_ (.RESET_B(net579),
    .D(_0516_),
    .Q(\vga_tetris.boardMem.board_15[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7050_ (.RESET_B(net578),
    .D(_0517_),
    .Q(\vga_tetris.boardMem.board_15[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _7051_ (.RESET_B(net577),
    .D(_0518_),
    .Q(\vga_tetris.boardMem.board_15[5] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _7052_ (.RESET_B(net576),
    .D(_0519_),
    .Q(\vga_tetris.boardMem.board_15[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _7053_ (.RESET_B(net575),
    .D(_0520_),
    .Q(\vga_tetris.boardMem.board_15[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7054_ (.RESET_B(net574),
    .D(_0521_),
    .Q(\vga_tetris.boardMem.board_15[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7055_ (.RESET_B(net573),
    .D(_0522_),
    .Q(\vga_tetris.boardMem.board_15[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _7056_ (.RESET_B(net572),
    .D(_0523_),
    .Q(\vga_tetris.boardMem.board_15[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7057_ (.RESET_B(net571),
    .D(_0524_),
    .Q(\vga_tetris.boardMem.board_15[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7058_ (.RESET_B(net570),
    .D(_0525_),
    .Q(\vga_tetris.boardMem.board_15[12] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _7059_ (.RESET_B(net569),
    .D(_0526_),
    .Q(\vga_tetris.boardMem.board_15[13] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _7060_ (.RESET_B(net568),
    .D(_0527_),
    .Q(\vga_tetris.boardMem.board_15[14] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7061_ (.RESET_B(net567),
    .D(_0528_),
    .Q(\vga_tetris.boardMem.board_15[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _7062_ (.RESET_B(net566),
    .D(net770),
    .Q(\vga_tetris.boardMem.board_15[16] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7063_ (.RESET_B(net565),
    .D(_0530_),
    .Q(\vga_tetris.boardMem.board_15[17] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7064_ (.RESET_B(net564),
    .D(_0531_),
    .Q(\vga_tetris.boardMem.board_15[18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7065_ (.RESET_B(net563),
    .D(_0532_),
    .Q(\vga_tetris.boardMem.board_15[19] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _7066_ (.RESET_B(net562),
    .D(net1592),
    .Q(\vga_tetris.boardMem.board_16[0] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _7067_ (.RESET_B(net561),
    .D(_0534_),
    .Q(\vga_tetris.boardMem.board_16[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _7068_ (.RESET_B(net560),
    .D(_0535_),
    .Q(\vga_tetris.boardMem.board_16[2] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _7069_ (.RESET_B(net559),
    .D(_0536_),
    .Q(\vga_tetris.boardMem.board_16[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7070_ (.RESET_B(net558),
    .D(_0537_),
    .Q(\vga_tetris.boardMem.board_16[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _7071_ (.RESET_B(net557),
    .D(_0538_),
    .Q(\vga_tetris.boardMem.board_16[5] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _7072_ (.RESET_B(net556),
    .D(_0539_),
    .Q(\vga_tetris.boardMem.board_16[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _7073_ (.RESET_B(net555),
    .D(_0540_),
    .Q(\vga_tetris.boardMem.board_16[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7074_ (.RESET_B(net554),
    .D(_0541_),
    .Q(\vga_tetris.boardMem.board_16[8] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7075_ (.RESET_B(net553),
    .D(_0542_),
    .Q(\vga_tetris.boardMem.board_16[9] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _7076_ (.RESET_B(net552),
    .D(_0543_),
    .Q(\vga_tetris.boardMem.board_16[10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7077_ (.RESET_B(net550),
    .D(_0544_),
    .Q(\vga_tetris.boardMem.board_16[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7078_ (.RESET_B(net548),
    .D(_0545_),
    .Q(\vga_tetris.boardMem.board_16[12] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _7079_ (.RESET_B(net519),
    .D(_0546_),
    .Q(\vga_tetris.boardMem.board_16[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _7080_ (.RESET_B(net517),
    .D(_0547_),
    .Q(\vga_tetris.boardMem.board_16[14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7081_ (.RESET_B(net515),
    .D(_0548_),
    .Q(\vga_tetris.boardMem.board_16[15] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _7082_ (.RESET_B(net513),
    .D(net1482),
    .Q(\vga_tetris.boardMem.board_16[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _7083_ (.RESET_B(net511),
    .D(_0550_),
    .Q(\vga_tetris.boardMem.board_16[17] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _7084_ (.RESET_B(net509),
    .D(_0551_),
    .Q(\vga_tetris.boardMem.board_16[18] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7085_ (.RESET_B(net507),
    .D(_0552_),
    .Q(\vga_tetris.boardMem.board_16[19] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _7086_ (.RESET_B(net505),
    .D(_0553_),
    .Q(\vga_tetris.boardMem.board_17[0] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _7087_ (.RESET_B(net503),
    .D(_0554_),
    .Q(\vga_tetris.boardMem.board_17[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _7088_ (.RESET_B(net501),
    .D(_0555_),
    .Q(\vga_tetris.boardMem.board_17[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7089_ (.RESET_B(net499),
    .D(_0556_),
    .Q(\vga_tetris.boardMem.board_17[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7090_ (.RESET_B(net497),
    .D(_0557_),
    .Q(\vga_tetris.boardMem.board_17[4] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _7091_ (.RESET_B(net487),
    .D(_0558_),
    .Q(\vga_tetris.boardMem.board_17[5] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _7092_ (.RESET_B(net485),
    .D(_0559_),
    .Q(\vga_tetris.boardMem.board_17[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7093_ (.RESET_B(net483),
    .D(_0560_),
    .Q(\vga_tetris.boardMem.board_17[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7094_ (.RESET_B(net481),
    .D(_0561_),
    .Q(\vga_tetris.boardMem.board_17[8] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _7095_ (.RESET_B(net479),
    .D(net1558),
    .Q(\vga_tetris.boardMem.board_17[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _7096_ (.RESET_B(net477),
    .D(net1419),
    .Q(\vga_tetris.boardMem.board_17[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7097_ (.RESET_B(net475),
    .D(_0564_),
    .Q(\vga_tetris.boardMem.board_17[11] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7098_ (.RESET_B(net473),
    .D(_0565_),
    .Q(\vga_tetris.boardMem.board_17[12] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _7099_ (.RESET_B(net471),
    .D(_0566_),
    .Q(\vga_tetris.boardMem.board_17[13] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _7100_ (.RESET_B(net469),
    .D(_0567_),
    .Q(\vga_tetris.boardMem.board_17[14] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _7101_ (.RESET_B(net467),
    .D(_0568_),
    .Q(\vga_tetris.boardMem.board_17[15] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _7102_ (.RESET_B(net465),
    .D(_0569_),
    .Q(\vga_tetris.boardMem.board_17[16] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _7103_ (.RESET_B(net463),
    .D(net1580),
    .Q(\vga_tetris.boardMem.board_17[17] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _7104_ (.RESET_B(net461),
    .D(net1444),
    .Q(\vga_tetris.boardMem.board_17[18] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7105_ (.RESET_B(net459),
    .D(_0572_),
    .Q(\vga_tetris.boardMem.board_17[19] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _7106_ (.RESET_B(net457),
    .D(net1545),
    .Q(\vga_tetris.boardMem.board_18[0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _7107_ (.RESET_B(net452),
    .D(net1434),
    .Q(\vga_tetris.boardMem.board_18[1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _7108_ (.RESET_B(net450),
    .D(_0575_),
    .Q(\vga_tetris.boardMem.board_18[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _7109_ (.RESET_B(net448),
    .D(_0576_),
    .Q(\vga_tetris.boardMem.board_18[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7110_ (.RESET_B(net446),
    .D(_0577_),
    .Q(\vga_tetris.boardMem.board_18[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7111_ (.RESET_B(net444),
    .D(_0578_),
    .Q(\vga_tetris.boardMem.board_18[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7112_ (.RESET_B(net442),
    .D(_0579_),
    .Q(\vga_tetris.boardMem.board_18[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7113_ (.RESET_B(net440),
    .D(_0580_),
    .Q(\vga_tetris.boardMem.board_18[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7114_ (.RESET_B(net438),
    .D(net1567),
    .Q(\vga_tetris.boardMem.board_18[8] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7115_ (.RESET_B(net436),
    .D(_0582_),
    .Q(\vga_tetris.boardMem.board_18[9] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7116_ (.RESET_B(net434),
    .D(net1465),
    .Q(\vga_tetris.boardMem.board_18[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7117_ (.RESET_B(net432),
    .D(_0584_),
    .Q(\vga_tetris.boardMem.board_18[11] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _7118_ (.RESET_B(net430),
    .D(_0585_),
    .Q(\vga_tetris.boardMem.board_18[12] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _7119_ (.RESET_B(net428),
    .D(_0586_),
    .Q(\vga_tetris.boardMem.board_18[13] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _7120_ (.RESET_B(net426),
    .D(_0587_),
    .Q(\vga_tetris.boardMem.board_18[14] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7121_ (.RESET_B(net424),
    .D(_0588_),
    .Q(\vga_tetris.boardMem.board_18[15] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7122_ (.RESET_B(net422),
    .D(_0589_),
    .Q(\vga_tetris.boardMem.board_18[16] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7123_ (.RESET_B(net420),
    .D(net1531),
    .Q(\vga_tetris.boardMem.board_18[17] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _7124_ (.RESET_B(net418),
    .D(_0591_),
    .Q(\vga_tetris.boardMem.board_18[18] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7125_ (.RESET_B(net416),
    .D(_0592_),
    .Q(\vga_tetris.boardMem.board_18[19] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _7126_ (.RESET_B(net414),
    .D(net1711),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _7127_ (.RESET_B(net412),
    .D(net1604),
    .Q(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7128_ (.RESET_B(net405),
    .D(_0595_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7129_ (.RESET_B(net390),
    .D(_0596_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7130_ (.RESET_B(net386),
    .D(net1600),
    .Q(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7131_ (.RESET_B(net382),
    .D(_0598_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7132_ (.RESET_B(net375),
    .D(_0599_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7133_ (.RESET_B(net371),
    .D(_0600_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7134_ (.RESET_B(net367),
    .D(_0601_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _7135_ (.RESET_B(net363),
    .D(net1691),
    .Q(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7136_ (.RESET_B(net359),
    .D(_0603_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7137_ (.RESET_B(net355),
    .D(_0604_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7138_ (.RESET_B(net351),
    .D(_0605_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _7139_ (.RESET_B(net347),
    .D(_0606_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7140_ (.RESET_B(net343),
    .D(net1820),
    .Q(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _7141_ (.RESET_B(net339),
    .D(_0608_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7142_ (.RESET_B(net331),
    .D(net1862),
    .Q(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7143_ (.RESET_B(net410),
    .D(_0610_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7144_ (.RESET_B(net388),
    .D(_0611_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _7145_ (.RESET_B(net377),
    .D(net1778),
    .Q(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7146_ (.RESET_B(net369),
    .D(_0613_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _7147_ (.RESET_B(net361),
    .D(_0614_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7148_ (.RESET_B(net353),
    .D(_0615_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7149_ (.RESET_B(net345),
    .D(_0616_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _7150_ (.RESET_B(net333),
    .D(_0617_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7151_ (.RESET_B(net403),
    .D(_0618_),
    .Q(\vga_tetris._tetrisDisplay_io_boardYCoord[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7152_ (.RESET_B(net373),
    .D(_0619_),
    .Q(\vga_tetris._tetrisDisplay_io_boardYCoord[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7153_ (.RESET_B(net357),
    .D(_0620_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7154_ (.RESET_B(net341),
    .D(net1758),
    .Q(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7155_ (.RESET_B(net384),
    .D(net1849),
    .Q(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _7156_ (.RESET_B(net349),
    .D(_0623_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7157_ (.RESET_B(net365),
    .D(_0624_),
    .Q(\vga_tetris.runningTetrisLogicQ ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_tiehi _6981__22 (.L_HI(net22));
 sg13g2_tiehi _6980__23 (.L_HI(net23));
 sg13g2_tiehi _6979__24 (.L_HI(net24));
 sg13g2_tiehi _6978__25 (.L_HI(net25));
 sg13g2_tiehi _6977__26 (.L_HI(net26));
 sg13g2_tiehi _6976__27 (.L_HI(net27));
 sg13g2_tiehi _6975__28 (.L_HI(net28));
 sg13g2_tiehi _6974__29 (.L_HI(net29));
 sg13g2_tiehi _6973__30 (.L_HI(net30));
 sg13g2_tiehi _6972__31 (.L_HI(net31));
 sg13g2_tiehi _6971__32 (.L_HI(net32));
 sg13g2_tiehi _6970__33 (.L_HI(net33));
 sg13g2_tiehi _6969__34 (.L_HI(net34));
 sg13g2_tiehi _6968__35 (.L_HI(net35));
 sg13g2_tiehi _6967__36 (.L_HI(net36));
 sg13g2_tiehi _6966__37 (.L_HI(net37));
 sg13g2_tiehi _6965__38 (.L_HI(net38));
 sg13g2_tiehi _6964__39 (.L_HI(net39));
 sg13g2_tiehi _6963__40 (.L_HI(net40));
 sg13g2_tiehi _6962__41 (.L_HI(net41));
 sg13g2_tiehi _6961__42 (.L_HI(net42));
 sg13g2_tiehi _6960__43 (.L_HI(net43));
 sg13g2_tiehi _6959__44 (.L_HI(net44));
 sg13g2_tiehi _6958__45 (.L_HI(net45));
 sg13g2_tiehi _6957__46 (.L_HI(net46));
 sg13g2_tiehi _6956__47 (.L_HI(net47));
 sg13g2_tiehi _6955__48 (.L_HI(net48));
 sg13g2_tiehi _6954__49 (.L_HI(net49));
 sg13g2_tiehi _6953__50 (.L_HI(net50));
 sg13g2_tiehi _6952__51 (.L_HI(net51));
 sg13g2_tiehi _6951__52 (.L_HI(net52));
 sg13g2_tiehi _6950__53 (.L_HI(net53));
 sg13g2_tiehi _6949__54 (.L_HI(net54));
 sg13g2_tiehi _6948__55 (.L_HI(net55));
 sg13g2_tiehi _6947__56 (.L_HI(net56));
 sg13g2_tiehi _6946__57 (.L_HI(net57));
 sg13g2_tiehi _6945__58 (.L_HI(net58));
 sg13g2_tiehi _6944__59 (.L_HI(net59));
 sg13g2_tiehi _6943__60 (.L_HI(net60));
 sg13g2_tiehi _6942__61 (.L_HI(net61));
 sg13g2_tiehi _6941__62 (.L_HI(net62));
 sg13g2_tiehi _6940__63 (.L_HI(net63));
 sg13g2_tiehi _6939__64 (.L_HI(net64));
 sg13g2_tiehi _6938__65 (.L_HI(net65));
 sg13g2_tiehi _6937__66 (.L_HI(net66));
 sg13g2_tiehi _6936__67 (.L_HI(net67));
 sg13g2_tiehi _6935__68 (.L_HI(net68));
 sg13g2_tiehi _6934__69 (.L_HI(net69));
 sg13g2_tiehi _6933__70 (.L_HI(net70));
 sg13g2_tiehi _6932__71 (.L_HI(net71));
 sg13g2_tiehi _6931__72 (.L_HI(net72));
 sg13g2_tiehi _6930__73 (.L_HI(net73));
 sg13g2_tiehi _6929__74 (.L_HI(net74));
 sg13g2_tiehi _6928__75 (.L_HI(net75));
 sg13g2_tiehi _6927__76 (.L_HI(net76));
 sg13g2_tiehi _6926__77 (.L_HI(net77));
 sg13g2_tiehi _6925__78 (.L_HI(net78));
 sg13g2_tiehi _6924__79 (.L_HI(net79));
 sg13g2_tiehi _6923__80 (.L_HI(net80));
 sg13g2_tiehi _6922__81 (.L_HI(net81));
 sg13g2_tiehi _6921__82 (.L_HI(net82));
 sg13g2_tiehi _6920__83 (.L_HI(net83));
 sg13g2_tiehi _6919__84 (.L_HI(net84));
 sg13g2_tiehi _6918__85 (.L_HI(net85));
 sg13g2_tiehi _6917__86 (.L_HI(net86));
 sg13g2_tiehi _6916__87 (.L_HI(net87));
 sg13g2_tiehi _6915__88 (.L_HI(net88));
 sg13g2_tiehi _6914__89 (.L_HI(net89));
 sg13g2_tiehi _6913__90 (.L_HI(net90));
 sg13g2_tiehi _6912__91 (.L_HI(net91));
 sg13g2_tiehi _6911__92 (.L_HI(net92));
 sg13g2_tiehi _6910__93 (.L_HI(net93));
 sg13g2_tiehi _6909__94 (.L_HI(net94));
 sg13g2_tiehi _6908__95 (.L_HI(net95));
 sg13g2_tiehi _6907__96 (.L_HI(net96));
 sg13g2_tiehi _6906__97 (.L_HI(net97));
 sg13g2_tiehi _6905__98 (.L_HI(net98));
 sg13g2_tiehi _6904__99 (.L_HI(net99));
 sg13g2_tiehi _6903__100 (.L_HI(net100));
 sg13g2_tiehi _6902__101 (.L_HI(net101));
 sg13g2_tiehi _6901__102 (.L_HI(net102));
 sg13g2_tiehi _6900__103 (.L_HI(net103));
 sg13g2_tiehi _6899__104 (.L_HI(net104));
 sg13g2_tiehi _6898__105 (.L_HI(net105));
 sg13g2_tiehi _6897__106 (.L_HI(net106));
 sg13g2_tiehi _6896__107 (.L_HI(net107));
 sg13g2_tiehi _6895__108 (.L_HI(net108));
 sg13g2_tiehi _6894__109 (.L_HI(net109));
 sg13g2_tiehi _6893__110 (.L_HI(net110));
 sg13g2_tiehi _6892__111 (.L_HI(net111));
 sg13g2_tiehi _6891__112 (.L_HI(net112));
 sg13g2_tiehi _6890__113 (.L_HI(net113));
 sg13g2_tiehi _6889__114 (.L_HI(net114));
 sg13g2_tiehi _6888__115 (.L_HI(net115));
 sg13g2_tiehi _6887__116 (.L_HI(net116));
 sg13g2_tiehi _6886__117 (.L_HI(net117));
 sg13g2_tiehi _6885__118 (.L_HI(net118));
 sg13g2_tiehi _6884__119 (.L_HI(net119));
 sg13g2_tiehi _6883__120 (.L_HI(net120));
 sg13g2_tiehi _6882__121 (.L_HI(net121));
 sg13g2_tiehi _6881__122 (.L_HI(net122));
 sg13g2_tiehi _6880__123 (.L_HI(net123));
 sg13g2_tiehi _6879__124 (.L_HI(net124));
 sg13g2_tiehi _6878__125 (.L_HI(net125));
 sg13g2_tiehi _6877__126 (.L_HI(net126));
 sg13g2_tiehi _6876__127 (.L_HI(net127));
 sg13g2_tiehi _6875__128 (.L_HI(net128));
 sg13g2_tiehi _6874__129 (.L_HI(net129));
 sg13g2_tiehi _6873__130 (.L_HI(net130));
 sg13g2_tiehi _6872__131 (.L_HI(net131));
 sg13g2_tiehi _6871__132 (.L_HI(net132));
 sg13g2_tiehi _6870__133 (.L_HI(net133));
 sg13g2_tiehi _6869__134 (.L_HI(net134));
 sg13g2_tiehi _6868__135 (.L_HI(net135));
 sg13g2_tiehi _6867__136 (.L_HI(net136));
 sg13g2_tiehi _6866__137 (.L_HI(net137));
 sg13g2_tiehi _6865__138 (.L_HI(net138));
 sg13g2_tiehi _6864__139 (.L_HI(net139));
 sg13g2_tiehi _6863__140 (.L_HI(net140));
 sg13g2_tiehi _6862__141 (.L_HI(net141));
 sg13g2_tiehi _6861__142 (.L_HI(net142));
 sg13g2_tiehi _6860__143 (.L_HI(net143));
 sg13g2_tiehi _6859__144 (.L_HI(net144));
 sg13g2_tiehi _6858__145 (.L_HI(net145));
 sg13g2_tiehi _6857__146 (.L_HI(net146));
 sg13g2_tiehi _6856__147 (.L_HI(net147));
 sg13g2_tiehi _6855__148 (.L_HI(net148));
 sg13g2_tiehi _6854__149 (.L_HI(net149));
 sg13g2_tiehi _6853__150 (.L_HI(net150));
 sg13g2_tiehi _6852__151 (.L_HI(net151));
 sg13g2_tiehi _6851__152 (.L_HI(net152));
 sg13g2_tiehi _6850__153 (.L_HI(net153));
 sg13g2_tiehi _6849__154 (.L_HI(net154));
 sg13g2_tiehi _6848__155 (.L_HI(net155));
 sg13g2_tiehi _6847__156 (.L_HI(net156));
 sg13g2_tiehi _6846__157 (.L_HI(net157));
 sg13g2_tiehi _6845__158 (.L_HI(net158));
 sg13g2_tiehi _6844__159 (.L_HI(net159));
 sg13g2_tiehi _6843__160 (.L_HI(net160));
 sg13g2_tiehi _6842__161 (.L_HI(net161));
 sg13g2_tiehi _6841__162 (.L_HI(net162));
 sg13g2_tiehi _6840__163 (.L_HI(net163));
 sg13g2_tiehi _6839__164 (.L_HI(net164));
 sg13g2_tiehi _6838__165 (.L_HI(net165));
 sg13g2_tiehi _6837__166 (.L_HI(net166));
 sg13g2_tiehi _6836__167 (.L_HI(net167));
 sg13g2_tiehi _6835__168 (.L_HI(net168));
 sg13g2_tiehi _6834__169 (.L_HI(net169));
 sg13g2_tiehi _6833__170 (.L_HI(net170));
 sg13g2_tiehi _6832__171 (.L_HI(net171));
 sg13g2_tiehi _6831__172 (.L_HI(net172));
 sg13g2_tiehi _6830__173 (.L_HI(net173));
 sg13g2_tiehi _6829__174 (.L_HI(net174));
 sg13g2_tiehi _6828__175 (.L_HI(net175));
 sg13g2_tiehi _6827__176 (.L_HI(net176));
 sg13g2_tiehi _6826__177 (.L_HI(net177));
 sg13g2_tiehi _6825__178 (.L_HI(net178));
 sg13g2_tiehi _6824__179 (.L_HI(net179));
 sg13g2_tiehi _6823__180 (.L_HI(net180));
 sg13g2_tiehi _6822__181 (.L_HI(net181));
 sg13g2_tiehi _6821__182 (.L_HI(net182));
 sg13g2_tiehi _6820__183 (.L_HI(net183));
 sg13g2_tiehi _6819__184 (.L_HI(net184));
 sg13g2_tiehi _6818__185 (.L_HI(net185));
 sg13g2_tiehi _6817__186 (.L_HI(net186));
 sg13g2_tiehi _6816__187 (.L_HI(net187));
 sg13g2_tiehi _6815__188 (.L_HI(net188));
 sg13g2_tiehi _6814__189 (.L_HI(net189));
 sg13g2_tiehi _6813__190 (.L_HI(net190));
 sg13g2_tiehi _6812__191 (.L_HI(net191));
 sg13g2_tiehi _6811__192 (.L_HI(net192));
 sg13g2_tiehi _6810__193 (.L_HI(net193));
 sg13g2_tiehi _6809__194 (.L_HI(net194));
 sg13g2_tiehi _6808__195 (.L_HI(net195));
 sg13g2_tiehi _6807__196 (.L_HI(net196));
 sg13g2_tiehi _6806__197 (.L_HI(net197));
 sg13g2_tiehi _6805__198 (.L_HI(net198));
 sg13g2_tiehi _6804__199 (.L_HI(net199));
 sg13g2_tiehi _6803__200 (.L_HI(net200));
 sg13g2_tiehi _6802__201 (.L_HI(net201));
 sg13g2_tiehi _6801__202 (.L_HI(net202));
 sg13g2_tiehi _6800__203 (.L_HI(net203));
 sg13g2_tiehi _6799__204 (.L_HI(net204));
 sg13g2_tiehi _6798__205 (.L_HI(net205));
 sg13g2_tiehi _6797__206 (.L_HI(net206));
 sg13g2_tiehi _6796__207 (.L_HI(net207));
 sg13g2_tiehi _6795__208 (.L_HI(net208));
 sg13g2_tiehi _6794__209 (.L_HI(net209));
 sg13g2_tiehi _6793__210 (.L_HI(net210));
 sg13g2_tiehi _6792__211 (.L_HI(net211));
 sg13g2_tiehi _6791__212 (.L_HI(net212));
 sg13g2_tiehi _6790__213 (.L_HI(net213));
 sg13g2_tiehi _6789__214 (.L_HI(net214));
 sg13g2_tiehi _6788__215 (.L_HI(net215));
 sg13g2_tiehi _6787__216 (.L_HI(net216));
 sg13g2_tiehi _6786__217 (.L_HI(net217));
 sg13g2_tiehi _6785__218 (.L_HI(net218));
 sg13g2_tiehi _6784__219 (.L_HI(net219));
 sg13g2_tiehi _6783__220 (.L_HI(net220));
 sg13g2_tiehi _6782__221 (.L_HI(net221));
 sg13g2_tiehi _6781__222 (.L_HI(net222));
 sg13g2_tiehi _6780__223 (.L_HI(net223));
 sg13g2_tiehi _6779__224 (.L_HI(net224));
 sg13g2_tiehi _6778__225 (.L_HI(net225));
 sg13g2_tiehi _6777__226 (.L_HI(net226));
 sg13g2_tiehi _6776__227 (.L_HI(net227));
 sg13g2_tiehi _6775__228 (.L_HI(net228));
 sg13g2_tiehi _6774__229 (.L_HI(net229));
 sg13g2_tiehi _6773__230 (.L_HI(net230));
 sg13g2_tiehi _6772__231 (.L_HI(net231));
 sg13g2_tiehi _6771__232 (.L_HI(net232));
 sg13g2_tiehi _6770__233 (.L_HI(net233));
 sg13g2_tiehi _6769__234 (.L_HI(net234));
 sg13g2_tiehi _6768__235 (.L_HI(net235));
 sg13g2_tiehi _6767__236 (.L_HI(net236));
 sg13g2_tiehi _6766__237 (.L_HI(net237));
 sg13g2_tiehi _6765__238 (.L_HI(net238));
 sg13g2_tiehi _6764__239 (.L_HI(net239));
 sg13g2_tiehi _6763__240 (.L_HI(net240));
 sg13g2_tiehi _6762__241 (.L_HI(net241));
 sg13g2_tiehi _6761__242 (.L_HI(net242));
 sg13g2_tiehi _6760__243 (.L_HI(net243));
 sg13g2_tiehi _6759__244 (.L_HI(net244));
 sg13g2_tiehi _6758__245 (.L_HI(net245));
 sg13g2_tiehi _6757__246 (.L_HI(net246));
 sg13g2_tiehi _6756__247 (.L_HI(net247));
 sg13g2_tiehi _6755__248 (.L_HI(net248));
 sg13g2_tiehi _6754__249 (.L_HI(net249));
 sg13g2_tiehi _6753__250 (.L_HI(net250));
 sg13g2_tiehi _6752__251 (.L_HI(net251));
 sg13g2_tiehi _6751__252 (.L_HI(net252));
 sg13g2_tiehi _6750__253 (.L_HI(net253));
 sg13g2_tiehi _6749__254 (.L_HI(net254));
 sg13g2_tiehi _6748__255 (.L_HI(net255));
 sg13g2_tiehi _6747__256 (.L_HI(net256));
 sg13g2_tiehi _6746__257 (.L_HI(net257));
 sg13g2_tiehi _6745__258 (.L_HI(net258));
 sg13g2_tiehi _6744__259 (.L_HI(net259));
 sg13g2_tiehi _6743__260 (.L_HI(net260));
 sg13g2_tiehi _6742__261 (.L_HI(net261));
 sg13g2_tiehi _6741__262 (.L_HI(net262));
 sg13g2_tiehi _6740__263 (.L_HI(net263));
 sg13g2_tiehi _6739__264 (.L_HI(net264));
 sg13g2_tiehi _6738__265 (.L_HI(net265));
 sg13g2_tiehi _6737__266 (.L_HI(net266));
 sg13g2_tiehi _6736__267 (.L_HI(net267));
 sg13g2_tiehi _6735__268 (.L_HI(net268));
 sg13g2_tiehi _6734__269 (.L_HI(net269));
 sg13g2_tiehi _6733__270 (.L_HI(net270));
 sg13g2_tiehi _6732__271 (.L_HI(net271));
 sg13g2_tiehi _6731__272 (.L_HI(net272));
 sg13g2_tiehi _6730__273 (.L_HI(net273));
 sg13g2_tiehi _6729__274 (.L_HI(net274));
 sg13g2_tiehi _6728__275 (.L_HI(net275));
 sg13g2_tiehi _6727__276 (.L_HI(net276));
 sg13g2_tiehi _6726__277 (.L_HI(net277));
 sg13g2_tiehi _6725__278 (.L_HI(net278));
 sg13g2_tiehi _6724__279 (.L_HI(net279));
 sg13g2_tiehi _6723__280 (.L_HI(net280));
 sg13g2_tiehi _6722__281 (.L_HI(net281));
 sg13g2_tiehi _6721__282 (.L_HI(net282));
 sg13g2_tiehi _6720__283 (.L_HI(net283));
 sg13g2_tiehi _6719__284 (.L_HI(net284));
 sg13g2_tiehi _6718__285 (.L_HI(net285));
 sg13g2_tiehi _6717__286 (.L_HI(net286));
 sg13g2_tiehi _6716__287 (.L_HI(net287));
 sg13g2_tiehi _6715__288 (.L_HI(net288));
 sg13g2_tiehi _6714__289 (.L_HI(net289));
 sg13g2_tiehi _6713__290 (.L_HI(net290));
 sg13g2_tiehi _6712__291 (.L_HI(net291));
 sg13g2_tiehi _6711__292 (.L_HI(net292));
 sg13g2_tiehi _6710__293 (.L_HI(net293));
 sg13g2_tiehi _6709__294 (.L_HI(net294));
 sg13g2_tiehi _6708__295 (.L_HI(net295));
 sg13g2_tiehi _6707__296 (.L_HI(net296));
 sg13g2_tiehi _6706__297 (.L_HI(net297));
 sg13g2_tiehi _6705__298 (.L_HI(net298));
 sg13g2_tiehi _6704__299 (.L_HI(net299));
 sg13g2_tiehi _6703__300 (.L_HI(net300));
 sg13g2_tiehi _6702__301 (.L_HI(net301));
 sg13g2_tiehi _6701__302 (.L_HI(net302));
 sg13g2_tiehi _6700__303 (.L_HI(net303));
 sg13g2_tiehi _6699__304 (.L_HI(net304));
 sg13g2_tiehi _6698__305 (.L_HI(net305));
 sg13g2_tiehi _6697__306 (.L_HI(net306));
 sg13g2_tiehi _6696__307 (.L_HI(net307));
 sg13g2_tiehi _6695__308 (.L_HI(net308));
 sg13g2_tiehi _6694__309 (.L_HI(net309));
 sg13g2_tiehi _6693__310 (.L_HI(net310));
 sg13g2_tiehi _6692__311 (.L_HI(net311));
 sg13g2_tiehi _6691__312 (.L_HI(net312));
 sg13g2_tiehi _6690__313 (.L_HI(net313));
 sg13g2_tiehi _6689__314 (.L_HI(net314));
 sg13g2_tiehi _6688__315 (.L_HI(net315));
 sg13g2_tiehi _6687__316 (.L_HI(net316));
 sg13g2_tiehi _6686__317 (.L_HI(net317));
 sg13g2_tiehi _6685__318 (.L_HI(net318));
 sg13g2_tiehi _6684__319 (.L_HI(net319));
 sg13g2_tiehi _6683__320 (.L_HI(net320));
 sg13g2_tiehi _6682__321 (.L_HI(net321));
 sg13g2_tiehi _6681__322 (.L_HI(net322));
 sg13g2_tiehi _6680__323 (.L_HI(net323));
 sg13g2_tiehi _6679__324 (.L_HI(net324));
 sg13g2_tiehi _6678__325 (.L_HI(net325));
 sg13g2_tiehi _6677__326 (.L_HI(net326));
 sg13g2_tiehi _6676__327 (.L_HI(net327));
 sg13g2_tiehi _6675__328 (.L_HI(net328));
 sg13g2_tiehi _6533__329 (.L_HI(net329));
 sg13g2_tiehi _6674__330 (.L_HI(net330));
 sg13g2_tiehi _7142__331 (.L_HI(net331));
 sg13g2_tiehi _6673__332 (.L_HI(net332));
 sg13g2_tiehi _7150__333 (.L_HI(net333));
 sg13g2_tiehi _6672__334 (.L_HI(net334));
 sg13g2_tiehi _6671__335 (.L_HI(net335));
 sg13g2_tiehi _6670__336 (.L_HI(net336));
 sg13g2_tiehi _6669__337 (.L_HI(net337));
 sg13g2_tiehi _6668__338 (.L_HI(net338));
 sg13g2_tiehi _7141__339 (.L_HI(net339));
 sg13g2_tiehi _6667__340 (.L_HI(net340));
 sg13g2_tiehi _7154__341 (.L_HI(net341));
 sg13g2_tiehi _6666__342 (.L_HI(net342));
 sg13g2_tiehi _7140__343 (.L_HI(net343));
 sg13g2_tiehi _6665__344 (.L_HI(net344));
 sg13g2_tiehi _7149__345 (.L_HI(net345));
 sg13g2_tiehi _6664__346 (.L_HI(net346));
 sg13g2_tiehi _7139__347 (.L_HI(net347));
 sg13g2_tiehi _6663__348 (.L_HI(net348));
 sg13g2_tiehi _7156__349 (.L_HI(net349));
 sg13g2_tiehi _6662__350 (.L_HI(net350));
 sg13g2_tiehi _7138__351 (.L_HI(net351));
 sg13g2_tiehi _6661__352 (.L_HI(net352));
 sg13g2_tiehi _7148__353 (.L_HI(net353));
 sg13g2_tiehi _6660__354 (.L_HI(net354));
 sg13g2_tiehi _7137__355 (.L_HI(net355));
 sg13g2_tiehi _6659__356 (.L_HI(net356));
 sg13g2_tiehi _7153__357 (.L_HI(net357));
 sg13g2_tiehi _6658__358 (.L_HI(net358));
 sg13g2_tiehi _7136__359 (.L_HI(net359));
 sg13g2_tiehi _6657__360 (.L_HI(net360));
 sg13g2_tiehi _7147__361 (.L_HI(net361));
 sg13g2_tiehi _6656__362 (.L_HI(net362));
 sg13g2_tiehi _7135__363 (.L_HI(net363));
 sg13g2_tiehi _6655__364 (.L_HI(net364));
 sg13g2_tiehi _7157__365 (.L_HI(net365));
 sg13g2_tiehi _6654__366 (.L_HI(net366));
 sg13g2_tiehi _7134__367 (.L_HI(net367));
 sg13g2_tiehi _6653__368 (.L_HI(net368));
 sg13g2_tiehi _7146__369 (.L_HI(net369));
 sg13g2_tiehi _6652__370 (.L_HI(net370));
 sg13g2_tiehi _7133__371 (.L_HI(net371));
 sg13g2_tiehi _6651__372 (.L_HI(net372));
 sg13g2_tiehi _7152__373 (.L_HI(net373));
 sg13g2_tiehi _6650__374 (.L_HI(net374));
 sg13g2_tiehi _7132__375 (.L_HI(net375));
 sg13g2_tiehi _6649__376 (.L_HI(net376));
 sg13g2_tiehi _7145__377 (.L_HI(net377));
 sg13g2_tiehi _6648__378 (.L_HI(net378));
 sg13g2_tiehi _6647__379 (.L_HI(net379));
 sg13g2_tiehi _6646__380 (.L_HI(net380));
 sg13g2_tiehi _6645__381 (.L_HI(net381));
 sg13g2_tiehi _7131__382 (.L_HI(net382));
 sg13g2_tiehi _6644__383 (.L_HI(net383));
 sg13g2_tiehi _7155__384 (.L_HI(net384));
 sg13g2_tiehi _6643__385 (.L_HI(net385));
 sg13g2_tiehi _7130__386 (.L_HI(net386));
 sg13g2_tiehi _6642__387 (.L_HI(net387));
 sg13g2_tiehi _7144__388 (.L_HI(net388));
 sg13g2_tiehi _6641__389 (.L_HI(net389));
 sg13g2_tiehi _7129__390 (.L_HI(net390));
 sg13g2_tiehi _6640__391 (.L_HI(net391));
 sg13g2_tiehi _6639__392 (.L_HI(net392));
 sg13g2_tiehi _6638__393 (.L_HI(net393));
 sg13g2_tiehi _6637__394 (.L_HI(net394));
 sg13g2_tiehi _6636__395 (.L_HI(net395));
 sg13g2_tiehi _6635__396 (.L_HI(net396));
 sg13g2_tiehi _6634__397 (.L_HI(net397));
 sg13g2_tiehi _6633__398 (.L_HI(net398));
 sg13g2_tiehi _6632__399 (.L_HI(net399));
 sg13g2_tiehi _6631__400 (.L_HI(net400));
 sg13g2_tiehi _6630__401 (.L_HI(net401));
 sg13g2_tiehi _6629__402 (.L_HI(net402));
 sg13g2_tiehi _7151__403 (.L_HI(net403));
 sg13g2_tiehi _6628__404 (.L_HI(net404));
 sg13g2_tiehi _7128__405 (.L_HI(net405));
 sg13g2_tiehi _6627__406 (.L_HI(net406));
 sg13g2_tiehi _6626__407 (.L_HI(net407));
 sg13g2_tiehi _6625__408 (.L_HI(net408));
 sg13g2_tiehi _6624__409 (.L_HI(net409));
 sg13g2_tiehi _7143__410 (.L_HI(net410));
 sg13g2_tiehi _6623__411 (.L_HI(net411));
 sg13g2_tiehi _7127__412 (.L_HI(net412));
 sg13g2_tiehi _6622__413 (.L_HI(net413));
 sg13g2_tiehi _7126__414 (.L_HI(net414));
 sg13g2_tiehi _6621__415 (.L_HI(net415));
 sg13g2_tiehi _7125__416 (.L_HI(net416));
 sg13g2_tiehi _6620__417 (.L_HI(net417));
 sg13g2_tiehi _7124__418 (.L_HI(net418));
 sg13g2_tiehi _6619__419 (.L_HI(net419));
 sg13g2_tiehi _7123__420 (.L_HI(net420));
 sg13g2_tiehi _6618__421 (.L_HI(net421));
 sg13g2_tiehi _7122__422 (.L_HI(net422));
 sg13g2_tiehi _6617__423 (.L_HI(net423));
 sg13g2_tiehi _7121__424 (.L_HI(net424));
 sg13g2_tiehi _6616__425 (.L_HI(net425));
 sg13g2_tiehi _7120__426 (.L_HI(net426));
 sg13g2_tiehi _6615__427 (.L_HI(net427));
 sg13g2_tiehi _7119__428 (.L_HI(net428));
 sg13g2_tiehi _6614__429 (.L_HI(net429));
 sg13g2_tiehi _7118__430 (.L_HI(net430));
 sg13g2_tiehi _6613__431 (.L_HI(net431));
 sg13g2_tiehi _7117__432 (.L_HI(net432));
 sg13g2_tiehi _6612__433 (.L_HI(net433));
 sg13g2_tiehi _7116__434 (.L_HI(net434));
 sg13g2_tiehi _6611__435 (.L_HI(net435));
 sg13g2_tiehi _7115__436 (.L_HI(net436));
 sg13g2_tiehi _6610__437 (.L_HI(net437));
 sg13g2_tiehi _7114__438 (.L_HI(net438));
 sg13g2_tiehi _6609__439 (.L_HI(net439));
 sg13g2_tiehi _7113__440 (.L_HI(net440));
 sg13g2_tiehi _6608__441 (.L_HI(net441));
 sg13g2_tiehi _7112__442 (.L_HI(net442));
 sg13g2_tiehi _6607__443 (.L_HI(net443));
 sg13g2_tiehi _7111__444 (.L_HI(net444));
 sg13g2_tiehi _6606__445 (.L_HI(net445));
 sg13g2_tiehi _7110__446 (.L_HI(net446));
 sg13g2_tiehi _6605__447 (.L_HI(net447));
 sg13g2_tiehi _7109__448 (.L_HI(net448));
 sg13g2_tiehi _6604__449 (.L_HI(net449));
 sg13g2_tiehi _7108__450 (.L_HI(net450));
 sg13g2_tiehi _6603__451 (.L_HI(net451));
 sg13g2_tiehi _7107__452 (.L_HI(net452));
 sg13g2_tiehi _6602__453 (.L_HI(net453));
 sg13g2_tiehi _6601__454 (.L_HI(net454));
 sg13g2_tiehi _6600__455 (.L_HI(net455));
 sg13g2_tiehi _6599__456 (.L_HI(net456));
 sg13g2_tiehi _7106__457 (.L_HI(net457));
 sg13g2_tiehi _6598__458 (.L_HI(net458));
 sg13g2_tiehi _7105__459 (.L_HI(net459));
 sg13g2_tiehi _6597__460 (.L_HI(net460));
 sg13g2_tiehi _7104__461 (.L_HI(net461));
 sg13g2_tiehi _6596__462 (.L_HI(net462));
 sg13g2_tiehi _7103__463 (.L_HI(net463));
 sg13g2_tiehi _6595__464 (.L_HI(net464));
 sg13g2_tiehi _7102__465 (.L_HI(net465));
 sg13g2_tiehi _6594__466 (.L_HI(net466));
 sg13g2_tiehi _7101__467 (.L_HI(net467));
 sg13g2_tiehi _6593__468 (.L_HI(net468));
 sg13g2_tiehi _7100__469 (.L_HI(net469));
 sg13g2_tiehi _6592__470 (.L_HI(net470));
 sg13g2_tiehi _7099__471 (.L_HI(net471));
 sg13g2_tiehi _6591__472 (.L_HI(net472));
 sg13g2_tiehi _7098__473 (.L_HI(net473));
 sg13g2_tiehi _6590__474 (.L_HI(net474));
 sg13g2_tiehi _7097__475 (.L_HI(net475));
 sg13g2_tiehi _6589__476 (.L_HI(net476));
 sg13g2_tiehi _7096__477 (.L_HI(net477));
 sg13g2_tiehi _6588__478 (.L_HI(net478));
 sg13g2_tiehi _7095__479 (.L_HI(net479));
 sg13g2_tiehi _6587__480 (.L_HI(net480));
 sg13g2_tiehi _7094__481 (.L_HI(net481));
 sg13g2_tiehi _6586__482 (.L_HI(net482));
 sg13g2_tiehi _7093__483 (.L_HI(net483));
 sg13g2_tiehi _6585__484 (.L_HI(net484));
 sg13g2_tiehi _7092__485 (.L_HI(net485));
 sg13g2_tiehi _6584__486 (.L_HI(net486));
 sg13g2_tiehi _7091__487 (.L_HI(net487));
 sg13g2_tiehi _6583__488 (.L_HI(net488));
 sg13g2_tiehi _6582__489 (.L_HI(net489));
 sg13g2_tiehi _6581__490 (.L_HI(net490));
 sg13g2_tiehi _6580__491 (.L_HI(net491));
 sg13g2_tiehi _6579__492 (.L_HI(net492));
 sg13g2_tiehi _6578__493 (.L_HI(net493));
 sg13g2_tiehi _6577__494 (.L_HI(net494));
 sg13g2_tiehi _6576__495 (.L_HI(net495));
 sg13g2_tiehi _6575__496 (.L_HI(net496));
 sg13g2_tiehi _7090__497 (.L_HI(net497));
 sg13g2_tiehi _6574__498 (.L_HI(net498));
 sg13g2_tiehi _7089__499 (.L_HI(net499));
 sg13g2_tiehi _6573__500 (.L_HI(net500));
 sg13g2_tiehi _7088__501 (.L_HI(net501));
 sg13g2_tiehi _6572__502 (.L_HI(net502));
 sg13g2_tiehi _7087__503 (.L_HI(net503));
 sg13g2_tiehi _6571__504 (.L_HI(net504));
 sg13g2_tiehi _7086__505 (.L_HI(net505));
 sg13g2_tiehi _6570__506 (.L_HI(net506));
 sg13g2_tiehi _7085__507 (.L_HI(net507));
 sg13g2_tiehi _6569__508 (.L_HI(net508));
 sg13g2_tiehi _7084__509 (.L_HI(net509));
 sg13g2_tiehi _6568__510 (.L_HI(net510));
 sg13g2_tiehi _7083__511 (.L_HI(net511));
 sg13g2_tiehi _6567__512 (.L_HI(net512));
 sg13g2_tiehi _7082__513 (.L_HI(net513));
 sg13g2_tiehi _6566__514 (.L_HI(net514));
 sg13g2_tiehi _7081__515 (.L_HI(net515));
 sg13g2_tiehi _6565__516 (.L_HI(net516));
 sg13g2_tiehi _7080__517 (.L_HI(net517));
 sg13g2_tiehi _6564__518 (.L_HI(net518));
 sg13g2_tiehi _7079__519 (.L_HI(net519));
 sg13g2_tiehi _6563__520 (.L_HI(net520));
 sg13g2_tiehi _6562__521 (.L_HI(net521));
 sg13g2_tiehi _6561__522 (.L_HI(net522));
 sg13g2_tiehi _6560__523 (.L_HI(net523));
 sg13g2_tiehi _6559__524 (.L_HI(net524));
 sg13g2_tiehi _6558__525 (.L_HI(net525));
 sg13g2_tiehi _6557__526 (.L_HI(net526));
 sg13g2_tiehi _6556__527 (.L_HI(net527));
 sg13g2_tiehi _6555__528 (.L_HI(net528));
 sg13g2_tiehi _6554__529 (.L_HI(net529));
 sg13g2_tiehi _6553__530 (.L_HI(net530));
 sg13g2_tiehi _6552__531 (.L_HI(net531));
 sg13g2_tiehi _6551__532 (.L_HI(net532));
 sg13g2_tiehi _6550__533 (.L_HI(net533));
 sg13g2_tiehi _6549__534 (.L_HI(net534));
 sg13g2_tiehi _6548__535 (.L_HI(net535));
 sg13g2_tiehi _6547__536 (.L_HI(net536));
 sg13g2_tiehi _6546__537 (.L_HI(net537));
 sg13g2_tiehi _6545__538 (.L_HI(net538));
 sg13g2_tiehi _6544__539 (.L_HI(net539));
 sg13g2_tiehi _6543__540 (.L_HI(net540));
 sg13g2_tiehi _6542__541 (.L_HI(net541));
 sg13g2_tiehi _6541__542 (.L_HI(net542));
 sg13g2_tiehi _6540__543 (.L_HI(net543));
 sg13g2_tiehi _6539__544 (.L_HI(net544));
 sg13g2_tiehi _6538__545 (.L_HI(net545));
 sg13g2_tiehi _6537__546 (.L_HI(net546));
 sg13g2_tiehi _6536__547 (.L_HI(net547));
 sg13g2_tiehi _7078__548 (.L_HI(net548));
 sg13g2_tiehi _6535__549 (.L_HI(net549));
 sg13g2_tiehi _7077__550 (.L_HI(net550));
 sg13g2_tiehi _6534__551 (.L_HI(net551));
 sg13g2_tiehi _7076__552 (.L_HI(net552));
 sg13g2_tiehi _7075__553 (.L_HI(net553));
 sg13g2_tiehi _7074__554 (.L_HI(net554));
 sg13g2_tiehi _7073__555 (.L_HI(net555));
 sg13g2_tiehi _7072__556 (.L_HI(net556));
 sg13g2_tiehi _7071__557 (.L_HI(net557));
 sg13g2_tiehi _7070__558 (.L_HI(net558));
 sg13g2_tiehi _7069__559 (.L_HI(net559));
 sg13g2_tiehi _7068__560 (.L_HI(net560));
 sg13g2_tiehi _7067__561 (.L_HI(net561));
 sg13g2_tiehi _7066__562 (.L_HI(net562));
 sg13g2_tiehi _7065__563 (.L_HI(net563));
 sg13g2_tiehi _7064__564 (.L_HI(net564));
 sg13g2_tiehi _7063__565 (.L_HI(net565));
 sg13g2_tiehi _7062__566 (.L_HI(net566));
 sg13g2_tiehi _7061__567 (.L_HI(net567));
 sg13g2_tiehi _7060__568 (.L_HI(net568));
 sg13g2_tiehi _7059__569 (.L_HI(net569));
 sg13g2_tiehi _7058__570 (.L_HI(net570));
 sg13g2_tiehi _7057__571 (.L_HI(net571));
 sg13g2_tiehi _7056__572 (.L_HI(net572));
 sg13g2_tiehi _7055__573 (.L_HI(net573));
 sg13g2_tiehi _7054__574 (.L_HI(net574));
 sg13g2_tiehi _7053__575 (.L_HI(net575));
 sg13g2_tiehi _7052__576 (.L_HI(net576));
 sg13g2_tiehi _7051__577 (.L_HI(net577));
 sg13g2_tiehi _7050__578 (.L_HI(net578));
 sg13g2_tiehi _7049__579 (.L_HI(net579));
 sg13g2_tiehi _7048__580 (.L_HI(net580));
 sg13g2_tiehi _7047__581 (.L_HI(net581));
 sg13g2_tiehi _7046__582 (.L_HI(net582));
 sg13g2_tiehi _7045__583 (.L_HI(net583));
 sg13g2_tiehi _7044__584 (.L_HI(net584));
 sg13g2_tiehi _7043__585 (.L_HI(net585));
 sg13g2_tiehi _7042__586 (.L_HI(net586));
 sg13g2_tiehi _7041__587 (.L_HI(net587));
 sg13g2_tiehi _7040__588 (.L_HI(net588));
 sg13g2_tiehi _7039__589 (.L_HI(net589));
 sg13g2_tiehi _7038__590 (.L_HI(net590));
 sg13g2_tiehi _7037__591 (.L_HI(net591));
 sg13g2_tiehi _7036__592 (.L_HI(net592));
 sg13g2_tiehi _7035__593 (.L_HI(net593));
 sg13g2_tiehi _7034__594 (.L_HI(net594));
 sg13g2_tiehi _7033__595 (.L_HI(net595));
 sg13g2_tiehi _7032__596 (.L_HI(net596));
 sg13g2_tiehi _7031__597 (.L_HI(net597));
 sg13g2_tiehi _7030__598 (.L_HI(net598));
 sg13g2_tiehi _7029__599 (.L_HI(net599));
 sg13g2_tiehi _7028__600 (.L_HI(net600));
 sg13g2_tiehi _7027__601 (.L_HI(net601));
 sg13g2_tiehi _7026__602 (.L_HI(net602));
 sg13g2_tiehi _7025__603 (.L_HI(net603));
 sg13g2_tiehi _7024__604 (.L_HI(net604));
 sg13g2_tiehi _7023__605 (.L_HI(net605));
 sg13g2_tiehi _7022__606 (.L_HI(net606));
 sg13g2_tiehi _7021__607 (.L_HI(net607));
 sg13g2_tiehi _7020__608 (.L_HI(net608));
 sg13g2_tiehi _7019__609 (.L_HI(net609));
 sg13g2_tiehi _7018__610 (.L_HI(net610));
 sg13g2_tiehi _7017__611 (.L_HI(net611));
 sg13g2_tiehi _7016__612 (.L_HI(net612));
 sg13g2_tiehi _7015__613 (.L_HI(net613));
 sg13g2_tiehi _7014__614 (.L_HI(net614));
 sg13g2_tiehi _7013__615 (.L_HI(net615));
 sg13g2_tiehi _7012__616 (.L_HI(net616));
 sg13g2_tiehi _7011__617 (.L_HI(net617));
 sg13g2_tiehi _7010__618 (.L_HI(net618));
 sg13g2_tiehi _7009__619 (.L_HI(net619));
 sg13g2_tiehi _7008__620 (.L_HI(net620));
 sg13g2_tiehi _7007__621 (.L_HI(net621));
 sg13g2_tiehi _7006__622 (.L_HI(net622));
 sg13g2_tiehi _7005__623 (.L_HI(net623));
 sg13g2_tiehi _7004__624 (.L_HI(net624));
 sg13g2_tiehi _7003__625 (.L_HI(net625));
 sg13g2_tiehi _7002__626 (.L_HI(net626));
 sg13g2_tiehi _7001__627 (.L_HI(net627));
 sg13g2_tiehi _7000__628 (.L_HI(net628));
 sg13g2_tiehi _6999__629 (.L_HI(net629));
 sg13g2_tiehi _6998__630 (.L_HI(net630));
 sg13g2_tiehi _6997__631 (.L_HI(net631));
 sg13g2_tiehi _6996__632 (.L_HI(net632));
 sg13g2_tiehi _6995__633 (.L_HI(net633));
 sg13g2_tiehi _6994__634 (.L_HI(net634));
 sg13g2_tiehi _6993__635 (.L_HI(net635));
 sg13g2_tiehi _6992__636 (.L_HI(net636));
 sg13g2_tiehi _6991__637 (.L_HI(net637));
 sg13g2_tiehi _6990__638 (.L_HI(net638));
 sg13g2_tiehi _6989__639 (.L_HI(net639));
 sg13g2_tiehi _6988__640 (.L_HI(net640));
 sg13g2_tiehi _6987__641 (.L_HI(net641));
 sg13g2_tiehi _6986__642 (.L_HI(net642));
 sg13g2_tiehi _6985__643 (.L_HI(net643));
 sg13g2_tiehi _6984__644 (.L_HI(net644));
 sg13g2_tiehi _6983__645 (.L_HI(net645));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_vga_tetris_6 (.L_LO(net6));
 sg13g2_tielo tt_um_vga_tetris_7 (.L_LO(net7));
 sg13g2_tielo tt_um_vga_tetris_8 (.L_LO(net8));
 sg13g2_tielo tt_um_vga_tetris_9 (.L_LO(net9));
 sg13g2_tielo tt_um_vga_tetris_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_tetris_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_tetris_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_tetris_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_tetris_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_tetris_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_tetris_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_tetris_17 (.L_LO(net17));
 sg13g2_tielo tt_um_vga_tetris_18 (.L_LO(net18));
 sg13g2_tielo tt_um_vga_tetris_19 (.L_LO(net19));
 sg13g2_tielo tt_um_vga_tetris_20 (.L_LO(net20));
 sg13g2_tiehi _6982__21 (.L_HI(net21));
 sg13g2_buf_1 _7799_ (.A(\vga_tetris._vgaController_io_vSync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7800_ (.A(vga_hs),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout842 (.A(_2144_),
    .X(net842));
 sg13g2_buf_8 fanout843 (.A(net847),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net847),
    .X(net844));
 sg13g2_buf_8 fanout845 (.A(net847),
    .X(net845));
 sg13g2_buf_8 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_8 fanout847 (.A(_0875_),
    .X(net847));
 sg13g2_buf_8 fanout848 (.A(net850),
    .X(net848));
 sg13g2_buf_1 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_8 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_8 fanout851 (.A(net855),
    .X(net851));
 sg13g2_buf_8 fanout852 (.A(net855),
    .X(net852));
 sg13g2_buf_1 fanout853 (.A(net855),
    .X(net853));
 sg13g2_buf_8 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_8 fanout855 (.A(_2851_),
    .X(net855));
 sg13g2_buf_8 fanout856 (.A(net858),
    .X(net856));
 sg13g2_buf_1 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_8 fanout858 (.A(net859),
    .X(net858));
 sg13g2_buf_8 fanout859 (.A(_2830_),
    .X(net859));
 sg13g2_buf_8 fanout860 (.A(net862),
    .X(net860));
 sg13g2_buf_1 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_8 fanout862 (.A(_2830_),
    .X(net862));
 sg13g2_buf_8 fanout863 (.A(net865),
    .X(net863));
 sg13g2_buf_1 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_8 fanout865 (.A(net869),
    .X(net865));
 sg13g2_buf_8 fanout866 (.A(net869),
    .X(net866));
 sg13g2_buf_1 fanout867 (.A(net869),
    .X(net867));
 sg13g2_buf_8 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_8 fanout869 (.A(_2809_),
    .X(net869));
 sg13g2_buf_8 fanout870 (.A(net872),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_8 fanout872 (.A(_2788_),
    .X(net872));
 sg13g2_buf_8 fanout873 (.A(net876),
    .X(net873));
 sg13g2_buf_8 fanout874 (.A(net876),
    .X(net874));
 sg13g2_buf_1 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_8 fanout876 (.A(_2788_),
    .X(net876));
 sg13g2_buf_8 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_8 fanout878 (.A(net883),
    .X(net878));
 sg13g2_buf_8 fanout879 (.A(net882),
    .X(net879));
 sg13g2_buf_8 fanout880 (.A(net882),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_8 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_8 fanout883 (.A(_2767_),
    .X(net883));
 sg13g2_buf_8 fanout884 (.A(net885),
    .X(net884));
 sg13g2_buf_8 fanout885 (.A(net890),
    .X(net885));
 sg13g2_buf_8 fanout886 (.A(net889),
    .X(net886));
 sg13g2_buf_8 fanout887 (.A(net889),
    .X(net887));
 sg13g2_buf_1 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_8 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_8 fanout890 (.A(_2746_),
    .X(net890));
 sg13g2_buf_8 fanout891 (.A(net893),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_8 fanout893 (.A(net897),
    .X(net893));
 sg13g2_buf_8 fanout894 (.A(net897),
    .X(net894));
 sg13g2_buf_8 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_8 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_8 fanout897 (.A(_2725_),
    .X(net897));
 sg13g2_buf_8 fanout898 (.A(net900),
    .X(net898));
 sg13g2_buf_1 fanout899 (.A(net900),
    .X(net899));
 sg13g2_buf_8 fanout900 (.A(net904),
    .X(net900));
 sg13g2_buf_8 fanout901 (.A(net903),
    .X(net901));
 sg13g2_buf_8 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_8 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_8 fanout904 (.A(_2703_),
    .X(net904));
 sg13g2_buf_8 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_8 fanout906 (.A(_2682_),
    .X(net906));
 sg13g2_buf_8 fanout907 (.A(net910),
    .X(net907));
 sg13g2_buf_8 fanout908 (.A(net910),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_8 fanout910 (.A(_2682_),
    .X(net910));
 sg13g2_buf_8 fanout911 (.A(net913),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_8 fanout913 (.A(_2661_),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(net916),
    .X(net914));
 sg13g2_buf_8 fanout915 (.A(net916),
    .X(net915));
 sg13g2_buf_8 fanout916 (.A(_2661_),
    .X(net916));
 sg13g2_buf_8 fanout917 (.A(net919),
    .X(net917));
 sg13g2_buf_1 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_8 fanout919 (.A(_2640_),
    .X(net919));
 sg13g2_buf_8 fanout920 (.A(net923),
    .X(net920));
 sg13g2_buf_8 fanout921 (.A(net923),
    .X(net921));
 sg13g2_buf_1 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_8 fanout923 (.A(_2640_),
    .X(net923));
 sg13g2_buf_8 fanout924 (.A(net926),
    .X(net924));
 sg13g2_buf_1 fanout925 (.A(net926),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(_2618_),
    .X(net926));
 sg13g2_buf_8 fanout927 (.A(net929),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_8 fanout929 (.A(_2618_),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(net932),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_8 fanout932 (.A(net936),
    .X(net932));
 sg13g2_buf_8 fanout933 (.A(net936),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net936),
    .X(net934));
 sg13g2_buf_8 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_8 fanout936 (.A(_2597_),
    .X(net936));
 sg13g2_buf_8 fanout937 (.A(net939),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_8 fanout939 (.A(net943),
    .X(net939));
 sg13g2_buf_8 fanout940 (.A(net942),
    .X(net940));
 sg13g2_buf_8 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_8 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_8 fanout943 (.A(_2576_),
    .X(net943));
 sg13g2_buf_8 fanout944 (.A(net946),
    .X(net944));
 sg13g2_buf_1 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_8 fanout946 (.A(net950),
    .X(net946));
 sg13g2_buf_8 fanout947 (.A(net950),
    .X(net947));
 sg13g2_buf_1 fanout948 (.A(net950),
    .X(net948));
 sg13g2_buf_8 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_8 fanout950 (.A(_2555_),
    .X(net950));
 sg13g2_buf_8 fanout951 (.A(net956),
    .X(net951));
 sg13g2_buf_8 fanout952 (.A(net956),
    .X(net952));
 sg13g2_buf_8 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_8 fanout954 (.A(net956),
    .X(net954));
 sg13g2_buf_8 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_8 fanout956 (.A(_2533_),
    .X(net956));
 sg13g2_buf_8 fanout957 (.A(net959),
    .X(net957));
 sg13g2_buf_1 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_8 fanout959 (.A(net963),
    .X(net959));
 sg13g2_buf_8 fanout960 (.A(net963),
    .X(net960));
 sg13g2_buf_1 fanout961 (.A(net963),
    .X(net961));
 sg13g2_buf_8 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_8 fanout963 (.A(_2511_),
    .X(net963));
 sg13g2_buf_8 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_8 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_8 fanout966 (.A(net970),
    .X(net966));
 sg13g2_buf_8 fanout967 (.A(net970),
    .X(net967));
 sg13g2_buf_1 fanout968 (.A(net970),
    .X(net968));
 sg13g2_buf_8 fanout969 (.A(net970),
    .X(net969));
 sg13g2_buf_8 fanout970 (.A(_2488_),
    .X(net970));
 sg13g2_buf_8 fanout971 (.A(net973),
    .X(net971));
 sg13g2_buf_1 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_8 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_8 fanout974 (.A(_2465_),
    .X(net974));
 sg13g2_buf_8 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_8 fanout977 (.A(_2465_),
    .X(net977));
 sg13g2_buf_8 fanout978 (.A(net980),
    .X(net978));
 sg13g2_buf_1 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_8 fanout980 (.A(net984),
    .X(net980));
 sg13g2_buf_8 fanout981 (.A(net983),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_8 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_8 fanout984 (.A(_2268_),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(_0874_),
    .X(net985));
 sg13g2_buf_8 fanout986 (.A(_0871_),
    .X(net986));
 sg13g2_buf_8 fanout987 (.A(_0877_),
    .X(net987));
 sg13g2_buf_8 fanout988 (.A(_0877_),
    .X(net988));
 sg13g2_buf_8 fanout989 (.A(_0870_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_0870_),
    .X(net990));
 sg13g2_buf_8 fanout991 (.A(_0868_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_0868_),
    .X(net992));
 sg13g2_buf_8 fanout993 (.A(_0867_),
    .X(net993));
 sg13g2_buf_8 fanout994 (.A(_0867_),
    .X(net994));
 sg13g2_buf_8 fanout995 (.A(_0866_),
    .X(net995));
 sg13g2_buf_8 fanout996 (.A(_0866_),
    .X(net996));
 sg13g2_buf_8 fanout997 (.A(_0864_),
    .X(net997));
 sg13g2_buf_8 fanout998 (.A(_0864_),
    .X(net998));
 sg13g2_buf_8 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_buf_8 fanout1000 (.A(_0863_),
    .X(net1000));
 sg13g2_buf_8 fanout1001 (.A(_0862_),
    .X(net1001));
 sg13g2_buf_8 fanout1002 (.A(_0862_),
    .X(net1002));
 sg13g2_buf_8 fanout1003 (.A(_0861_),
    .X(net1003));
 sg13g2_buf_8 fanout1004 (.A(_0861_),
    .X(net1004));
 sg13g2_buf_8 fanout1005 (.A(_0859_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_0859_),
    .X(net1006));
 sg13g2_buf_8 fanout1007 (.A(_0858_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_0858_),
    .X(net1008));
 sg13g2_buf_8 fanout1009 (.A(_0856_),
    .X(net1009));
 sg13g2_buf_8 fanout1010 (.A(_0856_),
    .X(net1010));
 sg13g2_buf_8 fanout1011 (.A(_0855_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_0855_),
    .X(net1012));
 sg13g2_buf_8 fanout1013 (.A(_0852_),
    .X(net1013));
 sg13g2_buf_8 fanout1014 (.A(_0852_),
    .X(net1014));
 sg13g2_buf_8 fanout1015 (.A(_0851_),
    .X(net1015));
 sg13g2_buf_8 fanout1016 (.A(_0851_),
    .X(net1016));
 sg13g2_buf_8 fanout1017 (.A(_0847_),
    .X(net1017));
 sg13g2_buf_8 fanout1018 (.A(_0847_),
    .X(net1018));
 sg13g2_buf_8 fanout1019 (.A(_0845_),
    .X(net1019));
 sg13g2_buf_8 fanout1020 (.A(_0845_),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(_0842_),
    .X(net1021));
 sg13g2_buf_8 fanout1022 (.A(_0842_),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(_0838_),
    .X(net1023));
 sg13g2_buf_8 fanout1024 (.A(_0838_),
    .X(net1024));
 sg13g2_buf_8 fanout1025 (.A(net1029),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1029),
    .X(net1026));
 sg13g2_buf_8 fanout1027 (.A(net1029),
    .X(net1027));
 sg13g2_buf_1 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_8 fanout1029 (.A(_0857_),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(_0857_),
    .X(net1030));
 sg13g2_buf_1 fanout1031 (.A(_0857_),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_8 fanout1033 (.A(net1038),
    .X(net1033));
 sg13g2_buf_8 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_8 fanout1035 (.A(net1038),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(net1038),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(_0854_),
    .X(net1038));
 sg13g2_buf_8 fanout1039 (.A(net1042),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(net1042),
    .X(net1040));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_8 fanout1042 (.A(_0850_),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(_0848_),
    .X(net1043));
 sg13g2_buf_8 fanout1044 (.A(net1048),
    .X(net1044));
 sg13g2_buf_1 fanout1045 (.A(net1048),
    .X(net1045));
 sg13g2_buf_8 fanout1046 (.A(net1048),
    .X(net1046));
 sg13g2_buf_1 fanout1047 (.A(net1048),
    .X(net1047));
 sg13g2_buf_8 fanout1048 (.A(_0846_),
    .X(net1048));
 sg13g2_buf_8 fanout1049 (.A(_0846_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_0846_),
    .X(net1050));
 sg13g2_buf_8 fanout1051 (.A(net1053),
    .X(net1051));
 sg13g2_buf_8 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_8 fanout1053 (.A(_0844_),
    .X(net1053));
 sg13g2_buf_8 fanout1054 (.A(net1056),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(net1056),
    .X(net1055));
 sg13g2_buf_1 fanout1056 (.A(_0844_),
    .X(net1056));
 sg13g2_buf_8 fanout1057 (.A(net1059),
    .X(net1057));
 sg13g2_buf_8 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_8 fanout1059 (.A(_0841_),
    .X(net1059));
 sg13g2_buf_8 fanout1060 (.A(net1061),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(_0841_),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(_0840_),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(_0840_),
    .X(net1063));
 sg13g2_buf_8 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_8 fanout1065 (.A(_0840_),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(net1069),
    .X(net1066));
 sg13g2_buf_8 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_8 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(net1072),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(net1072),
    .X(net1070));
 sg13g2_buf_1 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(_0837_),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(net1076),
    .X(net1073));
 sg13g2_buf_1 fanout1074 (.A(net1076),
    .X(net1074));
 sg13g2_buf_8 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_8 fanout1076 (.A(_0798_),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(net1079),
    .X(net1077));
 sg13g2_buf_1 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(_0798_),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(_2928_),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(_1630_),
    .X(net1081));
 sg13g2_buf_1 fanout1082 (.A(_1630_),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_buf_8 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(_0914_),
    .X(net1085));
 sg13g2_buf_8 fanout1086 (.A(_1640_),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(_1601_),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(_1790_),
    .X(net1088));
 sg13g2_buf_8 fanout1089 (.A(_1787_),
    .X(net1089));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(_1551_),
    .X(net1091));
 sg13g2_buf_8 fanout1092 (.A(_2421_),
    .X(net1092));
 sg13g2_buf_8 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_8 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_8 fanout1095 (.A(_2348_),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(net1098),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(_2344_),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net1101),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_8 fanout1101 (.A(_2340_),
    .X(net1101));
 sg13g2_buf_8 fanout1102 (.A(net1104),
    .X(net1102));
 sg13g2_buf_8 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_8 fanout1104 (.A(_2336_),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_8 fanout1106 (.A(_2332_),
    .X(net1106));
 sg13g2_buf_1 fanout1107 (.A(_2332_),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_8 fanout1110 (.A(_2328_),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(net1113),
    .X(net1111));
 sg13g2_buf_8 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_8 fanout1113 (.A(_2324_),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1116),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_8 fanout1116 (.A(_2320_),
    .X(net1116));
 sg13g2_buf_8 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_8 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(_2316_),
    .X(net1119));
 sg13g2_buf_8 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_8 fanout1122 (.A(_2312_),
    .X(net1122));
 sg13g2_buf_8 fanout1123 (.A(net1125),
    .X(net1123));
 sg13g2_buf_1 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_8 fanout1125 (.A(_2308_),
    .X(net1125));
 sg13g2_buf_8 fanout1126 (.A(net1128),
    .X(net1126));
 sg13g2_buf_8 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(_2304_),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_8 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(_2300_),
    .X(net1131));
 sg13g2_buf_8 fanout1132 (.A(net1134),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sg13g2_buf_8 fanout1134 (.A(_2296_),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_2292_),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(net1140),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(_2288_),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_2284_),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(_2284_),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(net1146),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(net1146),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(_2280_),
    .X(net1146));
 sg13g2_buf_8 fanout1147 (.A(net1149),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_8 fanout1149 (.A(_2276_),
    .X(net1149));
 sg13g2_buf_8 fanout1150 (.A(net1152),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_8 fanout1152 (.A(_2272_),
    .X(net1152));
 sg13g2_buf_8 fanout1153 (.A(_2216_),
    .X(net1153));
 sg13g2_buf_8 fanout1154 (.A(_2216_),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(_2142_),
    .X(net1155));
 sg13g2_buf_8 fanout1156 (.A(_2068_),
    .X(net1156));
 sg13g2_buf_1 fanout1157 (.A(_2068_),
    .X(net1157));
 sg13g2_buf_8 fanout1158 (.A(_1810_),
    .X(net1158));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(_2183_),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(_2066_),
    .X(net1161));
 sg13g2_buf_8 fanout1162 (.A(_1733_),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_8 fanout1164 (.A(_2182_),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(_2182_),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(_1954_),
    .X(net1166));
 sg13g2_buf_8 fanout1167 (.A(_1949_),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(net1171),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(net1171),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_8 fanout1171 (.A(_1539_),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1179),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(net1179),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(net1177),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(net1178),
    .X(net1177));
 sg13g2_buf_8 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_8 fanout1179 (.A(_0756_),
    .X(net1179));
 sg13g2_buf_8 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_1 fanout1181 (.A(_0731_),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_1 fanout1183 (.A(net1187),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_8 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_8 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_8 fanout1187 (.A(_1698_),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(_0723_),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(net1192),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(_0720_),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(_0719_),
    .X(net1193));
 sg13g2_buf_8 fanout1194 (.A(_1147_),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(net1196),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_8 fanout1197 (.A(_0889_),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(net1200),
    .X(net1198));
 sg13g2_buf_2 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(_0889_),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(net1202),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(_0672_),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(_0669_),
    .X(net1204));
 sg13g2_buf_8 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(net1771),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(net1848),
    .X(net1207));
 sg13g2_buf_8 fanout1208 (.A(net1899),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1911),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(net1907),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(net1215),
    .X(net1213));
 sg13g2_buf_1 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(net1890),
    .X(net1215));
 sg13g2_buf_8 fanout1216 (.A(net1217),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1884),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(net1901),
    .X(net1219));
 sg13g2_buf_8 fanout1220 (.A(net1860),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_2 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(net1912),
    .X(net1223));
 sg13g2_buf_8 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(net1872),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1723),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(net1228),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net1869),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(net1900),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(net1811),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .X(net1232));
 sg13g2_buf_8 fanout1233 (.A(net1234),
    .X(net1233));
 sg13g2_buf_1 fanout1234 (.A(net1894),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net1885),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net1655),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .X(net1240));
 sg13g2_buf_8 fanout1241 (.A(\vga_tetris.tetrisLogic.stateQ[1] ),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(net1781),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(net1244),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(net1258),
    .X(net1245));
 sg13g2_buf_8 fanout1246 (.A(net1250),
    .X(net1246));
 sg13g2_buf_8 fanout1247 (.A(net1250),
    .X(net1247));
 sg13g2_buf_8 fanout1248 (.A(net1250),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(net1250),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(net1258),
    .X(net1250));
 sg13g2_buf_8 fanout1251 (.A(net1258),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(net1258),
    .X(net1252));
 sg13g2_buf_8 fanout1253 (.A(net1257),
    .X(net1253));
 sg13g2_buf_1 fanout1254 (.A(net1257),
    .X(net1254));
 sg13g2_buf_8 fanout1255 (.A(net1257),
    .X(net1255));
 sg13g2_buf_1 fanout1256 (.A(net1257),
    .X(net1256));
 sg13g2_buf_8 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_8 fanout1258 (.A(_0703_),
    .X(net1258));
 sg13g2_buf_8 fanout1259 (.A(net1260),
    .X(net1259));
 sg13g2_buf_8 fanout1260 (.A(net1264),
    .X(net1260));
 sg13g2_buf_8 fanout1261 (.A(net1264),
    .X(net1261));
 sg13g2_buf_8 fanout1262 (.A(net1263),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(net1272),
    .X(net1264));
 sg13g2_buf_8 fanout1265 (.A(net1272),
    .X(net1265));
 sg13g2_buf_1 fanout1266 (.A(net1267),
    .X(net1266));
 sg13g2_buf_8 fanout1267 (.A(net1272),
    .X(net1267));
 sg13g2_buf_8 fanout1268 (.A(net1271),
    .X(net1268));
 sg13g2_buf_8 fanout1269 (.A(net1271),
    .X(net1269));
 sg13g2_buf_8 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_8 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(rst_n),
    .X(net1272));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_vga_tetris_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_2_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_90_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_84_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_85_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_89_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_11_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_82_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_83_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_14_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_18_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_23_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_25_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_32_clk));
 sg13g2_buf_1 clkload24 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_34_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_30_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_72_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_55_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_leaf_77_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_79_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_80_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_64_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_68_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_69_clk));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload38 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_39_clk));
 sg13g2_inv_8 clkload42 (.A(clknet_leaf_46_clk));
 sg13g2_buf_8 clkload43 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload44 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload46 (.A(clknet_leaf_41_clk));
 sg13g2_buf_8 clkload47 (.A(clknet_leaf_43_clk));
 sg13g2_buf_8 clkload48 (.A(clknet_leaf_45_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vga_tetris.vgaController.horizontalCounterQ[0] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vga_tetris.msTimer.msTimerQ[0] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0015_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold4 (.A(\vga_tetris.boardMem.board_8[7] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold5 (.A(\vga_tetris.boardMem.board_7[5] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vga_tetris.boardMem.board_10[3] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold7 (.A(\vga_tetris.boardMem.board_9[13] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold8 (.A(\vga_tetris.boardMem.board_13[4] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0477_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vga_tetris.boardMem.board_9[9] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold11 (.A(\vga_tetris.boardMem.board_5[5] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold12 (.A(\vga_tetris.boardMem.board_12[4] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold13 (.A(\vga_tetris.boardMem.board_15[11] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold14 (.A(\vga_tetris.boardMem.board_9[17] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold15 (.A(\vga_tetris.boardMem.board_10[2] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vga_tetris.boardMem.board_9[12] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold17 (.A(\vga_tetris.boardMem.board_13[1] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold18 (.A(\vga_tetris.boardMem.board_4[12] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold19 (.A(\vga_tetris.boardMem.board_12[0] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0453_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold21 (.A(\vga_tetris.boardMem.board_9[1] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold22 (.A(\vga_tetris.boardMem.board_4[14] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold23 (.A(\vga_tetris.boardMem.board_4[4] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold24 (.A(\vga_tetris.boardMem.board_13[16] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold25 (.A(\vga_tetris.boardMem.board_7[8] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold26 (.A(\vga_tetris.boardMem.board_7[3] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold27 (.A(\vga_tetris.boardMem.board_8[2] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0375_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold29 (.A(\vga_tetris.boardMem.board_15[10] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold30 (.A(\vga_tetris.boardMem.board_5[8] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold31 (.A(\vga_tetris.boardMem.board_11[6] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vga_tetris.boardMem.board_9[10] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0403_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold34 (.A(\vga_tetris.boardMem.board_12[11] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0464_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold36 (.A(\vga_tetris.boardMem.board_11[11] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vga_tetris.boardMem.board_11[18] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold38 (.A(\vga_tetris.boardMem.board_6[17] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vga_tetris.boardMem.board_9[8] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold40 (.A(\vga_tetris.boardMem.board_6[18] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold41 (.A(\vga_tetris.boardMem.board_4[11] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0304_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold43 (.A(\vga_tetris.boardMem.board_8[1] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold44 (.A(\vga_tetris.boardMem.board_13[15] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vga_tetris.boardMem.board_8[13] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold46 (.A(\vga_tetris.boardMem.board_11[13] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vga_tetris.boardMem.board_7[4] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold48 (.A(\vga_tetris.boardMem.board_12[3] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vga_tetris.boardMem.board_5[18] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vga_tetris.boardMem.board_11[12] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vga_tetris.boardMem.board_4[10] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0303_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold53 (.A(\vga_tetris.boardMem.board_7[13] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vga_tetris.boardMem.board_4[16] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold55 (.A(\vga_tetris.boardMem.board_7[18] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vga_tetris.boardMem.board_11[19] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0452_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold58 (.A(\vga_tetris.boardMem.board_5[17] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold59 (.A(\vga_tetris.boardMem.board_13[12] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vga_tetris.boardMem.board_12[13] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold61 (.A(\vga_tetris.boardMem.board_10[5] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold62 (.A(\vga_tetris.boardMem.board_6[15] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold63 (.A(\vga_tetris.boardMem.board_10[4] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold64 (.A(\vga_tetris.boardMem.board_9[15] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vga_tetris.boardMem.board_6[10] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0343_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold67 (.A(\vga_tetris.boardMem.board_12[1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold68 (.A(\vga_tetris.boardMem.board_9[18] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold69 (.A(\vga_tetris.boardMem.board_7[19] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold70 (.A(\vga_tetris.boardMem.board_15[8] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold71 (.A(\vga_tetris.boardMem.board_5[2] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold72 (.A(\vga_tetris.boardMem.board_8[11] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vga_tetris.boardMem.board_8[16] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold74 (.A(\vga_tetris.boardMem.board_8[12] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0385_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vga_tetris.boardMem.board_6[8] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold77 (.A(\vga_tetris.boardMem.board_10[10] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold78 (.A(\vga_tetris.boardMem.board_8[10] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold79 (.A(\vga_tetris.boardMem.board_12[2] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vga_tetris.boardMem.board_9[16] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vga_tetris.boardMem.board_12[10] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vga_tetris.boardMem.board_4[17] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0310_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold84 (.A(\vga_tetris.boardMem.board_11[9] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold85 (.A(\vga_tetris.boardMem.board_15[14] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vga_tetris.boardMem.board_11[4] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold87 (.A(\vga_tetris.boardMem.board_12[6] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold88 (.A(\vga_tetris.boardMem.board_9[4] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold89 (.A(\vga_tetris.boardMem.board_6[4] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vga_tetris.boardMem.board_15[3] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vga_tetris.boardMem.board_4[9] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold92 (.A(\vga_tetris.boardMem.board_15[6] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold93 (.A(\vga_tetris.vgaController.horizontalCounterQ[2] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold94 (.A(_1792_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0007_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vga_tetris.boardMem.board_10[14] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold97 (.A(\vga_tetris.boardMem.board_7[9] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold98 (.A(\vga_tetris.boardMem.board_10[15] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold99 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0068_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold101 (.A(\vga_tetris.boardMem.board_10[17] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0430_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vga_tetris.boardMem.board_15[17] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold104 (.A(\vga_tetris.boardMem.board_14[4] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold105 (.A(\vga_tetris.boardMem.board_13[17] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vga_tetris.boardMem.board_10[16] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold107 (.A(\vga_tetris.boardMem.board_13[0] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0473_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold109 (.A(\vga_tetris.boardMem.board_13[5] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold110 (.A(\vga_tetris.boardMem.board_6[16] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold111 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0122_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold113 (.A(\vga_tetris.boardMem.board_15[0] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vga_tetris.boardMem.board_4[6] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold115 (.A(\vga_tetris.boardMem.board_7[0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold116 (.A(\vga_tetris.boardMem.board_6[1] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vga_tetris.boardMem.board_12[16] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold118 (.A(\vga_tetris.boardMem.board_11[5] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold119 (.A(\vga_tetris.boardMem.board_13[2] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold120 (.A(\vga_tetris.boardMem.board_5[1] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold121 (.A(\vga_tetris.boardMem.board_8[9] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vga_tetris.boardMem.board_6[0] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold123 (.A(\vga_tetris.boardMem.board_12[14] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold124 (.A(\vga_tetris.boardMem.board_15[16] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0529_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold126 (.A(\vga_tetris.boardMem.board_10[8] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold127 (.A(\vga_tetris.boardMem.board_11[15] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold128 (.A(\vga_tetris.boardMem.board_7[1] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold129 (.A(\vga_tetris.boardMem.board_10[6] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold130 (.A(\vga_tetris.boardMem.board_9[6] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold131 (.A(\vga_tetris.boardMem.board_9[7] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0400_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold133 (.A(\vga_tetris.boardMem.board_8[17] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold134 (.A(\vga_tetris.boardMem.board_6[14] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vga_tetris.boardMem.board_13[13] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold136 (.A(\vga_tetris.boardMem.board_14[8] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold137 (.A(\vga_tetris.boardMem.board_15[18] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vga_tetris.boardMem.board_11[0] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold139 (.A(\vga_tetris.boardMem.board_13[18] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold140 (.A(\vga_tetris.boardMem.board_6[3] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold141 (.A(\vga_tetris.boardMem.board_14[10] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold142 (.A(\vga_tetris.boardMem.board_8[6] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vga_tetris.boardMem.board_8[4] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0377_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold145 (.A(\vga_tetris.boardMem.board_15[19] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold146 (.A(\vga_tetris.boardMem.board_14[14] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold147 (.A(\vga_tetris.boardMem.board_8[5] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vga_tetris.boardMem.board_5[11] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0324_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold150 (.A(\vga_tetris.boardMem.board_4[0] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold151 (.A(\vga_tetris.boardMem.board_12[8] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold152 (.A(\vga_tetris.boardMem.board_14[5] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold153 (.A(\vga_tetris.boardMem.board_14[9] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vga_tetris.boardMem.board_9[14] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold155 (.A(\vga_tetris.boardMem.board_12[5] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vga_tetris.boardMem.board_5[6] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold157 (.A(\vga_tetris.boardMem.board_8[3] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold158 (.A(\vga_tetris.boardMem.board_15[13] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vga_tetris.boardMem.board_7[17] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold160 (.A(\vga_tetris.boardMem.board_12[18] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold161 (.A(\vga_tetris.boardMem.board_13[6] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0479_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold163 (.A(\vga_tetris.boardMem.board_8[15] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold164 (.A(\vga_tetris.boardMem.board_5[19] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold165 (.A(\vga_tetris.boardMem.board_15[9] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold166 (.A(\vga_tetris.boardMem.board_10[9] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold167 (.A(\vga_tetris.boardMem.board_5[13] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold168 (.A(\vga_tetris.boardMem.board_14[17] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold169 (.A(\vga_tetris.boardMem.board_13[8] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold170 (.A(\vga_tetris.boardMem.board_9[19] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold171 (.A(\vga_tetris.boardMem.board_9[3] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vga_tetris.boardMem.board_13[10] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold173 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0119_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vga_tetris.boardMem.board_12[12] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold176 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0120_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold178 (.A(\vga_tetris.boardMem.board_11[10] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold179 (.A(\vga_tetris.boardMem.board_7[11] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold180 (.A(\vga_tetris.boardMem.board_5[10] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold181 (.A(\vga_tetris.boardMem.board_10[18] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold182 (.A(\vga_tetris.boardMem.board_12[9] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold183 (.A(\vga_tetris.boardMem.board_10[13] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vga_tetris.boardMem.board_12[17] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold185 (.A(\vga_tetris.boardMem.board_7[16] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold186 (.A(\vga_tetris.boardMem.board_11[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold187 (.A(\vga_tetris.boardMem.board_11[8] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold188 (.A(\vga_tetris.boardMem.board_5[9] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vga_tetris.boardMem.board_4[1] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold190 (.A(\vga_tetris.boardMem.board_4[2] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold191 (.A(\vga_tetris.boardMem.board_11[7] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0440_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold193 (.A(\vga_tetris.boardMem.board_5[3] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold194 (.A(\vga_tetris.boardMem.board_4[18] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold195 (.A(\vga_tetris.boardMem.board_7[15] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vga_tetris.boardMem.board_9[11] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold197 (.A(\vga_tetris.boardMem.board_12[19] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0472_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold199 (.A(\vga_tetris.boardMem.board_10[0] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold200 (.A(\vga_tetris.boardMem.board_13[9] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold201 (.A(\vga_tetris.boardMem.board_13[14] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vga_tetris.boardMem.board_11[17] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold203 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0134_),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold205 (.A(\vga_tetris.boardMem.board_5[15] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold206 (.A(\vga_tetris.boardMem.board_7[6] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold207 (.A(\vga_tetris.boardMem.board_10[19] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold208 (.A(\vga_tetris.boardMem.board_6[2] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold209 (.A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0094_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold211 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0127_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold213 (.A(\vga_tetris.boardMem.board_8[18] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vga_tetris.boardMem.board_9[0] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold215 (.A(\vga_tetris.boardMem.board_5[7] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold216 (.A(\vga_tetris.boardMem.board_11[3] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold217 (.A(\vga_tetris.boardMem.board_4[3] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold218 (.A(\vga_tetris.boardMem.board_8[8] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold219 (.A(\vga_tetris.boardMem.board_14[13] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold220 (.A(\vga_tetris.boardMem.board_14[0] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold221 (.A(\vga_tetris.boardMem.board_14[19] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold222 (.A(\vga_tetris.boardMem.board_7[7] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold223 (.A(\vga_tetris.boardMem.board_14[1] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold224 (.A(\vga_tetris.boardMem.board_14[3] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold225 (.A(\vga_tetris.boardMem.board_12[15] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold226 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0121_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vga_tetris.boardMem.board_14[2] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold229 (.A(\vga_tetris.boardMem.board_9[5] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold230 (.A(\vga_tetris.boardMem.board_4[8] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold231 (.A(\vga_tetris.boardMem.board_14[15] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vga_tetris.boardMem.board_10[12] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold233 (.A(\vga_tetris.boardMem.board_12[7] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold234 (.A(\vga_tetris.boardMem.board_11[2] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vga_tetris.boardMem.board_15[15] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold236 (.A(\vga_tetris.boardMem.board_14[11] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold237 (.A(\vga_tetris.boardMem.board_10[11] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold238 (.A(\vga_tetris.boardMem.board_15[7] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold239 (.A(\vga_tetris.boardMem.board_6[6] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold240 (.A(\vga_tetris.boardMem.board_10[7] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vga_tetris.boardMem.board_8[0] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold242 (.A(\vga_tetris.boardMem.board_7[2] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vga_tetris.boardMem.board_6[11] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold244 (.A(\vga_tetris.boardMem.board_6[5] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vga_tetris.boardMem.board_11[14] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold246 (.A(\vga_tetris.boardMem.board_8[19] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold247 (.A(\vga_tetris.boardMem.board_6[12] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold248 (.A(\vga_tetris.boardMem.board_4[7] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0300_),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold250 (.A(\vga_tetris.boardMem.board_5[16] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold251 (.A(\vga_tetris.boardMem.board_5[4] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold252 (.A(\vga_tetris.boardMem.board_6[13] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vga_tetris.boardMem.board_13[7] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold254 (.A(\vga_tetris.boardMem.board_13[3] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold255 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0053_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold257 (.A(\vga_tetris.boardMem.board_7[12] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0365_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold259 (.A(\vga_tetris.boardMem.board_15[1] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0514_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold261 (.A(\vga_tetris.boardMem.board_5[12] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold262 (.A(\vga_tetris.boardMem.board_10[1] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold263 (.A(\vga_tetris.boardMem.board_14[16] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0509_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold265 (.A(\vga_tetris.boardMem.board_4[13] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold266 (.A(\vga_tetris.boardMem.board_6[9] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vga_tetris.boardMem.board_8[14] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold268 (.A(\vga_tetris.boardMem.board_7[10] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold269 (.A(\vga_tetris.boardMem.board_5[0] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold270 (.A(\vga_tetris.msTimer.msTimerQ[13] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0028_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold272 (.A(\vga_tetris.boardMem.board_4[5] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold273 (.A(\vga_tetris.boardMem.board_15[5] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold274 (.A(\vga_tetris.boardMem.board_14[18] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold275 (.A(\vga_tetris.vgaController.horizontalCounterQ[1] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold276 (.A(\vga_tetris.boardMem.board_14[7] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold277 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold278 (.A(\vga_tetris.boardMem.board_13[11] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold279 (.A(\vga_tetris.msTimer.msTimerQ[2] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold280 (.A(_1814_),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0017_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold282 (.A(\vga_tetris.boardMem.board_13[19] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold283 (.A(\vga_tetris.boardMem.board_14[6] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold284 (.A(\vga_tetris.boardMem.board_4[19] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold285 (.A(\vga_tetris.inputs.buttonTimerQ_0[1] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold286 (.A(_2360_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0177_),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold288 (.A(\vga_tetris.boardMem.board_15[4] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold289 (.A(\vga_tetris.boardMem.board_6[7] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold290 (.A(\vga_tetris.boardMem.board_7[14] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold291 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0058_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold293 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0126_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold295 (.A(\vga_tetris.boardMem.board_11[16] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold296 (.A(\vga_tetris.boardMem.board_14[12] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0505_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold298 (.A(\vga_tetris.boardMem.board_15[12] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold299 (.A(\vga_tetris.boardMem.board_15[2] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold300 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold301 (.A(\vga_tetris.boardMem.board_5[14] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold302 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold303 (.A(\vga_tetris.boardMem.board_4[15] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold304 (.A(\vga_tetris.boardMem.board_9[2] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold305 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0080_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold307 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold308 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold309 (.A(\vga_tetris.msTimer.msTimerQ[14] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold310 (.A(_1836_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold311 (.A(\vga_tetris.boardMem.board_6[19] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold312 (.A(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold313 (.A(_2231_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0139_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold315 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0075_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold317 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold318 (.A(\vga_tetris.boardMem.board_2[11] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold319 (.A(\vga_tetris.boardMem.board_0[5] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0218_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold321 (.A(\vga_tetris.boardMem.board_2[8] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold323 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold324 (.A(\vga_tetris.boardMem.board_17[4] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold325 (.A(\vga_tetris.boardMem.board_17[7] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold326 (.A(\vga_tetris.boardMem.board_1[18] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold327 (.A(\vga_tetris.boardMem.board_17[12] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold328 (.A(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold329 (.A(_2252_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0150_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold331 (.A(\vga_tetris.boardMem.board_0[3] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0216_),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold333 (.A(\vga_tetris.boardMem.board_17[5] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold334 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0057_),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold336 (.A(\vga_tetris.boardMem.board_16[4] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vga_tetris.boardMem.board_16[14] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold339 (.A(\vga_tetris.boardMem.board_17[2] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold340 (.A(\vga_tetris.boardMem.board_0[16] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold341 (.A(\vga_tetris.boardMem.board_0[17] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold342 (.A(\vga_tetris.boardMem.board_17[10] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0563_),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold344 (.A(\vga_tetris.boardMem.board_17[14] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold345 (.A(\vga_tetris.boardMem.board_0[15] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0228_),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold347 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vga_tetris.inputs.buttonTimerQ_2[6] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold349 (.A(_2417_),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0198_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold351 (.A(\vga_tetris.boardMem.board_16[7] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold352 (.A(\vga_tetris.boardMem.board_19[12] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold353 (.A(\vga_tetris.boardMem.board_16[6] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold354 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0083_),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold356 (.A(\vga_tetris.boardMem.board_18[11] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold357 (.A(\vga_tetris.boardMem.board_18[1] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0574_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold359 (.A(\vga_tetris.boardMem.board_16[11] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold360 (.A(\vga_tetris.boardMem.board_19[16] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold361 (.A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0095_),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vga_tetris.boardMem.board_0[12] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold364 (.A(\vga_tetris.boardMem.board_0[7] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vga_tetris.boardMem.board_16[15] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold366 (.A(\vga_tetris.boardMem.board_3[6] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold367 (.A(\vga_tetris.boardMem.board_17[18] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0571_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0064_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold371 (.A(\vga_tetris.boardMem.board_0[11] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold372 (.A(\vga_tetris.boardMem.board_1[1] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0234_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold374 (.A(\vga_tetris.boardMem.board_17[0] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold375 (.A(\vga_tetris.boardMem.board_18[5] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold376 (.A(\vga_tetris.boardMem.board_18[16] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold378 (.A(_2243_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0146_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold380 (.A(\vga_tetris.boardMem.board_1[13] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold381 (.A(\vga_tetris.boardMem.board_18[13] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold382 (.A(\vga_tetris.boardMem.board_19[11] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold383 (.A(\vga_tetris.boardMem.board_18[4] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold384 (.A(\vga_tetris.boardMem.board_3[17] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold385 (.A(\vga_tetris.boardMem.board_2[16] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vga_tetris.boardMem.board_1[4] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold387 (.A(\vga_tetris.boardMem.board_18[19] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold388 (.A(\vga_tetris.boardMem.board_18[10] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0583_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0076_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold392 (.A(\vga_tetris.boardMem.board_16[3] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold393 (.A(\vga_tetris.boardMem.board_0[18] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold394 (.A(\vga_tetris.boardMem.board_17[1] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold395 (.A(\vga_tetris.boardMem.board_1[3] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold396 (.A(\vga_tetris.boardMem.board_16[8] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold397 (.A(\vga_tetris.boardMem.board_2[4] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold398 (.A(\vga_tetris.boardMem.board_17[8] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold399 (.A(\vga_tetris.boardMem.board_18[6] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold400 (.A(\vga_tetris.boardMem.board_17[19] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold401 (.A(\vga_tetris.boardMem.board_3[12] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold402 (.A(\vga_tetris.boardMem.board_2[0] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold403 (.A(\vga_tetris.boardMem.board_17[15] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold404 (.A(\vga_tetris.boardMem.board_16[2] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold405 (.A(\vga_tetris.boardMem.board_16[16] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0549_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold407 (.A(\vga_tetris.boardMem.board_16[5] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold408 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold409 (.A(\vga_tetris.boardMem.board_0[6] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vga_tetris.boardMem.board_19[10] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold411 (.A(\vga_tetris.boardMem.board_1[10] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold412 (.A(\vga_tetris.boardMem.board_17[16] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold413 (.A(\vga_tetris.boardMem.board_0[9] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0222_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vga_tetris.boardMem.board_18[9] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold416 (.A(\vga_tetris.boardMem.board_3[19] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold417 (.A(\vga_tetris.boardMem.board_2[6] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold418 (.A(\vga_tetris.boardMem.board_17[11] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vga_tetris.boardMem.board_16[19] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold420 (.A(\vga_tetris.boardMem.board_18[7] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold421 (.A(\vga_tetris.boardMem.board_1[11] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold422 (.A(\vga_tetris.boardMem.board_3[13] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold423 (.A(\vga_tetris.boardMem.board_18[12] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold424 (.A(\vga_tetris.boardMem.board_1[2] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold425 (.A(\vga_tetris.boardMem.board_0[0] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold426 (.A(\vga_tetris.boardMem.board_3[4] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold427 (.A(\vga_tetris.boardMem.board_19[14] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold428 (.A(\vga_tetris.boardMem.board_1[5] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold429 (.A(\vga_tetris.boardMem.board_2[1] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold430 (.A(\vga_tetris.boardMem.board_2[9] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold431 (.A(\vga_tetris.boardMem.board_3[14] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold432 (.A(\vga_tetris.boardMem.board_18[3] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold433 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold434 (.A(\vga_tetris.boardMem.board_2[2] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold435 (.A(\vga_tetris.boardMem.board_0[10] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0223_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold437 (.A(\vga_tetris.boardMem.board_16[18] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold438 (.A(\vga_tetris.boardMem.board_16[10] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold439 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold440 (.A(\vga_tetris.boardMem.board_16[12] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold441 (.A(\vga_tetris.boardMem.board_0[4] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold442 (.A(\vga_tetris.boardMem.board_19[5] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold443 (.A(\vga_tetris.boardMem.board_18[15] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold444 (.A(\vga_tetris.boardMem.board_3[5] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold445 (.A(\vga_tetris.boardMem.board_3[18] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold446 (.A(\vga_tetris.vgaController.horizontalCounterQ[3] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold447 (.A(\vga_tetris.boardMem.board_19[0] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold448 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold449 (.A(\vga_tetris.boardMem.board_1[12] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold450 (.A(\vga_tetris.boardMem.board_0[19] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold451 (.A(\vga_tetris.boardMem.board_0[8] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0221_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold453 (.A(\vga_tetris.boardMem.board_2[13] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold454 (.A(\vga_tetris.boardMem.board_18[17] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0590_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold456 (.A(\vga_tetris.boardMem.board_3[15] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold457 (.A(\vga_tetris.boardMem.board_2[10] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold458 (.A(\vga_tetris.boardMem.board_3[2] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold459 (.A(\vga_tetris.boardMem.board_3[3] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold460 (.A(\vga_tetris.boardMem.board_19[9] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold461 (.A(\vga_tetris.boardMem.board_0[1] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold462 (.A(\vga_tetris.boardMem.board_16[1] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold463 (.A(\vga_tetris.boardMem.board_0[14] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0227_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold465 (.A(\vga_tetris.boardMem.board_2[18] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold466 (.A(\vga_tetris.boardMem.board_1[17] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold467 (.A(\vga_tetris.boardMem.board_19[7] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold468 (.A(\vga_tetris.boardMem.board_18[0] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0573_),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold470 (.A(\vga_tetris.boardMem.board_0[13] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0226_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold472 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold473 (.A(_1908_),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0045_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold475 (.A(\vga_tetris.boardMem.board_16[9] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold476 (.A(\vga_tetris.boardMem.board_18[14] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold477 (.A(\vga_tetris.boardMem.board_1[19] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold478 (.A(\vga_tetris.boardMem.board_3[9] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold479 (.A(\vga_tetris.boardMem.board_2[7] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold480 (.A(\vga_tetris.boardMem.board_1[14] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold481 (.A(\vga_tetris.boardMem.board_17[9] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0562_),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold483 (.A(\vga_tetris.boardMem.board_1[9] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold484 (.A(\vga_tetris.boardMem.board_2[19] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold485 (.A(\vga_tetris.boardMem.board_2[15] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold486 (.A(\vga_tetris.boardMem.board_19[3] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold487 (.A(\vga_tetris.boardMem.board_3[7] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold488 (.A(\vga_tetris.boardMem.board_3[8] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0281_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold490 (.A(\vga_tetris.boardMem.board_18[8] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0581_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold492 (.A(\vga_tetris.boardMem.board_19[2] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold493 (.A(\vga_tetris.boardMem.board_1[7] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold494 (.A(\vga_tetris.boardMem.board_18[2] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold495 (.A(\vga_tetris.boardMem.board_18[18] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold496 (.A(\vga_tetris.boardMem.board_3[10] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold497 (.A(\vga_tetris.boardMem.board_3[16] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold498 (.A(\vga_tetris.boardMem.board_17[3] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold499 (.A(\vga_tetris.boardMem.board_3[1] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold500 (.A(\vga_tetris.boardMem.board_19[1] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold501 (.A(\vga_tetris.boardMem.board_19[18] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold502 (.A(\vga_tetris.boardMem.board_19[6] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold503 (.A(\vga_tetris.boardMem.board_17[17] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0570_),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold505 (.A(\vga_tetris.boardMem.board_1[15] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold506 (.A(\vga_tetris.boardMem.board_17[13] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold507 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold508 (.A(\vga_tetris.boardMem.board_19[15] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold509 (.A(\vga_tetris.boardMem.board_1[8] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold510 (.A(\vga_tetris.boardMem.board_16[17] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold511 (.A(\vga_tetris.boardMem.board_2[17] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold512 (.A(\vga_tetris.boardMem.board_19[4] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold513 (.A(\vga_tetris.boardMem.board_19[19] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold514 (.A(\vga_tetris.boardMem.board_19[17] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold515 (.A(\vga_tetris.boardMem.board_16[0] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0533_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold517 (.A(\vga_tetris.boardMem.board_2[5] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold518 (.A(\vga_tetris.boardMem.board_0[2] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0215_),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold520 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold521 (.A(_1952_),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold522 (.A(\vga_tetris.boardMem.board_2[14] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold523 (.A(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0597_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold525 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold526 (.A(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold527 (.A(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0594_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold529 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold530 (.A(\vga_tetris.boardMem.board_1[16] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0249_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold532 (.A(\vga_tetris.boardMem.board_3[0] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold533 (.A(\vga_tetris.boardMem.board_1[6] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold534 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0051_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold536 (.A(\vga_tetris.boardMem.board_1[0] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold537 (.A(\vga_tetris.boardMem.board_2[3] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold538 (.A(\vga_tetris.boardMem.board_19[13] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold539 (.A(\vga_tetris.boardMem.board_19[8] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0164_),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold541 (.A(\vga_tetris.boardMem.board_17[6] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold542 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold543 (.A(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold544 (.A(\vga_tetris.boardMem.board_2[12] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold545 (.A(\vga_tetris.boardMem.board_16[13] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold546 (.A(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold547 (.A(_2880_),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold548 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold549 (.A(_1867_),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold550 (.A(\vga_tetris.inputs.buttonTimerQ_0[7] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold551 (.A(_2373_),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0183_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold553 (.A(\vga_tetris.boardMem.board_3[11] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold554 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold555 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0062_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold557 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold558 (.A(_1989_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold559 (.A(\vga_tetris.inputs.buttonTimerQ_0[6] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold560 (.A(_2371_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0182_),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold562 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold563 (.A(_2026_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold564 (.A(\vga_tetris.msTimer.msTimerQ[6] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold565 (.A(_1822_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0021_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold567 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold568 (.A(_2011_),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold569 (.A(\vga_tetris.inputs.buttonTimerQ_2[0] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold570 (.A(_2402_),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0192_),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold572 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold573 (.A(_2020_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold574 (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold575 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold576 (.A(_2017_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold577 (.A(\vga_tetris.msTimer.msTimerQ[7] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold578 (.A(_1823_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold579 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold580 (.A(_1869_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold581 (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold582 (.A(\vga_tetris.msTimer.msTimerQ[3] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold583 (.A(_1816_),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0018_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold585 (.A(\vga_tetris._tetrisLogic_io_score_0[0] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold586 (.A(_2253_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold587 (.A(\vga_tetris.inputs.buttonTimerQ_1[0] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold588 (.A(_2379_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0184_),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold590 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold591 (.A(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold592 (.A(_2890_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold593 (.A(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold594 (.A(_1797_),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0011_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold596 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold597 (.A(\vga_tetris.inputs.buttonTimerQ_1[7] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold598 (.A(_2395_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold599 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold600 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold601 (.A(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold602 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold603 (.A(_1910_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0046_),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold605 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold606 (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold607 (.A(_1796_),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0010_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold609 (.A(\vga_tetris.msTimer.msTimerQ[5] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold610 (.A(_1820_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0020_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold612 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold613 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold614 (.A(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0602_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold616 (.A(\vga_tetris._inputs_io_downButtonActive ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0211_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold618 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold619 (.A(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold620 (.A(_1800_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold621 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0132_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold623 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold624 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold625 (.A(_1937_),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold626 (.A(_0066_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold627 (.A(\vga_tetris.msTimer.msTimerQ[4] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold628 (.A(_1818_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold629 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold630 (.A(\vga_tetris.inputs.buttonTimerQ_2[7] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold631 (.A(_2420_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0199_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold633 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold634 (.A(_2101_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold635 (.A(_0593_),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold636 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold637 (.A(_1912_),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold638 (.A(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold639 (.A(_2233_),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold640 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold641 (.A(\vga_tetris.inputs.buttonTimerQ_2[1] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold642 (.A(_0193_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold643 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold644 (.A(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold645 (.A(_2215_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold646 (.A(_0135_),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold647 (.A(\vga_tetris.startTetrisLogicQ ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0067_),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold649 (.A(\vga_tetris.inputs.buttonTimerQ_0[0] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold650 (.A(\vga_tetris.inputs.buttonTimerQ_1[1] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold651 (.A(_2381_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold652 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold653 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold654 (.A(\vga_tetris.inputs.buttonTimerQ_1[6] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold655 (.A(_2394_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold656 (.A(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[2] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold657 (.A(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold658 (.A(_2244_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold659 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold660 (.A(_1916_),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold661 (.A(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold662 (.A(_2226_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0137_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold664 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold665 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold666 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold667 (.A(\vga_tetris.msTimer.msTimerQ[8] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold668 (.A(\vga_tetris.msTimer.msTimerQ[1] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold669 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold670 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold671 (.A(\vga_tetris.msTimer.msTimerQ[12] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold672 (.A(_1834_),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold673 (.A(_0027_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold674 (.A(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold675 (.A(_2042_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold676 (.A(_0091_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold677 (.A(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold678 (.A(_2235_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold679 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold680 (.A(_1860_),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold681 (.A(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0621_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold683 (.A(\vga_tetris.msTimer.msTimerQ[9] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold684 (.A(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold685 (.A(_1803_),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold686 (.A(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold687 (.A(_2219_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold688 (.A(_2222_),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0136_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold690 (.A(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold691 (.A(\vga_tetris.inputs.buttonTimerQ_1[5] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold692 (.A(_2391_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0189_),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold694 (.A(\vga_tetris.msTimer.msTimerQ[10] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold695 (.A(\vga_tetris.runningTetrisLogicQ ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold696 (.A(_0212_),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold697 (.A(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold698 (.A(_2249_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold699 (.A(_0149_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold700 (.A(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold701 (.A(_2921_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold702 (.A(_0612_),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold703 (.A(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold704 (.A(\vga_tetris.msTimer.msTimerQ[11] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold705 (.A(\vga_tetris.tetrisLogic.stateQ[1] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold706 (.A(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold707 (.A(_2902_),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold708 (.A(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold709 (.A(_2240_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0145_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold711 (.A(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold712 (.A(\vga_tetris._vgaController_io_pixelPosX[1] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold713 (.A(\vga_tetris.tetrisLogic.stateQ[3] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold714 (.A(_1750_),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold715 (.A(\vga_tetris._tetrisLogic_io_score_0[2] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold716 (.A(_2257_),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold717 (.A(_0153_),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold718 (.A(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold719 (.A(_1802_),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold720 (.A(\vga_tetris.tetrisLogic.stateQ[2] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold721 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold722 (.A(\vga_tetris.inputs.buttonTimerQ_3[0] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold723 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold724 (.A(_2048_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold725 (.A(\vga_tetris.inputs.buttonTimerQ_3[3] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold726 (.A(_2433_),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold727 (.A(\vga_tetris.inputs.buttonTimerQ_3[7] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold728 (.A(_2445_),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold729 (.A(_2446_),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold730 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold731 (.A(_1943_),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold732 (.A(_0069_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold733 (.A(\vga_tetris._vgaController_io_pixelPosX[9] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold734 (.A(_2919_),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold735 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold736 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold737 (.A(\vga_tetris.inputs.buttonTimerQ_0[4] ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold738 (.A(_2368_),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold739 (.A(_0180_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold740 (.A(\vga_tetris.inputs.buttonTimerQ_2[4] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold741 (.A(_2413_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold742 (.A(_0196_),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold743 (.A(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold744 (.A(_0607_),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold745 (.A(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold746 (.A(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold747 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold748 (.A(\vga_tetris.inputs.buttonTimerQ_1[4] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold749 (.A(_2388_),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold750 (.A(_2390_),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold751 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold752 (.A(_2135_),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold753 (.A(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold754 (.A(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold755 (.A(_2211_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold756 (.A(_2247_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold757 (.A(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold758 (.A(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold759 (.A(_2435_),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold760 (.A(\vga_tetris.inputs.buttonTimerQ_2[2] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold761 (.A(_2408_),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold762 (.A(\vga_tetris.inputs.buttonTimerQ_1[2] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold763 (.A(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold764 (.A(_2238_),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold765 (.A(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold766 (.A(_2416_),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold767 (.A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold768 (.A(_0039_),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold769 (.A(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold770 (.A(_2366_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold771 (.A(\vga_tetris.inputs.buttonTimerQ_0[2] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold772 (.A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0622_),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold774 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold775 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold776 (.A(_0106_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold777 (.A(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold778 (.A(\vga_tetris._vgaController_io_vSync ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold779 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold780 (.A(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0187_),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold782 (.A(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold783 (.A(_2256_),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold784 (.A(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold785 (.A(_2914_),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold786 (.A(_0609_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold787 (.A(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold788 (.A(_1131_),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold789 (.A(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold790 (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold791 (.A(\vga_tetris.inputs.buttonTimerQ_3[6] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold792 (.A(_2442_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold793 (.A(\vga_tetris._tetrisLogic_io_gameOver ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold794 (.A(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold795 (.A(\vga_tetris._inputs_io_rightButtonActive ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold796 (.A(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold797 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold798 (.A(_2133_),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold799 (.A(_2134_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold800 (.A(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold801 (.A(_2411_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold802 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold803 (.A(_2052_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold804 (.A(\vga_tetris.tetrisLogic.stateQ[0] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold805 (.A(_0000_),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold806 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold807 (.A(_0098_),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold808 (.A(\vga_tetris._vgaController_io_pixelPosY[2] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold809 (.A(\vga_tetris.tetrisLogic.rotationQ[0] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold810 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold811 (.A(_0100_),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold812 (.A(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold813 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold814 (.A(\vga_tetris._vgaController_io_pixelPosY[3] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold815 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold816 (.A(_2128_),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold817 (.A(_0103_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold818 (.A(\vga_tetris.tetrisLogic.stateQ[4] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold819 (.A(_0041_),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold820 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold821 (.A(_0097_),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold822 (.A(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold823 (.A(\vga_tetris._vgaController_io_pixelPosY[6] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold824 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold825 (.A(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold826 (.A(_2915_),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold827 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold828 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold829 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold830 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold831 (.A(\vga_tetris._tetrisDisplay_io_boardYCoord[0] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold832 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold833 (.A(_0004_),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold834 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold835 (.A(\vga_tetris._tetrisDisplay_io_boardYCoord[1] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold836 (.A(\vga_tetris._vgaController_io_pixelPosX[4] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold837 (.A(\vga_tetris.msTimer.msTimerQ[12] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold838 (.A(_1804_),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold839 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold840 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold841 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold842 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold843 (.A(_2106_),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold844 (.A(\vga_tetris.boardMem.board_0[10] ),
    .X(net1920));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_4 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_512 ();
 sg13g2_decap_8 FILLER_4_519 ();
 sg13g2_decap_8 FILLER_4_526 ();
 sg13g2_decap_8 FILLER_4_533 ();
 sg13g2_decap_8 FILLER_4_540 ();
 sg13g2_decap_8 FILLER_4_547 ();
 sg13g2_fill_2 FILLER_4_554 ();
 sg13g2_fill_1 FILLER_4_556 ();
 sg13g2_decap_8 FILLER_4_561 ();
 sg13g2_decap_8 FILLER_4_568 ();
 sg13g2_decap_8 FILLER_4_575 ();
 sg13g2_decap_8 FILLER_4_582 ();
 sg13g2_decap_8 FILLER_4_589 ();
 sg13g2_decap_8 FILLER_4_596 ();
 sg13g2_decap_8 FILLER_4_603 ();
 sg13g2_decap_8 FILLER_4_610 ();
 sg13g2_decap_8 FILLER_4_617 ();
 sg13g2_decap_8 FILLER_4_624 ();
 sg13g2_decap_8 FILLER_4_631 ();
 sg13g2_decap_8 FILLER_4_638 ();
 sg13g2_decap_8 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_652 ();
 sg13g2_decap_8 FILLER_4_659 ();
 sg13g2_decap_8 FILLER_4_666 ();
 sg13g2_decap_8 FILLER_4_673 ();
 sg13g2_decap_8 FILLER_4_680 ();
 sg13g2_decap_8 FILLER_4_687 ();
 sg13g2_decap_8 FILLER_4_694 ();
 sg13g2_decap_8 FILLER_4_701 ();
 sg13g2_decap_8 FILLER_4_708 ();
 sg13g2_decap_8 FILLER_4_715 ();
 sg13g2_decap_8 FILLER_4_722 ();
 sg13g2_decap_8 FILLER_4_729 ();
 sg13g2_decap_8 FILLER_4_736 ();
 sg13g2_decap_8 FILLER_4_743 ();
 sg13g2_decap_8 FILLER_4_750 ();
 sg13g2_decap_8 FILLER_4_757 ();
 sg13g2_decap_8 FILLER_4_764 ();
 sg13g2_decap_8 FILLER_4_771 ();
 sg13g2_decap_8 FILLER_4_778 ();
 sg13g2_decap_8 FILLER_4_785 ();
 sg13g2_decap_8 FILLER_4_792 ();
 sg13g2_decap_8 FILLER_4_799 ();
 sg13g2_decap_8 FILLER_4_806 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_8 FILLER_4_834 ();
 sg13g2_decap_8 FILLER_4_841 ();
 sg13g2_decap_8 FILLER_4_848 ();
 sg13g2_decap_8 FILLER_4_855 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_4 FILLER_5_438 ();
 sg13g2_fill_1 FILLER_5_442 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_4 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_486 ();
 sg13g2_fill_1 FILLER_5_493 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_2 FILLER_5_612 ();
 sg13g2_fill_2 FILLER_5_628 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_635 ();
 sg13g2_decap_8 FILLER_5_642 ();
 sg13g2_decap_8 FILLER_5_649 ();
 sg13g2_decap_8 FILLER_5_656 ();
 sg13g2_decap_8 FILLER_5_663 ();
 sg13g2_decap_8 FILLER_5_670 ();
 sg13g2_decap_8 FILLER_5_677 ();
 sg13g2_decap_8 FILLER_5_684 ();
 sg13g2_decap_8 FILLER_5_691 ();
 sg13g2_decap_8 FILLER_5_698 ();
 sg13g2_decap_8 FILLER_5_705 ();
 sg13g2_decap_8 FILLER_5_712 ();
 sg13g2_decap_8 FILLER_5_719 ();
 sg13g2_decap_8 FILLER_5_726 ();
 sg13g2_decap_8 FILLER_5_733 ();
 sg13g2_decap_8 FILLER_5_740 ();
 sg13g2_decap_8 FILLER_5_747 ();
 sg13g2_decap_8 FILLER_5_754 ();
 sg13g2_decap_8 FILLER_5_761 ();
 sg13g2_decap_8 FILLER_5_768 ();
 sg13g2_decap_8 FILLER_5_775 ();
 sg13g2_decap_8 FILLER_5_782 ();
 sg13g2_decap_8 FILLER_5_789 ();
 sg13g2_decap_8 FILLER_5_796 ();
 sg13g2_decap_8 FILLER_5_803 ();
 sg13g2_decap_8 FILLER_5_810 ();
 sg13g2_decap_8 FILLER_5_817 ();
 sg13g2_decap_8 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_831 ();
 sg13g2_decap_8 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_845 ();
 sg13g2_decap_8 FILLER_5_852 ();
 sg13g2_fill_2 FILLER_5_859 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_fill_2 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_456 ();
 sg13g2_fill_1 FILLER_6_463 ();
 sg13g2_fill_1 FILLER_6_473 ();
 sg13g2_fill_2 FILLER_6_478 ();
 sg13g2_fill_1 FILLER_6_480 ();
 sg13g2_decap_4 FILLER_6_490 ();
 sg13g2_fill_2 FILLER_6_508 ();
 sg13g2_fill_1 FILLER_6_510 ();
 sg13g2_fill_2 FILLER_6_525 ();
 sg13g2_fill_1 FILLER_6_527 ();
 sg13g2_decap_4 FILLER_6_541 ();
 sg13g2_fill_2 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_587 ();
 sg13g2_fill_1 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_657 ();
 sg13g2_decap_8 FILLER_6_664 ();
 sg13g2_decap_8 FILLER_6_671 ();
 sg13g2_decap_8 FILLER_6_678 ();
 sg13g2_decap_4 FILLER_6_685 ();
 sg13g2_decap_8 FILLER_6_692 ();
 sg13g2_decap_8 FILLER_6_699 ();
 sg13g2_decap_8 FILLER_6_710 ();
 sg13g2_decap_8 FILLER_6_717 ();
 sg13g2_decap_4 FILLER_6_724 ();
 sg13g2_fill_2 FILLER_6_728 ();
 sg13g2_decap_4 FILLER_6_761 ();
 sg13g2_fill_2 FILLER_6_769 ();
 sg13g2_decap_8 FILLER_6_780 ();
 sg13g2_decap_8 FILLER_6_787 ();
 sg13g2_decap_8 FILLER_6_794 ();
 sg13g2_decap_8 FILLER_6_801 ();
 sg13g2_decap_8 FILLER_6_808 ();
 sg13g2_decap_8 FILLER_6_815 ();
 sg13g2_decap_8 FILLER_6_822 ();
 sg13g2_decap_8 FILLER_6_829 ();
 sg13g2_decap_8 FILLER_6_836 ();
 sg13g2_decap_8 FILLER_6_843 ();
 sg13g2_decap_8 FILLER_6_850 ();
 sg13g2_decap_4 FILLER_6_857 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_4 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_7_435 ();
 sg13g2_fill_1 FILLER_7_461 ();
 sg13g2_fill_1 FILLER_7_466 ();
 sg13g2_fill_1 FILLER_7_472 ();
 sg13g2_decap_8 FILLER_7_477 ();
 sg13g2_fill_1 FILLER_7_484 ();
 sg13g2_fill_2 FILLER_7_512 ();
 sg13g2_fill_2 FILLER_7_566 ();
 sg13g2_fill_2 FILLER_7_608 ();
 sg13g2_fill_1 FILLER_7_610 ();
 sg13g2_fill_2 FILLER_7_616 ();
 sg13g2_fill_2 FILLER_7_636 ();
 sg13g2_fill_1 FILLER_7_638 ();
 sg13g2_decap_8 FILLER_7_666 ();
 sg13g2_fill_1 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_732 ();
 sg13g2_fill_1 FILLER_7_734 ();
 sg13g2_fill_2 FILLER_7_748 ();
 sg13g2_fill_1 FILLER_7_759 ();
 sg13g2_decap_8 FILLER_7_787 ();
 sg13g2_decap_8 FILLER_7_794 ();
 sg13g2_decap_8 FILLER_7_801 ();
 sg13g2_decap_8 FILLER_7_808 ();
 sg13g2_decap_8 FILLER_7_815 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_decap_8 FILLER_7_829 ();
 sg13g2_decap_8 FILLER_7_836 ();
 sg13g2_decap_8 FILLER_7_843 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_decap_4 FILLER_7_857 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_fill_2 FILLER_8_392 ();
 sg13g2_fill_1 FILLER_8_394 ();
 sg13g2_fill_2 FILLER_8_400 ();
 sg13g2_fill_1 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_407 ();
 sg13g2_decap_4 FILLER_8_414 ();
 sg13g2_fill_2 FILLER_8_418 ();
 sg13g2_decap_4 FILLER_8_544 ();
 sg13g2_fill_1 FILLER_8_548 ();
 sg13g2_decap_4 FILLER_8_576 ();
 sg13g2_decap_4 FILLER_8_593 ();
 sg13g2_fill_1 FILLER_8_597 ();
 sg13g2_fill_2 FILLER_8_613 ();
 sg13g2_fill_1 FILLER_8_615 ();
 sg13g2_fill_2 FILLER_8_622 ();
 sg13g2_fill_1 FILLER_8_687 ();
 sg13g2_decap_8 FILLER_8_705 ();
 sg13g2_fill_1 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_8_727 ();
 sg13g2_fill_2 FILLER_8_743 ();
 sg13g2_fill_1 FILLER_8_755 ();
 sg13g2_decap_8 FILLER_8_789 ();
 sg13g2_fill_2 FILLER_8_796 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_4 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_4 FILLER_9_112 ();
 sg13g2_fill_2 FILLER_9_116 ();
 sg13g2_decap_4 FILLER_9_131 ();
 sg13g2_decap_4 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_decap_4 FILLER_9_184 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_4 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_fill_1 FILLER_9_384 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_433 ();
 sg13g2_decap_4 FILLER_9_438 ();
 sg13g2_fill_2 FILLER_9_442 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_4 FILLER_9_466 ();
 sg13g2_fill_1 FILLER_9_492 ();
 sg13g2_fill_2 FILLER_9_502 ();
 sg13g2_fill_1 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_fill_2 FILLER_9_532 ();
 sg13g2_fill_2 FILLER_9_540 ();
 sg13g2_fill_1 FILLER_9_542 ();
 sg13g2_decap_4 FILLER_9_574 ();
 sg13g2_decap_4 FILLER_9_586 ();
 sg13g2_decap_8 FILLER_9_632 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_decap_8 FILLER_9_646 ();
 sg13g2_fill_2 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_659 ();
 sg13g2_fill_2 FILLER_9_666 ();
 sg13g2_fill_1 FILLER_9_668 ();
 sg13g2_fill_2 FILLER_9_682 ();
 sg13g2_decap_8 FILLER_9_702 ();
 sg13g2_decap_4 FILLER_9_745 ();
 sg13g2_fill_2 FILLER_9_749 ();
 sg13g2_fill_2 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_832 ();
 sg13g2_decap_8 FILLER_9_839 ();
 sg13g2_decap_8 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_853 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_89 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_decap_4 FILLER_10_407 ();
 sg13g2_fill_2 FILLER_10_411 ();
 sg13g2_fill_1 FILLER_10_418 ();
 sg13g2_decap_4 FILLER_10_451 ();
 sg13g2_fill_1 FILLER_10_467 ();
 sg13g2_fill_2 FILLER_10_495 ();
 sg13g2_fill_2 FILLER_10_654 ();
 sg13g2_fill_2 FILLER_10_661 ();
 sg13g2_fill_1 FILLER_10_663 ();
 sg13g2_fill_2 FILLER_10_668 ();
 sg13g2_fill_2 FILLER_10_720 ();
 sg13g2_fill_1 FILLER_10_722 ();
 sg13g2_decap_4 FILLER_10_755 ();
 sg13g2_fill_2 FILLER_10_759 ();
 sg13g2_fill_2 FILLER_10_767 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_128 ();
 sg13g2_decap_4 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_233 ();
 sg13g2_fill_2 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_4 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_4 FILLER_11_432 ();
 sg13g2_fill_2 FILLER_11_436 ();
 sg13g2_decap_4 FILLER_11_442 ();
 sg13g2_fill_1 FILLER_11_459 ();
 sg13g2_decap_4 FILLER_11_469 ();
 sg13g2_fill_1 FILLER_11_473 ();
 sg13g2_decap_4 FILLER_11_478 ();
 sg13g2_decap_4 FILLER_11_486 ();
 sg13g2_fill_1 FILLER_11_503 ();
 sg13g2_fill_1 FILLER_11_514 ();
 sg13g2_decap_8 FILLER_11_561 ();
 sg13g2_decap_4 FILLER_11_568 ();
 sg13g2_fill_1 FILLER_11_585 ();
 sg13g2_fill_1 FILLER_11_599 ();
 sg13g2_decap_4 FILLER_11_604 ();
 sg13g2_fill_2 FILLER_11_608 ();
 sg13g2_fill_2 FILLER_11_625 ();
 sg13g2_fill_1 FILLER_11_627 ();
 sg13g2_decap_4 FILLER_11_636 ();
 sg13g2_decap_4 FILLER_11_702 ();
 sg13g2_fill_1 FILLER_11_706 ();
 sg13g2_fill_1 FILLER_11_720 ();
 sg13g2_fill_2 FILLER_11_725 ();
 sg13g2_fill_1 FILLER_11_727 ();
 sg13g2_fill_2 FILLER_11_742 ();
 sg13g2_fill_2 FILLER_11_759 ();
 sg13g2_fill_1 FILLER_11_761 ();
 sg13g2_decap_4 FILLER_11_781 ();
 sg13g2_fill_1 FILLER_11_785 ();
 sg13g2_fill_2 FILLER_11_795 ();
 sg13g2_fill_2 FILLER_11_802 ();
 sg13g2_fill_1 FILLER_11_804 ();
 sg13g2_fill_1 FILLER_11_810 ();
 sg13g2_fill_1 FILLER_11_820 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_43 ();
 sg13g2_fill_2 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_348 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_2 FILLER_12_366 ();
 sg13g2_fill_1 FILLER_12_368 ();
 sg13g2_decap_4 FILLER_12_378 ();
 sg13g2_decap_4 FILLER_12_386 ();
 sg13g2_fill_2 FILLER_12_403 ();
 sg13g2_fill_1 FILLER_12_405 ();
 sg13g2_fill_1 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_541 ();
 sg13g2_fill_1 FILLER_12_583 ();
 sg13g2_fill_2 FILLER_12_620 ();
 sg13g2_fill_2 FILLER_12_626 ();
 sg13g2_decap_4 FILLER_12_641 ();
 sg13g2_fill_2 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_651 ();
 sg13g2_fill_1 FILLER_12_657 ();
 sg13g2_decap_4 FILLER_12_662 ();
 sg13g2_fill_1 FILLER_12_666 ();
 sg13g2_fill_2 FILLER_12_768 ();
 sg13g2_fill_1 FILLER_12_775 ();
 sg13g2_fill_2 FILLER_12_803 ();
 sg13g2_fill_1 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_decap_4 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_decap_4 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_4 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_370 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_13_417 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_decap_8 FILLER_13_461 ();
 sg13g2_decap_8 FILLER_13_468 ();
 sg13g2_fill_1 FILLER_13_492 ();
 sg13g2_fill_1 FILLER_13_506 ();
 sg13g2_fill_2 FILLER_13_523 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_fill_2 FILLER_13_536 ();
 sg13g2_fill_1 FILLER_13_538 ();
 sg13g2_decap_8 FILLER_13_566 ();
 sg13g2_fill_1 FILLER_13_573 ();
 sg13g2_decap_4 FILLER_13_578 ();
 sg13g2_fill_1 FILLER_13_582 ();
 sg13g2_decap_4 FILLER_13_604 ();
 sg13g2_fill_1 FILLER_13_644 ();
 sg13g2_decap_4 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_710 ();
 sg13g2_fill_2 FILLER_13_726 ();
 sg13g2_fill_1 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_747 ();
 sg13g2_decap_8 FILLER_13_754 ();
 sg13g2_decap_4 FILLER_13_761 ();
 sg13g2_decap_4 FILLER_13_786 ();
 sg13g2_fill_2 FILLER_13_790 ();
 sg13g2_fill_2 FILLER_13_811 ();
 sg13g2_fill_1 FILLER_13_813 ();
 sg13g2_fill_1 FILLER_13_819 ();
 sg13g2_fill_1 FILLER_13_829 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_38 ();
 sg13g2_fill_1 FILLER_14_40 ();
 sg13g2_fill_2 FILLER_14_54 ();
 sg13g2_decap_8 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_86 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_100 ();
 sg13g2_decap_4 FILLER_14_111 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_decap_4 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_4 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_4 FILLER_14_434 ();
 sg13g2_decap_4 FILLER_14_514 ();
 sg13g2_fill_1 FILLER_14_545 ();
 sg13g2_fill_2 FILLER_14_616 ();
 sg13g2_decap_4 FILLER_14_622 ();
 sg13g2_fill_1 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_636 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_fill_1 FILLER_14_650 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_4 FILLER_14_662 ();
 sg13g2_fill_1 FILLER_14_666 ();
 sg13g2_fill_2 FILLER_14_699 ();
 sg13g2_fill_1 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_fill_1 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_799 ();
 sg13g2_fill_1 FILLER_14_806 ();
 sg13g2_fill_2 FILLER_14_826 ();
 sg13g2_fill_1 FILLER_14_828 ();
 sg13g2_fill_1 FILLER_14_834 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_285 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_fill_2 FILLER_15_409 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_decap_4 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_15_433 ();
 sg13g2_fill_2 FILLER_15_451 ();
 sg13g2_fill_1 FILLER_15_453 ();
 sg13g2_decap_8 FILLER_15_475 ();
 sg13g2_decap_4 FILLER_15_482 ();
 sg13g2_fill_2 FILLER_15_490 ();
 sg13g2_fill_2 FILLER_15_497 ();
 sg13g2_fill_1 FILLER_15_499 ();
 sg13g2_decap_8 FILLER_15_512 ();
 sg13g2_fill_2 FILLER_15_519 ();
 sg13g2_decap_4 FILLER_15_529 ();
 sg13g2_fill_2 FILLER_15_542 ();
 sg13g2_fill_1 FILLER_15_544 ();
 sg13g2_decap_4 FILLER_15_558 ();
 sg13g2_fill_2 FILLER_15_571 ();
 sg13g2_decap_4 FILLER_15_578 ();
 sg13g2_fill_1 FILLER_15_582 ();
 sg13g2_fill_2 FILLER_15_587 ();
 sg13g2_fill_1 FILLER_15_612 ();
 sg13g2_fill_1 FILLER_15_640 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_fill_2 FILLER_15_675 ();
 sg13g2_fill_1 FILLER_15_681 ();
 sg13g2_fill_2 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_706 ();
 sg13g2_fill_2 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_731 ();
 sg13g2_fill_1 FILLER_15_733 ();
 sg13g2_fill_2 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_853 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_10 ();
 sg13g2_decap_4 FILLER_16_17 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_41 ();
 sg13g2_decap_4 FILLER_16_46 ();
 sg13g2_fill_2 FILLER_16_50 ();
 sg13g2_decap_8 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_85 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_135 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_decap_4 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_4 FILLER_16_252 ();
 sg13g2_decap_4 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_400 ();
 sg13g2_decap_4 FILLER_16_433 ();
 sg13g2_fill_2 FILLER_16_510 ();
 sg13g2_fill_2 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_549 ();
 sg13g2_fill_1 FILLER_16_551 ();
 sg13g2_fill_2 FILLER_16_565 ();
 sg13g2_fill_1 FILLER_16_567 ();
 sg13g2_fill_1 FILLER_16_616 ();
 sg13g2_decap_4 FILLER_16_636 ();
 sg13g2_fill_2 FILLER_16_649 ();
 sg13g2_fill_2 FILLER_16_678 ();
 sg13g2_fill_1 FILLER_16_680 ();
 sg13g2_fill_2 FILLER_16_708 ();
 sg13g2_fill_1 FILLER_16_710 ();
 sg13g2_fill_1 FILLER_16_738 ();
 sg13g2_decap_4 FILLER_16_743 ();
 sg13g2_fill_2 FILLER_16_747 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_fill_2 FILLER_16_791 ();
 sg13g2_fill_1 FILLER_16_793 ();
 sg13g2_fill_2 FILLER_16_823 ();
 sg13g2_fill_1 FILLER_16_843 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_34 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_decap_8 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_decap_4 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_decap_4 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_4 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_4 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_358 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_decap_4 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_435 ();
 sg13g2_fill_2 FILLER_17_442 ();
 sg13g2_fill_1 FILLER_17_448 ();
 sg13g2_fill_2 FILLER_17_457 ();
 sg13g2_fill_1 FILLER_17_459 ();
 sg13g2_decap_8 FILLER_17_488 ();
 sg13g2_fill_2 FILLER_17_513 ();
 sg13g2_fill_2 FILLER_17_519 ();
 sg13g2_decap_4 FILLER_17_533 ();
 sg13g2_decap_4 FILLER_17_542 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_fill_1 FILLER_17_571 ();
 sg13g2_fill_1 FILLER_17_580 ();
 sg13g2_decap_4 FILLER_17_585 ();
 sg13g2_fill_1 FILLER_17_589 ();
 sg13g2_fill_2 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_607 ();
 sg13g2_decap_4 FILLER_17_641 ();
 sg13g2_decap_8 FILLER_17_653 ();
 sg13g2_decap_8 FILLER_17_660 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_2 FILLER_17_696 ();
 sg13g2_fill_1 FILLER_17_702 ();
 sg13g2_decap_4 FILLER_17_712 ();
 sg13g2_decap_8 FILLER_17_720 ();
 sg13g2_fill_2 FILLER_17_727 ();
 sg13g2_fill_1 FILLER_17_729 ();
 sg13g2_fill_2 FILLER_17_749 ();
 sg13g2_fill_1 FILLER_17_751 ();
 sg13g2_fill_1 FILLER_17_789 ();
 sg13g2_fill_2 FILLER_17_803 ();
 sg13g2_fill_1 FILLER_17_805 ();
 sg13g2_fill_1 FILLER_17_812 ();
 sg13g2_fill_2 FILLER_17_822 ();
 sg13g2_fill_1 FILLER_17_824 ();
 sg13g2_decap_8 FILLER_17_852 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_11 ();
 sg13g2_fill_2 FILLER_18_15 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_fill_1 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_decap_4 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_331 ();
 sg13g2_decap_4 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_fill_1 FILLER_18_414 ();
 sg13g2_fill_2 FILLER_18_460 ();
 sg13g2_fill_1 FILLER_18_462 ();
 sg13g2_fill_2 FILLER_18_540 ();
 sg13g2_fill_1 FILLER_18_569 ();
 sg13g2_fill_2 FILLER_18_608 ();
 sg13g2_fill_2 FILLER_18_627 ();
 sg13g2_fill_1 FILLER_18_629 ();
 sg13g2_fill_1 FILLER_18_639 ();
 sg13g2_fill_1 FILLER_18_667 ();
 sg13g2_fill_1 FILLER_18_685 ();
 sg13g2_fill_1 FILLER_18_705 ();
 sg13g2_decap_4 FILLER_18_710 ();
 sg13g2_fill_2 FILLER_18_714 ();
 sg13g2_fill_2 FILLER_18_769 ();
 sg13g2_fill_1 FILLER_18_812 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_41 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_92 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_4 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_fill_1 FILLER_19_444 ();
 sg13g2_fill_2 FILLER_19_489 ();
 sg13g2_fill_1 FILLER_19_491 ();
 sg13g2_decap_4 FILLER_19_501 ();
 sg13g2_fill_2 FILLER_19_505 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_fill_2 FILLER_19_532 ();
 sg13g2_fill_1 FILLER_19_592 ();
 sg13g2_fill_1 FILLER_19_603 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_fill_2 FILLER_19_657 ();
 sg13g2_fill_2 FILLER_19_684 ();
 sg13g2_fill_1 FILLER_19_686 ();
 sg13g2_fill_2 FILLER_19_699 ();
 sg13g2_fill_2 FILLER_19_742 ();
 sg13g2_fill_1 FILLER_19_744 ();
 sg13g2_decap_4 FILLER_19_795 ();
 sg13g2_decap_4 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_4 FILLER_19_858 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_10 ();
 sg13g2_fill_2 FILLER_20_17 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_decap_4 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_4 FILLER_20_431 ();
 sg13g2_fill_1 FILLER_20_435 ();
 sg13g2_decap_4 FILLER_20_462 ();
 sg13g2_decap_4 FILLER_20_470 ();
 sg13g2_fill_2 FILLER_20_474 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_fill_2 FILLER_20_511 ();
 sg13g2_fill_2 FILLER_20_526 ();
 sg13g2_fill_1 FILLER_20_528 ();
 sg13g2_fill_2 FILLER_20_646 ();
 sg13g2_fill_1 FILLER_20_648 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_fill_1 FILLER_20_707 ();
 sg13g2_fill_1 FILLER_20_758 ();
 sg13g2_fill_2 FILLER_20_803 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_fill_2 FILLER_20_833 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_4 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_decap_4 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_4 FILLER_21_375 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_decap_4 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_fill_2 FILLER_21_434 ();
 sg13g2_fill_1 FILLER_21_449 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_fill_2 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_490 ();
 sg13g2_fill_2 FILLER_21_518 ();
 sg13g2_decap_4 FILLER_21_525 ();
 sg13g2_fill_1 FILLER_21_533 ();
 sg13g2_fill_1 FILLER_21_613 ();
 sg13g2_fill_2 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_729 ();
 sg13g2_decap_4 FILLER_21_736 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_775 ();
 sg13g2_decap_4 FILLER_21_788 ();
 sg13g2_fill_1 FILLER_21_792 ();
 sg13g2_fill_1 FILLER_21_806 ();
 sg13g2_fill_1 FILLER_21_834 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_13 ();
 sg13g2_fill_1 FILLER_22_20 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_250 ();
 sg13g2_decap_4 FILLER_22_258 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_fill_1 FILLER_22_422 ();
 sg13g2_fill_2 FILLER_22_449 ();
 sg13g2_fill_1 FILLER_22_451 ();
 sg13g2_fill_1 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_fill_1 FILLER_22_513 ();
 sg13g2_fill_2 FILLER_22_541 ();
 sg13g2_fill_2 FILLER_22_576 ();
 sg13g2_fill_1 FILLER_22_578 ();
 sg13g2_fill_2 FILLER_22_607 ();
 sg13g2_fill_1 FILLER_22_658 ();
 sg13g2_fill_1 FILLER_22_706 ();
 sg13g2_fill_2 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_736 ();
 sg13g2_fill_1 FILLER_22_745 ();
 sg13g2_fill_2 FILLER_22_769 ();
 sg13g2_fill_2 FILLER_22_839 ();
 sg13g2_fill_1 FILLER_22_841 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_decap_4 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_decap_4 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_4 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_23_424 ();
 sg13g2_decap_4 FILLER_23_438 ();
 sg13g2_fill_2 FILLER_23_442 ();
 sg13g2_fill_2 FILLER_23_480 ();
 sg13g2_decap_4 FILLER_23_499 ();
 sg13g2_fill_2 FILLER_23_503 ();
 sg13g2_fill_1 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_523 ();
 sg13g2_fill_2 FILLER_23_533 ();
 sg13g2_fill_1 FILLER_23_535 ();
 sg13g2_fill_1 FILLER_23_555 ();
 sg13g2_fill_1 FILLER_23_578 ();
 sg13g2_fill_2 FILLER_23_588 ();
 sg13g2_fill_1 FILLER_23_600 ();
 sg13g2_decap_4 FILLER_23_614 ();
 sg13g2_fill_1 FILLER_23_618 ();
 sg13g2_fill_2 FILLER_23_725 ();
 sg13g2_fill_2 FILLER_23_731 ();
 sg13g2_fill_2 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_4 FILLER_23_777 ();
 sg13g2_decap_4 FILLER_23_785 ();
 sg13g2_fill_2 FILLER_23_789 ();
 sg13g2_fill_2 FILLER_23_800 ();
 sg13g2_decap_4 FILLER_23_812 ();
 sg13g2_fill_1 FILLER_23_816 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_27 ();
 sg13g2_fill_2 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_decap_4 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_decap_4 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_decap_4 FILLER_24_365 ();
 sg13g2_decap_4 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_400 ();
 sg13g2_fill_1 FILLER_24_433 ();
 sg13g2_fill_2 FILLER_24_461 ();
 sg13g2_fill_1 FILLER_24_476 ();
 sg13g2_fill_1 FILLER_24_483 ();
 sg13g2_decap_4 FILLER_24_511 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_fill_2 FILLER_24_521 ();
 sg13g2_fill_2 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_561 ();
 sg13g2_fill_2 FILLER_24_590 ();
 sg13g2_fill_1 FILLER_24_592 ();
 sg13g2_fill_2 FILLER_24_611 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_fill_2 FILLER_24_627 ();
 sg13g2_fill_1 FILLER_24_629 ();
 sg13g2_decap_4 FILLER_24_643 ();
 sg13g2_fill_1 FILLER_24_668 ();
 sg13g2_decap_4 FILLER_24_697 ();
 sg13g2_fill_1 FILLER_24_701 ();
 sg13g2_fill_2 FILLER_24_707 ();
 sg13g2_fill_2 FILLER_24_736 ();
 sg13g2_decap_4 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_fill_1 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_fill_1 FILLER_24_818 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_180 ();
 sg13g2_decap_4 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_4 FILLER_25_353 ();
 sg13g2_decap_4 FILLER_25_388 ();
 sg13g2_fill_2 FILLER_25_410 ();
 sg13g2_fill_2 FILLER_25_416 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_fill_1 FILLER_25_428 ();
 sg13g2_decap_4 FILLER_25_434 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_fill_2 FILLER_25_471 ();
 sg13g2_fill_1 FILLER_25_473 ();
 sg13g2_fill_1 FILLER_25_480 ();
 sg13g2_decap_4 FILLER_25_503 ();
 sg13g2_fill_2 FILLER_25_548 ();
 sg13g2_fill_1 FILLER_25_554 ();
 sg13g2_decap_4 FILLER_25_565 ();
 sg13g2_fill_2 FILLER_25_569 ();
 sg13g2_fill_1 FILLER_25_579 ();
 sg13g2_fill_2 FILLER_25_584 ();
 sg13g2_decap_4 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_612 ();
 sg13g2_decap_8 FILLER_25_619 ();
 sg13g2_fill_1 FILLER_25_626 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_fill_1 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_fill_2 FILLER_25_660 ();
 sg13g2_fill_1 FILLER_25_662 ();
 sg13g2_decap_4 FILLER_25_694 ();
 sg13g2_fill_1 FILLER_25_702 ();
 sg13g2_fill_2 FILLER_25_721 ();
 sg13g2_fill_1 FILLER_25_742 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_decap_4 FILLER_25_827 ();
 sg13g2_fill_2 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_decap_4 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_decap_4 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_460 ();
 sg13g2_fill_2 FILLER_26_518 ();
 sg13g2_fill_1 FILLER_26_562 ();
 sg13g2_decap_8 FILLER_26_601 ();
 sg13g2_fill_2 FILLER_26_608 ();
 sg13g2_decap_4 FILLER_26_637 ();
 sg13g2_fill_1 FILLER_26_667 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_fill_2 FILLER_26_679 ();
 sg13g2_fill_1 FILLER_26_681 ();
 sg13g2_fill_2 FILLER_26_687 ();
 sg13g2_fill_1 FILLER_26_689 ();
 sg13g2_fill_2 FILLER_26_699 ();
 sg13g2_fill_1 FILLER_26_701 ();
 sg13g2_fill_1 FILLER_26_759 ();
 sg13g2_fill_2 FILLER_26_766 ();
 sg13g2_fill_1 FILLER_26_768 ();
 sg13g2_fill_1 FILLER_26_777 ();
 sg13g2_fill_2 FILLER_26_800 ();
 sg13g2_fill_1 FILLER_26_802 ();
 sg13g2_fill_2 FILLER_26_829 ();
 sg13g2_fill_1 FILLER_26_831 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_decap_4 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_decap_4 FILLER_27_394 ();
 sg13g2_decap_4 FILLER_27_430 ();
 sg13g2_fill_1 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_fill_2 FILLER_27_452 ();
 sg13g2_fill_1 FILLER_27_454 ();
 sg13g2_fill_1 FILLER_27_480 ();
 sg13g2_decap_4 FILLER_27_496 ();
 sg13g2_fill_2 FILLER_27_513 ();
 sg13g2_fill_1 FILLER_27_515 ();
 sg13g2_fill_2 FILLER_27_583 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_fill_1 FILLER_27_608 ();
 sg13g2_fill_1 FILLER_27_614 ();
 sg13g2_fill_2 FILLER_27_623 ();
 sg13g2_fill_1 FILLER_27_693 ();
 sg13g2_fill_2 FILLER_27_727 ();
 sg13g2_fill_2 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_809 ();
 sg13g2_fill_2 FILLER_27_819 ();
 sg13g2_decap_4 FILLER_27_856 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_40 ();
 sg13g2_decap_4 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_decap_4 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_decap_4 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_28_434 ();
 sg13g2_fill_1 FILLER_28_491 ();
 sg13g2_fill_1 FILLER_28_546 ();
 sg13g2_fill_1 FILLER_28_569 ();
 sg13g2_decap_8 FILLER_28_597 ();
 sg13g2_fill_1 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_fill_2 FILLER_28_669 ();
 sg13g2_fill_1 FILLER_28_671 ();
 sg13g2_fill_1 FILLER_28_681 ();
 sg13g2_decap_4 FILLER_28_686 ();
 sg13g2_decap_4 FILLER_28_726 ();
 sg13g2_fill_1 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_fill_2 FILLER_28_788 ();
 sg13g2_fill_1 FILLER_28_790 ();
 sg13g2_fill_2 FILLER_28_832 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_13 ();
 sg13g2_fill_2 FILLER_29_17 ();
 sg13g2_decap_4 FILLER_29_29 ();
 sg13g2_fill_2 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_decap_8 FILLER_29_85 ();
 sg13g2_decap_8 FILLER_29_92 ();
 sg13g2_decap_4 FILLER_29_99 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_decap_4 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_428 ();
 sg13g2_fill_1 FILLER_29_437 ();
 sg13g2_decap_4 FILLER_29_453 ();
 sg13g2_fill_2 FILLER_29_467 ();
 sg13g2_fill_1 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_fill_2 FILLER_29_529 ();
 sg13g2_fill_2 FILLER_29_584 ();
 sg13g2_fill_1 FILLER_29_626 ();
 sg13g2_fill_1 FILLER_29_631 ();
 sg13g2_decap_4 FILLER_29_636 ();
 sg13g2_fill_1 FILLER_29_640 ();
 sg13g2_fill_1 FILLER_29_650 ();
 sg13g2_decap_4 FILLER_29_695 ();
 sg13g2_fill_2 FILLER_29_699 ();
 sg13g2_decap_4 FILLER_29_714 ();
 sg13g2_fill_2 FILLER_29_718 ();
 sg13g2_fill_2 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_792 ();
 sg13g2_decap_4 FILLER_29_799 ();
 sg13g2_fill_1 FILLER_29_809 ();
 sg13g2_fill_2 FILLER_29_815 ();
 sg13g2_fill_1 FILLER_29_817 ();
 sg13g2_decap_4 FILLER_29_822 ();
 sg13g2_fill_1 FILLER_29_830 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_decap_4 FILLER_30_185 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_409 ();
 sg13g2_decap_8 FILLER_30_452 ();
 sg13g2_fill_2 FILLER_30_491 ();
 sg13g2_fill_1 FILLER_30_493 ();
 sg13g2_fill_2 FILLER_30_507 ();
 sg13g2_fill_2 FILLER_30_559 ();
 sg13g2_fill_1 FILLER_30_561 ();
 sg13g2_fill_2 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_600 ();
 sg13g2_decap_8 FILLER_30_607 ();
 sg13g2_fill_2 FILLER_30_614 ();
 sg13g2_fill_1 FILLER_30_654 ();
 sg13g2_fill_1 FILLER_30_686 ();
 sg13g2_fill_2 FILLER_30_775 ();
 sg13g2_fill_1 FILLER_30_777 ();
 sg13g2_fill_2 FILLER_30_811 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_16 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_401 ();
 sg13g2_fill_2 FILLER_31_420 ();
 sg13g2_fill_2 FILLER_31_441 ();
 sg13g2_decap_4 FILLER_31_449 ();
 sg13g2_fill_1 FILLER_31_470 ();
 sg13g2_fill_2 FILLER_31_524 ();
 sg13g2_fill_1 FILLER_31_526 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_fill_2 FILLER_31_552 ();
 sg13g2_fill_2 FILLER_31_567 ();
 sg13g2_fill_2 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_624 ();
 sg13g2_fill_2 FILLER_31_678 ();
 sg13g2_fill_1 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_694 ();
 sg13g2_decap_4 FILLER_31_701 ();
 sg13g2_fill_1 FILLER_31_705 ();
 sg13g2_decap_4 FILLER_31_737 ();
 sg13g2_fill_2 FILLER_31_741 ();
 sg13g2_decap_4 FILLER_31_760 ();
 sg13g2_fill_1 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_fill_2 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_786 ();
 sg13g2_fill_2 FILLER_31_805 ();
 sg13g2_decap_4 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_4 FILLER_31_858 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_2 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_decap_4 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_197 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_decap_4 FILLER_32_213 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_decap_4 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_432 ();
 sg13g2_fill_1 FILLER_32_434 ();
 sg13g2_fill_2 FILLER_32_472 ();
 sg13g2_fill_2 FILLER_32_480 ();
 sg13g2_fill_1 FILLER_32_482 ();
 sg13g2_fill_1 FILLER_32_500 ();
 sg13g2_decap_8 FILLER_32_636 ();
 sg13g2_fill_2 FILLER_32_643 ();
 sg13g2_decap_4 FILLER_32_658 ();
 sg13g2_fill_2 FILLER_32_716 ();
 sg13g2_fill_1 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_fill_2 FILLER_32_755 ();
 sg13g2_fill_1 FILLER_32_771 ();
 sg13g2_fill_1 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_fill_1 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_decap_4 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_decap_4 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_420 ();
 sg13g2_fill_2 FILLER_33_448 ();
 sg13g2_fill_1 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_472 ();
 sg13g2_fill_1 FILLER_33_474 ();
 sg13g2_fill_2 FILLER_33_484 ();
 sg13g2_fill_1 FILLER_33_512 ();
 sg13g2_fill_1 FILLER_33_560 ();
 sg13g2_fill_1 FILLER_33_575 ();
 sg13g2_fill_1 FILLER_33_605 ();
 sg13g2_fill_1 FILLER_33_612 ();
 sg13g2_decap_8 FILLER_33_617 ();
 sg13g2_decap_8 FILLER_33_624 ();
 sg13g2_decap_8 FILLER_33_631 ();
 sg13g2_fill_2 FILLER_33_638 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_fill_2 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_666 ();
 sg13g2_decap_4 FILLER_33_671 ();
 sg13g2_fill_2 FILLER_33_675 ();
 sg13g2_decap_8 FILLER_33_681 ();
 sg13g2_fill_2 FILLER_33_688 ();
 sg13g2_fill_2 FILLER_33_716 ();
 sg13g2_fill_2 FILLER_33_758 ();
 sg13g2_fill_2 FILLER_33_791 ();
 sg13g2_fill_2 FILLER_33_799 ();
 sg13g2_fill_2 FILLER_33_842 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_29 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_4 FILLER_34_72 ();
 sg13g2_decap_4 FILLER_34_80 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_426 ();
 sg13g2_fill_2 FILLER_34_453 ();
 sg13g2_fill_1 FILLER_34_455 ();
 sg13g2_fill_2 FILLER_34_483 ();
 sg13g2_fill_1 FILLER_34_485 ();
 sg13g2_fill_2 FILLER_34_505 ();
 sg13g2_fill_2 FILLER_34_540 ();
 sg13g2_fill_1 FILLER_34_574 ();
 sg13g2_fill_2 FILLER_34_606 ();
 sg13g2_fill_2 FILLER_34_648 ();
 sg13g2_fill_2 FILLER_34_686 ();
 sg13g2_fill_1 FILLER_34_688 ();
 sg13g2_fill_2 FILLER_34_701 ();
 sg13g2_decap_4 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_743 ();
 sg13g2_fill_2 FILLER_34_753 ();
 sg13g2_fill_2 FILLER_34_773 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_fill_2 FILLER_34_833 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_9 ();
 sg13g2_fill_2 FILLER_35_16 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_decap_8 FILLER_35_36 ();
 sg13g2_decap_4 FILLER_35_43 ();
 sg13g2_fill_2 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_fill_2 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_decap_4 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_decap_4 FILLER_35_447 ();
 sg13g2_fill_2 FILLER_35_451 ();
 sg13g2_decap_4 FILLER_35_475 ();
 sg13g2_fill_1 FILLER_35_479 ();
 sg13g2_fill_1 FILLER_35_555 ();
 sg13g2_decap_4 FILLER_35_577 ();
 sg13g2_fill_1 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_586 ();
 sg13g2_fill_2 FILLER_35_593 ();
 sg13g2_fill_1 FILLER_35_595 ();
 sg13g2_fill_2 FILLER_35_614 ();
 sg13g2_fill_1 FILLER_35_634 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_670 ();
 sg13g2_fill_2 FILLER_35_677 ();
 sg13g2_decap_4 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_725 ();
 sg13g2_decap_4 FILLER_35_730 ();
 sg13g2_fill_2 FILLER_35_734 ();
 sg13g2_fill_1 FILLER_35_745 ();
 sg13g2_fill_2 FILLER_35_754 ();
 sg13g2_fill_1 FILLER_35_756 ();
 sg13g2_fill_2 FILLER_35_837 ();
 sg13g2_fill_1 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_165 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_decap_4 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_decap_4 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_fill_2 FILLER_36_411 ();
 sg13g2_fill_1 FILLER_36_413 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_fill_1 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_499 ();
 sg13g2_decap_8 FILLER_36_506 ();
 sg13g2_fill_1 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_4 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_640 ();
 sg13g2_fill_2 FILLER_36_701 ();
 sg13g2_fill_2 FILLER_36_707 ();
 sg13g2_fill_1 FILLER_36_709 ();
 sg13g2_fill_1 FILLER_36_719 ();
 sg13g2_decap_4 FILLER_36_733 ();
 sg13g2_decap_4 FILLER_36_746 ();
 sg13g2_fill_2 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_fill_1 FILLER_36_806 ();
 sg13g2_fill_2 FILLER_36_812 ();
 sg13g2_fill_1 FILLER_36_814 ();
 sg13g2_decap_4 FILLER_36_819 ();
 sg13g2_fill_2 FILLER_36_823 ();
 sg13g2_fill_2 FILLER_36_829 ();
 sg13g2_decap_4 FILLER_36_835 ();
 sg13g2_fill_1 FILLER_36_839 ();
 sg13g2_fill_2 FILLER_36_844 ();
 sg13g2_fill_1 FILLER_36_846 ();
 sg13g2_decap_4 FILLER_36_856 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_59 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_150 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_decap_4 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_decap_4 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_decap_4 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_37_414 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_1 FILLER_37_430 ();
 sg13g2_decap_8 FILLER_37_449 ();
 sg13g2_decap_4 FILLER_37_456 ();
 sg13g2_decap_4 FILLER_37_492 ();
 sg13g2_fill_2 FILLER_37_509 ();
 sg13g2_fill_1 FILLER_37_551 ();
 sg13g2_fill_2 FILLER_37_565 ();
 sg13g2_fill_2 FILLER_37_598 ();
 sg13g2_fill_2 FILLER_37_608 ();
 sg13g2_fill_1 FILLER_37_610 ();
 sg13g2_fill_2 FILLER_37_624 ();
 sg13g2_fill_1 FILLER_37_626 ();
 sg13g2_fill_2 FILLER_37_633 ();
 sg13g2_fill_1 FILLER_37_648 ();
 sg13g2_fill_2 FILLER_37_654 ();
 sg13g2_decap_4 FILLER_37_680 ();
 sg13g2_decap_4 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_752 ();
 sg13g2_fill_2 FILLER_37_758 ();
 sg13g2_fill_1 FILLER_37_760 ();
 sg13g2_fill_1 FILLER_37_819 ();
 sg13g2_fill_1 FILLER_37_825 ();
 sg13g2_fill_2 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_65 ();
 sg13g2_fill_1 FILLER_38_67 ();
 sg13g2_decap_4 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_decap_4 FILLER_38_128 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_153 ();
 sg13g2_decap_4 FILLER_38_168 ();
 sg13g2_decap_4 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_decap_4 FILLER_38_331 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_4 FILLER_38_445 ();
 sg13g2_fill_2 FILLER_38_449 ();
 sg13g2_fill_2 FILLER_38_464 ();
 sg13g2_fill_1 FILLER_38_466 ();
 sg13g2_decap_4 FILLER_38_489 ();
 sg13g2_fill_2 FILLER_38_493 ();
 sg13g2_fill_2 FILLER_38_521 ();
 sg13g2_fill_1 FILLER_38_523 ();
 sg13g2_fill_2 FILLER_38_537 ();
 sg13g2_fill_1 FILLER_38_539 ();
 sg13g2_fill_1 FILLER_38_553 ();
 sg13g2_fill_1 FILLER_38_564 ();
 sg13g2_fill_2 FILLER_38_604 ();
 sg13g2_fill_1 FILLER_38_606 ();
 sg13g2_decap_8 FILLER_38_634 ();
 sg13g2_fill_2 FILLER_38_702 ();
 sg13g2_fill_1 FILLER_38_704 ();
 sg13g2_fill_2 FILLER_38_714 ();
 sg13g2_fill_1 FILLER_38_716 ();
 sg13g2_fill_1 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_778 ();
 sg13g2_decap_4 FILLER_38_785 ();
 sg13g2_fill_2 FILLER_38_789 ();
 sg13g2_decap_4 FILLER_38_801 ();
 sg13g2_decap_4 FILLER_38_814 ();
 sg13g2_fill_1 FILLER_38_818 ();
 sg13g2_fill_2 FILLER_38_823 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_9 ();
 sg13g2_decap_8 FILLER_39_71 ();
 sg13g2_decap_8 FILLER_39_83 ();
 sg13g2_decap_8 FILLER_39_100 ();
 sg13g2_decap_8 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_138 ();
 sg13g2_fill_2 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_192 ();
 sg13g2_fill_1 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_282 ();
 sg13g2_fill_1 FILLER_39_284 ();
 sg13g2_decap_8 FILLER_39_290 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_318 ();
 sg13g2_decap_4 FILLER_39_365 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_4 FILLER_39_397 ();
 sg13g2_fill_1 FILLER_39_401 ();
 sg13g2_fill_2 FILLER_39_420 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_decap_8 FILLER_39_436 ();
 sg13g2_fill_2 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_489 ();
 sg13g2_fill_1 FILLER_39_496 ();
 sg13g2_fill_2 FILLER_39_510 ();
 sg13g2_fill_1 FILLER_39_512 ();
 sg13g2_fill_2 FILLER_39_526 ();
 sg13g2_fill_2 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_583 ();
 sg13g2_fill_2 FILLER_39_599 ();
 sg13g2_fill_2 FILLER_39_607 ();
 sg13g2_fill_2 FILLER_39_622 ();
 sg13g2_fill_2 FILLER_39_650 ();
 sg13g2_fill_2 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_663 ();
 sg13g2_decap_8 FILLER_39_670 ();
 sg13g2_decap_4 FILLER_39_677 ();
 sg13g2_fill_1 FILLER_39_713 ();
 sg13g2_fill_2 FILLER_39_726 ();
 sg13g2_fill_1 FILLER_39_728 ();
 sg13g2_fill_1 FILLER_39_755 ();
 sg13g2_fill_2 FILLER_39_765 ();
 sg13g2_fill_2 FILLER_39_788 ();
 sg13g2_decap_4 FILLER_39_806 ();
 sg13g2_fill_1 FILLER_39_819 ();
 sg13g2_fill_2 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_13 ();
 sg13g2_decap_8 FILLER_40_20 ();
 sg13g2_decap_8 FILLER_40_40 ();
 sg13g2_decap_4 FILLER_40_47 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_65 ();
 sg13g2_decap_8 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_78 ();
 sg13g2_fill_2 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_123 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_255 ();
 sg13g2_fill_1 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_288 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_decap_4 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_4 FILLER_40_362 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_4 FILLER_40_421 ();
 sg13g2_fill_1 FILLER_40_470 ();
 sg13g2_fill_2 FILLER_40_507 ();
 sg13g2_fill_1 FILLER_40_509 ();
 sg13g2_fill_2 FILLER_40_550 ();
 sg13g2_fill_1 FILLER_40_552 ();
 sg13g2_fill_2 FILLER_40_562 ();
 sg13g2_fill_1 FILLER_40_564 ();
 sg13g2_fill_2 FILLER_40_571 ();
 sg13g2_fill_1 FILLER_40_573 ();
 sg13g2_fill_1 FILLER_40_601 ();
 sg13g2_decap_4 FILLER_40_625 ();
 sg13g2_fill_2 FILLER_40_629 ();
 sg13g2_decap_4 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_644 ();
 sg13g2_decap_4 FILLER_40_702 ();
 sg13g2_fill_2 FILLER_40_706 ();
 sg13g2_decap_4 FILLER_40_717 ();
 sg13g2_fill_1 FILLER_40_721 ();
 sg13g2_fill_2 FILLER_40_824 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_111 ();
 sg13g2_fill_1 FILLER_41_113 ();
 sg13g2_fill_2 FILLER_41_127 ();
 sg13g2_fill_1 FILLER_41_129 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_fill_1 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_170 ();
 sg13g2_fill_1 FILLER_41_181 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_fill_1 FILLER_41_239 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_decap_4 FILLER_41_290 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_342 ();
 sg13g2_decap_4 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_386 ();
 sg13g2_fill_1 FILLER_41_388 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_492 ();
 sg13g2_fill_1 FILLER_41_542 ();
 sg13g2_fill_1 FILLER_41_588 ();
 sg13g2_fill_2 FILLER_41_609 ();
 sg13g2_decap_4 FILLER_41_647 ();
 sg13g2_decap_4 FILLER_41_655 ();
 sg13g2_fill_1 FILLER_41_659 ();
 sg13g2_fill_2 FILLER_41_674 ();
 sg13g2_decap_8 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_687 ();
 sg13g2_decap_8 FILLER_41_720 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_fill_1 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_fill_1 FILLER_41_784 ();
 sg13g2_fill_1 FILLER_41_816 ();
 sg13g2_fill_2 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_823 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_70 ();
 sg13g2_fill_2 FILLER_42_125 ();
 sg13g2_fill_2 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_213 ();
 sg13g2_fill_2 FILLER_42_220 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_258 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_decap_4 FILLER_42_271 ();
 sg13g2_fill_2 FILLER_42_275 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_decap_4 FILLER_42_320 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_decap_8 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_decap_4 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_decap_4 FILLER_42_397 ();
 sg13g2_fill_1 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_fill_1 FILLER_42_427 ();
 sg13g2_fill_2 FILLER_42_470 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_fill_2 FILLER_42_486 ();
 sg13g2_fill_2 FILLER_42_515 ();
 sg13g2_decap_8 FILLER_42_535 ();
 sg13g2_decap_4 FILLER_42_542 ();
 sg13g2_fill_1 FILLER_42_546 ();
 sg13g2_fill_2 FILLER_42_564 ();
 sg13g2_decap_4 FILLER_42_593 ();
 sg13g2_decap_4 FILLER_42_624 ();
 sg13g2_fill_2 FILLER_42_628 ();
 sg13g2_decap_8 FILLER_42_635 ();
 sg13g2_decap_4 FILLER_42_642 ();
 sg13g2_fill_2 FILLER_42_646 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_fill_2 FILLER_42_707 ();
 sg13g2_fill_1 FILLER_42_709 ();
 sg13g2_fill_1 FILLER_42_742 ();
 sg13g2_decap_4 FILLER_42_756 ();
 sg13g2_fill_2 FILLER_42_778 ();
 sg13g2_fill_1 FILLER_42_780 ();
 sg13g2_decap_4 FILLER_42_821 ();
 sg13g2_fill_1 FILLER_42_825 ();
 sg13g2_fill_2 FILLER_42_839 ();
 sg13g2_fill_1 FILLER_42_841 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_4 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_41 ();
 sg13g2_fill_2 FILLER_43_48 ();
 sg13g2_fill_1 FILLER_43_50 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_decap_8 FILLER_43_102 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_120 ();
 sg13g2_decap_4 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_decap_4 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_166 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_2 FILLER_43_213 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_280 ();
 sg13g2_decap_4 FILLER_43_290 ();
 sg13g2_fill_2 FILLER_43_294 ();
 sg13g2_decap_4 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_decap_4 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_decap_4 FILLER_43_334 ();
 sg13g2_fill_2 FILLER_43_338 ();
 sg13g2_fill_2 FILLER_43_352 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_4 FILLER_43_413 ();
 sg13g2_fill_1 FILLER_43_417 ();
 sg13g2_fill_2 FILLER_43_431 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_fill_2 FILLER_43_484 ();
 sg13g2_fill_1 FILLER_43_486 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_2 FILLER_43_510 ();
 sg13g2_fill_2 FILLER_43_521 ();
 sg13g2_fill_2 FILLER_43_550 ();
 sg13g2_fill_1 FILLER_43_552 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_4 FILLER_43_565 ();
 sg13g2_fill_2 FILLER_43_569 ();
 sg13g2_fill_2 FILLER_43_575 ();
 sg13g2_fill_1 FILLER_43_577 ();
 sg13g2_decap_4 FILLER_43_608 ();
 sg13g2_fill_2 FILLER_43_612 ();
 sg13g2_fill_1 FILLER_43_618 ();
 sg13g2_decap_4 FILLER_43_655 ();
 sg13g2_fill_1 FILLER_43_659 ();
 sg13g2_fill_2 FILLER_43_673 ();
 sg13g2_fill_1 FILLER_43_675 ();
 sg13g2_fill_1 FILLER_43_704 ();
 sg13g2_fill_2 FILLER_43_726 ();
 sg13g2_fill_1 FILLER_43_728 ();
 sg13g2_fill_2 FILLER_43_792 ();
 sg13g2_fill_1 FILLER_43_794 ();
 sg13g2_decap_4 FILLER_43_799 ();
 sg13g2_decap_8 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_850 ();
 sg13g2_decap_4 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_60 ();
 sg13g2_fill_1 FILLER_44_62 ();
 sg13g2_fill_1 FILLER_44_94 ();
 sg13g2_decap_4 FILLER_44_123 ();
 sg13g2_fill_2 FILLER_44_127 ();
 sg13g2_fill_2 FILLER_44_169 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_195 ();
 sg13g2_decap_8 FILLER_44_232 ();
 sg13g2_fill_1 FILLER_44_239 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_4 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_4 FILLER_44_392 ();
 sg13g2_decap_4 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_465 ();
 sg13g2_fill_2 FILLER_44_510 ();
 sg13g2_fill_1 FILLER_44_525 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_decap_4 FILLER_44_583 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_616 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_647 ();
 sg13g2_fill_1 FILLER_44_649 ();
 sg13g2_decap_4 FILLER_44_684 ();
 sg13g2_fill_1 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_fill_2 FILLER_44_732 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_decap_8 FILLER_44_748 ();
 sg13g2_fill_2 FILLER_44_755 ();
 sg13g2_fill_1 FILLER_44_757 ();
 sg13g2_fill_2 FILLER_44_776 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_4 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_36 ();
 sg13g2_decap_8 FILLER_45_43 ();
 sg13g2_decap_8 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_57 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_67 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_decap_4 FILLER_45_86 ();
 sg13g2_decap_4 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_143 ();
 sg13g2_fill_2 FILLER_45_150 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_304 ();
 sg13g2_fill_1 FILLER_45_310 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_410 ();
 sg13g2_fill_1 FILLER_45_412 ();
 sg13g2_fill_2 FILLER_45_422 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_fill_1 FILLER_45_442 ();
 sg13g2_fill_1 FILLER_45_456 ();
 sg13g2_decap_4 FILLER_45_467 ();
 sg13g2_fill_2 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_486 ();
 sg13g2_fill_2 FILLER_45_493 ();
 sg13g2_fill_1 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_500 ();
 sg13g2_decap_4 FILLER_45_521 ();
 sg13g2_decap_4 FILLER_45_528 ();
 sg13g2_fill_1 FILLER_45_532 ();
 sg13g2_decap_4 FILLER_45_560 ();
 sg13g2_fill_2 FILLER_45_564 ();
 sg13g2_decap_8 FILLER_45_575 ();
 sg13g2_fill_2 FILLER_45_582 ();
 sg13g2_fill_1 FILLER_45_602 ();
 sg13g2_fill_2 FILLER_45_648 ();
 sg13g2_fill_1 FILLER_45_650 ();
 sg13g2_fill_1 FILLER_45_678 ();
 sg13g2_fill_1 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_fill_2 FILLER_45_711 ();
 sg13g2_fill_1 FILLER_45_713 ();
 sg13g2_fill_2 FILLER_45_719 ();
 sg13g2_decap_4 FILLER_45_757 ();
 sg13g2_fill_1 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_53 ();
 sg13g2_fill_1 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_2 FILLER_46_111 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_126 ();
 sg13g2_fill_2 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_fill_2 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_353 ();
 sg13g2_fill_2 FILLER_46_367 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_decap_4 FILLER_46_383 ();
 sg13g2_fill_2 FILLER_46_403 ();
 sg13g2_fill_1 FILLER_46_405 ();
 sg13g2_decap_4 FILLER_46_414 ();
 sg13g2_fill_2 FILLER_46_418 ();
 sg13g2_fill_2 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_455 ();
 sg13g2_decap_4 FILLER_46_465 ();
 sg13g2_decap_4 FILLER_46_505 ();
 sg13g2_fill_2 FILLER_46_509 ();
 sg13g2_fill_2 FILLER_46_543 ();
 sg13g2_fill_1 FILLER_46_587 ();
 sg13g2_decap_8 FILLER_46_592 ();
 sg13g2_fill_2 FILLER_46_599 ();
 sg13g2_decap_8 FILLER_46_605 ();
 sg13g2_decap_4 FILLER_46_612 ();
 sg13g2_fill_2 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_622 ();
 sg13g2_fill_1 FILLER_46_629 ();
 sg13g2_fill_1 FILLER_46_643 ();
 sg13g2_fill_1 FILLER_46_667 ();
 sg13g2_fill_1 FILLER_46_686 ();
 sg13g2_fill_1 FILLER_46_728 ();
 sg13g2_fill_2 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_753 ();
 sg13g2_decap_4 FILLER_46_760 ();
 sg13g2_fill_2 FILLER_46_764 ();
 sg13g2_decap_4 FILLER_46_774 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_15 ();
 sg13g2_decap_8 FILLER_47_22 ();
 sg13g2_fill_1 FILLER_47_46 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_decap_4 FILLER_47_88 ();
 sg13g2_fill_2 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_102 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_fill_2 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_197 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_decap_8 FILLER_47_278 ();
 sg13g2_fill_2 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_fill_1 FILLER_47_299 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_fill_2 FILLER_47_342 ();
 sg13g2_fill_1 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_359 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_fill_1 FILLER_47_385 ();
 sg13g2_fill_1 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_440 ();
 sg13g2_fill_2 FILLER_47_447 ();
 sg13g2_fill_1 FILLER_47_449 ();
 sg13g2_fill_2 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_470 ();
 sg13g2_fill_1 FILLER_47_490 ();
 sg13g2_fill_2 FILLER_47_504 ();
 sg13g2_fill_1 FILLER_47_506 ();
 sg13g2_fill_1 FILLER_47_516 ();
 sg13g2_fill_1 FILLER_47_526 ();
 sg13g2_fill_2 FILLER_47_550 ();
 sg13g2_fill_1 FILLER_47_552 ();
 sg13g2_fill_1 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_621 ();
 sg13g2_fill_1 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_628 ();
 sg13g2_fill_1 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_decap_8 FILLER_47_647 ();
 sg13g2_fill_1 FILLER_47_654 ();
 sg13g2_fill_1 FILLER_47_691 ();
 sg13g2_fill_2 FILLER_47_698 ();
 sg13g2_fill_1 FILLER_47_736 ();
 sg13g2_decap_8 FILLER_47_764 ();
 sg13g2_decap_8 FILLER_47_771 ();
 sg13g2_decap_8 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_792 ();
 sg13g2_decap_8 FILLER_47_799 ();
 sg13g2_decap_8 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_decap_8 FILLER_47_834 ();
 sg13g2_decap_8 FILLER_47_841 ();
 sg13g2_decap_8 FILLER_47_848 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_45 ();
 sg13g2_fill_2 FILLER_48_54 ();
 sg13g2_fill_2 FILLER_48_68 ();
 sg13g2_decap_8 FILLER_48_92 ();
 sg13g2_decap_8 FILLER_48_99 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_fill_2 FILLER_48_141 ();
 sg13g2_fill_1 FILLER_48_143 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_209 ();
 sg13g2_fill_1 FILLER_48_211 ();
 sg13g2_decap_8 FILLER_48_276 ();
 sg13g2_decap_8 FILLER_48_283 ();
 sg13g2_fill_2 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_2 FILLER_48_320 ();
 sg13g2_fill_2 FILLER_48_412 ();
 sg13g2_fill_2 FILLER_48_441 ();
 sg13g2_fill_2 FILLER_48_475 ();
 sg13g2_fill_1 FILLER_48_481 ();
 sg13g2_fill_2 FILLER_48_522 ();
 sg13g2_fill_1 FILLER_48_524 ();
 sg13g2_decap_8 FILLER_48_530 ();
 sg13g2_decap_8 FILLER_48_537 ();
 sg13g2_decap_4 FILLER_48_544 ();
 sg13g2_fill_2 FILLER_48_557 ();
 sg13g2_fill_1 FILLER_48_559 ();
 sg13g2_fill_2 FILLER_48_570 ();
 sg13g2_fill_1 FILLER_48_612 ();
 sg13g2_decap_4 FILLER_48_646 ();
 sg13g2_fill_1 FILLER_48_650 ();
 sg13g2_fill_2 FILLER_48_656 ();
 sg13g2_fill_2 FILLER_48_679 ();
 sg13g2_decap_4 FILLER_48_685 ();
 sg13g2_fill_1 FILLER_48_692 ();
 sg13g2_fill_1 FILLER_48_724 ();
 sg13g2_fill_2 FILLER_48_734 ();
 sg13g2_fill_1 FILLER_48_736 ();
 sg13g2_fill_2 FILLER_48_746 ();
 sg13g2_decap_8 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_16 ();
 sg13g2_decap_8 FILLER_49_23 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_decap_4 FILLER_49_44 ();
 sg13g2_decap_4 FILLER_49_62 ();
 sg13g2_decap_4 FILLER_49_78 ();
 sg13g2_fill_1 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_fill_2 FILLER_49_144 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_173 ();
 sg13g2_fill_2 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_287 ();
 sg13g2_decap_4 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_4 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_330 ();
 sg13g2_fill_1 FILLER_49_344 ();
 sg13g2_decap_4 FILLER_49_360 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_2 FILLER_49_398 ();
 sg13g2_fill_1 FILLER_49_447 ();
 sg13g2_decap_4 FILLER_49_457 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_2 FILLER_49_481 ();
 sg13g2_fill_1 FILLER_49_483 ();
 sg13g2_decap_4 FILLER_49_505 ();
 sg13g2_decap_4 FILLER_49_513 ();
 sg13g2_fill_1 FILLER_49_517 ();
 sg13g2_decap_4 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_599 ();
 sg13g2_fill_2 FILLER_49_637 ();
 sg13g2_fill_1 FILLER_49_639 ();
 sg13g2_decap_4 FILLER_49_653 ();
 sg13g2_fill_2 FILLER_49_667 ();
 sg13g2_fill_1 FILLER_49_673 ();
 sg13g2_decap_8 FILLER_49_741 ();
 sg13g2_decap_8 FILLER_49_748 ();
 sg13g2_decap_8 FILLER_49_755 ();
 sg13g2_decap_8 FILLER_49_762 ();
 sg13g2_decap_8 FILLER_49_769 ();
 sg13g2_decap_8 FILLER_49_776 ();
 sg13g2_decap_8 FILLER_49_783 ();
 sg13g2_decap_8 FILLER_49_790 ();
 sg13g2_decap_8 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_804 ();
 sg13g2_decap_8 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_56 ();
 sg13g2_decap_4 FILLER_50_74 ();
 sg13g2_fill_2 FILLER_50_78 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_97 ();
 sg13g2_decap_8 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_4 FILLER_50_126 ();
 sg13g2_decap_4 FILLER_50_135 ();
 sg13g2_fill_1 FILLER_50_139 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_decap_4 FILLER_50_216 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_decap_4 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_decap_4 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_346 ();
 sg13g2_decap_4 FILLER_50_369 ();
 sg13g2_fill_2 FILLER_50_431 ();
 sg13g2_fill_1 FILLER_50_433 ();
 sg13g2_fill_1 FILLER_50_447 ();
 sg13g2_decap_8 FILLER_50_459 ();
 sg13g2_fill_2 FILLER_50_471 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_decap_4 FILLER_50_486 ();
 sg13g2_fill_2 FILLER_50_495 ();
 sg13g2_fill_1 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_508 ();
 sg13g2_fill_2 FILLER_50_515 ();
 sg13g2_fill_2 FILLER_50_522 ();
 sg13g2_decap_4 FILLER_50_536 ();
 sg13g2_decap_8 FILLER_50_549 ();
 sg13g2_decap_8 FILLER_50_556 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_fill_2 FILLER_50_616 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_fill_2 FILLER_50_625 ();
 sg13g2_fill_1 FILLER_50_627 ();
 sg13g2_fill_2 FILLER_50_668 ();
 sg13g2_fill_1 FILLER_50_670 ();
 sg13g2_fill_1 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_705 ();
 sg13g2_fill_1 FILLER_50_710 ();
 sg13g2_decap_8 FILLER_50_720 ();
 sg13g2_decap_4 FILLER_50_727 ();
 sg13g2_decap_8 FILLER_50_735 ();
 sg13g2_decap_8 FILLER_50_742 ();
 sg13g2_decap_8 FILLER_50_749 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_decap_8 FILLER_50_763 ();
 sg13g2_decap_8 FILLER_50_770 ();
 sg13g2_decap_8 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_784 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_fill_1 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_fill_2 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_232 ();
 sg13g2_fill_1 FILLER_51_234 ();
 sg13g2_decap_4 FILLER_51_284 ();
 sg13g2_decap_4 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_320 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_decap_8 FILLER_51_359 ();
 sg13g2_decap_8 FILLER_51_366 ();
 sg13g2_decap_4 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_386 ();
 sg13g2_fill_2 FILLER_51_424 ();
 sg13g2_decap_4 FILLER_51_440 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_fill_2 FILLER_51_468 ();
 sg13g2_fill_2 FILLER_51_481 ();
 sg13g2_decap_8 FILLER_51_503 ();
 sg13g2_fill_1 FILLER_51_510 ();
 sg13g2_fill_1 FILLER_51_521 ();
 sg13g2_decap_8 FILLER_51_533 ();
 sg13g2_fill_1 FILLER_51_540 ();
 sg13g2_decap_4 FILLER_51_547 ();
 sg13g2_fill_2 FILLER_51_577 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_decap_4 FILLER_51_651 ();
 sg13g2_decap_8 FILLER_51_669 ();
 sg13g2_fill_2 FILLER_51_691 ();
 sg13g2_fill_2 FILLER_51_707 ();
 sg13g2_fill_1 FILLER_51_709 ();
 sg13g2_decap_8 FILLER_51_723 ();
 sg13g2_decap_8 FILLER_51_730 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_decap_8 FILLER_51_744 ();
 sg13g2_decap_8 FILLER_51_751 ();
 sg13g2_decap_8 FILLER_51_758 ();
 sg13g2_decap_8 FILLER_51_765 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_786 ();
 sg13g2_decap_8 FILLER_51_793 ();
 sg13g2_decap_8 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_807 ();
 sg13g2_decap_8 FILLER_51_814 ();
 sg13g2_decap_8 FILLER_51_821 ();
 sg13g2_decap_8 FILLER_51_828 ();
 sg13g2_decap_8 FILLER_51_835 ();
 sg13g2_decap_8 FILLER_51_842 ();
 sg13g2_decap_8 FILLER_51_849 ();
 sg13g2_decap_4 FILLER_51_856 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_12 ();
 sg13g2_decap_8 FILLER_52_19 ();
 sg13g2_fill_1 FILLER_52_43 ();
 sg13g2_fill_1 FILLER_52_57 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_decap_4 FILLER_52_111 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_decap_4 FILLER_52_156 ();
 sg13g2_decap_4 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_222 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_decap_4 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_316 ();
 sg13g2_decap_8 FILLER_52_323 ();
 sg13g2_decap_8 FILLER_52_335 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_435 ();
 sg13g2_fill_1 FILLER_52_437 ();
 sg13g2_decap_8 FILLER_52_456 ();
 sg13g2_decap_4 FILLER_52_463 ();
 sg13g2_fill_1 FILLER_52_477 ();
 sg13g2_decap_8 FILLER_52_482 ();
 sg13g2_fill_2 FILLER_52_489 ();
 sg13g2_fill_2 FILLER_52_496 ();
 sg13g2_decap_4 FILLER_52_509 ();
 sg13g2_fill_2 FILLER_52_540 ();
 sg13g2_decap_8 FILLER_52_548 ();
 sg13g2_decap_4 FILLER_52_555 ();
 sg13g2_fill_2 FILLER_52_559 ();
 sg13g2_fill_2 FILLER_52_583 ();
 sg13g2_decap_4 FILLER_52_589 ();
 sg13g2_fill_1 FILLER_52_619 ();
 sg13g2_fill_1 FILLER_52_653 ();
 sg13g2_decap_4 FILLER_52_668 ();
 sg13g2_fill_1 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_727 ();
 sg13g2_decap_8 FILLER_52_734 ();
 sg13g2_decap_8 FILLER_52_741 ();
 sg13g2_decap_8 FILLER_52_748 ();
 sg13g2_decap_8 FILLER_52_755 ();
 sg13g2_decap_8 FILLER_52_762 ();
 sg13g2_decap_8 FILLER_52_769 ();
 sg13g2_decap_8 FILLER_52_776 ();
 sg13g2_decap_8 FILLER_52_783 ();
 sg13g2_decap_8 FILLER_52_790 ();
 sg13g2_decap_8 FILLER_52_797 ();
 sg13g2_decap_8 FILLER_52_804 ();
 sg13g2_decap_8 FILLER_52_811 ();
 sg13g2_decap_8 FILLER_52_818 ();
 sg13g2_decap_8 FILLER_52_825 ();
 sg13g2_decap_8 FILLER_52_832 ();
 sg13g2_decap_8 FILLER_52_839 ();
 sg13g2_decap_8 FILLER_52_846 ();
 sg13g2_decap_8 FILLER_52_853 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_4 ();
 sg13g2_fill_2 FILLER_53_42 ();
 sg13g2_fill_2 FILLER_53_48 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_1 FILLER_53_69 ();
 sg13g2_decap_8 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_89 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_118 ();
 sg13g2_decap_4 FILLER_53_133 ();
 sg13g2_decap_4 FILLER_53_148 ();
 sg13g2_decap_4 FILLER_53_167 ();
 sg13g2_decap_4 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_decap_4 FILLER_53_198 ();
 sg13g2_fill_1 FILLER_53_202 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_decap_8 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_decap_8 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_decap_4 FILLER_53_372 ();
 sg13g2_fill_1 FILLER_53_376 ();
 sg13g2_fill_1 FILLER_53_420 ();
 sg13g2_fill_2 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_432 ();
 sg13g2_decap_8 FILLER_53_461 ();
 sg13g2_fill_1 FILLER_53_468 ();
 sg13g2_fill_2 FILLER_53_481 ();
 sg13g2_fill_1 FILLER_53_483 ();
 sg13g2_fill_2 FILLER_53_489 ();
 sg13g2_fill_1 FILLER_53_491 ();
 sg13g2_decap_8 FILLER_53_513 ();
 sg13g2_fill_2 FILLER_53_520 ();
 sg13g2_fill_1 FILLER_53_533 ();
 sg13g2_decap_4 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_564 ();
 sg13g2_fill_1 FILLER_53_578 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_620 ();
 sg13g2_fill_2 FILLER_53_635 ();
 sg13g2_fill_1 FILLER_53_637 ();
 sg13g2_fill_2 FILLER_53_647 ();
 sg13g2_fill_1 FILLER_53_649 ();
 sg13g2_decap_8 FILLER_53_713 ();
 sg13g2_decap_8 FILLER_53_720 ();
 sg13g2_decap_8 FILLER_53_727 ();
 sg13g2_decap_8 FILLER_53_734 ();
 sg13g2_decap_8 FILLER_53_741 ();
 sg13g2_decap_8 FILLER_53_748 ();
 sg13g2_decap_8 FILLER_53_755 ();
 sg13g2_decap_8 FILLER_53_762 ();
 sg13g2_decap_8 FILLER_53_769 ();
 sg13g2_decap_8 FILLER_53_776 ();
 sg13g2_decap_8 FILLER_53_783 ();
 sg13g2_decap_8 FILLER_53_790 ();
 sg13g2_decap_8 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_804 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_decap_8 FILLER_53_818 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_15 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_99 ();
 sg13g2_fill_1 FILLER_54_101 ();
 sg13g2_fill_1 FILLER_54_136 ();
 sg13g2_decap_4 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_237 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_4 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_decap_8 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_284 ();
 sg13g2_decap_8 FILLER_54_289 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_fill_2 FILLER_54_316 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_decap_8 FILLER_54_324 ();
 sg13g2_decap_8 FILLER_54_331 ();
 sg13g2_decap_4 FILLER_54_338 ();
 sg13g2_fill_1 FILLER_54_342 ();
 sg13g2_decap_4 FILLER_54_359 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_418 ();
 sg13g2_decap_8 FILLER_54_433 ();
 sg13g2_decap_8 FILLER_54_458 ();
 sg13g2_decap_8 FILLER_54_465 ();
 sg13g2_fill_1 FILLER_54_472 ();
 sg13g2_fill_1 FILLER_54_494 ();
 sg13g2_decap_4 FILLER_54_509 ();
 sg13g2_fill_2 FILLER_54_513 ();
 sg13g2_decap_8 FILLER_54_528 ();
 sg13g2_fill_1 FILLER_54_535 ();
 sg13g2_fill_2 FILLER_54_569 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_2 FILLER_54_651 ();
 sg13g2_fill_1 FILLER_54_653 ();
 sg13g2_fill_2 FILLER_54_668 ();
 sg13g2_fill_1 FILLER_54_670 ();
 sg13g2_decap_4 FILLER_54_683 ();
 sg13g2_fill_2 FILLER_54_687 ();
 sg13g2_decap_8 FILLER_54_716 ();
 sg13g2_decap_8 FILLER_54_723 ();
 sg13g2_decap_8 FILLER_54_730 ();
 sg13g2_decap_8 FILLER_54_737 ();
 sg13g2_decap_8 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_758 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_8 FILLER_54_807 ();
 sg13g2_decap_8 FILLER_54_814 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_2 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_45 ();
 sg13g2_fill_2 FILLER_55_52 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_fill_2 FILLER_55_94 ();
 sg13g2_decap_4 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_fill_1 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_131 ();
 sg13g2_decap_4 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_142 ();
 sg13g2_decap_4 FILLER_55_158 ();
 sg13g2_fill_2 FILLER_55_182 ();
 sg13g2_decap_4 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_199 ();
 sg13g2_fill_1 FILLER_55_213 ();
 sg13g2_decap_4 FILLER_55_227 ();
 sg13g2_decap_4 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_decap_4 FILLER_55_274 ();
 sg13g2_decap_8 FILLER_55_323 ();
 sg13g2_decap_8 FILLER_55_330 ();
 sg13g2_decap_4 FILLER_55_337 ();
 sg13g2_fill_1 FILLER_55_341 ();
 sg13g2_fill_2 FILLER_55_362 ();
 sg13g2_fill_1 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_384 ();
 sg13g2_decap_8 FILLER_55_391 ();
 sg13g2_fill_2 FILLER_55_398 ();
 sg13g2_fill_1 FILLER_55_400 ();
 sg13g2_decap_4 FILLER_55_406 ();
 sg13g2_decap_4 FILLER_55_423 ();
 sg13g2_decap_8 FILLER_55_440 ();
 sg13g2_fill_1 FILLER_55_453 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_decap_8 FILLER_55_482 ();
 sg13g2_decap_4 FILLER_55_489 ();
 sg13g2_decap_8 FILLER_55_505 ();
 sg13g2_fill_2 FILLER_55_512 ();
 sg13g2_fill_1 FILLER_55_514 ();
 sg13g2_decap_4 FILLER_55_520 ();
 sg13g2_fill_2 FILLER_55_537 ();
 sg13g2_decap_8 FILLER_55_558 ();
 sg13g2_fill_2 FILLER_55_565 ();
 sg13g2_decap_4 FILLER_55_584 ();
 sg13g2_decap_8 FILLER_55_592 ();
 sg13g2_decap_8 FILLER_55_599 ();
 sg13g2_decap_4 FILLER_55_606 ();
 sg13g2_fill_1 FILLER_55_610 ();
 sg13g2_decap_4 FILLER_55_629 ();
 sg13g2_decap_8 FILLER_55_687 ();
 sg13g2_decap_8 FILLER_55_694 ();
 sg13g2_decap_8 FILLER_55_701 ();
 sg13g2_decap_8 FILLER_55_708 ();
 sg13g2_decap_8 FILLER_55_715 ();
 sg13g2_decap_8 FILLER_55_722 ();
 sg13g2_decap_8 FILLER_55_729 ();
 sg13g2_decap_8 FILLER_55_736 ();
 sg13g2_decap_8 FILLER_55_743 ();
 sg13g2_decap_8 FILLER_55_750 ();
 sg13g2_decap_8 FILLER_55_757 ();
 sg13g2_decap_8 FILLER_55_764 ();
 sg13g2_decap_8 FILLER_55_771 ();
 sg13g2_decap_8 FILLER_55_778 ();
 sg13g2_decap_8 FILLER_55_785 ();
 sg13g2_decap_8 FILLER_55_792 ();
 sg13g2_decap_8 FILLER_55_799 ();
 sg13g2_decap_8 FILLER_55_806 ();
 sg13g2_decap_8 FILLER_55_813 ();
 sg13g2_decap_8 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_827 ();
 sg13g2_decap_8 FILLER_55_834 ();
 sg13g2_decap_8 FILLER_55_841 ();
 sg13g2_decap_8 FILLER_55_848 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_17 ();
 sg13g2_fill_2 FILLER_56_33 ();
 sg13g2_fill_1 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_45 ();
 sg13g2_decap_8 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_61 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_78 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_2 FILLER_56_85 ();
 sg13g2_fill_1 FILLER_56_87 ();
 sg13g2_fill_2 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_141 ();
 sg13g2_decap_4 FILLER_56_162 ();
 sg13g2_fill_2 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_decap_4 FILLER_56_287 ();
 sg13g2_fill_1 FILLER_56_291 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_decap_4 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_369 ();
 sg13g2_decap_8 FILLER_56_386 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_4 FILLER_56_404 ();
 sg13g2_fill_2 FILLER_56_408 ();
 sg13g2_decap_4 FILLER_56_436 ();
 sg13g2_fill_2 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_473 ();
 sg13g2_fill_2 FILLER_56_488 ();
 sg13g2_fill_2 FILLER_56_508 ();
 sg13g2_fill_1 FILLER_56_510 ();
 sg13g2_fill_2 FILLER_56_520 ();
 sg13g2_fill_1 FILLER_56_522 ();
 sg13g2_decap_8 FILLER_56_536 ();
 sg13g2_decap_8 FILLER_56_549 ();
 sg13g2_decap_8 FILLER_56_556 ();
 sg13g2_fill_1 FILLER_56_563 ();
 sg13g2_fill_2 FILLER_56_581 ();
 sg13g2_decap_8 FILLER_56_610 ();
 sg13g2_decap_8 FILLER_56_617 ();
 sg13g2_decap_8 FILLER_56_624 ();
 sg13g2_decap_4 FILLER_56_649 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_1 FILLER_56_659 ();
 sg13g2_fill_1 FILLER_56_664 ();
 sg13g2_decap_8 FILLER_56_669 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_decap_8 FILLER_56_691 ();
 sg13g2_decap_8 FILLER_56_698 ();
 sg13g2_decap_8 FILLER_56_705 ();
 sg13g2_decap_8 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_8 FILLER_56_726 ();
 sg13g2_decap_8 FILLER_56_733 ();
 sg13g2_decap_8 FILLER_56_740 ();
 sg13g2_decap_8 FILLER_56_747 ();
 sg13g2_decap_8 FILLER_56_754 ();
 sg13g2_decap_8 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_768 ();
 sg13g2_decap_8 FILLER_56_775 ();
 sg13g2_decap_8 FILLER_56_782 ();
 sg13g2_decap_8 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_46 ();
 sg13g2_fill_2 FILLER_57_54 ();
 sg13g2_fill_2 FILLER_57_61 ();
 sg13g2_decap_4 FILLER_57_92 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_125 ();
 sg13g2_fill_1 FILLER_57_129 ();
 sg13g2_decap_8 FILLER_57_134 ();
 sg13g2_decap_8 FILLER_57_159 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_decap_4 FILLER_57_243 ();
 sg13g2_fill_1 FILLER_57_247 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_decap_8 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_4 FILLER_57_379 ();
 sg13g2_fill_1 FILLER_57_383 ();
 sg13g2_decap_4 FILLER_57_422 ();
 sg13g2_fill_2 FILLER_57_426 ();
 sg13g2_fill_2 FILLER_57_467 ();
 sg13g2_fill_1 FILLER_57_469 ();
 sg13g2_decap_4 FILLER_57_484 ();
 sg13g2_fill_2 FILLER_57_488 ();
 sg13g2_decap_4 FILLER_57_516 ();
 sg13g2_fill_2 FILLER_57_520 ();
 sg13g2_decap_8 FILLER_57_533 ();
 sg13g2_decap_4 FILLER_57_540 ();
 sg13g2_fill_1 FILLER_57_544 ();
 sg13g2_fill_2 FILLER_57_581 ();
 sg13g2_decap_4 FILLER_57_592 ();
 sg13g2_fill_1 FILLER_57_596 ();
 sg13g2_fill_2 FILLER_57_608 ();
 sg13g2_decap_4 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_617 ();
 sg13g2_decap_4 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_636 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_decap_8 FILLER_57_653 ();
 sg13g2_fill_2 FILLER_57_660 ();
 sg13g2_fill_1 FILLER_57_668 ();
 sg13g2_decap_8 FILLER_57_673 ();
 sg13g2_decap_8 FILLER_57_680 ();
 sg13g2_decap_8 FILLER_57_687 ();
 sg13g2_decap_8 FILLER_57_694 ();
 sg13g2_decap_8 FILLER_57_701 ();
 sg13g2_decap_8 FILLER_57_708 ();
 sg13g2_decap_8 FILLER_57_715 ();
 sg13g2_decap_8 FILLER_57_722 ();
 sg13g2_decap_8 FILLER_57_729 ();
 sg13g2_decap_8 FILLER_57_736 ();
 sg13g2_decap_8 FILLER_57_743 ();
 sg13g2_decap_8 FILLER_57_750 ();
 sg13g2_decap_8 FILLER_57_757 ();
 sg13g2_decap_8 FILLER_57_764 ();
 sg13g2_decap_8 FILLER_57_771 ();
 sg13g2_decap_8 FILLER_57_778 ();
 sg13g2_decap_8 FILLER_57_785 ();
 sg13g2_decap_8 FILLER_57_792 ();
 sg13g2_decap_8 FILLER_57_799 ();
 sg13g2_decap_8 FILLER_57_806 ();
 sg13g2_decap_8 FILLER_57_813 ();
 sg13g2_decap_8 FILLER_57_820 ();
 sg13g2_decap_8 FILLER_57_827 ();
 sg13g2_decap_8 FILLER_57_834 ();
 sg13g2_decap_8 FILLER_57_841 ();
 sg13g2_decap_8 FILLER_57_848 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_fill_1 FILLER_58_13 ();
 sg13g2_fill_2 FILLER_58_63 ();
 sg13g2_fill_1 FILLER_58_65 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_4 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_100 ();
 sg13g2_decap_4 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_111 ();
 sg13g2_decap_8 FILLER_58_130 ();
 sg13g2_decap_8 FILLER_58_137 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_fill_2 FILLER_58_158 ();
 sg13g2_fill_1 FILLER_58_160 ();
 sg13g2_decap_4 FILLER_58_202 ();
 sg13g2_fill_2 FILLER_58_224 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_264 ();
 sg13g2_fill_2 FILLER_58_293 ();
 sg13g2_fill_1 FILLER_58_295 ();
 sg13g2_decap_4 FILLER_58_300 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_decap_8 FILLER_58_333 ();
 sg13g2_decap_4 FILLER_58_340 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_358 ();
 sg13g2_decap_8 FILLER_58_367 ();
 sg13g2_fill_2 FILLER_58_400 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_457 ();
 sg13g2_fill_2 FILLER_58_472 ();
 sg13g2_decap_4 FILLER_58_487 ();
 sg13g2_fill_2 FILLER_58_491 ();
 sg13g2_fill_1 FILLER_58_506 ();
 sg13g2_decap_8 FILLER_58_524 ();
 sg13g2_fill_2 FILLER_58_544 ();
 sg13g2_fill_2 FILLER_58_564 ();
 sg13g2_fill_1 FILLER_58_566 ();
 sg13g2_fill_1 FILLER_58_580 ();
 sg13g2_fill_1 FILLER_58_596 ();
 sg13g2_decap_4 FILLER_58_619 ();
 sg13g2_fill_1 FILLER_58_623 ();
 sg13g2_fill_1 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_640 ();
 sg13g2_fill_1 FILLER_58_651 ();
 sg13g2_fill_2 FILLER_58_657 ();
 sg13g2_fill_1 FILLER_58_659 ();
 sg13g2_decap_8 FILLER_58_683 ();
 sg13g2_decap_8 FILLER_58_690 ();
 sg13g2_decap_8 FILLER_58_697 ();
 sg13g2_decap_8 FILLER_58_704 ();
 sg13g2_decap_8 FILLER_58_711 ();
 sg13g2_decap_8 FILLER_58_718 ();
 sg13g2_decap_8 FILLER_58_725 ();
 sg13g2_decap_8 FILLER_58_732 ();
 sg13g2_decap_8 FILLER_58_739 ();
 sg13g2_decap_8 FILLER_58_746 ();
 sg13g2_decap_8 FILLER_58_753 ();
 sg13g2_decap_8 FILLER_58_760 ();
 sg13g2_decap_8 FILLER_58_767 ();
 sg13g2_decap_8 FILLER_58_774 ();
 sg13g2_decap_8 FILLER_58_781 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_decap_8 FILLER_58_795 ();
 sg13g2_decap_8 FILLER_58_802 ();
 sg13g2_decap_8 FILLER_58_809 ();
 sg13g2_decap_8 FILLER_58_816 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_830 ();
 sg13g2_decap_8 FILLER_58_837 ();
 sg13g2_decap_8 FILLER_58_844 ();
 sg13g2_decap_8 FILLER_58_851 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_60 ();
 sg13g2_fill_2 FILLER_59_75 ();
 sg13g2_decap_8 FILLER_59_81 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_decap_8 FILLER_59_108 ();
 sg13g2_fill_2 FILLER_59_115 ();
 sg13g2_fill_1 FILLER_59_117 ();
 sg13g2_decap_4 FILLER_59_140 ();
 sg13g2_fill_2 FILLER_59_144 ();
 sg13g2_decap_8 FILLER_59_151 ();
 sg13g2_decap_8 FILLER_59_158 ();
 sg13g2_decap_8 FILLER_59_165 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_fill_1 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_282 ();
 sg13g2_decap_4 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_379 ();
 sg13g2_fill_2 FILLER_59_394 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_414 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_fill_2 FILLER_59_432 ();
 sg13g2_fill_2 FILLER_59_441 ();
 sg13g2_fill_1 FILLER_59_443 ();
 sg13g2_fill_2 FILLER_59_453 ();
 sg13g2_decap_4 FILLER_59_464 ();
 sg13g2_decap_8 FILLER_59_477 ();
 sg13g2_decap_8 FILLER_59_484 ();
 sg13g2_decap_4 FILLER_59_491 ();
 sg13g2_decap_8 FILLER_59_508 ();
 sg13g2_decap_4 FILLER_59_515 ();
 sg13g2_fill_2 FILLER_59_519 ();
 sg13g2_decap_8 FILLER_59_590 ();
 sg13g2_decap_4 FILLER_59_597 ();
 sg13g2_fill_1 FILLER_59_601 ();
 sg13g2_fill_2 FILLER_59_618 ();
 sg13g2_fill_1 FILLER_59_620 ();
 sg13g2_decap_8 FILLER_59_692 ();
 sg13g2_decap_8 FILLER_59_699 ();
 sg13g2_decap_8 FILLER_59_706 ();
 sg13g2_decap_8 FILLER_59_713 ();
 sg13g2_decap_8 FILLER_59_720 ();
 sg13g2_decap_8 FILLER_59_727 ();
 sg13g2_decap_8 FILLER_59_734 ();
 sg13g2_decap_8 FILLER_59_741 ();
 sg13g2_decap_8 FILLER_59_748 ();
 sg13g2_decap_8 FILLER_59_755 ();
 sg13g2_decap_8 FILLER_59_762 ();
 sg13g2_decap_8 FILLER_59_769 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_8 FILLER_59_797 ();
 sg13g2_decap_8 FILLER_59_804 ();
 sg13g2_decap_8 FILLER_59_811 ();
 sg13g2_decap_8 FILLER_59_818 ();
 sg13g2_decap_8 FILLER_59_825 ();
 sg13g2_decap_8 FILLER_59_832 ();
 sg13g2_decap_8 FILLER_59_839 ();
 sg13g2_decap_8 FILLER_59_846 ();
 sg13g2_decap_8 FILLER_59_853 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_11 ();
 sg13g2_fill_1 FILLER_60_15 ();
 sg13g2_fill_1 FILLER_60_47 ();
 sg13g2_fill_1 FILLER_60_61 ();
 sg13g2_decap_4 FILLER_60_115 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_150 ();
 sg13g2_decap_8 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_fill_2 FILLER_60_204 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_289 ();
 sg13g2_fill_1 FILLER_60_320 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_decap_4 FILLER_60_382 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_fill_2 FILLER_60_430 ();
 sg13g2_fill_1 FILLER_60_432 ();
 sg13g2_fill_1 FILLER_60_488 ();
 sg13g2_fill_2 FILLER_60_516 ();
 sg13g2_fill_1 FILLER_60_518 ();
 sg13g2_fill_1 FILLER_60_572 ();
 sg13g2_fill_2 FILLER_60_596 ();
 sg13g2_decap_8 FILLER_60_620 ();
 sg13g2_decap_8 FILLER_60_627 ();
 sg13g2_decap_4 FILLER_60_634 ();
 sg13g2_fill_2 FILLER_60_643 ();
 sg13g2_fill_1 FILLER_60_645 ();
 sg13g2_decap_8 FILLER_60_662 ();
 sg13g2_fill_1 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_680 ();
 sg13g2_decap_8 FILLER_60_687 ();
 sg13g2_decap_4 FILLER_60_694 ();
 sg13g2_fill_2 FILLER_60_698 ();
 sg13g2_decap_4 FILLER_60_704 ();
 sg13g2_fill_1 FILLER_60_708 ();
 sg13g2_decap_8 FILLER_60_714 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_decap_8 FILLER_60_725 ();
 sg13g2_decap_8 FILLER_60_732 ();
 sg13g2_decap_8 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_746 ();
 sg13g2_decap_8 FILLER_60_753 ();
 sg13g2_decap_8 FILLER_60_760 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_795 ();
 sg13g2_decap_8 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_decap_8 FILLER_60_851 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_30 ();
 sg13g2_fill_1 FILLER_61_71 ();
 sg13g2_fill_1 FILLER_61_82 ();
 sg13g2_decap_8 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_99 ();
 sg13g2_fill_1 FILLER_61_101 ();
 sg13g2_decap_4 FILLER_61_109 ();
 sg13g2_fill_2 FILLER_61_151 ();
 sg13g2_fill_1 FILLER_61_153 ();
 sg13g2_decap_8 FILLER_61_159 ();
 sg13g2_decap_4 FILLER_61_166 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_decap_8 FILLER_61_176 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_211 ();
 sg13g2_fill_2 FILLER_61_245 ();
 sg13g2_fill_2 FILLER_61_254 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_decap_8 FILLER_61_275 ();
 sg13g2_decap_8 FILLER_61_282 ();
 sg13g2_decap_4 FILLER_61_289 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_fill_1 FILLER_61_307 ();
 sg13g2_fill_2 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_decap_8 FILLER_61_339 ();
 sg13g2_decap_8 FILLER_61_346 ();
 sg13g2_decap_4 FILLER_61_375 ();
 sg13g2_fill_2 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_2 FILLER_61_422 ();
 sg13g2_fill_1 FILLER_61_424 ();
 sg13g2_decap_8 FILLER_61_456 ();
 sg13g2_fill_2 FILLER_61_463 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_decap_4 FILLER_61_492 ();
 sg13g2_fill_2 FILLER_61_512 ();
 sg13g2_fill_1 FILLER_61_524 ();
 sg13g2_fill_2 FILLER_61_581 ();
 sg13g2_fill_1 FILLER_61_583 ();
 sg13g2_fill_1 FILLER_61_611 ();
 sg13g2_fill_1 FILLER_61_625 ();
 sg13g2_decap_4 FILLER_61_643 ();
 sg13g2_decap_8 FILLER_61_652 ();
 sg13g2_decap_4 FILLER_61_659 ();
 sg13g2_fill_1 FILLER_61_663 ();
 sg13g2_fill_2 FILLER_61_668 ();
 sg13g2_decap_8 FILLER_61_674 ();
 sg13g2_decap_4 FILLER_61_681 ();
 sg13g2_decap_8 FILLER_61_740 ();
 sg13g2_decap_8 FILLER_61_747 ();
 sg13g2_decap_8 FILLER_61_754 ();
 sg13g2_decap_8 FILLER_61_761 ();
 sg13g2_decap_8 FILLER_61_768 ();
 sg13g2_decap_8 FILLER_61_775 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_decap_8 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_8 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_4 ();
 sg13g2_decap_8 FILLER_62_10 ();
 sg13g2_fill_2 FILLER_62_30 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_159 ();
 sg13g2_decap_8 FILLER_62_166 ();
 sg13g2_decap_8 FILLER_62_173 ();
 sg13g2_decap_8 FILLER_62_180 ();
 sg13g2_fill_2 FILLER_62_187 ();
 sg13g2_decap_4 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_fill_2 FILLER_62_235 ();
 sg13g2_decap_4 FILLER_62_255 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_decap_8 FILLER_62_281 ();
 sg13g2_decap_4 FILLER_62_288 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_decap_4 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_fill_1 FILLER_62_383 ();
 sg13g2_fill_1 FILLER_62_431 ();
 sg13g2_decap_4 FILLER_62_440 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_4 FILLER_62_464 ();
 sg13g2_decap_8 FILLER_62_484 ();
 sg13g2_decap_4 FILLER_62_491 ();
 sg13g2_fill_2 FILLER_62_495 ();
 sg13g2_fill_2 FILLER_62_512 ();
 sg13g2_decap_8 FILLER_62_541 ();
 sg13g2_fill_2 FILLER_62_548 ();
 sg13g2_fill_1 FILLER_62_550 ();
 sg13g2_fill_1 FILLER_62_600 ();
 sg13g2_decap_8 FILLER_62_621 ();
 sg13g2_decap_4 FILLER_62_628 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_decap_4 FILLER_62_648 ();
 sg13g2_fill_1 FILLER_62_652 ();
 sg13g2_fill_2 FILLER_62_657 ();
 sg13g2_decap_4 FILLER_62_717 ();
 sg13g2_decap_8 FILLER_62_748 ();
 sg13g2_decap_8 FILLER_62_755 ();
 sg13g2_decap_8 FILLER_62_762 ();
 sg13g2_decap_8 FILLER_62_769 ();
 sg13g2_decap_8 FILLER_62_776 ();
 sg13g2_decap_8 FILLER_62_783 ();
 sg13g2_decap_8 FILLER_62_790 ();
 sg13g2_decap_8 FILLER_62_797 ();
 sg13g2_decap_8 FILLER_62_804 ();
 sg13g2_decap_8 FILLER_62_811 ();
 sg13g2_decap_8 FILLER_62_818 ();
 sg13g2_decap_8 FILLER_62_825 ();
 sg13g2_decap_8 FILLER_62_832 ();
 sg13g2_decap_8 FILLER_62_839 ();
 sg13g2_decap_8 FILLER_62_846 ();
 sg13g2_decap_8 FILLER_62_853 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_fill_2 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_107 ();
 sg13g2_decap_4 FILLER_63_111 ();
 sg13g2_fill_1 FILLER_63_115 ();
 sg13g2_fill_1 FILLER_63_131 ();
 sg13g2_fill_2 FILLER_63_142 ();
 sg13g2_decap_8 FILLER_63_153 ();
 sg13g2_decap_8 FILLER_63_160 ();
 sg13g2_fill_2 FILLER_63_167 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_fill_2 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_decap_4 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_342 ();
 sg13g2_decap_4 FILLER_63_350 ();
 sg13g2_fill_1 FILLER_63_354 ();
 sg13g2_decap_4 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_388 ();
 sg13g2_decap_4 FILLER_63_393 ();
 sg13g2_decap_8 FILLER_63_411 ();
 sg13g2_decap_4 FILLER_63_418 ();
 sg13g2_fill_1 FILLER_63_422 ();
 sg13g2_fill_2 FILLER_63_435 ();
 sg13g2_fill_1 FILLER_63_437 ();
 sg13g2_fill_2 FILLER_63_443 ();
 sg13g2_fill_2 FILLER_63_464 ();
 sg13g2_fill_1 FILLER_63_466 ();
 sg13g2_decap_8 FILLER_63_488 ();
 sg13g2_fill_2 FILLER_63_495 ();
 sg13g2_fill_1 FILLER_63_501 ();
 sg13g2_decap_4 FILLER_63_508 ();
 sg13g2_fill_2 FILLER_63_512 ();
 sg13g2_decap_4 FILLER_63_537 ();
 sg13g2_fill_2 FILLER_63_541 ();
 sg13g2_decap_4 FILLER_63_547 ();
 sg13g2_fill_1 FILLER_63_551 ();
 sg13g2_fill_2 FILLER_63_561 ();
 sg13g2_fill_1 FILLER_63_572 ();
 sg13g2_fill_1 FILLER_63_595 ();
 sg13g2_decap_4 FILLER_63_602 ();
 sg13g2_fill_1 FILLER_63_625 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_730 ();
 sg13g2_decap_8 FILLER_63_737 ();
 sg13g2_decap_8 FILLER_63_744 ();
 sg13g2_decap_8 FILLER_63_751 ();
 sg13g2_decap_8 FILLER_63_758 ();
 sg13g2_decap_8 FILLER_63_765 ();
 sg13g2_decap_8 FILLER_63_772 ();
 sg13g2_decap_8 FILLER_63_779 ();
 sg13g2_decap_8 FILLER_63_786 ();
 sg13g2_decap_8 FILLER_63_793 ();
 sg13g2_decap_8 FILLER_63_800 ();
 sg13g2_decap_8 FILLER_63_807 ();
 sg13g2_decap_8 FILLER_63_814 ();
 sg13g2_decap_8 FILLER_63_821 ();
 sg13g2_decap_8 FILLER_63_828 ();
 sg13g2_decap_8 FILLER_63_835 ();
 sg13g2_decap_8 FILLER_63_842 ();
 sg13g2_decap_8 FILLER_63_849 ();
 sg13g2_decap_4 FILLER_63_856 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_12 ();
 sg13g2_fill_1 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_132 ();
 sg13g2_decap_8 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_193 ();
 sg13g2_fill_2 FILLER_64_212 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_fill_2 FILLER_64_228 ();
 sg13g2_fill_2 FILLER_64_243 ();
 sg13g2_fill_1 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_258 ();
 sg13g2_fill_2 FILLER_64_277 ();
 sg13g2_decap_4 FILLER_64_287 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_309 ();
 sg13g2_fill_1 FILLER_64_319 ();
 sg13g2_decap_4 FILLER_64_325 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_391 ();
 sg13g2_decap_8 FILLER_64_402 ();
 sg13g2_fill_2 FILLER_64_409 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_decap_8 FILLER_64_435 ();
 sg13g2_decap_8 FILLER_64_447 ();
 sg13g2_fill_1 FILLER_64_454 ();
 sg13g2_fill_1 FILLER_64_464 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_fill_1 FILLER_64_478 ();
 sg13g2_decap_4 FILLER_64_487 ();
 sg13g2_fill_2 FILLER_64_491 ();
 sg13g2_decap_8 FILLER_64_515 ();
 sg13g2_decap_4 FILLER_64_533 ();
 sg13g2_fill_1 FILLER_64_570 ();
 sg13g2_decap_4 FILLER_64_601 ();
 sg13g2_fill_1 FILLER_64_605 ();
 sg13g2_decap_4 FILLER_64_611 ();
 sg13g2_decap_4 FILLER_64_619 ();
 sg13g2_fill_2 FILLER_64_627 ();
 sg13g2_fill_1 FILLER_64_629 ();
 sg13g2_fill_1 FILLER_64_640 ();
 sg13g2_fill_2 FILLER_64_650 ();
 sg13g2_fill_1 FILLER_64_652 ();
 sg13g2_fill_1 FILLER_64_681 ();
 sg13g2_fill_1 FILLER_64_701 ();
 sg13g2_fill_1 FILLER_64_711 ();
 sg13g2_decap_8 FILLER_64_730 ();
 sg13g2_decap_8 FILLER_64_737 ();
 sg13g2_decap_8 FILLER_64_744 ();
 sg13g2_decap_8 FILLER_64_751 ();
 sg13g2_decap_8 FILLER_64_758 ();
 sg13g2_decap_8 FILLER_64_765 ();
 sg13g2_decap_8 FILLER_64_772 ();
 sg13g2_decap_8 FILLER_64_779 ();
 sg13g2_decap_8 FILLER_64_786 ();
 sg13g2_decap_8 FILLER_64_793 ();
 sg13g2_decap_8 FILLER_64_800 ();
 sg13g2_decap_8 FILLER_64_807 ();
 sg13g2_decap_8 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_828 ();
 sg13g2_decap_8 FILLER_64_835 ();
 sg13g2_decap_8 FILLER_64_842 ();
 sg13g2_decap_8 FILLER_64_849 ();
 sg13g2_decap_4 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_78 ();
 sg13g2_decap_8 FILLER_65_93 ();
 sg13g2_fill_1 FILLER_65_100 ();
 sg13g2_fill_2 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_116 ();
 sg13g2_fill_2 FILLER_65_121 ();
 sg13g2_fill_1 FILLER_65_123 ();
 sg13g2_fill_2 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_130 ();
 sg13g2_decap_4 FILLER_65_135 ();
 sg13g2_fill_2 FILLER_65_139 ();
 sg13g2_decap_8 FILLER_65_155 ();
 sg13g2_fill_2 FILLER_65_162 ();
 sg13g2_decap_8 FILLER_65_185 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_2 FILLER_65_265 ();
 sg13g2_decap_4 FILLER_65_272 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_297 ();
 sg13g2_decap_4 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_4 FILLER_65_339 ();
 sg13g2_decap_8 FILLER_65_347 ();
 sg13g2_fill_1 FILLER_65_354 ();
 sg13g2_fill_2 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_442 ();
 sg13g2_fill_1 FILLER_65_468 ();
 sg13g2_decap_4 FILLER_65_490 ();
 sg13g2_fill_2 FILLER_65_494 ();
 sg13g2_decap_8 FILLER_65_512 ();
 sg13g2_decap_4 FILLER_65_539 ();
 sg13g2_fill_2 FILLER_65_543 ();
 sg13g2_fill_1 FILLER_65_575 ();
 sg13g2_decap_8 FILLER_65_580 ();
 sg13g2_fill_2 FILLER_65_587 ();
 sg13g2_decap_8 FILLER_65_593 ();
 sg13g2_fill_2 FILLER_65_638 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_fill_1 FILLER_65_651 ();
 sg13g2_decap_4 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_667 ();
 sg13g2_fill_1 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_751 ();
 sg13g2_decap_8 FILLER_65_758 ();
 sg13g2_decap_8 FILLER_65_765 ();
 sg13g2_decap_8 FILLER_65_772 ();
 sg13g2_decap_8 FILLER_65_779 ();
 sg13g2_decap_8 FILLER_65_786 ();
 sg13g2_decap_8 FILLER_65_793 ();
 sg13g2_decap_8 FILLER_65_800 ();
 sg13g2_decap_8 FILLER_65_807 ();
 sg13g2_decap_8 FILLER_65_814 ();
 sg13g2_decap_8 FILLER_65_821 ();
 sg13g2_decap_8 FILLER_65_828 ();
 sg13g2_decap_8 FILLER_65_835 ();
 sg13g2_decap_8 FILLER_65_842 ();
 sg13g2_decap_8 FILLER_65_849 ();
 sg13g2_decap_4 FILLER_65_856 ();
 sg13g2_fill_2 FILLER_65_860 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_9 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_18 ();
 sg13g2_fill_2 FILLER_66_44 ();
 sg13g2_decap_8 FILLER_66_101 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_fill_2 FILLER_66_144 ();
 sg13g2_fill_1 FILLER_66_146 ();
 sg13g2_decap_4 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_184 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_2 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_276 ();
 sg13g2_decap_4 FILLER_66_287 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_fill_2 FILLER_66_300 ();
 sg13g2_fill_2 FILLER_66_334 ();
 sg13g2_fill_1 FILLER_66_336 ();
 sg13g2_fill_1 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_decap_4 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_395 ();
 sg13g2_decap_4 FILLER_66_417 ();
 sg13g2_decap_8 FILLER_66_432 ();
 sg13g2_fill_2 FILLER_66_439 ();
 sg13g2_decap_8 FILLER_66_446 ();
 sg13g2_decap_8 FILLER_66_453 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_fill_1 FILLER_66_468 ();
 sg13g2_decap_8 FILLER_66_485 ();
 sg13g2_fill_2 FILLER_66_492 ();
 sg13g2_decap_8 FILLER_66_509 ();
 sg13g2_decap_8 FILLER_66_516 ();
 sg13g2_fill_2 FILLER_66_523 ();
 sg13g2_fill_2 FILLER_66_529 ();
 sg13g2_fill_2 FILLER_66_544 ();
 sg13g2_fill_1 FILLER_66_546 ();
 sg13g2_fill_2 FILLER_66_584 ();
 sg13g2_fill_1 FILLER_66_586 ();
 sg13g2_fill_1 FILLER_66_626 ();
 sg13g2_fill_1 FILLER_66_660 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_729 ();
 sg13g2_decap_8 FILLER_66_756 ();
 sg13g2_decap_8 FILLER_66_763 ();
 sg13g2_decap_8 FILLER_66_770 ();
 sg13g2_decap_8 FILLER_66_777 ();
 sg13g2_decap_8 FILLER_66_784 ();
 sg13g2_decap_8 FILLER_66_791 ();
 sg13g2_decap_8 FILLER_66_798 ();
 sg13g2_decap_8 FILLER_66_805 ();
 sg13g2_decap_8 FILLER_66_812 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_854 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_4 ();
 sg13g2_fill_1 FILLER_67_32 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_fill_2 FILLER_67_71 ();
 sg13g2_decap_8 FILLER_67_86 ();
 sg13g2_decap_8 FILLER_67_93 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_fill_2 FILLER_67_221 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_decap_4 FILLER_67_249 ();
 sg13g2_decap_4 FILLER_67_258 ();
 sg13g2_fill_1 FILLER_67_262 ();
 sg13g2_fill_2 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_278 ();
 sg13g2_decap_8 FILLER_67_289 ();
 sg13g2_fill_1 FILLER_67_346 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_fill_1 FILLER_67_373 ();
 sg13g2_fill_2 FILLER_67_378 ();
 sg13g2_fill_1 FILLER_67_380 ();
 sg13g2_fill_2 FILLER_67_405 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_fill_1 FILLER_67_430 ();
 sg13g2_fill_2 FILLER_67_441 ();
 sg13g2_fill_2 FILLER_67_457 ();
 sg13g2_decap_8 FILLER_67_478 ();
 sg13g2_decap_8 FILLER_67_485 ();
 sg13g2_decap_4 FILLER_67_492 ();
 sg13g2_fill_1 FILLER_67_496 ();
 sg13g2_decap_8 FILLER_67_512 ();
 sg13g2_fill_1 FILLER_67_519 ();
 sg13g2_fill_2 FILLER_67_525 ();
 sg13g2_fill_1 FILLER_67_544 ();
 sg13g2_fill_2 FILLER_67_554 ();
 sg13g2_fill_2 FILLER_67_583 ();
 sg13g2_fill_1 FILLER_67_585 ();
 sg13g2_fill_1 FILLER_67_628 ();
 sg13g2_decap_4 FILLER_67_642 ();
 sg13g2_decap_8 FILLER_67_750 ();
 sg13g2_decap_8 FILLER_67_757 ();
 sg13g2_decap_8 FILLER_67_764 ();
 sg13g2_decap_8 FILLER_67_771 ();
 sg13g2_decap_8 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_785 ();
 sg13g2_decap_8 FILLER_67_792 ();
 sg13g2_decap_8 FILLER_67_799 ();
 sg13g2_decap_8 FILLER_67_806 ();
 sg13g2_decap_8 FILLER_67_813 ();
 sg13g2_decap_8 FILLER_67_820 ();
 sg13g2_decap_8 FILLER_67_827 ();
 sg13g2_decap_8 FILLER_67_834 ();
 sg13g2_decap_8 FILLER_67_841 ();
 sg13g2_decap_8 FILLER_67_848 ();
 sg13g2_decap_8 FILLER_67_855 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_4 FILLER_68_10 ();
 sg13g2_fill_1 FILLER_68_38 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_92 ();
 sg13g2_fill_1 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_decap_8 FILLER_68_163 ();
 sg13g2_decap_8 FILLER_68_174 ();
 sg13g2_fill_2 FILLER_68_181 ();
 sg13g2_decap_4 FILLER_68_248 ();
 sg13g2_fill_1 FILLER_68_252 ();
 sg13g2_fill_2 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_decap_4 FILLER_68_263 ();
 sg13g2_fill_1 FILLER_68_275 ();
 sg13g2_decap_8 FILLER_68_293 ();
 sg13g2_decap_4 FILLER_68_337 ();
 sg13g2_fill_2 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_fill_2 FILLER_68_431 ();
 sg13g2_fill_2 FILLER_68_456 ();
 sg13g2_fill_2 FILLER_68_463 ();
 sg13g2_fill_1 FILLER_68_465 ();
 sg13g2_decap_8 FILLER_68_479 ();
 sg13g2_decap_4 FILLER_68_486 ();
 sg13g2_fill_1 FILLER_68_490 ();
 sg13g2_decap_8 FILLER_68_509 ();
 sg13g2_fill_2 FILLER_68_521 ();
 sg13g2_fill_2 FILLER_68_528 ();
 sg13g2_fill_1 FILLER_68_551 ();
 sg13g2_decap_4 FILLER_68_587 ();
 sg13g2_decap_8 FILLER_68_595 ();
 sg13g2_decap_4 FILLER_68_602 ();
 sg13g2_fill_1 FILLER_68_618 ();
 sg13g2_fill_2 FILLER_68_647 ();
 sg13g2_fill_1 FILLER_68_649 ();
 sg13g2_fill_1 FILLER_68_672 ();
 sg13g2_fill_2 FILLER_68_695 ();
 sg13g2_fill_2 FILLER_68_706 ();
 sg13g2_fill_1 FILLER_68_737 ();
 sg13g2_decap_8 FILLER_68_755 ();
 sg13g2_decap_8 FILLER_68_762 ();
 sg13g2_decap_8 FILLER_68_769 ();
 sg13g2_decap_8 FILLER_68_776 ();
 sg13g2_decap_8 FILLER_68_783 ();
 sg13g2_decap_8 FILLER_68_790 ();
 sg13g2_decap_8 FILLER_68_797 ();
 sg13g2_decap_8 FILLER_68_804 ();
 sg13g2_decap_8 FILLER_68_811 ();
 sg13g2_decap_8 FILLER_68_818 ();
 sg13g2_decap_8 FILLER_68_825 ();
 sg13g2_decap_8 FILLER_68_832 ();
 sg13g2_decap_8 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_fill_2 FILLER_68_860 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_fill_1 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_56 ();
 sg13g2_fill_2 FILLER_69_66 ();
 sg13g2_fill_1 FILLER_69_68 ();
 sg13g2_fill_2 FILLER_69_85 ();
 sg13g2_fill_1 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_116 ();
 sg13g2_fill_2 FILLER_69_122 ();
 sg13g2_decap_4 FILLER_69_151 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_205 ();
 sg13g2_decap_4 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_229 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_decap_4 FILLER_69_249 ();
 sg13g2_decap_8 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_289 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_305 ();
 sg13g2_fill_1 FILLER_69_322 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_decap_4 FILLER_69_364 ();
 sg13g2_fill_1 FILLER_69_368 ();
 sg13g2_fill_2 FILLER_69_402 ();
 sg13g2_fill_2 FILLER_69_428 ();
 sg13g2_fill_1 FILLER_69_430 ();
 sg13g2_decap_4 FILLER_69_435 ();
 sg13g2_fill_2 FILLER_69_439 ();
 sg13g2_decap_8 FILLER_69_453 ();
 sg13g2_decap_8 FILLER_69_481 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_506 ();
 sg13g2_fill_1 FILLER_69_508 ();
 sg13g2_fill_2 FILLER_69_575 ();
 sg13g2_fill_1 FILLER_69_618 ();
 sg13g2_fill_1 FILLER_69_632 ();
 sg13g2_decap_4 FILLER_69_642 ();
 sg13g2_fill_2 FILLER_69_659 ();
 sg13g2_decap_4 FILLER_69_696 ();
 sg13g2_fill_1 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_758 ();
 sg13g2_decap_8 FILLER_69_765 ();
 sg13g2_decap_8 FILLER_69_772 ();
 sg13g2_decap_8 FILLER_69_779 ();
 sg13g2_decap_8 FILLER_69_786 ();
 sg13g2_decap_8 FILLER_69_793 ();
 sg13g2_decap_8 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_807 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_26 ();
 sg13g2_fill_2 FILLER_70_36 ();
 sg13g2_fill_1 FILLER_70_103 ();
 sg13g2_decap_4 FILLER_70_136 ();
 sg13g2_decap_8 FILLER_70_153 ();
 sg13g2_fill_2 FILLER_70_160 ();
 sg13g2_fill_1 FILLER_70_162 ();
 sg13g2_decap_4 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_decap_4 FILLER_70_229 ();
 sg13g2_fill_1 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_296 ();
 sg13g2_fill_2 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_303 ();
 sg13g2_decap_4 FILLER_70_322 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_347 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_1 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_401 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_fill_1 FILLER_70_423 ();
 sg13g2_fill_2 FILLER_70_429 ();
 sg13g2_fill_1 FILLER_70_431 ();
 sg13g2_decap_4 FILLER_70_445 ();
 sg13g2_decap_4 FILLER_70_462 ();
 sg13g2_fill_2 FILLER_70_511 ();
 sg13g2_fill_2 FILLER_70_553 ();
 sg13g2_fill_1 FILLER_70_555 ();
 sg13g2_fill_1 FILLER_70_560 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_604 ();
 sg13g2_decap_8 FILLER_70_637 ();
 sg13g2_fill_2 FILLER_70_644 ();
 sg13g2_fill_1 FILLER_70_646 ();
 sg13g2_decap_4 FILLER_70_685 ();
 sg13g2_decap_8 FILLER_70_748 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_813 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_4 ();
 sg13g2_decap_4 FILLER_71_78 ();
 sg13g2_fill_2 FILLER_71_95 ();
 sg13g2_fill_2 FILLER_71_106 ();
 sg13g2_decap_4 FILLER_71_144 ();
 sg13g2_decap_4 FILLER_71_156 ();
 sg13g2_fill_1 FILLER_71_177 ();
 sg13g2_fill_2 FILLER_71_206 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_fill_2 FILLER_71_250 ();
 sg13g2_decap_8 FILLER_71_261 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_decap_4 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_fill_1 FILLER_71_297 ();
 sg13g2_fill_2 FILLER_71_311 ();
 sg13g2_fill_1 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_437 ();
 sg13g2_fill_1 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_537 ();
 sg13g2_decap_4 FILLER_71_542 ();
 sg13g2_fill_1 FILLER_71_546 ();
 sg13g2_fill_2 FILLER_71_568 ();
 sg13g2_fill_2 FILLER_71_579 ();
 sg13g2_fill_1 FILLER_71_598 ();
 sg13g2_decap_8 FILLER_71_608 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_fill_1 FILLER_71_630 ();
 sg13g2_fill_1 FILLER_71_645 ();
 sg13g2_decap_4 FILLER_71_681 ();
 sg13g2_fill_2 FILLER_71_685 ();
 sg13g2_fill_1 FILLER_71_714 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_21 ();
 sg13g2_fill_2 FILLER_72_134 ();
 sg13g2_fill_1 FILLER_72_136 ();
 sg13g2_fill_2 FILLER_72_156 ();
 sg13g2_decap_4 FILLER_72_164 ();
 sg13g2_decap_8 FILLER_72_239 ();
 sg13g2_fill_1 FILLER_72_267 ();
 sg13g2_decap_8 FILLER_72_277 ();
 sg13g2_decap_8 FILLER_72_284 ();
 sg13g2_fill_2 FILLER_72_291 ();
 sg13g2_fill_1 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_decap_4 FILLER_72_303 ();
 sg13g2_fill_2 FILLER_72_307 ();
 sg13g2_decap_4 FILLER_72_323 ();
 sg13g2_fill_2 FILLER_72_327 ();
 sg13g2_fill_2 FILLER_72_338 ();
 sg13g2_fill_2 FILLER_72_361 ();
 sg13g2_fill_1 FILLER_72_363 ();
 sg13g2_decap_4 FILLER_72_373 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_fill_1 FILLER_72_386 ();
 sg13g2_fill_2 FILLER_72_409 ();
 sg13g2_fill_1 FILLER_72_411 ();
 sg13g2_fill_2 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_427 ();
 sg13g2_fill_2 FILLER_72_437 ();
 sg13g2_fill_1 FILLER_72_439 ();
 sg13g2_fill_2 FILLER_72_453 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_475 ();
 sg13g2_decap_8 FILLER_72_482 ();
 sg13g2_fill_2 FILLER_72_489 ();
 sg13g2_decap_4 FILLER_72_495 ();
 sg13g2_fill_2 FILLER_72_507 ();
 sg13g2_decap_8 FILLER_72_513 ();
 sg13g2_fill_1 FILLER_72_601 ();
 sg13g2_fill_2 FILLER_72_629 ();
 sg13g2_decap_8 FILLER_72_667 ();
 sg13g2_decap_4 FILLER_72_674 ();
 sg13g2_fill_2 FILLER_72_678 ();
 sg13g2_fill_2 FILLER_72_737 ();
 sg13g2_decap_8 FILLER_72_775 ();
 sg13g2_decap_8 FILLER_72_782 ();
 sg13g2_decap_8 FILLER_72_789 ();
 sg13g2_decap_8 FILLER_72_796 ();
 sg13g2_decap_8 FILLER_72_803 ();
 sg13g2_decap_8 FILLER_72_810 ();
 sg13g2_decap_8 FILLER_72_817 ();
 sg13g2_decap_8 FILLER_72_824 ();
 sg13g2_decap_8 FILLER_72_831 ();
 sg13g2_decap_8 FILLER_72_838 ();
 sg13g2_decap_8 FILLER_72_845 ();
 sg13g2_decap_8 FILLER_72_852 ();
 sg13g2_fill_2 FILLER_72_859 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_52 ();
 sg13g2_fill_1 FILLER_73_54 ();
 sg13g2_decap_8 FILLER_73_64 ();
 sg13g2_fill_1 FILLER_73_71 ();
 sg13g2_fill_2 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_fill_2 FILLER_73_146 ();
 sg13g2_decap_8 FILLER_73_157 ();
 sg13g2_fill_1 FILLER_73_164 ();
 sg13g2_fill_2 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_222 ();
 sg13g2_fill_1 FILLER_73_224 ();
 sg13g2_fill_2 FILLER_73_235 ();
 sg13g2_decap_4 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_291 ();
 sg13g2_fill_1 FILLER_73_364 ();
 sg13g2_fill_2 FILLER_73_373 ();
 sg13g2_fill_1 FILLER_73_375 ();
 sg13g2_fill_1 FILLER_73_412 ();
 sg13g2_decap_8 FILLER_73_417 ();
 sg13g2_fill_2 FILLER_73_424 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_decap_4 FILLER_73_431 ();
 sg13g2_fill_2 FILLER_73_478 ();
 sg13g2_fill_1 FILLER_73_480 ();
 sg13g2_fill_2 FILLER_73_494 ();
 sg13g2_fill_1 FILLER_73_496 ();
 sg13g2_decap_4 FILLER_73_525 ();
 sg13g2_decap_8 FILLER_73_542 ();
 sg13g2_decap_4 FILLER_73_549 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_fill_2 FILLER_73_595 ();
 sg13g2_fill_1 FILLER_73_597 ();
 sg13g2_fill_1 FILLER_73_611 ();
 sg13g2_fill_2 FILLER_73_636 ();
 sg13g2_decap_8 FILLER_73_651 ();
 sg13g2_fill_1 FILLER_73_658 ();
 sg13g2_decap_8 FILLER_73_663 ();
 sg13g2_decap_4 FILLER_73_670 ();
 sg13g2_fill_2 FILLER_73_674 ();
 sg13g2_fill_1 FILLER_73_718 ();
 sg13g2_fill_2 FILLER_73_736 ();
 sg13g2_fill_2 FILLER_73_769 ();
 sg13g2_decap_8 FILLER_73_788 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_4 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_11 ();
 sg13g2_decap_8 FILLER_74_17 ();
 sg13g2_fill_2 FILLER_74_24 ();
 sg13g2_fill_1 FILLER_74_132 ();
 sg13g2_fill_2 FILLER_74_192 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_fill_2 FILLER_74_217 ();
 sg13g2_fill_2 FILLER_74_260 ();
 sg13g2_decap_4 FILLER_74_271 ();
 sg13g2_fill_1 FILLER_74_275 ();
 sg13g2_decap_8 FILLER_74_304 ();
 sg13g2_decap_8 FILLER_74_311 ();
 sg13g2_fill_2 FILLER_74_318 ();
 sg13g2_fill_1 FILLER_74_320 ();
 sg13g2_fill_2 FILLER_74_347 ();
 sg13g2_fill_1 FILLER_74_349 ();
 sg13g2_fill_2 FILLER_74_378 ();
 sg13g2_fill_2 FILLER_74_405 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_fill_2 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_fill_1 FILLER_74_456 ();
 sg13g2_fill_2 FILLER_74_483 ();
 sg13g2_fill_1 FILLER_74_485 ();
 sg13g2_fill_1 FILLER_74_529 ();
 sg13g2_decap_4 FILLER_74_557 ();
 sg13g2_fill_1 FILLER_74_596 ();
 sg13g2_fill_2 FILLER_74_608 ();
 sg13g2_fill_1 FILLER_74_610 ();
 sg13g2_decap_8 FILLER_74_656 ();
 sg13g2_decap_4 FILLER_74_663 ();
 sg13g2_fill_1 FILLER_74_667 ();
 sg13g2_fill_2 FILLER_74_677 ();
 sg13g2_fill_1 FILLER_74_679 ();
 sg13g2_fill_1 FILLER_74_702 ();
 sg13g2_fill_2 FILLER_74_721 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_55 ();
 sg13g2_decap_8 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_73 ();
 sg13g2_fill_2 FILLER_75_97 ();
 sg13g2_fill_2 FILLER_75_143 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_fill_1 FILLER_75_251 ();
 sg13g2_fill_1 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_381 ();
 sg13g2_fill_1 FILLER_75_383 ();
 sg13g2_fill_2 FILLER_75_412 ();
 sg13g2_fill_1 FILLER_75_414 ();
 sg13g2_decap_8 FILLER_75_423 ();
 sg13g2_fill_2 FILLER_75_430 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_457 ();
 sg13g2_fill_1 FILLER_75_459 ();
 sg13g2_fill_2 FILLER_75_474 ();
 sg13g2_fill_1 FILLER_75_476 ();
 sg13g2_fill_1 FILLER_75_531 ();
 sg13g2_fill_2 FILLER_75_537 ();
 sg13g2_fill_1 FILLER_75_539 ();
 sg13g2_fill_1 FILLER_75_572 ();
 sg13g2_fill_2 FILLER_75_741 ();
 sg13g2_fill_2 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_18 ();
 sg13g2_decap_8 FILLER_76_23 ();
 sg13g2_decap_4 FILLER_76_30 ();
 sg13g2_fill_1 FILLER_76_34 ();
 sg13g2_decap_8 FILLER_76_57 ();
 sg13g2_decap_8 FILLER_76_64 ();
 sg13g2_decap_8 FILLER_76_71 ();
 sg13g2_decap_4 FILLER_76_78 ();
 sg13g2_fill_2 FILLER_76_82 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_122 ();
 sg13g2_fill_2 FILLER_76_132 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_fill_2 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_255 ();
 sg13g2_decap_8 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_318 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_391 ();
 sg13g2_fill_1 FILLER_76_401 ();
 sg13g2_fill_2 FILLER_76_429 ();
 sg13g2_fill_1 FILLER_76_431 ();
 sg13g2_decap_4 FILLER_76_435 ();
 sg13g2_fill_1 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_467 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_fill_1 FILLER_76_515 ();
 sg13g2_fill_2 FILLER_76_544 ();
 sg13g2_decap_4 FILLER_76_550 ();
 sg13g2_fill_2 FILLER_76_554 ();
 sg13g2_fill_2 FILLER_76_565 ();
 sg13g2_fill_2 FILLER_76_612 ();
 sg13g2_fill_1 FILLER_76_614 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_662 ();
 sg13g2_fill_2 FILLER_76_669 ();
 sg13g2_fill_1 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_fill_2 FILLER_76_683 ();
 sg13g2_fill_1 FILLER_76_716 ();
 sg13g2_fill_1 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_47 ();
 sg13g2_decap_8 FILLER_77_54 ();
 sg13g2_decap_8 FILLER_77_61 ();
 sg13g2_decap_8 FILLER_77_68 ();
 sg13g2_decap_8 FILLER_77_75 ();
 sg13g2_decap_8 FILLER_77_82 ();
 sg13g2_fill_2 FILLER_77_89 ();
 sg13g2_fill_1 FILLER_77_121 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_fill_2 FILLER_77_295 ();
 sg13g2_fill_2 FILLER_77_344 ();
 sg13g2_fill_1 FILLER_77_346 ();
 sg13g2_fill_2 FILLER_77_412 ();
 sg13g2_fill_1 FILLER_77_435 ();
 sg13g2_fill_1 FILLER_77_469 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_fill_2 FILLER_77_501 ();
 sg13g2_fill_1 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_526 ();
 sg13g2_decap_4 FILLER_77_554 ();
 sg13g2_fill_1 FILLER_77_558 ();
 sg13g2_fill_2 FILLER_77_567 ();
 sg13g2_fill_2 FILLER_77_575 ();
 sg13g2_fill_1 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_656 ();
 sg13g2_decap_4 FILLER_77_663 ();
 sg13g2_fill_2 FILLER_77_704 ();
 sg13g2_fill_1 FILLER_77_724 ();
 sg13g2_fill_2 FILLER_77_739 ();
 sg13g2_fill_1 FILLER_77_741 ();
 sg13g2_fill_1 FILLER_77_756 ();
 sg13g2_fill_2 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_775 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_decap_4 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_163 ();
 sg13g2_decap_8 FILLER_78_206 ();
 sg13g2_decap_4 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_244 ();
 sg13g2_fill_2 FILLER_78_259 ();
 sg13g2_fill_1 FILLER_78_274 ();
 sg13g2_decap_4 FILLER_78_290 ();
 sg13g2_fill_1 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_394 ();
 sg13g2_fill_1 FILLER_78_396 ();
 sg13g2_fill_2 FILLER_78_410 ();
 sg13g2_fill_2 FILLER_78_572 ();
 sg13g2_fill_2 FILLER_78_593 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_8 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_fill_2 FILLER_78_678 ();
 sg13g2_fill_1 FILLER_78_680 ();
 sg13g2_fill_1 FILLER_78_734 ();
 sg13g2_fill_2 FILLER_78_744 ();
 sg13g2_fill_1 FILLER_78_746 ();
 sg13g2_fill_2 FILLER_78_756 ();
 sg13g2_fill_2 FILLER_78_777 ();
 sg13g2_fill_1 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_fill_2 FILLER_79_119 ();
 sg13g2_fill_2 FILLER_79_264 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_371 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_fill_2 FILLER_79_445 ();
 sg13g2_fill_2 FILLER_79_461 ();
 sg13g2_fill_1 FILLER_79_476 ();
 sg13g2_fill_2 FILLER_79_499 ();
 sg13g2_fill_1 FILLER_79_501 ();
 sg13g2_fill_1 FILLER_79_540 ();
 sg13g2_fill_2 FILLER_79_560 ();
 sg13g2_fill_1 FILLER_79_562 ();
 sg13g2_fill_2 FILLER_79_568 ();
 sg13g2_fill_1 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_4 FILLER_79_686 ();
 sg13g2_fill_2 FILLER_79_707 ();
 sg13g2_fill_1 FILLER_79_709 ();
 sg13g2_fill_2 FILLER_79_724 ();
 sg13g2_fill_1 FILLER_79_726 ();
 sg13g2_fill_2 FILLER_79_768 ();
 sg13g2_fill_1 FILLER_79_770 ();
 sg13g2_fill_2 FILLER_79_780 ();
 sg13g2_fill_1 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_4 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_170 ();
 sg13g2_decap_4 FILLER_80_183 ();
 sg13g2_fill_2 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_decap_4 FILLER_80_209 ();
 sg13g2_fill_1 FILLER_80_213 ();
 sg13g2_fill_2 FILLER_80_248 ();
 sg13g2_fill_2 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_fill_2 FILLER_80_492 ();
 sg13g2_fill_1 FILLER_80_494 ();
 sg13g2_fill_2 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_fill_2 FILLER_80_791 ();
 sg13g2_fill_1 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule
