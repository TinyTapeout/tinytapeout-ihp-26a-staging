module tt_um_phsauter_vga_maze (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire clknet_0_clk;
 wire \ent_x[0] ;
 wire \ent_x[1] ;
 wire \ent_y[0] ;
 wire \ent_y[1] ;
 wire \filled_width[1] ;
 wire \gamepad.decoder.data_reg[0] ;
 wire \gamepad.decoder.data_reg[10] ;
 wire \gamepad.decoder.data_reg[11] ;
 wire \gamepad.decoder.data_reg[1] ;
 wire \gamepad.decoder.data_reg[2] ;
 wire \gamepad.decoder.data_reg[3] ;
 wire \gamepad.decoder.data_reg[4] ;
 wire \gamepad.decoder.data_reg[5] ;
 wire \gamepad.decoder.data_reg[6] ;
 wire \gamepad.decoder.data_reg[7] ;
 wire \gamepad.decoder.data_reg[8] ;
 wire \gamepad.decoder.data_reg[9] ;
 wire \gamepad.driver.pmod_clk_prev ;
 wire \gamepad.driver.pmod_clk_sync[0] ;
 wire \gamepad.driver.pmod_clk_sync[1] ;
 wire \gamepad.driver.pmod_data_sync[0] ;
 wire \gamepad.driver.pmod_data_sync[1] ;
 wire \gamepad.driver.pmod_latch_prev ;
 wire \gamepad.driver.pmod_latch_sync[0] ;
 wire \gamepad.driver.pmod_latch_sync[1] ;
 wire \gamepad.driver.shift_reg[0] ;
 wire \gamepad.driver.shift_reg[10] ;
 wire \gamepad.driver.shift_reg[11] ;
 wire \gamepad.driver.shift_reg[1] ;
 wire \gamepad.driver.shift_reg[2] ;
 wire \gamepad.driver.shift_reg[3] ;
 wire \gamepad.driver.shift_reg[4] ;
 wire \gamepad.driver.shift_reg[5] ;
 wire \gamepad.driver.shift_reg[6] ;
 wire \gamepad.driver.shift_reg[7] ;
 wire \gamepad.driver.shift_reg[8] ;
 wire \gamepad.driver.shift_reg[9] ;
 wire \gen_frame_count[0] ;
 wire \gen_frame_count[1] ;
 wire \gen_frame_count[2] ;
 wire \gen_frame_count[3] ;
 wire \gen_row[0] ;
 wire \gen_row[1] ;
 wire \gen_row[2] ;
 wire generating;
 wire hsync;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire inp_a_prev;
 wire inp_b_prev;
 wire inp_down_prev;
 wire inp_l_prev;
 wire inp_left_prev;
 wire inp_r_prev;
 wire inp_right_prev;
 wire inp_select_prev;
 wire inp_start_prev;
 wire inp_up_prev;
 wire inp_x_prev;
 wire inp_y_prev;
 wire \lfsr[0] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[5] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \maze_seed[0] ;
 wire \maze_seed[1] ;
 wire \maze_seed[2] ;
 wire \maze_seed[3] ;
 wire \maze_seed[4] ;
 wire player_won;
 wire \player_x[0] ;
 wire \player_x[1] ;
 wire \player_x[2] ;
 wire \player_y[0] ;
 wire \player_y[1] ;
 wire \player_y[2] ;
 wire single_step_mode;
 wire \solver_frame_count[0] ;
 wire \solver_frame_count[1] ;
 wire \solver_frame_count[2] ;
 wire \solver_frame_count[3] ;
 wire \solver_l_dir[0] ;
 wire \solver_l_dir[1] ;
 wire \solver_l_dir[2] ;
 wire \solver_l_dir[3] ;
 wire solver_l_won;
 wire \solver_l_x[0] ;
 wire \solver_l_x[1] ;
 wire \solver_l_x[2] ;
 wire \solver_l_y[0] ;
 wire \solver_l_y[1] ;
 wire \solver_l_y[2] ;
 wire \solver_r_dir[0] ;
 wire \solver_r_dir[1] ;
 wire \solver_r_dir[2] ;
 wire \solver_r_dir[3] ;
 wire solver_r_won;
 wire \solver_r_x[0] ;
 wire \solver_r_x[1] ;
 wire \solver_r_x[2] ;
 wire \solver_r_y[0] ;
 wire \solver_r_y[1] ;
 wire \solver_r_y[2] ;
 wire \solver_speed[1] ;
 wire \solver_speed[2] ;
 wire \solver_speed[3] ;
 wire solvers_active;
 wire step_requested;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire vsync_prev;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;

 sg13g2_inv_1 _1105_ (.Y(_0297_),
    .A(net238));
 sg13g2_inv_1 _1106_ (.Y(_0298_),
    .A(net242));
 sg13g2_inv_1 _1107_ (.Y(_0299_),
    .A(net271));
 sg13g2_inv_1 _1108_ (.Y(_0300_),
    .A(net248));
 sg13g2_inv_1 _1109_ (.Y(_0301_),
    .A(net266));
 sg13g2_inv_1 _1110_ (.Y(_0302_),
    .A(net269));
 sg13g2_inv_1 _1111_ (.Y(_0303_),
    .A(net264));
 sg13g2_inv_1 _1112_ (.Y(_0304_),
    .A(net262));
 sg13g2_inv_1 _1113_ (.Y(_0305_),
    .A(net268));
 sg13g2_inv_1 _1114_ (.Y(_0306_),
    .A(net250));
 sg13g2_inv_1 _1115_ (.Y(_0307_),
    .A(net258));
 sg13g2_inv_1 _1116_ (.Y(_0308_),
    .A(net265));
 sg13g2_inv_1 _1117_ (.Y(_0309_),
    .A(\solver_speed[3] ));
 sg13g2_inv_1 _1118_ (.Y(_0310_),
    .A(net348));
 sg13g2_inv_1 _1119_ (.Y(_0311_),
    .A(net224));
 sg13g2_inv_2 _1120_ (.Y(_0312_),
    .A(generating));
 sg13g2_inv_1 _1121_ (.Y(_0313_),
    .A(solvers_active));
 sg13g2_inv_2 _1122_ (.Y(_0314_),
    .A(net184));
 sg13g2_inv_1 _1123_ (.Y(_0315_),
    .A(net255));
 sg13g2_inv_1 _1124_ (.Y(_0316_),
    .A(\maze_seed[2] ));
 sg13g2_inv_1 _1125_ (.Y(_0317_),
    .A(net240));
 sg13g2_inv_2 _1126_ (.Y(_0318_),
    .A(\maze_seed[0] ));
 sg13g2_inv_1 _1127_ (.Y(_0319_),
    .A(net288));
 sg13g2_inv_1 _1128_ (.Y(_0320_),
    .A(net228));
 sg13g2_inv_1 _1129_ (.Y(_0321_),
    .A(net292));
 sg13g2_inv_1 _1130_ (.Y(_0322_),
    .A(net200));
 sg13g2_inv_1 _1131_ (.Y(_0323_),
    .A(solver_l_won));
 sg13g2_inv_2 _1132_ (.Y(_0324_),
    .A(player_won));
 sg13g2_inv_2 _1133_ (.Y(_0325_),
    .A(solver_r_won));
 sg13g2_inv_4 _1134_ (.A(\solver_l_x[0] ),
    .Y(_0326_));
 sg13g2_inv_1 _1135_ (.Y(_0327_),
    .A(net186));
 sg13g2_inv_1 _1136_ (.Y(_0328_),
    .A(net187));
 sg13g2_inv_1 _1137_ (.Y(_0329_),
    .A(net189));
 sg13g2_inv_1 _1138_ (.Y(_0330_),
    .A(net185));
 sg13g2_inv_1 _1139_ (.Y(_0331_),
    .A(\solver_r_y[2] ));
 sg13g2_inv_2 _1140_ (.Y(_0332_),
    .A(net172));
 sg13g2_inv_1 _1141_ (.Y(_0333_),
    .A(net338));
 sg13g2_inv_2 _1142_ (.Y(_0334_),
    .A(net359));
 sg13g2_inv_2 _1143_ (.Y(_0335_),
    .A(net326));
 sg13g2_inv_2 _1144_ (.Y(_0336_),
    .A(net295));
 sg13g2_inv_2 _1145_ (.Y(_0337_),
    .A(net290));
 sg13g2_inv_1 _1146_ (.Y(_0338_),
    .A(net300));
 sg13g2_inv_1 _1147_ (.Y(_0339_),
    .A(net339));
 sg13g2_inv_2 _1148_ (.Y(_0340_),
    .A(\hvsync_gen.hpos[4] ));
 sg13g2_inv_1 _1149_ (.Y(_0341_),
    .A(net174));
 sg13g2_inv_2 _1150_ (.Y(_0342_),
    .A(net180));
 sg13g2_inv_1 _1151_ (.Y(_0343_),
    .A(net179));
 sg13g2_inv_2 _1152_ (.Y(_0344_),
    .A(\player_x[0] ));
 sg13g2_nor2b_2 _1153_ (.A(net281),
    .B_N(net247),
    .Y(_0345_));
 sg13g2_nand2b_2 _1154_ (.Y(_0346_),
    .B(net247),
    .A_N(net281));
 sg13g2_or3_1 _1155_ (.A(net282),
    .B(net302),
    .C(net163),
    .X(_0347_));
 sg13g2_nor3_2 _1156_ (.A(net304),
    .B(\solver_frame_count[2] ),
    .C(_0347_),
    .Y(_0348_));
 sg13g2_nor2b_1 _1157_ (.A(step_requested),
    .B_N(single_step_mode),
    .Y(_0349_));
 sg13g2_nand2_1 _1158_ (.Y(_0350_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_nand4_1 _1159_ (.B(_0323_),
    .C(_0324_),
    .A(_0312_),
    .Y(_0351_),
    .D(_0325_));
 sg13g2_nor2_1 _1160_ (.A(_0313_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor3_1 _1161_ (.A(_0313_),
    .B(_0349_),
    .C(_0351_),
    .Y(_0353_));
 sg13g2_o21ai_1 _1162_ (.B1(_0353_),
    .Y(_0354_),
    .A1(single_step_mode),
    .A2(_0348_));
 sg13g2_nand3_1 _1163_ (.B(\gamepad.decoder.data_reg[1] ),
    .C(\gamepad.decoder.data_reg[0] ),
    .A(\gamepad.decoder.data_reg[2] ),
    .Y(_0355_));
 sg13g2_nand4_1 _1164_ (.B(\gamepad.decoder.data_reg[5] ),
    .C(\gamepad.decoder.data_reg[4] ),
    .A(\gamepad.decoder.data_reg[6] ),
    .Y(_0356_),
    .D(\gamepad.decoder.data_reg[3] ));
 sg13g2_nand4_1 _1165_ (.B(\gamepad.decoder.data_reg[9] ),
    .C(\gamepad.decoder.data_reg[8] ),
    .A(\gamepad.decoder.data_reg[11] ),
    .Y(_0357_),
    .D(\gamepad.decoder.data_reg[7] ));
 sg13g2_nor3_1 _1166_ (.A(_0355_),
    .B(_0356_),
    .C(_0357_),
    .Y(_0358_));
 sg13g2_nand2_1 _1167_ (.Y(_0359_),
    .A(net237),
    .B(_0358_));
 sg13g2_nand2_1 _1168_ (.Y(_0360_),
    .A(net272),
    .B(net156));
 sg13g2_nor3_2 _1169_ (.A(generating),
    .B(inp_b_prev),
    .C(_0360_),
    .Y(_0361_));
 sg13g2_inv_1 _1170_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_nand2_1 _1171_ (.Y(_0363_),
    .A(net270),
    .B(net156));
 sg13g2_nor2_2 _1172_ (.A(inp_select_prev),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_or2_1 _1173_ (.X(_0365_),
    .B(_0363_),
    .A(inp_select_prev));
 sg13g2_nor2_2 _1174_ (.A(net193),
    .B(_0364_),
    .Y(_0366_));
 sg13g2_nand2_2 _1175_ (.Y(_0367_),
    .A(net202),
    .B(_0365_));
 sg13g2_nor2_1 _1176_ (.A(_0361_),
    .B(_0364_),
    .Y(_0368_));
 sg13g2_nor2_2 _1177_ (.A(_0361_),
    .B(_0367_),
    .Y(_0369_));
 sg13g2_and2_1 _1178_ (.A(net153),
    .B(_0369_),
    .X(_0370_));
 sg13g2_nor2_2 _1179_ (.A(net197),
    .B(net153),
    .Y(_0371_));
 sg13g2_nor3_2 _1180_ (.A(\solver_l_y[2] ),
    .B(net170),
    .C(\solver_l_y[1] ),
    .Y(_0372_));
 sg13g2_o21ai_1 _1181_ (.B1(_0372_),
    .Y(_0373_),
    .A1(\solver_l_x[2] ),
    .A2(\solver_l_x[1] ));
 sg13g2_nand2_2 _1182_ (.Y(_0374_),
    .A(_0326_),
    .B(_0373_));
 sg13g2_and2_1 _1183_ (.A(net188),
    .B(_0374_),
    .X(_0375_));
 sg13g2_nand2_1 _1184_ (.Y(_0376_),
    .A(net188),
    .B(_0374_));
 sg13g2_a22oi_1 _1185_ (.Y(_0377_),
    .B1(net151),
    .B2(_0375_),
    .A2(_0370_),
    .A1(net186));
 sg13g2_and2_1 _1186_ (.A(net170),
    .B(\solver_l_y[1] ),
    .X(_0378_));
 sg13g2_nand2_1 _1187_ (.Y(_0379_),
    .A(\solver_l_y[2] ),
    .B(_0378_));
 sg13g2_xnor2_1 _1188_ (.Y(_0380_),
    .A(\solver_l_y[1] ),
    .B(\solver_l_x[2] ));
 sg13g2_xnor2_1 _1189_ (.Y(_0381_),
    .A(\maze_seed[1] ),
    .B(_0380_));
 sg13g2_xor2_1 _1190_ (.B(_0381_),
    .A(net170),
    .X(_0382_));
 sg13g2_xnor2_1 _1191_ (.Y(_0383_),
    .A(\maze_seed[2] ),
    .B(\solver_l_y[2] ));
 sg13g2_xor2_1 _1192_ (.B(_0383_),
    .A(_0378_),
    .X(_0384_));
 sg13g2_a21oi_1 _1193_ (.A1(net182),
    .A2(_0382_),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_xor2_1 _1194_ (.B(\solver_l_x[1] ),
    .A(\maze_seed[0] ),
    .X(_0386_));
 sg13g2_xnor2_1 _1195_ (.Y(_0387_),
    .A(net170),
    .B(_0386_));
 sg13g2_or2_1 _1196_ (.X(_0388_),
    .B(_0387_),
    .A(net182));
 sg13g2_nand4_1 _1197_ (.B(_0382_),
    .C(_0384_),
    .A(net182),
    .Y(_0389_),
    .D(_0387_));
 sg13g2_o21ai_1 _1198_ (.B1(_0389_),
    .Y(_0390_),
    .A1(_0382_),
    .A2(_0388_));
 sg13g2_nor2_1 _1199_ (.A(_0385_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_xnor2_1 _1200_ (.Y(_0392_),
    .A(\maze_seed[4] ),
    .B(\solver_l_x[0] ));
 sg13g2_xnor2_1 _1201_ (.Y(_0393_),
    .A(_0381_),
    .B(_0392_));
 sg13g2_xnor2_1 _1202_ (.Y(_0394_),
    .A(_0387_),
    .B(_0393_));
 sg13g2_xnor2_1 _1203_ (.Y(_0395_),
    .A(_0391_),
    .B(_0394_));
 sg13g2_and2_1 _1204_ (.A(_0379_),
    .B(_0395_),
    .X(_0396_));
 sg13g2_nand2_2 _1205_ (.Y(_0397_),
    .A(_0379_),
    .B(_0395_));
 sg13g2_nor2_1 _1206_ (.A(net154),
    .B(_0361_),
    .Y(_0398_));
 sg13g2_nand4_1 _1207_ (.B(_0374_),
    .C(net143),
    .A(net399),
    .Y(_0399_),
    .D(_0398_));
 sg13g2_o21ai_1 _1208_ (.B1(_0377_),
    .Y(_0400_),
    .A1(_0367_),
    .A2(_0399_));
 sg13g2_o21ai_1 _1209_ (.B1(_0388_),
    .Y(_0401_),
    .A1(_0314_),
    .A2(_0381_));
 sg13g2_nand2_1 _1210_ (.Y(_0402_),
    .A(_0381_),
    .B(_0388_));
 sg13g2_a21oi_1 _1211_ (.A1(net182),
    .A2(_0387_),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_mux2_1 _1212_ (.A0(_0401_),
    .A1(_0403_),
    .S(_0383_),
    .X(_0404_));
 sg13g2_nor2_1 _1213_ (.A(net183),
    .B(net170),
    .Y(_0405_));
 sg13g2_a21oi_1 _1214_ (.A1(net183),
    .A2(_0386_),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_xnor2_1 _1215_ (.Y(_0407_),
    .A(_0393_),
    .B(_0406_));
 sg13g2_xnor2_1 _1216_ (.Y(_0408_),
    .A(_0404_),
    .B(_0407_));
 sg13g2_nor2_2 _1217_ (.A(_0372_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_or2_1 _1218_ (.X(_0410_),
    .B(_0408_),
    .A(_0372_));
 sg13g2_a21oi_1 _1219_ (.A1(net189),
    .A2(_0410_),
    .Y(_0411_),
    .B1(net187));
 sg13g2_inv_1 _1220_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_nand2_1 _1221_ (.Y(_0413_),
    .A(net151),
    .B(net143));
 sg13g2_and2_1 _1222_ (.A(\solver_l_x[0] ),
    .B(\solver_l_x[1] ),
    .X(_0414_));
 sg13g2_nor2_1 _1223_ (.A(_0326_),
    .B(_0372_),
    .Y(_0415_));
 sg13g2_a21oi_2 _1224_ (.B1(_0415_),
    .Y(_0416_),
    .A2(_0414_),
    .A1(\solver_l_x[2] ));
 sg13g2_nand2b_2 _1225_ (.Y(_0417_),
    .B(net187),
    .A_N(_0416_));
 sg13g2_nor3_1 _1226_ (.A(_0329_),
    .B(_0409_),
    .C(_0416_),
    .Y(_0418_));
 sg13g2_nor3_1 _1227_ (.A(_0411_),
    .B(_0413_),
    .C(_0416_),
    .Y(_0419_));
 sg13g2_nand2_1 _1228_ (.Y(_0420_),
    .A(_0374_),
    .B(net143));
 sg13g2_or2_1 _1229_ (.X(_0003_),
    .B(_0419_),
    .A(_0400_));
 sg13g2_nor3_1 _1230_ (.A(_0327_),
    .B(_0374_),
    .C(_0396_),
    .Y(_0421_));
 sg13g2_nand2_1 _1231_ (.Y(_0422_),
    .A(net394),
    .B(_0416_));
 sg13g2_nand2_1 _1232_ (.Y(_0423_),
    .A(net151),
    .B(_0422_));
 sg13g2_a21oi_1 _1233_ (.A1(_0410_),
    .A2(_0421_),
    .Y(_0424_),
    .B1(_0423_));
 sg13g2_nand2_2 _1234_ (.Y(_0425_),
    .A(_0410_),
    .B(_0416_));
 sg13g2_nand2b_1 _1235_ (.Y(_0426_),
    .B(_0425_),
    .A_N(net153));
 sg13g2_nand3_1 _1236_ (.B(\solver_l_dir[0] ),
    .C(_0426_),
    .A(net204),
    .Y(_0427_));
 sg13g2_o21ai_1 _1237_ (.B1(_0425_),
    .Y(_0428_),
    .A1(_0362_),
    .A2(_0410_));
 sg13g2_and3_2 _1238_ (.X(_0429_),
    .A(_0326_),
    .B(net188),
    .C(_0373_));
 sg13g2_nand3_1 _1239_ (.B(_0428_),
    .C(_0429_),
    .A(net151),
    .Y(_0430_));
 sg13g2_nand2_1 _1240_ (.Y(_0431_),
    .A(_0427_),
    .B(_0430_));
 sg13g2_nor2_1 _1241_ (.A(net191),
    .B(_0363_),
    .Y(_0080_));
 sg13g2_nor2_2 _1242_ (.A(net193),
    .B(_0365_),
    .Y(_0432_));
 sg13g2_nand3_1 _1243_ (.B(_0409_),
    .C(_0429_),
    .A(_0398_),
    .Y(_0433_));
 sg13g2_nor4_1 _1244_ (.A(net153),
    .B(_0361_),
    .C(net143),
    .D(_0417_),
    .Y(_0434_));
 sg13g2_or4_1 _1245_ (.A(net154),
    .B(_0361_),
    .C(net143),
    .D(_0417_),
    .X(_0435_));
 sg13g2_nand3_1 _1246_ (.B(_0433_),
    .C(_0435_),
    .A(_0399_),
    .Y(_0436_));
 sg13g2_nand2_1 _1247_ (.Y(_0437_),
    .A(_0371_),
    .B(_0396_));
 sg13g2_nand4_1 _1248_ (.B(_0371_),
    .C(_0374_),
    .A(\solver_l_dir[3] ),
    .Y(_0438_),
    .D(_0397_));
 sg13g2_o21ai_1 _1249_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0417_),
    .A2(_0437_));
 sg13g2_a221oi_1 _1250_ (.B2(_0361_),
    .C1(_0431_),
    .B1(_0439_),
    .A1(_0432_),
    .Y(_0440_),
    .A2(_0436_));
 sg13g2_o21ai_1 _1251_ (.B1(_0440_),
    .Y(_0000_),
    .A1(_0370_),
    .A2(_0424_));
 sg13g2_and2_1 _1252_ (.A(\solver_r_x[1] ),
    .B(net172),
    .X(_0441_));
 sg13g2_nand2_1 _1253_ (.Y(_0442_),
    .A(\solver_r_x[2] ),
    .B(_0441_));
 sg13g2_nor3_2 _1254_ (.A(net171),
    .B(\solver_r_y[1] ),
    .C(\solver_r_y[2] ),
    .Y(_0443_));
 sg13g2_nor2_1 _1255_ (.A(_0332_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_2 _1256_ (.B1(_0444_),
    .Y(_0445_),
    .A2(_0441_),
    .A1(\solver_r_x[2] ));
 sg13g2_inv_1 _1257_ (.Y(_0446_),
    .A(_0445_));
 sg13g2_xnor2_1 _1258_ (.Y(_0447_),
    .A(\solver_r_x[1] ),
    .B(net171));
 sg13g2_xnor2_1 _1259_ (.Y(_0448_),
    .A(\maze_seed[0] ),
    .B(_0447_));
 sg13g2_nor2_1 _1260_ (.A(_0314_),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_nand2_1 _1261_ (.Y(_0450_),
    .A(net183),
    .B(_0448_));
 sg13g2_xnor2_1 _1262_ (.Y(_0451_),
    .A(net183),
    .B(_0448_));
 sg13g2_xnor2_1 _1263_ (.Y(_0452_),
    .A(\maze_seed[1] ),
    .B(\solver_r_x[2] ));
 sg13g2_xnor2_1 _1264_ (.Y(_0453_),
    .A(\solver_r_y[1] ),
    .B(_0452_));
 sg13g2_xnor2_1 _1265_ (.Y(_0454_),
    .A(\maze_seed[2] ),
    .B(\solver_r_y[2] ));
 sg13g2_nor2_1 _1266_ (.A(_0448_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_nor2_1 _1267_ (.A(_0451_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nor2_1 _1268_ (.A(net183),
    .B(_0453_),
    .Y(_0457_));
 sg13g2_a22oi_1 _1269_ (.Y(_0458_),
    .B1(_0457_),
    .B2(_0455_),
    .A2(_0456_),
    .A1(_0453_));
 sg13g2_xnor2_1 _1270_ (.Y(_0459_),
    .A(\maze_seed[4] ),
    .B(net171));
 sg13g2_xnor2_1 _1271_ (.Y(_0460_),
    .A(net172),
    .B(_0459_));
 sg13g2_xnor2_1 _1272_ (.Y(_0461_),
    .A(_0454_),
    .B(_0460_));
 sg13g2_xnor2_1 _1273_ (.Y(_0462_),
    .A(_0449_),
    .B(_0461_));
 sg13g2_xor2_1 _1274_ (.B(_0462_),
    .A(_0458_),
    .X(_0463_));
 sg13g2_nor2_2 _1275_ (.A(_0443_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_nor3_2 _1276_ (.A(_0332_),
    .B(_0443_),
    .C(_0463_),
    .Y(_0465_));
 sg13g2_nor2_1 _1277_ (.A(net153),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_nand2_1 _1278_ (.Y(_0467_),
    .A(net279),
    .B(_0369_));
 sg13g2_nand2_1 _1279_ (.Y(_0468_),
    .A(net171),
    .B(\solver_r_y[1] ));
 sg13g2_nand3_1 _1280_ (.B(\solver_r_y[1] ),
    .C(\solver_r_y[2] ),
    .A(net171),
    .Y(_0469_));
 sg13g2_xor2_1 _1281_ (.B(\solver_r_y[1] ),
    .A(net171),
    .X(_0470_));
 sg13g2_xor2_1 _1282_ (.B(_0470_),
    .A(_0452_),
    .X(_0471_));
 sg13g2_xor2_1 _1283_ (.B(_0468_),
    .A(_0454_),
    .X(_0472_));
 sg13g2_nor2_1 _1284_ (.A(_0451_),
    .B(_0471_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1285_ (.A1(_0448_),
    .A2(_0472_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_a21oi_1 _1286_ (.A1(net183),
    .A2(_0471_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_xnor2_1 _1287_ (.Y(_0476_),
    .A(net172),
    .B(_0475_));
 sg13g2_xnor2_1 _1288_ (.Y(_0477_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_xnor2_1 _1289_ (.Y(_0478_),
    .A(_0450_),
    .B(_0459_));
 sg13g2_xnor2_1 _1290_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_xnor2_1 _1291_ (.Y(_0480_),
    .A(_0476_),
    .B(_0479_));
 sg13g2_nand2_2 _1292_ (.Y(_0481_),
    .A(_0469_),
    .B(_0480_));
 sg13g2_nand3_1 _1293_ (.B(_0446_),
    .C(_0481_),
    .A(\solver_r_dir[0] ),
    .Y(_0482_));
 sg13g2_nand2_1 _1294_ (.Y(_0483_),
    .A(_0334_),
    .B(_0482_));
 sg13g2_nand3_1 _1295_ (.B(_0464_),
    .C(_0483_),
    .A(net151),
    .Y(_0484_));
 sg13g2_o21ai_1 _1296_ (.B1(_0484_),
    .Y(_0005_),
    .A1(_0466_),
    .A2(_0467_));
 sg13g2_or2_1 _1297_ (.X(_0485_),
    .B(_0421_),
    .A(net189));
 sg13g2_nand3_1 _1298_ (.B(_0409_),
    .C(_0485_),
    .A(_0371_),
    .Y(_0486_));
 sg13g2_nand2_1 _1299_ (.Y(_0487_),
    .A(net313),
    .B(_0370_));
 sg13g2_or2_1 _1300_ (.X(_0488_),
    .B(_0433_),
    .A(_0367_));
 sg13g2_nand3_1 _1301_ (.B(_0487_),
    .C(_0488_),
    .A(_0486_),
    .Y(_0001_));
 sg13g2_nor2_1 _1302_ (.A(\solver_r_x[1] ),
    .B(\solver_r_x[2] ),
    .Y(_0489_));
 sg13g2_nor2b_1 _1303_ (.A(_0489_),
    .B_N(_0443_),
    .Y(_0490_));
 sg13g2_nor2_2 _1304_ (.A(net172),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_inv_1 _1305_ (.Y(_0492_),
    .A(_0491_));
 sg13g2_nor2_2 _1306_ (.A(_0334_),
    .B(_0464_),
    .Y(_0493_));
 sg13g2_nand2_1 _1307_ (.Y(_0494_),
    .A(\solver_r_dir[3] ),
    .B(_0491_));
 sg13g2_nand2_1 _1308_ (.Y(_0495_),
    .A(_0491_),
    .B(_0493_));
 sg13g2_and2_1 _1309_ (.A(\solver_r_dir[2] ),
    .B(_0491_),
    .X(_0496_));
 sg13g2_a221oi_1 _1310_ (.B2(net146),
    .C1(\solver_r_dir[0] ),
    .B1(_0496_),
    .A1(_0491_),
    .Y(_0497_),
    .A2(_0493_));
 sg13g2_nor4_1 _1311_ (.A(net197),
    .B(net153),
    .C(_0481_),
    .D(_0497_),
    .Y(_0498_));
 sg13g2_a21o_1 _1312_ (.A2(_0370_),
    .A1(net320),
    .B1(_0498_),
    .X(_0006_));
 sg13g2_nor2_1 _1313_ (.A(net186),
    .B(_0418_),
    .Y(_0499_));
 sg13g2_a22oi_1 _1314_ (.Y(_0500_),
    .B1(_0434_),
    .B2(_0366_),
    .A2(_0370_),
    .A1(net187));
 sg13g2_o21ai_1 _1315_ (.B1(_0500_),
    .Y(_0002_),
    .A1(_0437_),
    .A2(_0499_));
 sg13g2_nand3_1 _1316_ (.B(_0480_),
    .C(_0496_),
    .A(_0469_),
    .Y(_0501_));
 sg13g2_a22oi_1 _1317_ (.Y(_0502_),
    .B1(_0492_),
    .B2(_0493_),
    .A2(_0465_),
    .A1(net185));
 sg13g2_a21oi_1 _1318_ (.A1(_0501_),
    .A2(_0502_),
    .Y(_0503_),
    .B1(net146));
 sg13g2_nor2_2 _1319_ (.A(net338),
    .B(_0496_),
    .Y(_0504_));
 sg13g2_o21ai_1 _1320_ (.B1(_0495_),
    .Y(_0505_),
    .A1(_0446_),
    .A2(_0504_));
 sg13g2_a221oi_1 _1321_ (.B2(_0505_),
    .C1(_0503_),
    .B1(_0481_),
    .A1(net185),
    .Y(_0506_),
    .A2(_0445_));
 sg13g2_a22oi_1 _1322_ (.Y(_0004_),
    .B1(net151),
    .B2(_0506_),
    .A2(_0370_),
    .A1(_0333_));
 sg13g2_nand2_2 _1323_ (.Y(_0507_),
    .A(net320),
    .B(_0492_));
 sg13g2_a21oi_1 _1324_ (.A1(net338),
    .A2(_0481_),
    .Y(_0508_),
    .B1(net185));
 sg13g2_or2_1 _1325_ (.X(_0509_),
    .B(_0508_),
    .A(_0445_));
 sg13g2_o21ai_1 _1326_ (.B1(_0507_),
    .Y(_0510_),
    .A1(_0464_),
    .A2(_0509_));
 sg13g2_nand2_1 _1327_ (.Y(_0511_),
    .A(net151),
    .B(_0510_));
 sg13g2_nor2_2 _1328_ (.A(_0464_),
    .B(_0491_),
    .Y(_0512_));
 sg13g2_o21ai_1 _1329_ (.B1(_0369_),
    .Y(_0513_),
    .A1(net153),
    .A2(_0512_));
 sg13g2_o21ai_1 _1330_ (.B1(_0511_),
    .Y(_0007_),
    .A1(_0334_),
    .A2(_0513_));
 sg13g2_nand4_1 _1331_ (.B(_0337_),
    .C(net167),
    .A(net295),
    .Y(_0514_),
    .D(\hvsync_gen.vpos[6] ));
 sg13g2_nand2_1 _1332_ (.Y(_0515_),
    .A(net300),
    .B(_0339_));
 sg13g2_nand2_1 _1333_ (.Y(_0516_),
    .A(net300),
    .B(net166));
 sg13g2_nand2_1 _1334_ (.Y(_0517_),
    .A(net168),
    .B(_0335_));
 sg13g2_nor4_1 _1335_ (.A(_0514_),
    .B(_0515_),
    .C(_0516_),
    .D(_0517_),
    .Y(_0009_));
 sg13g2_and3_1 _1336_ (.X(_0518_),
    .A(net175),
    .B(net176),
    .C(net178));
 sg13g2_nor3_1 _1337_ (.A(net175),
    .B(net176),
    .C(net178),
    .Y(_0519_));
 sg13g2_nand2_1 _1338_ (.Y(_0520_),
    .A(net276),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_nor4_1 _1339_ (.A(net174),
    .B(_0518_),
    .C(_0519_),
    .D(net277),
    .Y(_0008_));
 sg13g2_o21ai_1 _1340_ (.B1(\hvsync_gen.vpos[8] ),
    .Y(_0521_),
    .A1(net166),
    .A2(\hvsync_gen.vpos[6] ));
 sg13g2_nor2_1 _1341_ (.A(\hvsync_gen.vpos[9] ),
    .B(\hvsync_gen.hpos[9] ),
    .Y(_0522_));
 sg13g2_nand2_1 _1342_ (.Y(_0523_),
    .A(\hvsync_gen.hpos[6] ),
    .B(net174));
 sg13g2_o21ai_1 _1343_ (.B1(net174),
    .Y(_0524_),
    .A1(\hvsync_gen.hpos[7] ),
    .A2(\hvsync_gen.hpos[6] ));
 sg13g2_nand3_1 _1344_ (.B(_0522_),
    .C(_0524_),
    .A(_0521_),
    .Y(_0525_));
 sg13g2_nand2b_1 _1345_ (.Y(_0526_),
    .B(net166),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_nor2b_2 _1346_ (.A(\hvsync_gen.vpos[6] ),
    .B_N(\hvsync_gen.vpos[8] ),
    .Y(_0527_));
 sg13g2_nor2b_2 _1347_ (.A(net166),
    .B_N(\hvsync_gen.vpos[9] ),
    .Y(_0528_));
 sg13g2_nor2b_1 _1348_ (.A(\hvsync_gen.vpos[8] ),
    .B_N(\hvsync_gen.vpos[6] ),
    .Y(_0529_));
 sg13g2_nand2b_1 _1349_ (.Y(_0530_),
    .B(_0528_),
    .A_N(_0529_));
 sg13g2_o21ai_1 _1350_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0526_),
    .A2(_0527_));
 sg13g2_or3_1 _1351_ (.A(_0527_),
    .B(_0528_),
    .C(_0529_),
    .X(_0532_));
 sg13g2_a22oi_1 _1352_ (.Y(_0533_),
    .B1(_0528_),
    .B2(_0529_),
    .A2(_0527_),
    .A1(_0526_));
 sg13g2_and2_1 _1353_ (.A(_0532_),
    .B(_0533_),
    .X(_0534_));
 sg13g2_a21o_2 _1354_ (.A2(_0533_),
    .A1(_0532_),
    .B1(net167),
    .X(_0535_));
 sg13g2_nand2_1 _1355_ (.Y(_0536_),
    .A(_0531_),
    .B(_0535_));
 sg13g2_a21o_1 _1356_ (.A2(_0527_),
    .A1(_0526_),
    .B1(_0528_),
    .X(_0537_));
 sg13g2_and2_1 _1357_ (.A(_0530_),
    .B(_0537_),
    .X(_0538_));
 sg13g2_a21oi_2 _1358_ (.B1(_0538_),
    .Y(_0539_),
    .A2(_0535_),
    .A1(_0531_));
 sg13g2_xor2_1 _1359_ (.B(net152),
    .A(net167),
    .X(_0540_));
 sg13g2_xnor2_1 _1360_ (.Y(_0541_),
    .A(net167),
    .B(_0539_));
 sg13g2_a21o_1 _1361_ (.A2(_0537_),
    .A1(_0535_),
    .B1(_0531_),
    .X(_0542_));
 sg13g2_and2_1 _1362_ (.A(_0536_),
    .B(_0542_),
    .X(_0543_));
 sg13g2_nand2_1 _1363_ (.Y(_0544_),
    .A(_0536_),
    .B(_0542_));
 sg13g2_o21ai_1 _1364_ (.B1(_0534_),
    .Y(_0545_),
    .A1(net167),
    .A2(net152));
 sg13g2_nand2b_1 _1365_ (.Y(_0546_),
    .B(_0538_),
    .A_N(_0535_));
 sg13g2_a22oi_1 _1366_ (.Y(_0547_),
    .B1(_0545_),
    .B2(_0546_),
    .A2(_0540_),
    .A1(_0337_));
 sg13g2_nor2_2 _1367_ (.A(_0543_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_o21ai_1 _1368_ (.B1(_0337_),
    .Y(_0549_),
    .A1(_0543_),
    .A2(_0547_));
 sg13g2_nor3_1 _1369_ (.A(\hvsync_gen.vpos[4] ),
    .B(_0541_),
    .C(_0544_),
    .Y(_0550_));
 sg13g2_and3_1 _1370_ (.X(_0551_),
    .A(_0544_),
    .B(_0545_),
    .C(_0546_));
 sg13g2_nor3_1 _1371_ (.A(_0547_),
    .B(_0550_),
    .C(_0551_),
    .Y(_0552_));
 sg13g2_nand4_1 _1372_ (.B(_0544_),
    .C(_0545_),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_0553_),
    .D(_0546_));
 sg13g2_nand2_1 _1373_ (.Y(_0554_),
    .A(_0549_),
    .B(_0553_));
 sg13g2_nand3_1 _1374_ (.B(_0549_),
    .C(_0553_),
    .A(_0336_),
    .Y(_0555_));
 sg13g2_xnor2_1 _1375_ (.Y(_0556_),
    .A(_0541_),
    .B(_0549_));
 sg13g2_a21oi_1 _1376_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0557_),
    .B1(_0552_));
 sg13g2_or2_1 _1377_ (.X(_0558_),
    .B(net140),
    .A(\gen_row[0] ));
 sg13g2_nand2_1 _1378_ (.Y(_0559_),
    .A(\gen_row[2] ),
    .B(net152));
 sg13g2_or2_1 _1379_ (.X(_0560_),
    .B(net152),
    .A(\gen_row[2] ));
 sg13g2_o21ai_1 _1380_ (.B1(_0560_),
    .Y(_0561_),
    .A1(\gen_row[1] ),
    .A2(net144));
 sg13g2_xnor2_1 _1381_ (.Y(_0562_),
    .A(\gen_row[1] ),
    .B(net144));
 sg13g2_a21oi_1 _1382_ (.A1(\gen_row[0] ),
    .A2(net140),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_nand4_1 _1383_ (.B(_0559_),
    .C(_0560_),
    .A(_0558_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_or2_1 _1384_ (.X(_0565_),
    .B(_0563_),
    .A(_0561_));
 sg13g2_nand4_1 _1385_ (.B(_0559_),
    .C(_0564_),
    .A(generating),
    .Y(_0566_),
    .D(_0565_));
 sg13g2_inv_1 _1386_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_nand2b_2 _1387_ (.Y(_0568_),
    .B(\hvsync_gen.hpos[9] ),
    .A_N(\hvsync_gen.hpos[7] ));
 sg13g2_and2_1 _1388_ (.A(net174),
    .B(_0568_),
    .X(_0569_));
 sg13g2_nor2b_1 _1389_ (.A(\hvsync_gen.hpos[9] ),
    .B_N(\hvsync_gen.hpos[7] ),
    .Y(_0570_));
 sg13g2_or2_1 _1390_ (.X(_0571_),
    .B(_0570_),
    .A(net175));
 sg13g2_nor2_1 _1391_ (.A(net174),
    .B(_0568_),
    .Y(_0572_));
 sg13g2_a21oi_1 _1392_ (.A1(_0569_),
    .A2(_0571_),
    .Y(_0573_),
    .B1(_0572_));
 sg13g2_a22oi_1 _1393_ (.Y(_0574_),
    .B1(_0573_),
    .B2(_0569_),
    .A2(_0572_),
    .A1(net175));
 sg13g2_a21oi_1 _1394_ (.A1(net175),
    .A2(_0341_),
    .Y(_0575_),
    .B1(_0568_));
 sg13g2_nand2b_1 _1395_ (.Y(_0576_),
    .B(net174),
    .A_N(net175));
 sg13g2_a21oi_1 _1396_ (.A1(_0570_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0575_));
 sg13g2_inv_1 _1397_ (.Y(_0578_),
    .A(_0577_));
 sg13g2_xnor2_1 _1398_ (.Y(_0579_),
    .A(net175),
    .B(_0573_));
 sg13g2_nor2_1 _1399_ (.A(net176),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_o21ai_1 _1400_ (.B1(_0578_),
    .Y(_0581_),
    .A1(net176),
    .A2(_0579_));
 sg13g2_and2_1 _1401_ (.A(_0574_),
    .B(_0581_),
    .X(_0582_));
 sg13g2_a21o_1 _1402_ (.A2(_0581_),
    .A1(_0574_),
    .B1(net176),
    .X(_0583_));
 sg13g2_nand3_1 _1403_ (.B(_0574_),
    .C(_0581_),
    .A(net176),
    .Y(_0584_));
 sg13g2_nand2_1 _1404_ (.Y(_0585_),
    .A(_0583_),
    .B(_0584_));
 sg13g2_nand3_1 _1405_ (.B(_0583_),
    .C(_0584_),
    .A(_0340_),
    .Y(_0586_));
 sg13g2_xnor2_1 _1406_ (.Y(_0587_),
    .A(_0579_),
    .B(_0583_));
 sg13g2_nand2_1 _1407_ (.Y(_0588_),
    .A(_0586_),
    .B(_0587_));
 sg13g2_o21ai_1 _1408_ (.B1(_0577_),
    .Y(_0589_),
    .A1(_0574_),
    .A2(_0580_));
 sg13g2_nand2_1 _1409_ (.Y(_0590_),
    .A(_0581_),
    .B(_0589_));
 sg13g2_or2_1 _1410_ (.X(_0591_),
    .B(_0590_),
    .A(_0586_));
 sg13g2_nand2b_1 _1411_ (.Y(_0592_),
    .B(_0586_),
    .A_N(_0590_));
 sg13g2_nand2b_1 _1412_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0587_));
 sg13g2_and2_1 _1413_ (.A(_0588_),
    .B(_0593_),
    .X(_0594_));
 sg13g2_nand2_1 _1414_ (.Y(_0595_),
    .A(_0588_),
    .B(_0593_));
 sg13g2_a22oi_1 _1415_ (.Y(_0596_),
    .B1(_0589_),
    .B2(_0581_),
    .A2(_0587_),
    .A1(_0586_));
 sg13g2_o21ai_1 _1416_ (.B1(_0585_),
    .Y(_0597_),
    .A1(\hvsync_gen.hpos[4] ),
    .A2(net142));
 sg13g2_and2_1 _1417_ (.A(_0591_),
    .B(_0597_),
    .X(_0598_));
 sg13g2_xnor2_1 _1418_ (.Y(_0599_),
    .A(_0340_),
    .B(net142));
 sg13g2_xnor2_1 _1419_ (.Y(_0600_),
    .A(net178),
    .B(net142));
 sg13g2_nor2_1 _1420_ (.A(net179),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_a22oi_1 _1421_ (.Y(_0602_),
    .B1(_0599_),
    .B2(_0343_),
    .A2(_0597_),
    .A1(_0591_));
 sg13g2_nor2_2 _1422_ (.A(_0594_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1423_ (.Y(_0604_),
    .A(\solver_r_y[2] ),
    .B(_0539_));
 sg13g2_xnor2_1 _1424_ (.Y(_0605_),
    .A(\solver_r_x[2] ),
    .B(_0582_));
 sg13g2_xnor2_1 _1425_ (.Y(_0606_),
    .A(\solver_r_y[1] ),
    .B(net144));
 sg13g2_xnor2_1 _1426_ (.Y(_0607_),
    .A(\solver_r_x[1] ),
    .B(net142));
 sg13g2_nor4_1 _1427_ (.A(_0604_),
    .B(_0605_),
    .C(_0606_),
    .D(_0607_),
    .Y(_0608_));
 sg13g2_xor2_1 _1428_ (.B(net141),
    .A(net171),
    .X(_0609_));
 sg13g2_xnor2_1 _1429_ (.Y(_0610_),
    .A(_0332_),
    .B(_0603_));
 sg13g2_nand3_1 _1430_ (.B(_0609_),
    .C(_0610_),
    .A(_0608_),
    .Y(_0611_));
 sg13g2_inv_1 _1431_ (.Y(_0612_),
    .A(_0611_));
 sg13g2_xnor2_1 _1432_ (.Y(_0613_),
    .A(_0344_),
    .B(_0603_));
 sg13g2_xnor2_1 _1433_ (.Y(_0614_),
    .A(\player_y[2] ),
    .B(net152));
 sg13g2_a21oi_1 _1434_ (.A1(\player_x[2] ),
    .A2(_0582_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_o21ai_1 _1435_ (.B1(_0615_),
    .Y(_0616_),
    .A1(\player_x[2] ),
    .A2(_0582_));
 sg13g2_xnor2_1 _1436_ (.Y(_0617_),
    .A(\player_x[1] ),
    .B(net142));
 sg13g2_xnor2_1 _1437_ (.Y(_0618_),
    .A(\player_y[1] ),
    .B(net144));
 sg13g2_nor3_1 _1438_ (.A(_0616_),
    .B(_0617_),
    .C(_0618_),
    .Y(_0619_));
 sg13g2_xor2_1 _1439_ (.B(net140),
    .A(net173),
    .X(_0620_));
 sg13g2_nand3_1 _1440_ (.B(_0619_),
    .C(_0620_),
    .A(_0613_),
    .Y(_0621_));
 sg13g2_nor2_1 _1441_ (.A(_0611_),
    .B(_0621_),
    .Y(_0622_));
 sg13g2_or2_1 _1442_ (.X(_0623_),
    .B(_0621_),
    .A(_0611_));
 sg13g2_o21ai_1 _1443_ (.B1(_0343_),
    .Y(_0624_),
    .A1(_0594_),
    .A2(_0602_));
 sg13g2_nand3_1 _1444_ (.B(_0595_),
    .C(_0598_),
    .A(net179),
    .Y(_0625_));
 sg13g2_a21oi_2 _1445_ (.B1(_0342_),
    .Y(_0626_),
    .A2(_0625_),
    .A1(_0624_));
 sg13g2_and3_1 _1446_ (.X(_0627_),
    .A(_0342_),
    .B(_0624_),
    .C(_0625_));
 sg13g2_nor2_1 _1447_ (.A(\hvsync_gen.vpos[3] ),
    .B(net141),
    .Y(_0628_));
 sg13g2_xnor2_1 _1448_ (.Y(_0629_),
    .A(\hvsync_gen.vpos[3] ),
    .B(net141));
 sg13g2_nor2_1 _1449_ (.A(\hvsync_gen.vpos[2] ),
    .B(_0629_),
    .Y(_0630_));
 sg13g2_nand2_1 _1450_ (.Y(_0631_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_0629_));
 sg13g2_nand2b_2 _1451_ (.Y(_0632_),
    .B(_0631_),
    .A_N(_0630_));
 sg13g2_nor3_1 _1452_ (.A(_0626_),
    .B(_0627_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_or3_1 _1453_ (.A(_0626_),
    .B(_0627_),
    .C(_0632_),
    .X(_0634_));
 sg13g2_xor2_1 _1454_ (.B(net180),
    .A(\hvsync_gen.vpos[2] ),
    .X(_0635_));
 sg13g2_nand2_1 _1455_ (.Y(_0636_),
    .A(\ent_x[0] ),
    .B(net169));
 sg13g2_xor2_1 _1456_ (.B(net181),
    .A(net168),
    .X(_0637_));
 sg13g2_nor2b_1 _1457_ (.A(_0636_),
    .B_N(_0637_),
    .Y(_0638_));
 sg13g2_a21o_1 _1458_ (.A2(net181),
    .A1(net168),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_nand2_1 _1459_ (.Y(_0640_),
    .A(_0635_),
    .B(_0639_));
 sg13g2_o21ai_1 _1460_ (.B1(_0640_),
    .Y(_0641_),
    .A1(\hvsync_gen.vpos[2] ),
    .A2(net180));
 sg13g2_o21ai_1 _1461_ (.B1(_0632_),
    .Y(_0642_),
    .A1(_0626_),
    .A2(_0627_));
 sg13g2_nand3_1 _1462_ (.B(_0641_),
    .C(_0642_),
    .A(_0634_),
    .Y(_0643_));
 sg13g2_a21o_2 _1463_ (.A2(_0642_),
    .A1(_0641_),
    .B1(_0633_),
    .X(_0644_));
 sg13g2_xor2_1 _1464_ (.B(_0639_),
    .A(_0635_),
    .X(_0645_));
 sg13g2_a21o_1 _1465_ (.A2(_0642_),
    .A1(_0634_),
    .B1(_0641_),
    .X(_0646_));
 sg13g2_a21o_1 _1466_ (.A2(_0646_),
    .A1(_0643_),
    .B1(_0645_),
    .X(_0647_));
 sg13g2_nand3_1 _1467_ (.B(_0644_),
    .C(_0647_),
    .A(_0622_),
    .Y(_0648_));
 sg13g2_or2_1 _1468_ (.X(_0649_),
    .B(net169),
    .A(\ent_x[0] ));
 sg13g2_and2_1 _1469_ (.A(_0636_),
    .B(_0637_),
    .X(_0650_));
 sg13g2_and3_1 _1470_ (.X(_0651_),
    .A(_0645_),
    .B(_0649_),
    .C(_0650_));
 sg13g2_a21oi_2 _1471_ (.B1(_0644_),
    .Y(_0652_),
    .A2(_0651_),
    .A1(_0646_));
 sg13g2_nand2_1 _1472_ (.Y(_0653_),
    .A(_0611_),
    .B(_0621_));
 sg13g2_o21ai_1 _1473_ (.B1(_0653_),
    .Y(_0654_),
    .A1(_0622_),
    .A2(_0652_));
 sg13g2_nand2b_1 _1474_ (.Y(_0655_),
    .B(_0648_),
    .A_N(_0654_));
 sg13g2_xnor2_1 _1475_ (.Y(_0656_),
    .A(_0326_),
    .B(_0603_));
 sg13g2_xor2_1 _1476_ (.B(net141),
    .A(net170),
    .X(_0657_));
 sg13g2_xnor2_1 _1477_ (.Y(_0658_),
    .A(\solver_l_y[1] ),
    .B(_0548_));
 sg13g2_xnor2_1 _1478_ (.Y(_0659_),
    .A(\solver_l_y[2] ),
    .B(_0539_));
 sg13g2_xnor2_1 _1479_ (.Y(_0660_),
    .A(\solver_l_x[2] ),
    .B(_0582_));
 sg13g2_xnor2_1 _1480_ (.Y(_0661_),
    .A(\solver_l_x[1] ),
    .B(net142));
 sg13g2_nor4_1 _1481_ (.A(_0658_),
    .B(_0659_),
    .C(_0660_),
    .D(_0661_),
    .Y(_0662_));
 sg13g2_nand3_1 _1482_ (.B(_0657_),
    .C(_0662_),
    .A(_0656_),
    .Y(_0663_));
 sg13g2_inv_1 _1483_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_xnor2_1 _1484_ (.Y(_0665_),
    .A(_0600_),
    .B(_0624_));
 sg13g2_xnor2_1 _1485_ (.Y(_0666_),
    .A(_0554_),
    .B(_0628_));
 sg13g2_mux2_1 _1486_ (.A0(_0595_),
    .A1(_0598_),
    .S(_0601_),
    .X(_0667_));
 sg13g2_a21oi_1 _1487_ (.A1(_0552_),
    .A2(_0555_),
    .Y(_0668_),
    .B1(_0556_));
 sg13g2_a21o_1 _1488_ (.A2(_0556_),
    .A1(_0555_),
    .B1(_0668_),
    .X(_0669_));
 sg13g2_nand3_1 _1489_ (.B(_0667_),
    .C(_0669_),
    .A(_0312_),
    .Y(_0670_));
 sg13g2_xnor2_1 _1490_ (.Y(_0671_),
    .A(_0631_),
    .B(_0666_));
 sg13g2_xnor2_1 _1491_ (.Y(_0672_),
    .A(_0626_),
    .B(_0665_));
 sg13g2_nor3_1 _1492_ (.A(_0670_),
    .B(_0671_),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_nor2_1 _1493_ (.A(net144),
    .B(net140),
    .Y(_0674_));
 sg13g2_xnor2_1 _1494_ (.Y(_0675_),
    .A(\maze_seed[2] ),
    .B(net152));
 sg13g2_xnor2_1 _1495_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_or3_1 _1496_ (.A(\maze_seed[4] ),
    .B(_0594_),
    .C(_0602_),
    .X(_0677_));
 sg13g2_o21ai_1 _1497_ (.B1(\maze_seed[4] ),
    .Y(_0678_),
    .A1(_0594_),
    .A2(_0602_));
 sg13g2_xnor2_1 _1498_ (.Y(_0679_),
    .A(_0318_),
    .B(net142));
 sg13g2_nand3_1 _1499_ (.B(_0678_),
    .C(_0679_),
    .A(_0677_),
    .Y(_0680_));
 sg13g2_a21o_1 _1500_ (.A2(_0678_),
    .A1(_0677_),
    .B1(_0679_),
    .X(_0681_));
 sg13g2_a21o_1 _1501_ (.A2(_0681_),
    .A1(_0680_),
    .B1(_0676_),
    .X(_0682_));
 sg13g2_nand3_1 _1502_ (.B(_0680_),
    .C(_0681_),
    .A(_0676_),
    .Y(_0683_));
 sg13g2_xnor2_1 _1503_ (.Y(_0684_),
    .A(\maze_seed[1] ),
    .B(_0582_));
 sg13g2_xnor2_1 _1504_ (.Y(_0685_),
    .A(net144),
    .B(_0684_));
 sg13g2_xor2_1 _1505_ (.B(_0685_),
    .A(net140),
    .X(_0686_));
 sg13g2_nand2_1 _1506_ (.Y(_0687_),
    .A(net182),
    .B(_0686_));
 sg13g2_xor2_1 _1507_ (.B(_0679_),
    .A(net140),
    .X(_0688_));
 sg13g2_nand2_1 _1508_ (.Y(_0689_),
    .A(_0676_),
    .B(_0688_));
 sg13g2_o21ai_1 _1509_ (.B1(_0689_),
    .Y(_0690_),
    .A1(net182),
    .A2(_0686_));
 sg13g2_and4_1 _1510_ (.A(_0682_),
    .B(_0683_),
    .C(_0687_),
    .D(_0690_),
    .X(_0691_));
 sg13g2_nor3_1 _1511_ (.A(net152),
    .B(net144),
    .C(net140),
    .Y(_0692_));
 sg13g2_a22oi_1 _1512_ (.Y(_0693_),
    .B1(_0687_),
    .B2(_0690_),
    .A2(_0683_),
    .A1(_0682_));
 sg13g2_nor3_1 _1513_ (.A(_0691_),
    .B(_0692_),
    .C(_0693_),
    .Y(_0694_));
 sg13g2_o21ai_1 _1514_ (.B1(\hvsync_gen.vpos[2] ),
    .Y(_0695_),
    .A1(net169),
    .A2(net168));
 sg13g2_nor2_1 _1515_ (.A(_0554_),
    .B(_0629_),
    .Y(_0696_));
 sg13g2_a21o_1 _1516_ (.A2(_0696_),
    .A1(_0695_),
    .B1(_0669_),
    .X(_0697_));
 sg13g2_xor2_1 _1517_ (.B(_0686_),
    .A(_0675_),
    .X(_0698_));
 sg13g2_nand3_1 _1518_ (.B(_0678_),
    .C(_0698_),
    .A(_0677_),
    .Y(_0699_));
 sg13g2_a21o_1 _1519_ (.A2(_0678_),
    .A1(_0677_),
    .B1(_0698_),
    .X(_0700_));
 sg13g2_and2_1 _1520_ (.A(net182),
    .B(_0685_),
    .X(_0701_));
 sg13g2_nor3_1 _1521_ (.A(net182),
    .B(_0675_),
    .C(_0685_),
    .Y(_0702_));
 sg13g2_a21oi_1 _1522_ (.A1(_0675_),
    .A2(_0701_),
    .Y(_0703_),
    .B1(_0702_));
 sg13g2_mux2_1 _1523_ (.A0(_0703_),
    .A1(_0701_),
    .S(_0688_),
    .X(_0704_));
 sg13g2_nand3_1 _1524_ (.B(_0700_),
    .C(_0704_),
    .A(_0699_),
    .Y(_0705_));
 sg13g2_nand3_1 _1525_ (.B(net144),
    .C(net140),
    .A(net152),
    .Y(_0706_));
 sg13g2_a21o_1 _1526_ (.A2(_0700_),
    .A1(_0699_),
    .B1(_0704_),
    .X(_0707_));
 sg13g2_nand3_1 _1527_ (.B(_0706_),
    .C(_0707_),
    .A(_0705_),
    .Y(_0708_));
 sg13g2_nand2_1 _1528_ (.Y(_0709_),
    .A(net169),
    .B(net168));
 sg13g2_and4_1 _1529_ (.A(_0630_),
    .B(_0666_),
    .C(_0669_),
    .D(_0709_),
    .X(_0710_));
 sg13g2_and2_1 _1530_ (.A(net223),
    .B(net181),
    .X(_0711_));
 sg13g2_nor2_1 _1531_ (.A(net180),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_nor3_1 _1532_ (.A(net180),
    .B(net179),
    .C(_0711_),
    .Y(_0713_));
 sg13g2_a21oi_1 _1533_ (.A1(_0582_),
    .A2(net142),
    .Y(_0714_),
    .B1(_0706_));
 sg13g2_nand3_1 _1534_ (.B(_0598_),
    .C(_0713_),
    .A(_0595_),
    .Y(_0715_));
 sg13g2_nor3_1 _1535_ (.A(_0665_),
    .B(_0714_),
    .C(_0715_),
    .Y(_0716_));
 sg13g2_nor2_1 _1536_ (.A(_0582_),
    .B(_0596_),
    .Y(_0717_));
 sg13g2_or2_1 _1537_ (.X(_0718_),
    .B(_0717_),
    .A(_0706_));
 sg13g2_nor2_1 _1538_ (.A(net223),
    .B(net181),
    .Y(_0719_));
 sg13g2_o21ai_1 _1539_ (.B1(net180),
    .Y(_0720_),
    .A1(\ent_x[0] ),
    .A2(\ent_x[1] ));
 sg13g2_and2_1 _1540_ (.A(_0599_),
    .B(_0720_),
    .X(_0721_));
 sg13g2_a221oi_1 _1541_ (.B2(net179),
    .C1(_0595_),
    .B1(_0721_),
    .A1(_0598_),
    .Y(_0722_),
    .A2(_0601_));
 sg13g2_a221oi_1 _1542_ (.B2(_0722_),
    .C1(_0716_),
    .B1(_0718_),
    .A1(_0708_),
    .Y(_0723_),
    .A2(_0710_));
 sg13g2_o21ai_1 _1543_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0694_),
    .A2(_0697_));
 sg13g2_nor2_1 _1544_ (.A(_0312_),
    .B(_0564_),
    .Y(_0725_));
 sg13g2_inv_1 _1545_ (.Y(_0726_),
    .A(_0725_));
 sg13g2_nand2_1 _1546_ (.Y(_0727_),
    .A(_0621_),
    .B(_0663_));
 sg13g2_o21ai_1 _1547_ (.B1(_0673_),
    .Y(_0728_),
    .A1(_0653_),
    .A2(_0664_));
 sg13g2_nor2_1 _1548_ (.A(_0663_),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_a221oi_1 _1549_ (.B2(_0655_),
    .C1(solver_l_won),
    .B1(_0729_),
    .A1(_0724_),
    .Y(_0730_),
    .A2(_0726_));
 sg13g2_nand2_1 _1550_ (.Y(_0731_),
    .A(_0692_),
    .B(_0717_));
 sg13g2_nor4_1 _1551_ (.A(_0603_),
    .B(_0653_),
    .C(_0664_),
    .D(_0731_),
    .Y(_0732_));
 sg13g2_and2_1 _1552_ (.A(_0673_),
    .B(_0732_),
    .X(_0733_));
 sg13g2_or2_1 _1553_ (.X(_0734_),
    .B(_0733_),
    .A(_0725_));
 sg13g2_nor3_1 _1554_ (.A(_0724_),
    .B(_0725_),
    .C(_0733_),
    .Y(_0735_));
 sg13g2_nand2_1 _1555_ (.Y(_0736_),
    .A(_0728_),
    .B(_0735_));
 sg13g2_a21o_1 _1556_ (.A2(_0736_),
    .A1(_0730_),
    .B1(_0350_),
    .X(_0737_));
 sg13g2_a21o_1 _1557_ (.A2(_0737_),
    .A1(_0566_),
    .B1(_0525_),
    .X(_0738_));
 sg13g2_nor4_1 _1558_ (.A(\hvsync_gen.vpos[4] ),
    .B(net166),
    .C(net167),
    .D(\hvsync_gen.vpos[6] ),
    .Y(_0739_));
 sg13g2_nand3_1 _1559_ (.B(_0339_),
    .C(_0739_),
    .A(_0338_),
    .Y(_0740_));
 sg13g2_nor4_1 _1560_ (.A(net169),
    .B(net168),
    .C(_0335_),
    .D(_0336_),
    .Y(_0741_));
 sg13g2_nor3_1 _1561_ (.A(net168),
    .B(_0335_),
    .C(\hvsync_gen.vpos[3] ),
    .Y(_0742_));
 sg13g2_a21oi_1 _1562_ (.A1(\ent_y[0] ),
    .A2(_0742_),
    .Y(_0743_),
    .B1(_0741_));
 sg13g2_nor3_1 _1563_ (.A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[9] ),
    .C(_0523_),
    .Y(_0744_));
 sg13g2_nor3_1 _1564_ (.A(\ent_x[0] ),
    .B(net180),
    .C(net179),
    .Y(_0745_));
 sg13g2_and4_1 _1565_ (.A(net177),
    .B(_0340_),
    .C(\ent_x[1] ),
    .D(_0745_),
    .X(_0746_));
 sg13g2_nor3_1 _1566_ (.A(net177),
    .B(net178),
    .C(net179),
    .Y(_0747_));
 sg13g2_nor2_1 _1567_ (.A(_0342_),
    .B(net181),
    .Y(_0748_));
 sg13g2_and3_1 _1568_ (.X(_0749_),
    .A(\ent_x[0] ),
    .B(_0747_),
    .C(_0748_));
 sg13g2_o21ai_1 _1569_ (.B1(_0744_),
    .Y(_0750_),
    .A1(_0746_),
    .A2(_0749_));
 sg13g2_o21ai_1 _1570_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0740_),
    .A2(_0743_));
 sg13g2_a22oi_1 _1571_ (.Y(_0752_),
    .B1(_0720_),
    .B2(_0747_),
    .A2(net178),
    .A1(net177));
 sg13g2_nand2_1 _1572_ (.Y(_0753_),
    .A(_0744_),
    .B(_0752_));
 sg13g2_xnor2_1 _1573_ (.Y(_0754_),
    .A(_0336_),
    .B(_0695_));
 sg13g2_nor2b_1 _1574_ (.A(_0713_),
    .B_N(net177),
    .Y(_0755_));
 sg13g2_nor4_1 _1575_ (.A(_0740_),
    .B(_0753_),
    .C(_0754_),
    .D(_0755_),
    .Y(_0756_));
 sg13g2_nand2_2 _1576_ (.Y(_0757_),
    .A(_0751_),
    .B(_0756_));
 sg13g2_o21ai_1 _1577_ (.B1(_0738_),
    .Y(uo_out[6]),
    .A1(single_step_mode),
    .A2(_0757_));
 sg13g2_o21ai_1 _1578_ (.B1(_0730_),
    .Y(_0758_),
    .A1(_0724_),
    .A2(_0726_));
 sg13g2_nand2b_1 _1579_ (.Y(_0759_),
    .B(_0566_),
    .A_N(_0525_));
 sg13g2_nor2_1 _1580_ (.A(_0350_),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_nand2_1 _1581_ (.Y(_0761_),
    .A(_0758_),
    .B(_0760_));
 sg13g2_o21ai_1 _1582_ (.B1(_0761_),
    .Y(uo_out[2]),
    .A1(single_step_mode),
    .A2(_0757_));
 sg13g2_nand2_1 _1583_ (.Y(_0762_),
    .A(_0612_),
    .B(_0664_));
 sg13g2_mux2_1 _1584_ (.A0(_0623_),
    .A1(_0762_),
    .S(_0652_),
    .X(_0763_));
 sg13g2_nor2_1 _1585_ (.A(_0623_),
    .B(_0663_),
    .Y(_0764_));
 sg13g2_nor2_1 _1586_ (.A(_0645_),
    .B(_0650_),
    .Y(_0765_));
 sg13g2_o21ai_1 _1587_ (.B1(_0765_),
    .Y(_0766_),
    .A1(_0636_),
    .A2(_0637_));
 sg13g2_a21oi_1 _1588_ (.A1(_0646_),
    .A2(_0766_),
    .Y(_0767_),
    .B1(_0644_));
 sg13g2_a21oi_1 _1589_ (.A1(_0644_),
    .A2(_0647_),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_a21o_1 _1590_ (.A2(_0647_),
    .A1(_0644_),
    .B1(_0767_),
    .X(_0769_));
 sg13g2_a22oi_1 _1591_ (.Y(_0770_),
    .B1(_0764_),
    .B2(_0769_),
    .A2(_0763_),
    .A1(_0727_));
 sg13g2_nor2_1 _1592_ (.A(solver_l_won),
    .B(_0724_),
    .Y(_0771_));
 sg13g2_o21ai_1 _1593_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0728_),
    .A2(_0770_));
 sg13g2_o21ai_1 _1594_ (.B1(_0325_),
    .Y(_0773_),
    .A1(_0734_),
    .A2(_0772_));
 sg13g2_nor2_1 _1595_ (.A(player_won),
    .B(_0567_),
    .Y(_0774_));
 sg13g2_a21oi_1 _1596_ (.A1(_0773_),
    .A2(_0774_),
    .Y(_0775_),
    .B1(_0525_));
 sg13g2_nor2_1 _1597_ (.A(\solver_speed[1] ),
    .B(\filled_width[1] ),
    .Y(_0776_));
 sg13g2_nor3_1 _1598_ (.A(\solver_speed[2] ),
    .B(\solver_speed[1] ),
    .C(\filled_width[1] ),
    .Y(_0777_));
 sg13g2_xnor2_1 _1599_ (.Y(_0778_),
    .A(net386),
    .B(_0777_));
 sg13g2_a21oi_1 _1600_ (.A1(net180),
    .A2(net181),
    .Y(_0779_),
    .B1(net179));
 sg13g2_xnor2_1 _1601_ (.Y(_0780_),
    .A(net178),
    .B(_0779_));
 sg13g2_nand3_1 _1602_ (.B(net181),
    .C(\hvsync_gen.hpos[3] ),
    .A(\hvsync_gen.hpos[2] ),
    .Y(_0781_));
 sg13g2_nor2b_1 _1603_ (.A(_0779_),
    .B_N(_0781_),
    .Y(_0782_));
 sg13g2_xnor2_1 _1604_ (.Y(_0783_),
    .A(net328),
    .B(_0776_));
 sg13g2_or2_1 _1605_ (.X(_0784_),
    .B(net181),
    .A(\filled_width[1] ));
 sg13g2_nand3_1 _1606_ (.B(_0342_),
    .C(_0784_),
    .A(\solver_speed[1] ),
    .Y(_0785_));
 sg13g2_o21ai_1 _1607_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0782_),
    .A2(_0783_));
 sg13g2_nor3_1 _1608_ (.A(_0748_),
    .B(_0776_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_a221oi_1 _1609_ (.B2(_0783_),
    .C1(_0787_),
    .B1(_0782_),
    .A1(_0778_),
    .Y(_0788_),
    .A2(_0780_));
 sg13g2_nor2_1 _1610_ (.A(_0778_),
    .B(_0780_),
    .Y(_0789_));
 sg13g2_nand2b_1 _1611_ (.Y(_0790_),
    .B(_0756_),
    .A_N(_0788_));
 sg13g2_o21ai_1 _1612_ (.B1(_0757_),
    .Y(_0791_),
    .A1(_0789_),
    .A2(_0790_));
 sg13g2_or2_1 _1613_ (.X(uo_out[5]),
    .B(_0791_),
    .A(_0775_));
 sg13g2_o21ai_1 _1614_ (.B1(_0325_),
    .Y(_0792_),
    .A1(_0733_),
    .A2(_0772_));
 sg13g2_a21oi_1 _1615_ (.A1(_0324_),
    .A2(_0792_),
    .Y(_0793_),
    .B1(_0759_));
 sg13g2_or2_1 _1616_ (.X(uo_out[1]),
    .B(_0793_),
    .A(_0791_));
 sg13g2_mux2_1 _1617_ (.A0(_0663_),
    .A1(_0621_),
    .S(_0652_),
    .X(_0794_));
 sg13g2_a22oi_1 _1618_ (.Y(_0795_),
    .B1(_0794_),
    .B2(_0612_),
    .A2(_0768_),
    .A1(_0764_));
 sg13g2_nor2_1 _1619_ (.A(_0724_),
    .B(_0733_),
    .Y(_0796_));
 sg13g2_o21ai_1 _1620_ (.B1(_0796_),
    .Y(_0797_),
    .A1(_0728_),
    .A2(_0795_));
 sg13g2_a21o_1 _1621_ (.A2(_0797_),
    .A1(_0323_),
    .B1(solver_r_won),
    .X(_0798_));
 sg13g2_nand2_1 _1622_ (.Y(_0799_),
    .A(_0324_),
    .B(_0798_));
 sg13g2_a21oi_1 _1623_ (.A1(_0324_),
    .A2(_0798_),
    .Y(_0800_),
    .B1(_0567_));
 sg13g2_o21ai_1 _1624_ (.B1(_0757_),
    .Y(uo_out[4]),
    .A1(_0525_),
    .A2(_0800_));
 sg13g2_o21ai_1 _1625_ (.B1(_0757_),
    .Y(uo_out[0]),
    .A1(_0759_),
    .A2(_0799_));
 sg13g2_and2_1 _1626_ (.A(net247),
    .B(net201),
    .X(_0010_));
 sg13g2_xnor2_1 _1627_ (.Y(_0801_),
    .A(net273),
    .B(net255));
 sg13g2_xnor2_1 _1628_ (.Y(_0802_),
    .A(net234),
    .B(net292));
 sg13g2_a21oi_1 _1629_ (.A1(_0801_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0346_));
 sg13g2_o21ai_1 _1630_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0801_),
    .A2(_0802_));
 sg13g2_a21oi_1 _1631_ (.A1(net288),
    .A2(_0346_),
    .Y(_0805_),
    .B1(net196));
 sg13g2_nand2_1 _1632_ (.Y(_0011_),
    .A(_0804_),
    .B(_0805_));
 sg13g2_o21ai_1 _1633_ (.B1(net202),
    .Y(_0806_),
    .A1(net245),
    .A2(net164));
 sg13g2_a21oi_1 _1634_ (.A1(_0319_),
    .A2(net164),
    .Y(_0012_),
    .B1(_0806_));
 sg13g2_a21oi_1 _1635_ (.A1(net245),
    .A2(net164),
    .Y(_0807_),
    .B1(net193));
 sg13g2_o21ai_1 _1636_ (.B1(_0807_),
    .Y(_0013_),
    .A1(_0317_),
    .A2(net164));
 sg13g2_o21ai_1 _1637_ (.B1(net202),
    .Y(_0808_),
    .A1(net255),
    .A2(net164));
 sg13g2_a21oi_1 _1638_ (.A1(_0317_),
    .A2(net164),
    .Y(_0014_),
    .B1(net256));
 sg13g2_o21ai_1 _1639_ (.B1(net201),
    .Y(_0809_),
    .A1(net273),
    .A2(net165));
 sg13g2_a21oi_1 _1640_ (.A1(_0315_),
    .A2(net165),
    .Y(_0015_),
    .B1(net274));
 sg13g2_a21oi_1 _1641_ (.A1(net273),
    .A2(net165),
    .Y(_0810_),
    .B1(net196));
 sg13g2_o21ai_1 _1642_ (.B1(_0810_),
    .Y(_0016_),
    .A1(_0321_),
    .A2(net165));
 sg13g2_o21ai_1 _1643_ (.B1(net200),
    .Y(_0811_),
    .A1(\lfsr[5] ),
    .A2(net163));
 sg13g2_a21oi_1 _1644_ (.A1(_0320_),
    .A2(net163),
    .Y(_0017_),
    .B1(_0811_));
 sg13g2_a21oi_1 _1645_ (.A1(net234),
    .A2(net163),
    .Y(_0812_),
    .B1(net194));
 sg13g2_o21ai_1 _1646_ (.B1(net235),
    .Y(_0018_),
    .A1(_0320_),
    .A2(net163));
 sg13g2_a22oi_1 _1647_ (.Y(_0019_),
    .B1(_0432_),
    .B2(_0319_),
    .A2(net149),
    .A1(_0318_));
 sg13g2_a22oi_1 _1648_ (.Y(_0813_),
    .B1(_0432_),
    .B2(net245),
    .A2(net149),
    .A1(\maze_seed[1] ));
 sg13g2_inv_1 _1649_ (.Y(_0020_),
    .A(net246));
 sg13g2_a22oi_1 _1650_ (.Y(_0021_),
    .B1(_0432_),
    .B2(_0317_),
    .A2(net149),
    .A1(_0316_));
 sg13g2_a22oi_1 _1651_ (.Y(_0814_),
    .B1(_0432_),
    .B2(net255),
    .A2(net149),
    .A1(net184));
 sg13g2_inv_1 _1652_ (.Y(_0022_),
    .A(_0814_));
 sg13g2_a22oi_1 _1653_ (.Y(_0815_),
    .B1(_0432_),
    .B2(net273),
    .A2(net149),
    .A1(net299));
 sg13g2_inv_1 _1654_ (.Y(_0023_),
    .A(_0815_));
 sg13g2_and2_1 _1655_ (.A(net347),
    .B(_0711_),
    .X(_0816_));
 sg13g2_and2_1 _1656_ (.A(net332),
    .B(_0816_),
    .X(_0817_));
 sg13g2_nand2_1 _1657_ (.Y(_0818_),
    .A(net178),
    .B(_0817_));
 sg13g2_inv_2 _1658_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_nor4_2 _1659_ (.A(net176),
    .B(_0568_),
    .C(_0576_),
    .Y(_0820_),
    .D(_0818_));
 sg13g2_nor2_2 _1660_ (.A(net198),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_nand2b_2 _1661_ (.Y(_0822_),
    .B(net203),
    .A_N(_0820_));
 sg13g2_nor2_1 _1662_ (.A(net223),
    .B(_0822_),
    .Y(_0024_));
 sg13g2_nor3_1 _1663_ (.A(_0711_),
    .B(_0719_),
    .C(_0822_),
    .Y(_0025_));
 sg13g2_nor3_1 _1664_ (.A(net198),
    .B(_0712_),
    .C(_0816_),
    .Y(_0026_));
 sg13g2_o21ai_1 _1665_ (.B1(net203),
    .Y(_0823_),
    .A1(net332),
    .A2(_0816_));
 sg13g2_nor2_1 _1666_ (.A(net333),
    .B(_0823_),
    .Y(_0027_));
 sg13g2_o21ai_1 _1667_ (.B1(net203),
    .Y(_0824_),
    .A1(net178),
    .A2(_0817_));
 sg13g2_nor2_1 _1668_ (.A(_0819_),
    .B(_0824_),
    .Y(_0028_));
 sg13g2_o21ai_1 _1669_ (.B1(net145),
    .Y(_0825_),
    .A1(net176),
    .A2(_0819_));
 sg13g2_a21oi_1 _1670_ (.A1(net177),
    .A2(_0819_),
    .Y(_0029_),
    .B1(_0825_));
 sg13g2_a21oi_1 _1671_ (.A1(net177),
    .A2(_0819_),
    .Y(_0826_),
    .B1(net175));
 sg13g2_and2_1 _1672_ (.A(_0518_),
    .B(_0817_),
    .X(_0827_));
 sg13g2_nor3_1 _1673_ (.A(_0822_),
    .B(_0826_),
    .C(_0827_),
    .Y(_0030_));
 sg13g2_nor2_1 _1674_ (.A(net276),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_and2_1 _1675_ (.A(net276),
    .B(_0827_),
    .X(_0829_));
 sg13g2_nor3_1 _1676_ (.A(_0822_),
    .B(_0828_),
    .C(_0829_),
    .Y(_0031_));
 sg13g2_or2_1 _1677_ (.X(_0830_),
    .B(_0829_),
    .A(net174));
 sg13g2_nand2_1 _1678_ (.Y(_0831_),
    .A(net377),
    .B(_0829_));
 sg13g2_nand3_1 _1679_ (.B(_0830_),
    .C(_0831_),
    .A(_0821_),
    .Y(_0832_));
 sg13g2_inv_1 _1680_ (.Y(_0032_),
    .A(_0832_));
 sg13g2_xor2_1 _1681_ (.B(_0831_),
    .A(net352),
    .X(_0833_));
 sg13g2_nor2_1 _1682_ (.A(_0822_),
    .B(net353),
    .Y(_0033_));
 sg13g2_nor3_2 _1683_ (.A(\player_y[2] ),
    .B(\player_y[1] ),
    .C(net173),
    .Y(_0834_));
 sg13g2_and2_1 _1684_ (.A(\player_x[1] ),
    .B(net286),
    .X(_0835_));
 sg13g2_nand2_1 _1685_ (.Y(_0836_),
    .A(\player_x[2] ),
    .B(_0835_));
 sg13g2_o21ai_1 _1686_ (.B1(_0836_),
    .Y(_0837_),
    .A1(_0344_),
    .A2(_0834_));
 sg13g2_nor2_1 _1687_ (.A(inp_right_prev),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_nand3_1 _1688_ (.B(net155),
    .C(_0838_),
    .A(net226),
    .Y(_0839_));
 sg13g2_o21ai_1 _1689_ (.B1(_0834_),
    .Y(_0840_),
    .A1(\player_x[2] ),
    .A2(\player_x[1] ));
 sg13g2_nor2_1 _1690_ (.A(net342),
    .B(net286),
    .Y(_0841_));
 sg13g2_a21oi_1 _1691_ (.A1(_0344_),
    .A2(_0840_),
    .Y(_0842_),
    .B1(inp_left_prev));
 sg13g2_nand3_1 _1692_ (.B(net155),
    .C(_0842_),
    .A(net227),
    .Y(_0843_));
 sg13g2_a21oi_2 _1693_ (.B1(_0351_),
    .Y(_0844_),
    .A2(_0843_),
    .A1(_0839_));
 sg13g2_nand2_1 _1694_ (.Y(_0845_),
    .A(net202),
    .B(_0844_));
 sg13g2_nand2_1 _1695_ (.Y(_0846_),
    .A(net286),
    .B(_0369_));
 sg13g2_a22oi_1 _1696_ (.Y(_0034_),
    .B1(_0845_),
    .B2(_0846_),
    .A2(_0844_),
    .A1(net286));
 sg13g2_nand2_1 _1697_ (.Y(_0847_),
    .A(net342),
    .B(_0369_));
 sg13g2_nor2_1 _1698_ (.A(_0835_),
    .B(_0841_),
    .Y(_0848_));
 sg13g2_xnor2_1 _1699_ (.Y(_0849_),
    .A(_0839_),
    .B(_0848_));
 sg13g2_a22oi_1 _1700_ (.Y(_0035_),
    .B1(_0849_),
    .B2(_0844_),
    .A2(_0847_),
    .A1(_0845_));
 sg13g2_nand2_1 _1701_ (.Y(_0850_),
    .A(net350),
    .B(_0369_));
 sg13g2_mux2_1 _1702_ (.A0(_0835_),
    .A1(_0841_),
    .S(_0839_),
    .X(_0851_));
 sg13g2_xnor2_1 _1703_ (.Y(_0852_),
    .A(net350),
    .B(_0851_));
 sg13g2_a22oi_1 _1704_ (.Y(_0036_),
    .B1(_0852_),
    .B2(_0844_),
    .A2(_0850_),
    .A1(_0845_));
 sg13g2_and2_1 _1705_ (.A(\player_y[1] ),
    .B(net173),
    .X(_0853_));
 sg13g2_xnor2_1 _1706_ (.Y(_0854_),
    .A(\maze_seed[2] ),
    .B(\player_y[2] ));
 sg13g2_xnor2_1 _1707_ (.Y(_0855_),
    .A(_0853_),
    .B(_0854_));
 sg13g2_inv_1 _1708_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_xnor2_1 _1709_ (.Y(_0857_),
    .A(\player_x[1] ),
    .B(net173));
 sg13g2_xnor2_1 _1710_ (.Y(_0858_),
    .A(_0318_),
    .B(_0857_));
 sg13g2_xnor2_1 _1711_ (.Y(_0859_),
    .A(\player_x[2] ),
    .B(\player_y[1] ));
 sg13g2_xnor2_1 _1712_ (.Y(_0860_),
    .A(\maze_seed[1] ),
    .B(_0859_));
 sg13g2_xnor2_1 _1713_ (.Y(_0861_),
    .A(\player_y[0] ),
    .B(_0860_));
 sg13g2_o21ai_1 _1714_ (.B1(net184),
    .Y(_0862_),
    .A1(_0856_),
    .A2(_0858_));
 sg13g2_mux2_1 _1715_ (.A0(_0862_),
    .A1(_0858_),
    .S(_0861_),
    .X(_0863_));
 sg13g2_nor3_1 _1716_ (.A(_0314_),
    .B(_0856_),
    .C(_0863_),
    .Y(_0864_));
 sg13g2_a21oi_1 _1717_ (.A1(_0856_),
    .A2(_0863_),
    .Y(_0865_),
    .B1(_0864_));
 sg13g2_nor2_1 _1718_ (.A(net184),
    .B(_0858_),
    .Y(_0866_));
 sg13g2_xnor2_1 _1719_ (.Y(_0867_),
    .A(\maze_seed[4] ),
    .B(\player_x[0] ));
 sg13g2_xnor2_1 _1720_ (.Y(_0868_),
    .A(_0860_),
    .B(_0867_));
 sg13g2_xnor2_1 _1721_ (.Y(_0869_),
    .A(_0866_),
    .B(_0868_));
 sg13g2_nand2_1 _1722_ (.Y(_0870_),
    .A(\player_y[2] ),
    .B(_0853_));
 sg13g2_a21oi_1 _1723_ (.A1(\player_y[2] ),
    .A2(_0853_),
    .Y(_0871_),
    .B1(inp_down_prev));
 sg13g2_xnor2_1 _1724_ (.Y(_0872_),
    .A(_0865_),
    .B(_0869_));
 sg13g2_and4_1 _1725_ (.A(\gamepad.decoder.data_reg[6] ),
    .B(net155),
    .C(_0871_),
    .D(_0872_),
    .X(_0873_));
 sg13g2_xor2_1 _1726_ (.B(_0861_),
    .A(\maze_seed[4] ),
    .X(_0874_));
 sg13g2_and3_1 _1727_ (.X(_0875_),
    .A(net184),
    .B(_0854_),
    .C(_0858_));
 sg13g2_nor2_1 _1728_ (.A(net184),
    .B(_0854_),
    .Y(_0876_));
 sg13g2_nor2_1 _1729_ (.A(_0860_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_nor3_1 _1730_ (.A(_0866_),
    .B(_0875_),
    .C(_0877_),
    .Y(_0878_));
 sg13g2_a21oi_1 _1731_ (.A1(net184),
    .A2(_0858_),
    .Y(_0879_),
    .B1(_0854_));
 sg13g2_or2_1 _1732_ (.X(_0880_),
    .B(_0879_),
    .A(_0875_));
 sg13g2_nand2_1 _1733_ (.Y(_0881_),
    .A(net260),
    .B(net155));
 sg13g2_nor3_1 _1734_ (.A(inp_up_prev),
    .B(_0834_),
    .C(_0881_),
    .Y(_0882_));
 sg13g2_xnor2_1 _1735_ (.Y(_0883_),
    .A(_0874_),
    .B(_0880_));
 sg13g2_xnor2_1 _1736_ (.Y(_0884_),
    .A(_0344_),
    .B(_0878_));
 sg13g2_xnor2_1 _1737_ (.Y(_0885_),
    .A(_0883_),
    .B(_0884_));
 sg13g2_a21oi_1 _1738_ (.A1(_0882_),
    .A2(_0885_),
    .Y(_0886_),
    .B1(_0873_));
 sg13g2_nor2_2 _1739_ (.A(_0351_),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_a21oi_1 _1740_ (.A1(net173),
    .A2(net148),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_a21oi_1 _1741_ (.A1(net173),
    .A2(_0887_),
    .Y(_0889_),
    .B1(net193));
 sg13g2_nor2b_1 _1742_ (.A(net385),
    .B_N(_0889_),
    .Y(_0037_));
 sg13g2_a21oi_1 _1743_ (.A1(net371),
    .A2(net148),
    .Y(_0890_),
    .B1(_0887_));
 sg13g2_xor2_1 _1744_ (.B(net173),
    .A(\player_y[1] ),
    .X(_0891_));
 sg13g2_xnor2_1 _1745_ (.Y(_0892_),
    .A(_0873_),
    .B(_0891_));
 sg13g2_nor3_1 _1746_ (.A(_0351_),
    .B(_0886_),
    .C(_0892_),
    .Y(_0893_));
 sg13g2_nor3_1 _1747_ (.A(net193),
    .B(net372),
    .C(_0893_),
    .Y(_0038_));
 sg13g2_nor2_1 _1748_ (.A(\player_y[2] ),
    .B(_0853_),
    .Y(_0894_));
 sg13g2_o21ai_1 _1749_ (.B1(\player_y[2] ),
    .Y(_0895_),
    .A1(\player_y[1] ),
    .A2(net173));
 sg13g2_nor2b_1 _1750_ (.A(_0834_),
    .B_N(_0895_),
    .Y(_0896_));
 sg13g2_mux2_1 _1751_ (.A0(_0896_),
    .A1(_0894_),
    .S(_0873_),
    .X(_0897_));
 sg13g2_and2_1 _1752_ (.A(_0887_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_a21oi_1 _1753_ (.A1(net367),
    .A2(net148),
    .Y(_0899_),
    .B1(_0887_));
 sg13g2_nor3_1 _1754_ (.A(net193),
    .B(_0898_),
    .C(net368),
    .Y(_0039_));
 sg13g2_nand2_1 _1755_ (.Y(_0900_),
    .A(net172),
    .B(net146));
 sg13g2_nand2_2 _1756_ (.Y(_0901_),
    .A(_0445_),
    .B(_0481_));
 sg13g2_a21oi_1 _1757_ (.A1(_0900_),
    .A2(_0901_),
    .Y(_0902_),
    .B1(_0504_));
 sg13g2_o21ai_1 _1758_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0332_),
    .A2(_0901_));
 sg13g2_nand2_1 _1759_ (.Y(_0904_),
    .A(_0330_),
    .B(_0333_));
 sg13g2_nor2_1 _1760_ (.A(net185),
    .B(net359),
    .Y(_0905_));
 sg13g2_nor3_1 _1761_ (.A(\solver_r_dir[3] ),
    .B(\solver_r_dir[2] ),
    .C(_0904_),
    .Y(_0906_));
 sg13g2_or2_1 _1762_ (.X(_0907_),
    .B(_0906_),
    .A(net153));
 sg13g2_nand3_1 _1763_ (.B(net146),
    .C(_0464_),
    .A(net172),
    .Y(_0908_));
 sg13g2_nor2_1 _1764_ (.A(net185),
    .B(_0490_),
    .Y(_0909_));
 sg13g2_o21ai_1 _1765_ (.B1(_0908_),
    .Y(_0910_),
    .A1(net172),
    .A2(_0909_));
 sg13g2_o21ai_1 _1766_ (.B1(_0905_),
    .Y(_0911_),
    .A1(net401),
    .A2(_0507_));
 sg13g2_a21oi_1 _1767_ (.A1(_0910_),
    .A2(_0911_),
    .Y(_0912_),
    .B1(net150));
 sg13g2_a221oi_1 _1768_ (.B2(_0903_),
    .C1(net197),
    .B1(_0912_),
    .A1(_0900_),
    .Y(_0040_),
    .A2(net150));
 sg13g2_xor2_1 _1769_ (.B(net403),
    .A(\solver_r_x[1] ),
    .X(_0913_));
 sg13g2_nand2_1 _1770_ (.Y(_0914_),
    .A(net392),
    .B(net146));
 sg13g2_a21oi_1 _1771_ (.A1(_0901_),
    .A2(_0914_),
    .Y(_0915_),
    .B1(_0504_));
 sg13g2_o21ai_1 _1772_ (.B1(_0915_),
    .Y(_0916_),
    .A1(_0901_),
    .A2(_0913_));
 sg13g2_or2_1 _1773_ (.X(_0917_),
    .B(_0914_),
    .A(_0512_));
 sg13g2_o21ai_1 _1774_ (.B1(_0913_),
    .Y(_0918_),
    .A1(_0330_),
    .A2(_0446_));
 sg13g2_o21ai_1 _1775_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0512_),
    .A2(_0913_));
 sg13g2_nor2_1 _1776_ (.A(\solver_r_dir[3] ),
    .B(_0913_),
    .Y(_0920_));
 sg13g2_a221oi_1 _1777_ (.B2(_0445_),
    .C1(_0905_),
    .B1(_0920_),
    .A1(_0917_),
    .Y(_0921_),
    .A2(_0919_));
 sg13g2_nor2_1 _1778_ (.A(_0507_),
    .B(_0913_),
    .Y(_0922_));
 sg13g2_nor3_1 _1779_ (.A(net150),
    .B(_0921_),
    .C(_0922_),
    .Y(_0923_));
 sg13g2_a221oi_1 _1780_ (.B2(_0923_),
    .C1(net197),
    .B1(_0916_),
    .A1(net150),
    .Y(_0041_),
    .A2(_0914_));
 sg13g2_nand2_1 _1781_ (.Y(_0924_),
    .A(net383),
    .B(net146));
 sg13g2_or3_1 _1782_ (.A(\solver_r_x[2] ),
    .B(_0441_),
    .C(_0444_),
    .X(_0925_));
 sg13g2_nand2b_1 _1783_ (.Y(_0926_),
    .B(_0481_),
    .A_N(_0925_));
 sg13g2_a21oi_1 _1784_ (.A1(_0901_),
    .A2(_0924_),
    .Y(_0927_),
    .B1(_0504_));
 sg13g2_nand2_1 _1785_ (.Y(_0928_),
    .A(_0926_),
    .B(_0927_));
 sg13g2_nor2b_1 _1786_ (.A(_0512_),
    .B_N(_0924_),
    .Y(_0929_));
 sg13g2_nand2_1 _1787_ (.Y(_0930_),
    .A(net185),
    .B(_0925_));
 sg13g2_o21ai_1 _1788_ (.B1(\solver_r_x[2] ),
    .Y(_0931_),
    .A1(\solver_r_x[1] ),
    .A2(\solver_r_x[0] ));
 sg13g2_a221oi_1 _1789_ (.B2(_0512_),
    .C1(_0929_),
    .B1(_0931_),
    .A1(_0334_),
    .Y(_0932_),
    .A2(_0930_));
 sg13g2_nand3_1 _1790_ (.B(_0445_),
    .C(_0925_),
    .A(net185),
    .Y(_0933_));
 sg13g2_o21ai_1 _1791_ (.B1(_0933_),
    .Y(_0934_),
    .A1(_0507_),
    .A2(_0931_));
 sg13g2_nor3_1 _1792_ (.A(net150),
    .B(_0932_),
    .C(_0934_),
    .Y(_0935_));
 sg13g2_a221oi_1 _1793_ (.B2(_0935_),
    .C1(net197),
    .B1(_0928_),
    .A1(net150),
    .Y(_0042_),
    .A2(_0924_));
 sg13g2_nand3_1 _1794_ (.B(_0480_),
    .C(_0491_),
    .A(_0469_),
    .Y(_0936_));
 sg13g2_nor2_1 _1795_ (.A(net320),
    .B(_0493_),
    .Y(_0937_));
 sg13g2_o21ai_1 _1796_ (.B1(_0936_),
    .Y(_0938_),
    .A1(net320),
    .A2(_0493_));
 sg13g2_o21ai_1 _1797_ (.B1(_0938_),
    .Y(_0939_),
    .A1(_0465_),
    .A2(_0508_));
 sg13g2_or2_1 _1798_ (.X(_0940_),
    .B(_0939_),
    .A(net150));
 sg13g2_nand3_1 _1799_ (.B(_0369_),
    .C(_0940_),
    .A(net171),
    .Y(_0941_));
 sg13g2_a21oi_1 _1800_ (.A1(_0494_),
    .A2(_0504_),
    .Y(_0942_),
    .B1(_0481_));
 sg13g2_a221oi_1 _1801_ (.B2(_0904_),
    .C1(_0942_),
    .B1(_0465_),
    .A1(\solver_r_dir[3] ),
    .Y(_0943_),
    .A2(_0464_));
 sg13g2_nand2b_1 _1802_ (.Y(_0944_),
    .B(net151),
    .A_N(net345));
 sg13g2_o21ai_1 _1803_ (.B1(_0941_),
    .Y(_0043_),
    .A1(_0943_),
    .A2(_0944_));
 sg13g2_nand2_1 _1804_ (.Y(_0945_),
    .A(net374),
    .B(net146));
 sg13g2_nand2b_1 _1805_ (.Y(_0946_),
    .B(_0939_),
    .A_N(_0945_));
 sg13g2_nand2_1 _1806_ (.Y(_0947_),
    .A(_0334_),
    .B(_0509_));
 sg13g2_nor3_1 _1807_ (.A(_0443_),
    .B(_0463_),
    .C(_0470_),
    .Y(_0948_));
 sg13g2_nand2_1 _1808_ (.Y(_0949_),
    .A(net338),
    .B(_0480_));
 sg13g2_o21ai_1 _1809_ (.B1(_0949_),
    .Y(_0950_),
    .A1(_0936_),
    .A2(_0937_));
 sg13g2_a221oi_1 _1810_ (.B2(_0470_),
    .C1(net150),
    .B1(_0950_),
    .A1(_0947_),
    .Y(_0951_),
    .A2(_0948_));
 sg13g2_a221oi_1 _1811_ (.B2(_0951_),
    .C1(net197),
    .B1(_0946_),
    .A1(_0907_),
    .Y(_0044_),
    .A2(_0945_));
 sg13g2_o21ai_1 _1812_ (.B1(\solver_r_y[2] ),
    .Y(_0952_),
    .A1(\solver_r_y[0] ),
    .A2(\solver_r_y[1] ));
 sg13g2_nor2_1 _1813_ (.A(_0463_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_a221oi_1 _1814_ (.B2(_0504_),
    .C1(_0481_),
    .B1(_0495_),
    .A1(_0331_),
    .Y(_0954_),
    .A2(_0468_));
 sg13g2_a21oi_1 _1815_ (.A1(_0947_),
    .A2(_0953_),
    .Y(_0955_),
    .B1(_0954_));
 sg13g2_nand3_1 _1816_ (.B(net146),
    .C(_0940_),
    .A(net402),
    .Y(_0956_));
 sg13g2_o21ai_1 _1817_ (.B1(_0956_),
    .Y(_0957_),
    .A1(_0907_),
    .A2(_0955_));
 sg13g2_and2_1 _1818_ (.A(net204),
    .B(_0957_),
    .X(_0045_));
 sg13g2_nand2_1 _1819_ (.Y(_0958_),
    .A(net379),
    .B(net147));
 sg13g2_a21oi_1 _1820_ (.A1(_0326_),
    .A2(net188),
    .Y(_0959_),
    .B1(net189));
 sg13g2_a221oi_1 _1821_ (.B2(_0958_),
    .C1(_0959_),
    .B1(_0425_),
    .A1(net379),
    .Y(_0960_),
    .A2(_0416_));
 sg13g2_and2_1 _1822_ (.A(_0396_),
    .B(_0958_),
    .X(_0961_));
 sg13g2_nand2_1 _1823_ (.Y(_0962_),
    .A(_0327_),
    .B(_0417_));
 sg13g2_nor2_1 _1824_ (.A(\solver_l_x[0] ),
    .B(_0373_),
    .Y(_0963_));
 sg13g2_o21ai_1 _1825_ (.B1(_0962_),
    .Y(_0964_),
    .A1(_0396_),
    .A2(_0963_));
 sg13g2_nor4_1 _1826_ (.A(net188),
    .B(net186),
    .C(net187),
    .D(net189),
    .Y(_0965_));
 sg13g2_nor2_1 _1827_ (.A(net154),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_or2_1 _1828_ (.X(_0967_),
    .B(_0965_),
    .A(net154));
 sg13g2_a21oi_1 _1829_ (.A1(_0326_),
    .A2(net187),
    .Y(_0968_),
    .B1(_0967_));
 sg13g2_o21ai_1 _1830_ (.B1(_0968_),
    .Y(_0969_),
    .A1(_0961_),
    .A2(_0964_));
 sg13g2_o21ai_1 _1831_ (.B1(net204),
    .Y(_0970_),
    .A1(_0960_),
    .A2(_0969_));
 sg13g2_a21oi_1 _1832_ (.A1(_0958_),
    .A2(_0967_),
    .Y(_0046_),
    .B1(_0970_));
 sg13g2_nor2_1 _1833_ (.A(\solver_l_x[0] ),
    .B(\solver_l_x[1] ),
    .Y(_0971_));
 sg13g2_nor2_2 _1834_ (.A(_0414_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_or2_1 _1835_ (.X(_0973_),
    .B(_0429_),
    .A(net189));
 sg13g2_nand2_1 _1836_ (.Y(_0974_),
    .A(net381),
    .B(net147));
 sg13g2_o21ai_1 _1837_ (.B1(_0973_),
    .Y(_0975_),
    .A1(_0425_),
    .A2(_0972_));
 sg13g2_a21oi_1 _1838_ (.A1(_0425_),
    .A2(_0974_),
    .Y(_0976_),
    .B1(_0975_));
 sg13g2_nand3_1 _1839_ (.B(net143),
    .C(_0972_),
    .A(_0374_),
    .Y(_0128_));
 sg13g2_a21oi_1 _1840_ (.A1(net187),
    .A2(_0972_),
    .Y(_0129_),
    .B1(_0962_));
 sg13g2_a21oi_1 _1841_ (.A1(_0420_),
    .A2(_0974_),
    .Y(_0130_),
    .B1(_0129_));
 sg13g2_nand2_1 _1842_ (.Y(_0131_),
    .A(_0128_),
    .B(_0130_));
 sg13g2_nand3_1 _1843_ (.B(_0416_),
    .C(_0972_),
    .A(net187),
    .Y(_0132_));
 sg13g2_o21ai_1 _1844_ (.B1(_0132_),
    .Y(_0133_),
    .A1(_0376_),
    .A2(_0972_));
 sg13g2_nor3_1 _1845_ (.A(_0967_),
    .B(_0976_),
    .C(_0133_),
    .Y(_0134_));
 sg13g2_a221oi_1 _1846_ (.B2(_0134_),
    .C1(net197),
    .B1(_0131_),
    .A1(_0967_),
    .Y(_0047_),
    .A2(_0974_));
 sg13g2_nor2b_2 _1847_ (.A(_0971_),
    .B_N(net390),
    .Y(_0135_));
 sg13g2_nor3_1 _1848_ (.A(\solver_l_x[2] ),
    .B(_0414_),
    .C(_0415_),
    .Y(_0136_));
 sg13g2_nand2b_1 _1849_ (.Y(_0137_),
    .B(\solver_l_dir[2] ),
    .A_N(_0136_));
 sg13g2_nand2_1 _1850_ (.Y(_0138_),
    .A(net390),
    .B(net147));
 sg13g2_a22oi_1 _1851_ (.Y(_0139_),
    .B1(_0138_),
    .B2(_0420_),
    .A2(_0137_),
    .A1(_0327_));
 sg13g2_o21ai_1 _1852_ (.B1(_0139_),
    .Y(_0140_),
    .A1(_0420_),
    .A2(_0135_));
 sg13g2_a21oi_1 _1853_ (.A1(net188),
    .A2(_0135_),
    .Y(_0141_),
    .B1(_0973_));
 sg13g2_a221oi_1 _1854_ (.B2(_0425_),
    .C1(_0141_),
    .B1(_0138_),
    .A1(_0410_),
    .Y(_0142_),
    .A2(_0136_));
 sg13g2_nand2_1 _1855_ (.Y(_0143_),
    .A(_0375_),
    .B(_0135_));
 sg13g2_o21ai_1 _1856_ (.B1(_0143_),
    .Y(_0144_),
    .A1(_0422_),
    .A2(_0136_));
 sg13g2_nor3_1 _1857_ (.A(_0967_),
    .B(_0142_),
    .C(_0144_),
    .Y(_0145_));
 sg13g2_a221oi_1 _1858_ (.B2(_0145_),
    .C1(net198),
    .B1(_0140_),
    .A1(_0967_),
    .Y(_0048_),
    .A2(_0138_));
 sg13g2_nand2_1 _1859_ (.Y(_0146_),
    .A(net231),
    .B(net155));
 sg13g2_nor3_1 _1860_ (.A(net307),
    .B(_0351_),
    .C(_0146_),
    .Y(_0147_));
 sg13g2_a21oi_1 _1861_ (.A1(solvers_active),
    .A2(_0365_),
    .Y(_0148_),
    .B1(_0147_));
 sg13g2_and2_1 _1862_ (.A(solvers_active),
    .B(_0147_),
    .X(_0149_));
 sg13g2_nor4_1 _1863_ (.A(net192),
    .B(_0361_),
    .C(net308),
    .D(_0149_),
    .Y(_0049_));
 sg13g2_nand2b_1 _1864_ (.Y(_0150_),
    .B(_0396_),
    .A_N(_0416_));
 sg13g2_nor2_1 _1865_ (.A(\solver_l_x[0] ),
    .B(_0410_),
    .Y(_0151_));
 sg13g2_a21oi_1 _1866_ (.A1(net186),
    .A2(net143),
    .Y(_0152_),
    .B1(net188));
 sg13g2_o21ai_1 _1867_ (.B1(_0966_),
    .Y(_0153_),
    .A1(_0151_),
    .A2(_0152_));
 sg13g2_a21oi_1 _1868_ (.A1(_0412_),
    .A2(_0150_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_nor2b_1 _1869_ (.A(_0154_),
    .B_N(net147),
    .Y(_0155_));
 sg13g2_inv_1 _1870_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_o21ai_1 _1871_ (.B1(_0151_),
    .Y(_0157_),
    .A1(net188),
    .A2(net186));
 sg13g2_a21oi_1 _1872_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0158_),
    .B1(_0150_));
 sg13g2_a221oi_1 _1873_ (.B2(net189),
    .C1(_0158_),
    .B1(_0409_),
    .A1(net186),
    .Y(_0159_),
    .A2(_0396_));
 sg13g2_a21oi_1 _1874_ (.A1(_0157_),
    .A2(_0159_),
    .Y(_0160_),
    .B1(_0967_));
 sg13g2_o21ai_1 _1875_ (.B1(net204),
    .Y(_0161_),
    .A1(net170),
    .A2(_0160_));
 sg13g2_a21oi_1 _1876_ (.A1(net170),
    .A2(_0156_),
    .Y(_0050_),
    .B1(_0161_));
 sg13g2_nand2b_1 _1877_ (.Y(_0162_),
    .B(_0151_),
    .A_N(_0152_));
 sg13g2_xor2_1 _1878_ (.B(net360),
    .A(\solver_l_y[0] ),
    .X(_0163_));
 sg13g2_a21oi_1 _1879_ (.A1(net189),
    .A2(_0409_),
    .Y(_0164_),
    .B1(_0163_));
 sg13g2_nor2_1 _1880_ (.A(_0411_),
    .B(_0150_),
    .Y(_0165_));
 sg13g2_a21oi_1 _1881_ (.A1(net186),
    .A2(_0395_),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_a221oi_1 _1882_ (.B2(_0163_),
    .C1(_0967_),
    .B1(_0166_),
    .A1(_0162_),
    .Y(_0167_),
    .A2(_0164_));
 sg13g2_a21oi_1 _1883_ (.A1(net360),
    .A2(_0155_),
    .Y(_0168_),
    .B1(_0167_));
 sg13g2_nor2_1 _1884_ (.A(net198),
    .B(net361),
    .Y(_0051_));
 sg13g2_o21ai_1 _1885_ (.B1(\solver_l_y[2] ),
    .Y(_0169_),
    .A1(\solver_l_y[0] ),
    .A2(\solver_l_y[1] ));
 sg13g2_nor2_1 _1886_ (.A(_0408_),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_o21ai_1 _1887_ (.B1(_0170_),
    .Y(_0171_),
    .A1(_0421_),
    .A2(_0973_));
 sg13g2_nand2_1 _1888_ (.Y(_0172_),
    .A(_0417_),
    .B(_0499_));
 sg13g2_o21ai_1 _1889_ (.B1(_0172_),
    .Y(_0173_),
    .A1(net376),
    .A2(_0378_));
 sg13g2_o21ai_1 _1890_ (.B1(_0171_),
    .Y(_0174_),
    .A1(net143),
    .A2(_0173_));
 sg13g2_a22oi_1 _1891_ (.Y(_0175_),
    .B1(_0174_),
    .B2(_0966_),
    .A2(_0155_),
    .A1(net376));
 sg13g2_nor2_1 _1892_ (.A(net197),
    .B(_0175_),
    .Y(_0052_));
 sg13g2_nor3_1 _1893_ (.A(_0351_),
    .B(_0836_),
    .C(_0870_),
    .Y(_0176_));
 sg13g2_a21oi_1 _1894_ (.A1(net297),
    .A2(net148),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_nor2_1 _1895_ (.A(net193),
    .B(net298),
    .Y(_0053_));
 sg13g2_nor2_1 _1896_ (.A(_0442_),
    .B(_0469_),
    .Y(_0178_));
 sg13g2_a22oi_1 _1897_ (.Y(_0179_),
    .B1(_0178_),
    .B2(_0352_),
    .A2(net148),
    .A1(net315));
 sg13g2_nor2_1 _1898_ (.A(net196),
    .B(net316),
    .Y(_0054_));
 sg13g2_and2_1 _1899_ (.A(net369),
    .B(net156),
    .X(_0180_));
 sg13g2_nand3b_1 _1900_ (.B(_0180_),
    .C(generating),
    .Y(_0181_),
    .A_N(net396));
 sg13g2_inv_1 _1901_ (.Y(_0182_),
    .A(_0181_));
 sg13g2_nand3_1 _1902_ (.B(\gen_row[1] ),
    .C(\gen_row[0] ),
    .A(net324),
    .Y(_0183_));
 sg13g2_or2_1 _1903_ (.X(_0184_),
    .B(net218),
    .A(net216));
 sg13g2_a21oi_1 _1904_ (.A1(net224),
    .A2(\gen_frame_count[0] ),
    .Y(_0185_),
    .B1(_0184_));
 sg13g2_nand2_2 _1905_ (.Y(_0186_),
    .A(generating),
    .B(net164));
 sg13g2_nand2_1 _1906_ (.Y(_0187_),
    .A(_0181_),
    .B(_0186_));
 sg13g2_o21ai_1 _1907_ (.B1(_0187_),
    .Y(_0188_),
    .A1(_0183_),
    .A2(_0185_));
 sg13g2_nand2_1 _1908_ (.Y(_0189_),
    .A(_0365_),
    .B(_0188_));
 sg13g2_nor3_1 _1909_ (.A(_0312_),
    .B(net165),
    .C(_0364_),
    .Y(_0190_));
 sg13g2_o21ai_1 _1910_ (.B1(net397),
    .Y(_0191_),
    .A1(_0189_),
    .A2(_0190_));
 sg13g2_nand2_1 _1911_ (.Y(_0055_),
    .A(net200),
    .B(net398));
 sg13g2_nand4_1 _1912_ (.B(_0365_),
    .C(_0181_),
    .A(generating),
    .Y(_0192_),
    .D(_0185_));
 sg13g2_and2_1 _1913_ (.A(_0189_),
    .B(_0192_),
    .X(_0193_));
 sg13g2_o21ai_1 _1914_ (.B1(_0181_),
    .Y(_0194_),
    .A1(net365),
    .A2(_0364_));
 sg13g2_inv_1 _1915_ (.Y(_0195_),
    .A(_0194_));
 sg13g2_o21ai_1 _1916_ (.B1(net201),
    .Y(_0196_),
    .A1(net365),
    .A2(_0193_));
 sg13g2_a21oi_1 _1917_ (.A1(_0193_),
    .A2(_0195_),
    .Y(_0056_),
    .B1(_0196_));
 sg13g2_xor2_1 _1918_ (.B(\gen_row[0] ),
    .A(net363),
    .X(_0197_));
 sg13g2_a21oi_1 _1919_ (.A1(_0365_),
    .A2(_0197_),
    .Y(_0198_),
    .B1(_0182_));
 sg13g2_o21ai_1 _1920_ (.B1(net201),
    .Y(_0199_),
    .A1(net363),
    .A2(_0193_));
 sg13g2_a21oi_1 _1921_ (.A1(_0193_),
    .A2(_0198_),
    .Y(_0057_),
    .B1(_0199_));
 sg13g2_a21o_1 _1922_ (.A2(\gen_row[0] ),
    .A1(\gen_row[1] ),
    .B1(net324),
    .X(_0200_));
 sg13g2_and2_1 _1923_ (.A(_0183_),
    .B(_0200_),
    .X(_0201_));
 sg13g2_a21oi_1 _1924_ (.A1(_0365_),
    .A2(_0201_),
    .Y(_0202_),
    .B1(_0182_));
 sg13g2_o21ai_1 _1925_ (.B1(net201),
    .Y(_0203_),
    .A1(net324),
    .A2(_0193_));
 sg13g2_a21oi_1 _1926_ (.A1(_0193_),
    .A2(_0202_),
    .Y(_0058_),
    .B1(_0203_));
 sg13g2_nor2_1 _1927_ (.A(_0184_),
    .B(_0186_),
    .Y(_0204_));
 sg13g2_nand3_1 _1928_ (.B(generating),
    .C(net164),
    .A(net322),
    .Y(_0205_));
 sg13g2_o21ai_1 _1929_ (.B1(_0205_),
    .Y(_0206_),
    .A1(net322),
    .A2(_0204_));
 sg13g2_nor2_1 _1930_ (.A(_0367_),
    .B(net323),
    .Y(_0059_));
 sg13g2_o21ai_1 _1931_ (.B1(net149),
    .Y(_0207_),
    .A1(_0185_),
    .A2(_0186_));
 sg13g2_a21oi_1 _1932_ (.A1(_0311_),
    .A2(_0205_),
    .Y(_0060_),
    .B1(_0207_));
 sg13g2_and3_1 _1933_ (.X(_0061_),
    .A(net218),
    .B(net149),
    .C(_0186_));
 sg13g2_and3_1 _1934_ (.X(_0062_),
    .A(net216),
    .B(net149),
    .C(_0186_));
 sg13g2_nand2_1 _1935_ (.Y(_0208_),
    .A(net263),
    .B(net156));
 sg13g2_nor3_1 _1936_ (.A(\solver_speed[3] ),
    .B(\solver_speed[2] ),
    .C(\solver_speed[1] ),
    .Y(_0209_));
 sg13g2_nor3_2 _1937_ (.A(inp_r_prev),
    .B(_0208_),
    .C(_0209_),
    .Y(_0210_));
 sg13g2_and2_1 _1938_ (.A(net362),
    .B(net156),
    .X(_0211_));
 sg13g2_nand3_1 _1939_ (.B(net354),
    .C(net348),
    .A(net328),
    .Y(_0212_));
 sg13g2_nor2b_1 _1940_ (.A(inp_l_prev),
    .B_N(_0211_),
    .Y(_0213_));
 sg13g2_o21ai_1 _1941_ (.B1(_0213_),
    .Y(_0214_),
    .A1(_0309_),
    .A2(_0212_));
 sg13g2_nor2b_2 _1942_ (.A(_0210_),
    .B_N(_0214_),
    .Y(_0215_));
 sg13g2_o21ai_1 _1943_ (.B1(net201),
    .Y(_0216_),
    .A1(_0310_),
    .A2(_0215_));
 sg13g2_a21oi_1 _1944_ (.A1(_0310_),
    .A2(_0215_),
    .Y(_0063_),
    .B1(_0216_));
 sg13g2_xnor2_1 _1945_ (.Y(_0217_),
    .A(\solver_speed[1] ),
    .B(net348));
 sg13g2_inv_1 _1946_ (.Y(_0218_),
    .A(_0217_));
 sg13g2_nand2b_1 _1947_ (.Y(_0219_),
    .B(_0217_),
    .A_N(_0210_));
 sg13g2_o21ai_1 _1948_ (.B1(_0218_),
    .Y(_0220_),
    .A1(_0210_),
    .A2(_0214_));
 sg13g2_a22oi_1 _1949_ (.Y(_0221_),
    .B1(_0219_),
    .B2(_0220_),
    .A2(_0215_),
    .A1(net354));
 sg13g2_nor2_1 _1950_ (.A(net196),
    .B(net355),
    .Y(_0064_));
 sg13g2_xnor2_1 _1951_ (.Y(_0222_),
    .A(_0783_),
    .B(_0219_));
 sg13g2_a21oi_1 _1952_ (.A1(net328),
    .A2(_0215_),
    .Y(_0223_),
    .B1(net196));
 sg13g2_o21ai_1 _1953_ (.B1(net329),
    .Y(_0065_),
    .A1(_0215_),
    .A2(_0222_));
 sg13g2_nor2_1 _1954_ (.A(net386),
    .B(_0210_),
    .Y(_0224_));
 sg13g2_o21ai_1 _1955_ (.B1(net387),
    .Y(_0225_),
    .A1(_0212_),
    .A2(_0214_));
 sg13g2_a21oi_1 _1956_ (.A1(_0778_),
    .A2(_0210_),
    .Y(_0226_),
    .B1(net196));
 sg13g2_and2_1 _1957_ (.A(net388),
    .B(_0226_),
    .X(_0066_));
 sg13g2_nor4_1 _1958_ (.A(\solver_frame_count[3] ),
    .B(\solver_frame_count[2] ),
    .C(net282),
    .D(_0310_),
    .Y(_0227_));
 sg13g2_nor3_1 _1959_ (.A(net302),
    .B(net163),
    .C(_0227_),
    .Y(_0228_));
 sg13g2_a21oi_1 _1960_ (.A1(net302),
    .A2(net163),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_nor2_1 _1961_ (.A(net194),
    .B(net303),
    .Y(_0067_));
 sg13g2_o21ai_1 _1962_ (.B1(net282),
    .Y(_0230_),
    .A1(\solver_frame_count[0] ),
    .A2(net163));
 sg13g2_a221oi_1 _1963_ (.B2(_0347_),
    .C1(net194),
    .B1(net283),
    .A1(_0348_),
    .Y(_0068_),
    .A2(_0218_));
 sg13g2_nor2b_1 _1964_ (.A(net304),
    .B_N(_0783_),
    .Y(_0231_));
 sg13g2_nor3_1 _1965_ (.A(net312),
    .B(_0347_),
    .C(_0231_),
    .Y(_0232_));
 sg13g2_a21oi_1 _1966_ (.A1(net312),
    .A2(_0347_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_nor2_1 _1967_ (.A(net195),
    .B(_0233_),
    .Y(_0069_));
 sg13g2_o21ai_1 _1968_ (.B1(net304),
    .Y(_0234_),
    .A1(\solver_frame_count[2] ),
    .A2(_0347_));
 sg13g2_nand2b_1 _1969_ (.Y(_0235_),
    .B(_0348_),
    .A_N(_0778_));
 sg13g2_a21oi_1 _1970_ (.A1(net305),
    .A2(_0235_),
    .Y(_0070_),
    .B1(net199));
 sg13g2_nand2_1 _1971_ (.Y(_0236_),
    .A(net232),
    .B(net156));
 sg13g2_nor2_1 _1972_ (.A(inp_x_prev),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_o21ai_1 _1973_ (.B1(net356),
    .Y(_0238_),
    .A1(_0364_),
    .A2(_0237_));
 sg13g2_o21ai_1 _1974_ (.B1(net200),
    .Y(_0239_),
    .A1(net356),
    .A2(_0237_));
 sg13g2_nor2b_1 _1975_ (.A(net357),
    .B_N(_0238_),
    .Y(_0071_));
 sg13g2_nand2_1 _1976_ (.Y(_0240_),
    .A(single_step_mode),
    .B(solvers_active));
 sg13g2_nand2_1 _1977_ (.Y(_0241_),
    .A(step_requested),
    .B(_0240_));
 sg13g2_nor3_1 _1978_ (.A(_0367_),
    .B(_0237_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_and3_1 _1979_ (.X(_0083_),
    .A(net237),
    .B(net200),
    .C(net156));
 sg13g2_nor3_1 _1980_ (.A(net317),
    .B(_0351_),
    .C(_0240_),
    .Y(_0243_));
 sg13g2_a21o_1 _1981_ (.A2(net318),
    .A1(_0083_),
    .B1(_0242_),
    .X(_0072_));
 sg13g2_and4_1 _1982_ (.A(\solver_l_y[2] ),
    .B(\solver_l_x[2] ),
    .C(_0378_),
    .D(_0414_),
    .X(_0244_));
 sg13g2_a22oi_1 _1983_ (.Y(_0245_),
    .B1(_0244_),
    .B2(_0352_),
    .A2(net148),
    .A1(net310));
 sg13g2_nor2_1 _1984_ (.A(net196),
    .B(net311),
    .Y(_0073_));
 sg13g2_nor2_1 _1985_ (.A(net192),
    .B(_0881_),
    .Y(_0074_));
 sg13g2_and3_1 _1986_ (.X(_0075_),
    .A(net230),
    .B(net202),
    .C(net155));
 sg13g2_and3_1 _1987_ (.X(_0076_),
    .A(net227),
    .B(net202),
    .C(net155));
 sg13g2_and3_1 _1988_ (.X(_0077_),
    .A(net226),
    .B(net202),
    .C(net155));
 sg13g2_nor2_1 _1989_ (.A(net192),
    .B(_0146_),
    .Y(_0078_));
 sg13g2_nor2_1 _1990_ (.A(net192),
    .B(_0360_),
    .Y(_0079_));
 sg13g2_and2_1 _1991_ (.A(net202),
    .B(_0180_),
    .X(_0081_));
 sg13g2_nor2_1 _1992_ (.A(net195),
    .B(net233),
    .Y(_0082_));
 sg13g2_and2_1 _1993_ (.A(net200),
    .B(_0211_),
    .X(_0084_));
 sg13g2_nor2_1 _1994_ (.A(net195),
    .B(_0208_),
    .Y(_0085_));
 sg13g2_and2_1 _1995_ (.A(net203),
    .B(net1),
    .X(_0086_));
 sg13g2_and2_1 _1996_ (.A(net203),
    .B(net214),
    .X(_0087_));
 sg13g2_nand4_1 _1997_ (.B(\hvsync_gen.vpos[9] ),
    .C(_0739_),
    .A(_0338_),
    .Y(_0246_),
    .D(_0741_));
 sg13g2_nand3_1 _1998_ (.B(_0820_),
    .C(_0246_),
    .A(net203),
    .Y(_0247_));
 sg13g2_inv_2 _1999_ (.Y(_0248_),
    .A(_0247_));
 sg13g2_mux2_1 _2000_ (.A0(_0248_),
    .A1(net145),
    .S(net169),
    .X(_0088_));
 sg13g2_nand2_1 _2001_ (.Y(_0249_),
    .A(net168),
    .B(net145));
 sg13g2_xnor2_1 _2002_ (.Y(_0250_),
    .A(net169),
    .B(net340));
 sg13g2_o21ai_1 _2003_ (.B1(_0249_),
    .Y(_0089_),
    .A1(_0247_),
    .A2(net341));
 sg13g2_nand2_1 _2004_ (.Y(_0251_),
    .A(net326),
    .B(net145));
 sg13g2_nand3_1 _2005_ (.B(\ent_y[1] ),
    .C(\hvsync_gen.vpos[2] ),
    .A(net169),
    .Y(_0252_));
 sg13g2_xnor2_1 _2006_ (.Y(_0253_),
    .A(_0335_),
    .B(_0709_));
 sg13g2_o21ai_1 _2007_ (.B1(_0251_),
    .Y(_0090_),
    .A1(_0247_),
    .A2(_0253_));
 sg13g2_nand2_1 _2008_ (.Y(_0254_),
    .A(net295),
    .B(net145));
 sg13g2_or2_1 _2009_ (.X(_0255_),
    .B(_0252_),
    .A(_0336_));
 sg13g2_xnor2_1 _2010_ (.Y(_0256_),
    .A(_0336_),
    .B(_0252_));
 sg13g2_o21ai_1 _2011_ (.B1(_0254_),
    .Y(_0091_),
    .A1(_0247_),
    .A2(_0256_));
 sg13g2_nand2_1 _2012_ (.Y(_0257_),
    .A(net290),
    .B(net145));
 sg13g2_nor2_1 _2013_ (.A(_0337_),
    .B(_0255_),
    .Y(_0258_));
 sg13g2_xnor2_1 _2014_ (.Y(_0259_),
    .A(_0337_),
    .B(_0255_));
 sg13g2_o21ai_1 _2015_ (.B1(_0257_),
    .Y(_0092_),
    .A1(_0247_),
    .A2(_0259_));
 sg13g2_nand2_1 _2016_ (.Y(_0260_),
    .A(net167),
    .B(net145));
 sg13g2_xnor2_1 _2017_ (.Y(_0261_),
    .A(net167),
    .B(_0258_));
 sg13g2_o21ai_1 _2018_ (.B1(_0260_),
    .Y(_0093_),
    .A1(_0247_),
    .A2(_0261_));
 sg13g2_a21oi_1 _2019_ (.A1(net336),
    .A2(_0258_),
    .Y(_0262_),
    .B1(net344));
 sg13g2_and3_2 _2020_ (.X(_0263_),
    .A(net336),
    .B(\hvsync_gen.vpos[6] ),
    .C(_0258_));
 sg13g2_nor3_1 _2021_ (.A(_0247_),
    .B(_0262_),
    .C(_0263_),
    .Y(_0264_));
 sg13g2_a21o_1 _2022_ (.A2(_0821_),
    .A1(net344),
    .B1(_0264_),
    .X(_0094_));
 sg13g2_o21ai_1 _2023_ (.B1(_0248_),
    .Y(_0265_),
    .A1(net166),
    .A2(_0263_));
 sg13g2_a21oi_1 _2024_ (.A1(net166),
    .A2(_0263_),
    .Y(_0266_),
    .B1(_0265_));
 sg13g2_a21o_1 _2025_ (.A2(net145),
    .A1(net293),
    .B1(_0266_),
    .X(_0095_));
 sg13g2_nand2b_1 _2026_ (.Y(_0267_),
    .B(_0263_),
    .A_N(_0516_));
 sg13g2_nand2_1 _2027_ (.Y(_0268_),
    .A(_0248_),
    .B(_0267_));
 sg13g2_nand3_1 _2028_ (.B(_0248_),
    .C(net337),
    .A(net166),
    .Y(_0269_));
 sg13g2_a22oi_1 _2029_ (.Y(_0096_),
    .B1(_0269_),
    .B2(_0338_),
    .A2(_0268_),
    .A1(_0822_));
 sg13g2_a21o_1 _2030_ (.A2(_0268_),
    .A1(_0822_),
    .B1(_0339_),
    .X(_0270_));
 sg13g2_o21ai_1 _2031_ (.B1(_0270_),
    .Y(_0097_),
    .A1(_0515_),
    .A2(_0269_));
 sg13g2_nand2b_2 _2032_ (.Y(_0271_),
    .B(net222),
    .A_N(net261));
 sg13g2_a21oi_1 _2033_ (.A1(net263),
    .A2(net162),
    .Y(_0272_),
    .B1(net194));
 sg13g2_o21ai_1 _2034_ (.B1(_0272_),
    .Y(_0098_),
    .A1(_0308_),
    .A2(net162));
 sg13g2_a21oi_1 _2035_ (.A1(\gamepad.decoder.data_reg[1] ),
    .A2(net162),
    .Y(_0273_),
    .B1(net194));
 sg13g2_o21ai_1 _2036_ (.B1(_0273_),
    .Y(_0099_),
    .A1(_0307_),
    .A2(net162));
 sg13g2_a21oi_1 _2037_ (.A1(net232),
    .A2(net162),
    .Y(_0274_),
    .B1(net195));
 sg13g2_o21ai_1 _2038_ (.B1(_0274_),
    .Y(_0100_),
    .A1(_0306_),
    .A2(_0271_));
 sg13g2_a21oi_1 _2039_ (.A1(net231),
    .A2(net160),
    .Y(_0275_),
    .B1(net190));
 sg13g2_o21ai_1 _2040_ (.B1(_0275_),
    .Y(_0101_),
    .A1(_0305_),
    .A2(net161));
 sg13g2_a21oi_1 _2041_ (.A1(net226),
    .A2(net160),
    .Y(_0276_),
    .B1(net190));
 sg13g2_o21ai_1 _2042_ (.B1(_0276_),
    .Y(_0102_),
    .A1(_0304_),
    .A2(net160));
 sg13g2_a21oi_1 _2043_ (.A1(net227),
    .A2(net160),
    .Y(_0277_),
    .B1(net190));
 sg13g2_o21ai_1 _2044_ (.B1(_0277_),
    .Y(_0103_),
    .A1(_0303_),
    .A2(net160));
 sg13g2_a21oi_1 _2045_ (.A1(net230),
    .A2(net160),
    .Y(_0278_),
    .B1(net190));
 sg13g2_o21ai_1 _2046_ (.B1(_0278_),
    .Y(_0104_),
    .A1(_0302_),
    .A2(net160));
 sg13g2_a21oi_1 _2047_ (.A1(net260),
    .A2(net161),
    .Y(_0279_),
    .B1(net191));
 sg13g2_o21ai_1 _2048_ (.B1(_0279_),
    .Y(_0105_),
    .A1(_0301_),
    .A2(net160));
 sg13g2_a21oi_1 _2049_ (.A1(\gamepad.decoder.data_reg[8] ),
    .A2(net161),
    .Y(_0280_),
    .B1(net191));
 sg13g2_o21ai_1 _2050_ (.B1(_0280_),
    .Y(_0106_),
    .A1(_0300_),
    .A2(net161));
 sg13g2_a21oi_1 _2051_ (.A1(net270),
    .A2(net162),
    .Y(_0281_),
    .B1(net191));
 sg13g2_o21ai_1 _2052_ (.B1(_0281_),
    .Y(_0107_),
    .A1(_0299_),
    .A2(net161));
 sg13g2_a21oi_1 _2053_ (.A1(net237),
    .A2(net162),
    .Y(_0282_),
    .B1(net195));
 sg13g2_o21ai_1 _2054_ (.B1(_0282_),
    .Y(_0108_),
    .A1(_0298_),
    .A2(_0271_));
 sg13g2_a21oi_1 _2055_ (.A1(\gamepad.decoder.data_reg[11] ),
    .A2(net161),
    .Y(_0283_),
    .B1(net191));
 sg13g2_o21ai_1 _2056_ (.B1(_0283_),
    .Y(_0109_),
    .A1(_0297_),
    .A2(net161));
 sg13g2_and2_1 _2057_ (.A(net200),
    .B(net221),
    .X(_0110_));
 sg13g2_nor2b_2 _2058_ (.A(net267),
    .B_N(net221),
    .Y(_0284_));
 sg13g2_a21oi_1 _2059_ (.A1(net252),
    .A2(_0284_),
    .Y(_0285_),
    .B1(net194));
 sg13g2_o21ai_1 _2060_ (.B1(net253),
    .Y(_0111_),
    .A1(_0308_),
    .A2(net159));
 sg13g2_a21oi_1 _2061_ (.A1(net265),
    .A2(net159),
    .Y(_0286_),
    .B1(net194));
 sg13g2_o21ai_1 _2062_ (.B1(_0286_),
    .Y(_0112_),
    .A1(_0307_),
    .A2(net159));
 sg13g2_a21oi_1 _2063_ (.A1(net258),
    .A2(net159),
    .Y(_0287_),
    .B1(net194));
 sg13g2_o21ai_1 _2064_ (.B1(_0287_),
    .Y(_0113_),
    .A1(_0306_),
    .A2(net159));
 sg13g2_a21oi_1 _2065_ (.A1(net250),
    .A2(net159),
    .Y(_0288_),
    .B1(net195));
 sg13g2_o21ai_1 _2066_ (.B1(_0288_),
    .Y(_0114_),
    .A1(_0305_),
    .A2(net157));
 sg13g2_a21oi_1 _2067_ (.A1(net268),
    .A2(net157),
    .Y(_0289_),
    .B1(net190));
 sg13g2_o21ai_1 _2068_ (.B1(_0289_),
    .Y(_0115_),
    .A1(_0304_),
    .A2(net157));
 sg13g2_a21oi_1 _2069_ (.A1(net262),
    .A2(net157),
    .Y(_0290_),
    .B1(net190));
 sg13g2_o21ai_1 _2070_ (.B1(_0290_),
    .Y(_0116_),
    .A1(_0303_),
    .A2(net157));
 sg13g2_a21oi_1 _2071_ (.A1(net264),
    .A2(net157),
    .Y(_0291_),
    .B1(net190));
 sg13g2_o21ai_1 _2072_ (.B1(_0291_),
    .Y(_0117_),
    .A1(_0302_),
    .A2(net157));
 sg13g2_a21oi_1 _2073_ (.A1(net269),
    .A2(net157),
    .Y(_0292_),
    .B1(net190));
 sg13g2_o21ai_1 _2074_ (.B1(_0292_),
    .Y(_0118_),
    .A1(_0301_),
    .A2(net158));
 sg13g2_a21oi_1 _2075_ (.A1(net266),
    .A2(net158),
    .Y(_0293_),
    .B1(net191));
 sg13g2_o21ai_1 _2076_ (.B1(_0293_),
    .Y(_0119_),
    .A1(_0300_),
    .A2(net158));
 sg13g2_a21oi_1 _2077_ (.A1(net248),
    .A2(net158),
    .Y(_0294_),
    .B1(net191));
 sg13g2_o21ai_1 _2078_ (.B1(_0294_),
    .Y(_0120_),
    .A1(_0299_),
    .A2(net158));
 sg13g2_a21oi_1 _2079_ (.A1(net271),
    .A2(net158),
    .Y(_0295_),
    .B1(net191));
 sg13g2_o21ai_1 _2080_ (.B1(_0295_),
    .Y(_0121_),
    .A1(_0298_),
    .A2(net159));
 sg13g2_a21oi_1 _2081_ (.A1(net242),
    .A2(net159),
    .Y(_0296_),
    .B1(net195));
 sg13g2_o21ai_1 _2082_ (.B1(net243),
    .Y(_0122_),
    .A1(_0297_),
    .A2(net158));
 sg13g2_and2_1 _2083_ (.A(net204),
    .B(net222),
    .X(_0123_));
 sg13g2_and2_1 _2084_ (.A(net203),
    .B(net3),
    .X(_0124_));
 sg13g2_and2_1 _2085_ (.A(net200),
    .B(net215),
    .X(_0125_));
 sg13g2_and2_1 _2086_ (.A(net203),
    .B(net2),
    .X(_0126_));
 sg13g2_and2_1 _2087_ (.A(net201),
    .B(net220),
    .X(_0127_));
 sg13g2_dfrbpq_1 _2088_ (.RESET_B(net22),
    .D(_0010_),
    .Q(vsync_prev),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _2089_ (.RESET_B(net23),
    .D(net395),
    .Q(\solver_l_dir[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _2090_ (.RESET_B(net24),
    .D(net314),
    .Q(\solver_l_dir[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _2091_ (.RESET_B(net25),
    .D(_0002_),
    .Q(\solver_l_dir[2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _2092_ (.RESET_B(net26),
    .D(_0003_),
    .Q(\solver_l_dir[3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _2093_ (.RESET_B(net27),
    .D(_0004_),
    .Q(\solver_r_dir[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _2094_ (.RESET_B(net28),
    .D(net280),
    .Q(\solver_r_dir[1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _2095_ (.RESET_B(net106),
    .D(net321),
    .Q(\solver_r_dir[2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _2096_ (.RESET_B(net21),
    .D(_0007_),
    .Q(\solver_r_dir[3] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _2097_ (.RESET_B(net32),
    .D(_0011_),
    .Q(\lfsr[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _2098_ (.RESET_B(net30),
    .D(_0012_),
    .Q(\lfsr[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _2099_ (.RESET_B(net20),
    .D(_0013_),
    .Q(\lfsr[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _2100_ (.RESET_B(net212),
    .D(net257),
    .Q(\lfsr[3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _2101_ (.RESET_B(net210),
    .D(net275),
    .Q(\lfsr[4] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _2102_ (.RESET_B(net208),
    .D(_0016_),
    .Q(\lfsr[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _2103_ (.RESET_B(net206),
    .D(net229),
    .Q(\lfsr[6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _2104_ (.RESET_B(net138),
    .D(net236),
    .Q(\lfsr[7] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _2105_ (.RESET_B(net136),
    .D(net289),
    .Q(\maze_seed[0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _2106_ (.RESET_B(net134),
    .D(_0020_),
    .Q(\maze_seed[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _2107_ (.RESET_B(net132),
    .D(net241),
    .Q(\maze_seed[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _2108_ (.RESET_B(net130),
    .D(_0022_),
    .Q(\maze_seed[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _2109_ (.RESET_B(net128),
    .D(_0023_),
    .Q(\maze_seed[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _2110_ (.RESET_B(net126),
    .D(_0024_),
    .Q(\ent_x[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _2111_ (.RESET_B(net125),
    .D(_0025_),
    .Q(\ent_x[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _2112_ (.RESET_B(net124),
    .D(_0026_),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _2113_ (.RESET_B(net123),
    .D(_0027_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _2114_ (.RESET_B(net122),
    .D(_0028_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _2115_ (.RESET_B(net121),
    .D(net335),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _2116_ (.RESET_B(net120),
    .D(_0030_),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _2117_ (.RESET_B(net119),
    .D(_0031_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _2118_ (.RESET_B(net118),
    .D(_0032_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _2119_ (.RESET_B(net116),
    .D(_0033_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _2120_ (.RESET_B(net115),
    .D(net287),
    .Q(\player_x[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _2121_ (.RESET_B(net114),
    .D(net343),
    .Q(\player_x[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _2122_ (.RESET_B(net113),
    .D(net351),
    .Q(\player_x[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _2123_ (.RESET_B(net112),
    .D(_0037_),
    .Q(\player_y[0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _2124_ (.RESET_B(net111),
    .D(net373),
    .Q(\player_y[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _2125_ (.RESET_B(net110),
    .D(_0039_),
    .Q(\player_y[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _2126_ (.RESET_B(net109),
    .D(_0040_),
    .Q(\solver_r_x[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _2127_ (.RESET_B(net108),
    .D(_0041_),
    .Q(\solver_r_x[1] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _2128_ (.RESET_B(net107),
    .D(_0042_),
    .Q(\solver_r_x[2] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _2129_ (.RESET_B(net105),
    .D(net346),
    .Q(\solver_r_y[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _2130_ (.RESET_B(net104),
    .D(net375),
    .Q(\solver_r_y[1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _2131_ (.RESET_B(net103),
    .D(_0045_),
    .Q(\solver_r_y[2] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _2132_ (.RESET_B(net102),
    .D(net380),
    .Q(\solver_l_x[0] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _2133_ (.RESET_B(net101),
    .D(net382),
    .Q(\solver_l_x[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _2134_ (.RESET_B(net100),
    .D(net391),
    .Q(\solver_l_x[2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _2135_ (.RESET_B(net99),
    .D(net309),
    .Q(solvers_active),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _2136_ (.RESET_B(net97),
    .D(_0050_),
    .Q(\solver_l_y[0] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _2137_ (.RESET_B(net96),
    .D(_0051_),
    .Q(\solver_l_y[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _2138_ (.RESET_B(net95),
    .D(_0052_),
    .Q(\solver_l_y[2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _2139_ (.RESET_B(net94),
    .D(_0053_),
    .Q(player_won),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _2140_ (.RESET_B(net93),
    .D(_0054_),
    .Q(solver_r_won),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _2141_ (.RESET_B(net92),
    .D(_0055_),
    .Q(generating),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _2142_ (.RESET_B(net90),
    .D(net366),
    .Q(\gen_row[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _2143_ (.RESET_B(net88),
    .D(net364),
    .Q(\gen_row[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _2144_ (.RESET_B(net86),
    .D(net325),
    .Q(\gen_row[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _2145_ (.RESET_B(net84),
    .D(_0059_),
    .Q(\gen_frame_count[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _2146_ (.RESET_B(net82),
    .D(net225),
    .Q(\gen_frame_count[1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _2147_ (.RESET_B(net80),
    .D(net219),
    .Q(\gen_frame_count[2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _2148_ (.RESET_B(net78),
    .D(net217),
    .Q(\gen_frame_count[3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _2149_ (.RESET_B(net76),
    .D(net349),
    .Q(\filled_width[1] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _2150_ (.RESET_B(net74),
    .D(_0064_),
    .Q(\solver_speed[1] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _2151_ (.RESET_B(net72),
    .D(net330),
    .Q(\solver_speed[2] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _2152_ (.RESET_B(net70),
    .D(net389),
    .Q(\solver_speed[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _2153_ (.RESET_B(net68),
    .D(_0067_),
    .Q(\solver_frame_count[0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _2154_ (.RESET_B(net66),
    .D(net284),
    .Q(\solver_frame_count[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _2155_ (.RESET_B(net64),
    .D(_0069_),
    .Q(\solver_frame_count[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _2156_ (.RESET_B(net62),
    .D(net306),
    .Q(\solver_frame_count[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _2157_ (.RESET_B(net60),
    .D(net358),
    .Q(single_step_mode),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _2158_ (.RESET_B(net58),
    .D(net319),
    .Q(step_requested),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _2159_ (.RESET_B(net56),
    .D(_0073_),
    .Q(solver_l_won),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _2160_ (.RESET_B(net55),
    .D(_0074_),
    .Q(inp_up_prev),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _2161_ (.RESET_B(net54),
    .D(_0075_),
    .Q(inp_down_prev),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _2162_ (.RESET_B(net53),
    .D(_0076_),
    .Q(inp_left_prev),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _2163_ (.RESET_B(net52),
    .D(_0077_),
    .Q(inp_right_prev),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _2164_ (.RESET_B(net51),
    .D(_0078_),
    .Q(inp_a_prev),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _2165_ (.RESET_B(net50),
    .D(_0079_),
    .Q(inp_b_prev),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _2166_ (.RESET_B(net49),
    .D(_0080_),
    .Q(inp_select_prev),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _2167_ (.RESET_B(net48),
    .D(_0081_),
    .Q(inp_start_prev),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _2168_ (.RESET_B(net47),
    .D(_0082_),
    .Q(inp_x_prev),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _2169_ (.RESET_B(net46),
    .D(_0083_),
    .Q(inp_y_prev),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _2170_ (.RESET_B(net45),
    .D(_0084_),
    .Q(inp_l_prev),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _2171_ (.RESET_B(net44),
    .D(_0085_),
    .Q(inp_r_prev),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _2172_ (.RESET_B(net43),
    .D(_0086_),
    .Q(\gamepad.driver.pmod_latch_sync[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _2173_ (.RESET_B(net117),
    .D(_0087_),
    .Q(\gamepad.driver.pmod_latch_sync[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _2174_ (.RESET_B(net42),
    .D(net278),
    .Q(hsync),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _2175_ (.RESET_B(net41),
    .D(_0088_),
    .Q(\ent_y[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _2176_ (.RESET_B(net39),
    .D(_0089_),
    .Q(\ent_y[1] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _2177_ (.RESET_B(net37),
    .D(net327),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _2178_ (.RESET_B(net35),
    .D(net296),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _2179_ (.RESET_B(net33),
    .D(net291),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _2180_ (.RESET_B(net29),
    .D(_0093_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _2181_ (.RESET_B(net211),
    .D(_0094_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _2182_ (.RESET_B(net207),
    .D(net294),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _2183_ (.RESET_B(net137),
    .D(_0096_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _2184_ (.RESET_B(net75),
    .D(_0097_),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _2185_ (.RESET_B(net133),
    .D(net301),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _2186_ (.RESET_B(net129),
    .D(_0098_),
    .Q(\gamepad.decoder.data_reg[0] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _2187_ (.RESET_B(net98),
    .D(net259),
    .Q(\gamepad.decoder.data_reg[1] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _2188_ (.RESET_B(net89),
    .D(net251),
    .Q(\gamepad.decoder.data_reg[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _2189_ (.RESET_B(net85),
    .D(_0101_),
    .Q(\gamepad.decoder.data_reg[3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _2190_ (.RESET_B(net81),
    .D(_0102_),
    .Q(\gamepad.decoder.data_reg[4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _2191_ (.RESET_B(net77),
    .D(_0103_),
    .Q(\gamepad.decoder.data_reg[5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _2192_ (.RESET_B(net73),
    .D(_0104_),
    .Q(\gamepad.decoder.data_reg[6] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _2193_ (.RESET_B(net69),
    .D(_0105_),
    .Q(\gamepad.decoder.data_reg[7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _2194_ (.RESET_B(net65),
    .D(net249),
    .Q(\gamepad.decoder.data_reg[8] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _2195_ (.RESET_B(net61),
    .D(_0107_),
    .Q(\gamepad.decoder.data_reg[9] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _2196_ (.RESET_B(net57),
    .D(_0108_),
    .Q(\gamepad.decoder.data_reg[10] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _2197_ (.RESET_B(net38),
    .D(net239),
    .Q(\gamepad.decoder.data_reg[11] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _2198_ (.RESET_B(net34),
    .D(_0110_),
    .Q(\gamepad.driver.pmod_clk_prev ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _2199_ (.RESET_B(net31),
    .D(net254),
    .Q(\gamepad.driver.shift_reg[0] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _2200_ (.RESET_B(net209),
    .D(_0112_),
    .Q(\gamepad.driver.shift_reg[1] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _2201_ (.RESET_B(net135),
    .D(_0113_),
    .Q(\gamepad.driver.shift_reg[2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _2202_ (.RESET_B(net127),
    .D(_0114_),
    .Q(\gamepad.driver.shift_reg[3] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _2203_ (.RESET_B(net87),
    .D(_0115_),
    .Q(\gamepad.driver.shift_reg[4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _2204_ (.RESET_B(net79),
    .D(_0116_),
    .Q(\gamepad.driver.shift_reg[5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _2205_ (.RESET_B(net71),
    .D(_0117_),
    .Q(\gamepad.driver.shift_reg[6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _2206_ (.RESET_B(net63),
    .D(_0118_),
    .Q(\gamepad.driver.shift_reg[7] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _2207_ (.RESET_B(net40),
    .D(_0119_),
    .Q(\gamepad.driver.shift_reg[8] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _2208_ (.RESET_B(net213),
    .D(_0120_),
    .Q(\gamepad.driver.shift_reg[9] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _2209_ (.RESET_B(net131),
    .D(_0121_),
    .Q(\gamepad.driver.shift_reg[10] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _2210_ (.RESET_B(net83),
    .D(net244),
    .Q(\gamepad.driver.shift_reg[11] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _2211_ (.RESET_B(net67),
    .D(_0123_),
    .Q(\gamepad.driver.pmod_latch_prev ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _2212_ (.RESET_B(net59),
    .D(_0124_),
    .Q(\gamepad.driver.pmod_data_sync[0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _2213_ (.RESET_B(net36),
    .D(_0125_),
    .Q(\gamepad.driver.pmod_data_sync[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _2214_ (.RESET_B(net139),
    .D(_0126_),
    .Q(\gamepad.driver.pmod_clk_sync[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _2215_ (.RESET_B(net91),
    .D(_0127_),
    .Q(\gamepad.driver.pmod_clk_sync[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_tiehi _2096__21 (.L_HI(net21));
 sg13g2_tiehi _2088__22 (.L_HI(net22));
 sg13g2_tiehi _2089__23 (.L_HI(net23));
 sg13g2_tiehi _2090__24 (.L_HI(net24));
 sg13g2_tiehi _2091__25 (.L_HI(net25));
 sg13g2_tiehi _2092__26 (.L_HI(net26));
 sg13g2_tiehi _2093__27 (.L_HI(net27));
 sg13g2_tiehi _2094__28 (.L_HI(net28));
 sg13g2_tiehi _2180__29 (.L_HI(net29));
 sg13g2_tiehi _2098__30 (.L_HI(net30));
 sg13g2_tiehi _2199__31 (.L_HI(net31));
 sg13g2_tiehi _2097__32 (.L_HI(net32));
 sg13g2_tiehi _2179__33 (.L_HI(net33));
 sg13g2_tiehi _2198__34 (.L_HI(net34));
 sg13g2_tiehi _2178__35 (.L_HI(net35));
 sg13g2_tiehi _2213__36 (.L_HI(net36));
 sg13g2_tiehi _2177__37 (.L_HI(net37));
 sg13g2_tiehi _2197__38 (.L_HI(net38));
 sg13g2_tiehi _2176__39 (.L_HI(net39));
 sg13g2_tiehi _2207__40 (.L_HI(net40));
 sg13g2_tiehi _2175__41 (.L_HI(net41));
 sg13g2_tiehi _2174__42 (.L_HI(net42));
 sg13g2_tiehi _2172__43 (.L_HI(net43));
 sg13g2_tiehi _2171__44 (.L_HI(net44));
 sg13g2_tiehi _2170__45 (.L_HI(net45));
 sg13g2_tiehi _2169__46 (.L_HI(net46));
 sg13g2_tiehi _2168__47 (.L_HI(net47));
 sg13g2_tiehi _2167__48 (.L_HI(net48));
 sg13g2_tiehi _2166__49 (.L_HI(net49));
 sg13g2_tiehi _2165__50 (.L_HI(net50));
 sg13g2_tiehi _2164__51 (.L_HI(net51));
 sg13g2_tiehi _2163__52 (.L_HI(net52));
 sg13g2_tiehi _2162__53 (.L_HI(net53));
 sg13g2_tiehi _2161__54 (.L_HI(net54));
 sg13g2_tiehi _2160__55 (.L_HI(net55));
 sg13g2_tiehi _2159__56 (.L_HI(net56));
 sg13g2_tiehi _2196__57 (.L_HI(net57));
 sg13g2_tiehi _2158__58 (.L_HI(net58));
 sg13g2_tiehi _2212__59 (.L_HI(net59));
 sg13g2_tiehi _2157__60 (.L_HI(net60));
 sg13g2_tiehi _2195__61 (.L_HI(net61));
 sg13g2_tiehi _2156__62 (.L_HI(net62));
 sg13g2_tiehi _2206__63 (.L_HI(net63));
 sg13g2_tiehi _2155__64 (.L_HI(net64));
 sg13g2_tiehi _2194__65 (.L_HI(net65));
 sg13g2_tiehi _2154__66 (.L_HI(net66));
 sg13g2_tiehi _2211__67 (.L_HI(net67));
 sg13g2_tiehi _2153__68 (.L_HI(net68));
 sg13g2_tiehi _2193__69 (.L_HI(net69));
 sg13g2_tiehi _2152__70 (.L_HI(net70));
 sg13g2_tiehi _2205__71 (.L_HI(net71));
 sg13g2_tiehi _2151__72 (.L_HI(net72));
 sg13g2_tiehi _2192__73 (.L_HI(net73));
 sg13g2_tiehi _2150__74 (.L_HI(net74));
 sg13g2_tiehi _2184__75 (.L_HI(net75));
 sg13g2_tiehi _2149__76 (.L_HI(net76));
 sg13g2_tiehi _2191__77 (.L_HI(net77));
 sg13g2_tiehi _2148__78 (.L_HI(net78));
 sg13g2_tiehi _2204__79 (.L_HI(net79));
 sg13g2_tiehi _2147__80 (.L_HI(net80));
 sg13g2_tiehi _2190__81 (.L_HI(net81));
 sg13g2_tiehi _2146__82 (.L_HI(net82));
 sg13g2_tiehi _2210__83 (.L_HI(net83));
 sg13g2_tiehi _2145__84 (.L_HI(net84));
 sg13g2_tiehi _2189__85 (.L_HI(net85));
 sg13g2_tiehi _2144__86 (.L_HI(net86));
 sg13g2_tiehi _2203__87 (.L_HI(net87));
 sg13g2_tiehi _2143__88 (.L_HI(net88));
 sg13g2_tiehi _2188__89 (.L_HI(net89));
 sg13g2_tiehi _2142__90 (.L_HI(net90));
 sg13g2_tiehi _2215__91 (.L_HI(net91));
 sg13g2_tiehi _2141__92 (.L_HI(net92));
 sg13g2_tiehi _2140__93 (.L_HI(net93));
 sg13g2_tiehi _2139__94 (.L_HI(net94));
 sg13g2_tiehi _2138__95 (.L_HI(net95));
 sg13g2_tiehi _2137__96 (.L_HI(net96));
 sg13g2_tiehi _2136__97 (.L_HI(net97));
 sg13g2_tiehi _2187__98 (.L_HI(net98));
 sg13g2_tiehi _2135__99 (.L_HI(net99));
 sg13g2_tiehi _2134__100 (.L_HI(net100));
 sg13g2_tiehi _2133__101 (.L_HI(net101));
 sg13g2_tiehi _2132__102 (.L_HI(net102));
 sg13g2_tiehi _2131__103 (.L_HI(net103));
 sg13g2_tiehi _2130__104 (.L_HI(net104));
 sg13g2_tiehi _2129__105 (.L_HI(net105));
 sg13g2_tiehi _2095__106 (.L_HI(net106));
 sg13g2_tiehi _2128__107 (.L_HI(net107));
 sg13g2_tiehi _2127__108 (.L_HI(net108));
 sg13g2_tiehi _2126__109 (.L_HI(net109));
 sg13g2_tiehi _2125__110 (.L_HI(net110));
 sg13g2_tiehi _2124__111 (.L_HI(net111));
 sg13g2_tiehi _2123__112 (.L_HI(net112));
 sg13g2_tiehi _2122__113 (.L_HI(net113));
 sg13g2_tiehi _2121__114 (.L_HI(net114));
 sg13g2_tiehi _2120__115 (.L_HI(net115));
 sg13g2_tiehi _2119__116 (.L_HI(net116));
 sg13g2_tiehi _2173__117 (.L_HI(net117));
 sg13g2_tiehi _2118__118 (.L_HI(net118));
 sg13g2_tiehi _2117__119 (.L_HI(net119));
 sg13g2_tiehi _2116__120 (.L_HI(net120));
 sg13g2_tiehi _2115__121 (.L_HI(net121));
 sg13g2_tiehi _2114__122 (.L_HI(net122));
 sg13g2_tiehi _2113__123 (.L_HI(net123));
 sg13g2_tiehi _2112__124 (.L_HI(net124));
 sg13g2_tiehi _2111__125 (.L_HI(net125));
 sg13g2_tiehi _2110__126 (.L_HI(net126));
 sg13g2_tiehi _2202__127 (.L_HI(net127));
 sg13g2_tiehi _2109__128 (.L_HI(net128));
 sg13g2_tiehi _2186__129 (.L_HI(net129));
 sg13g2_tiehi _2108__130 (.L_HI(net130));
 sg13g2_tiehi _2209__131 (.L_HI(net131));
 sg13g2_tiehi _2107__132 (.L_HI(net132));
 sg13g2_tiehi _2185__133 (.L_HI(net133));
 sg13g2_tiehi _2106__134 (.L_HI(net134));
 sg13g2_tiehi _2201__135 (.L_HI(net135));
 sg13g2_tiehi _2105__136 (.L_HI(net136));
 sg13g2_tiehi _2183__137 (.L_HI(net137));
 sg13g2_tiehi _2104__138 (.L_HI(net138));
 sg13g2_tiehi _2214__139 (.L_HI(net139));
 sg13g2_tiehi _2103__140 (.L_HI(net206));
 sg13g2_tiehi _2182__141 (.L_HI(net207));
 sg13g2_tiehi _2102__142 (.L_HI(net208));
 sg13g2_tiehi _2200__143 (.L_HI(net209));
 sg13g2_tiehi _2101__144 (.L_HI(net210));
 sg13g2_tiehi _2181__145 (.L_HI(net211));
 sg13g2_tiehi _2100__146 (.L_HI(net212));
 sg13g2_tiehi _2208__147 (.L_HI(net213));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_phsauter_vga_maze_5 (.L_LO(net5));
 sg13g2_tielo tt_um_phsauter_vga_maze_6 (.L_LO(net6));
 sg13g2_tielo tt_um_phsauter_vga_maze_7 (.L_LO(net7));
 sg13g2_tielo tt_um_phsauter_vga_maze_8 (.L_LO(net8));
 sg13g2_tielo tt_um_phsauter_vga_maze_9 (.L_LO(net9));
 sg13g2_tielo tt_um_phsauter_vga_maze_10 (.L_LO(net10));
 sg13g2_tielo tt_um_phsauter_vga_maze_11 (.L_LO(net11));
 sg13g2_tielo tt_um_phsauter_vga_maze_12 (.L_LO(net12));
 sg13g2_tielo tt_um_phsauter_vga_maze_13 (.L_LO(net13));
 sg13g2_tielo tt_um_phsauter_vga_maze_14 (.L_LO(net14));
 sg13g2_tielo tt_um_phsauter_vga_maze_15 (.L_LO(net15));
 sg13g2_tielo tt_um_phsauter_vga_maze_16 (.L_LO(net16));
 sg13g2_tielo tt_um_phsauter_vga_maze_17 (.L_LO(net17));
 sg13g2_tielo tt_um_phsauter_vga_maze_18 (.L_LO(net18));
 sg13g2_tielo tt_um_phsauter_vga_maze_19 (.L_LO(net19));
 sg13g2_tiehi _2099__20 (.L_HI(net20));
 sg13g2_buf_1 _2360_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2361_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout140 (.A(_0557_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0557_),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(_0596_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(_0397_),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0548_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0821_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(_0368_),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(_0366_),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0907_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(_0371_),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(_0539_),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(_0354_),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(_0354_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(_0359_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(_0284_),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(_0284_),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(_0271_),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(_0346_),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_0345_),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(_0345_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net293),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net336),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net340),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net393),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net370),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net345),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net401),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net384),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net377),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net378),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net334),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net400),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(\hvsync_gen.hpos[3] ),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(net347),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(net331),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(net285),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(net279),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(net399),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(net394),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(\solver_l_dir[1] ),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(\solver_l_dir[0] ),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(net199),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net199),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(_0322_),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net205),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(net205),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(net205),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_8 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(rst_n),
    .X(net205));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_tielo tt_um_phsauter_vga_maze_4 (.L_LO(net4));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad.driver.pmod_latch_sync[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad.driver.pmod_data_sync[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold3 (.A(\gen_frame_count[3] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0062_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold5 (.A(\gen_frame_count[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0061_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold7 (.A(\gamepad.driver.pmod_clk_sync[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold8 (.A(\gamepad.driver.pmod_clk_sync[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold9 (.A(\gamepad.driver.pmod_latch_sync[1] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ent_x[0] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold11 (.A(\gen_frame_count[1] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0060_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold13 (.A(\gamepad.decoder.data_reg[4] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold14 (.A(\gamepad.decoder.data_reg[5] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold15 (.A(\lfsr[6] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0017_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold17 (.A(\gamepad.decoder.data_reg[6] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold18 (.A(\gamepad.decoder.data_reg[3] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold19 (.A(\gamepad.decoder.data_reg[2] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0236_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold21 (.A(\lfsr[7] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0812_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0018_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold24 (.A(\gamepad.decoder.data_reg[10] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold25 (.A(\gamepad.driver.shift_reg[11] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0109_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold27 (.A(\lfsr[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0021_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold29 (.A(\gamepad.driver.shift_reg[10] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0296_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0122_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold32 (.A(\lfsr[1] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0813_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.vsync ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold35 (.A(\gamepad.driver.shift_reg[8] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0106_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold37 (.A(\gamepad.driver.shift_reg[2] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0100_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold39 (.A(\gamepad.driver.pmod_data_sync[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0285_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0111_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold42 (.A(\lfsr[3] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0808_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0014_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold45 (.A(\gamepad.driver.shift_reg[1] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0099_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold47 (.A(\gamepad.decoder.data_reg[7] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold48 (.A(\gamepad.driver.pmod_latch_prev ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold49 (.A(\gamepad.driver.shift_reg[4] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold50 (.A(\gamepad.decoder.data_reg[0] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold51 (.A(\gamepad.driver.shift_reg[5] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold52 (.A(\gamepad.driver.shift_reg[0] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold53 (.A(\gamepad.driver.shift_reg[7] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold54 (.A(\gamepad.driver.pmod_clk_prev ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold55 (.A(\gamepad.driver.shift_reg[3] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold56 (.A(\gamepad.driver.shift_reg[6] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold57 (.A(\gamepad.decoder.data_reg[9] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold58 (.A(\gamepad.driver.shift_reg[9] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold59 (.A(\gamepad.decoder.data_reg[11] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold60 (.A(\lfsr[4] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0809_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0015_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold63 (.A(\hvsync_gen.hpos[7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0520_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0008_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold66 (.A(\solver_r_dir[1] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0005_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold68 (.A(vsync_prev),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold69 (.A(\solver_frame_count[1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0230_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0068_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold72 (.A(\maze_seed[3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold73 (.A(\player_x[0] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0034_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold75 (.A(\lfsr[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0019_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold77 (.A(\hvsync_gen.vpos[4] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0092_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold79 (.A(\lfsr[5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold80 (.A(\hvsync_gen.vpos[7] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0095_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold82 (.A(\hvsync_gen.vpos[3] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0091_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold84 (.A(player_won),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0177_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold86 (.A(\maze_seed[4] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold87 (.A(\hvsync_gen.vpos[8] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0009_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold89 (.A(\solver_frame_count[0] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0229_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold91 (.A(\solver_frame_count[3] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0234_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0070_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold94 (.A(inp_a_prev),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0148_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0049_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold97 (.A(solver_l_won),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0245_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold99 (.A(\solver_frame_count[2] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold100 (.A(\solver_l_dir[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0001_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold102 (.A(solver_r_won),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0179_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold104 (.A(inp_y_prev),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0243_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0072_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold107 (.A(\solver_r_dir[2] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0006_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold109 (.A(\gen_frame_count[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0206_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold111 (.A(\gen_row[2] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0058_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold113 (.A(\hvsync_gen.vpos[2] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0090_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold115 (.A(\solver_speed[2] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0223_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0065_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ent_x[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold119 (.A(\hvsync_gen.hpos[3] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0817_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold121 (.A(\hvsync_gen.hpos[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0029_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold123 (.A(\hvsync_gen.vpos[5] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0263_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold125 (.A(\solver_r_dir[0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold126 (.A(\hvsync_gen.vpos[9] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold127 (.A(\ent_y[1] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0250_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold129 (.A(\player_x[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0035_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold131 (.A(\hvsync_gen.vpos[6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold132 (.A(\solver_r_y[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0043_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold134 (.A(\hvsync_gen.hpos[2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold135 (.A(\filled_width[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0063_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold137 (.A(\player_x[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0036_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold139 (.A(\hvsync_gen.hpos[9] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0833_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold141 (.A(\solver_speed[1] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0221_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold143 (.A(single_step_mode),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0239_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0071_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold146 (.A(\solver_r_dir[3] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold147 (.A(\solver_l_y[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0168_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold149 (.A(\gamepad.decoder.data_reg[1] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold150 (.A(\gen_row[1] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0057_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold152 (.A(\gen_row[0] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0056_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold154 (.A(\player_y[2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0899_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold156 (.A(\gamepad.decoder.data_reg[8] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold157 (.A(\solver_l_y[0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold158 (.A(\player_y[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0890_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0038_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold161 (.A(\solver_r_y[1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0044_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold163 (.A(\solver_l_y[2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold164 (.A(\hvsync_gen.hpos[8] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold165 (.A(\hvsync_gen.hpos[6] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold166 (.A(\solver_l_x[0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0046_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold168 (.A(\solver_l_x[1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0047_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold170 (.A(\solver_r_x[2] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold171 (.A(\player_y[0] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0888_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold173 (.A(\solver_speed[3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0224_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0225_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0066_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold177 (.A(\solver_l_x[2] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0048_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold179 (.A(\solver_r_x[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold180 (.A(\ent_y[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold181 (.A(\solver_l_dir[2] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0000_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold183 (.A(inp_start_prev),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0181_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0191_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold186 (.A(\solver_l_dir[3] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold187 (.A(\hvsync_gen.hpos[4] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold188 (.A(\solver_r_x[0] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold189 (.A(\solver_r_y[2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold190 (.A(\solver_r_x[0] ),
    .X(net403));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_135 ();
 sg13g2_fill_2 FILLER_0_152 ();
 sg13g2_fill_1 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_4 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_4 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_4 FILLER_0_252 ();
 sg13g2_fill_1 FILLER_0_269 ();
 sg13g2_fill_2 FILLER_0_288 ();
 sg13g2_fill_1 FILLER_0_295 ();
 sg13g2_decap_4 FILLER_0_305 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_fill_2 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_fill_2 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_4 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_4 FILLER_1_208 ();
 sg13g2_fill_2 FILLER_1_212 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_1 FILLER_1_298 ();
 sg13g2_fill_1 FILLER_1_307 ();
 sg13g2_decap_4 FILLER_1_330 ();
 sg13g2_fill_1 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_4 FILLER_1_351 ();
 sg13g2_decap_4 FILLER_1_368 ();
 sg13g2_fill_1 FILLER_1_372 ();
 sg13g2_fill_2 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_37 ();
 sg13g2_fill_1 FILLER_2_43 ();
 sg13g2_decap_4 FILLER_2_72 ();
 sg13g2_fill_2 FILLER_2_76 ();
 sg13g2_fill_2 FILLER_2_94 ();
 sg13g2_decap_8 FILLER_2_100 ();
 sg13g2_decap_8 FILLER_2_107 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_decap_4 FILLER_2_121 ();
 sg13g2_fill_1 FILLER_2_125 ();
 sg13g2_fill_1 FILLER_2_155 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_232 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_2 FILLER_2_260 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_decap_4 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_4 FILLER_2_319 ();
 sg13g2_fill_1 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_fill_2 FILLER_2_344 ();
 sg13g2_fill_1 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_4 ();
 sg13g2_fill_2 FILLER_3_10 ();
 sg13g2_fill_1 FILLER_3_12 ();
 sg13g2_decap_4 FILLER_3_17 ();
 sg13g2_fill_2 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_33 ();
 sg13g2_fill_1 FILLER_3_48 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_fill_2 FILLER_3_67 ();
 sg13g2_decap_4 FILLER_3_85 ();
 sg13g2_fill_2 FILLER_3_89 ();
 sg13g2_fill_2 FILLER_3_118 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_163 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_fill_2 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_222 ();
 sg13g2_decap_8 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_310 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_356 ();
 sg13g2_decap_4 FILLER_3_376 ();
 sg13g2_fill_2 FILLER_3_380 ();
 sg13g2_fill_2 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_fill_2 FILLER_4_77 ();
 sg13g2_fill_2 FILLER_4_106 ();
 sg13g2_fill_1 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_136 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_decap_4 FILLER_4_229 ();
 sg13g2_fill_2 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_263 ();
 sg13g2_fill_2 FILLER_4_273 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_fill_2 FILLER_4_305 ();
 sg13g2_fill_1 FILLER_4_307 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_fill_1 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_364 ();
 sg13g2_fill_2 FILLER_4_375 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_16 ();
 sg13g2_fill_2 FILLER_5_44 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_fill_2 FILLER_5_74 ();
 sg13g2_fill_1 FILLER_5_76 ();
 sg13g2_fill_1 FILLER_5_81 ();
 sg13g2_fill_1 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_135 ();
 sg13g2_fill_2 FILLER_5_153 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_178 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_fill_2 FILLER_5_218 ();
 sg13g2_fill_2 FILLER_5_257 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_fill_1 FILLER_5_369 ();
 sg13g2_fill_2 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_120 ();
 sg13g2_decap_4 FILLER_6_127 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_4 FILLER_6_142 ();
 sg13g2_fill_2 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_decap_4 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_223 ();
 sg13g2_fill_2 FILLER_6_229 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_decap_4 FILLER_6_240 ();
 sg13g2_fill_2 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_266 ();
 sg13g2_decap_4 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_308 ();
 sg13g2_fill_1 FILLER_6_329 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_decap_4 FILLER_7_10 ();
 sg13g2_fill_2 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_61 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_123 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_166 ();
 sg13g2_decap_4 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_decap_4 FILLER_7_194 ();
 sg13g2_fill_2 FILLER_7_198 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_decap_4 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_decap_4 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_decap_4 FILLER_7_335 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_2 FILLER_7_365 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_8_27 ();
 sg13g2_fill_1 FILLER_8_60 ();
 sg13g2_decap_4 FILLER_8_126 ();
 sg13g2_decap_4 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_180 ();
 sg13g2_decap_8 FILLER_8_187 ();
 sg13g2_decap_8 FILLER_8_215 ();
 sg13g2_decap_8 FILLER_8_222 ();
 sg13g2_decap_4 FILLER_8_241 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_292 ();
 sg13g2_fill_2 FILLER_8_308 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_decap_4 FILLER_9_9 ();
 sg13g2_fill_1 FILLER_9_13 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_81 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_decap_4 FILLER_9_139 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_decap_4 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_decap_4 FILLER_9_219 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_293 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_fill_1 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_9 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_78 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_decap_4 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_245 ();
 sg13g2_fill_2 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_264 ();
 sg13g2_decap_4 FILLER_10_271 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_4 FILLER_10_297 ();
 sg13g2_fill_2 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_311 ();
 sg13g2_fill_1 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_342 ();
 sg13g2_fill_2 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_27 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_195 ();
 sg13g2_decap_4 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_11_370 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_132 ();
 sg13g2_decap_4 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_204 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_246 ();
 sg13g2_fill_2 FILLER_12_253 ();
 sg13g2_decap_4 FILLER_12_271 ();
 sg13g2_decap_4 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_fill_2 FILLER_12_365 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_27 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_fill_2 FILLER_13_235 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_257 ();
 sg13g2_decap_4 FILLER_13_264 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_24 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_decap_4 FILLER_14_74 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_2 FILLER_14_197 ();
 sg13g2_decap_4 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_decap_4 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_365 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_386 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_4 FILLER_15_368 ();
 sg13g2_fill_2 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_10 ();
 sg13g2_fill_2 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_fill_2 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_83 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_4 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_99 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_345 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_397 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_decap_4 FILLER_17_9 ();
 sg13g2_decap_4 FILLER_17_48 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_decap_4 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_decap_4 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_374 ();
 sg13g2_decap_4 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_27 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_decap_4 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_132 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_decap_8 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_decap_4 FILLER_18_335 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_decap_4 FILLER_18_375 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_50 ();
 sg13g2_fill_2 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_80 ();
 sg13g2_decap_4 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_4 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_fill_2 FILLER_20_51 ();
 sg13g2_decap_4 FILLER_20_62 ();
 sg13g2_fill_1 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_4 FILLER_20_274 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_4 FILLER_20_285 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_9 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_decap_4 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_4 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_decap_4 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_decap_4 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_4 FILLER_22_271 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_decap_4 FILLER_22_344 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_9 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_68 ();
 sg13g2_decap_4 FILLER_23_75 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_decap_8 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_229 ();
 sg13g2_decap_8 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_decap_4 FILLER_24_9 ();
 sg13g2_fill_2 FILLER_24_13 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_25_27 ();
 sg13g2_fill_2 FILLER_25_100 ();
 sg13g2_fill_1 FILLER_25_125 ();
 sg13g2_decap_4 FILLER_25_143 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_4 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_decap_4 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_4 FILLER_25_393 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_fill_2 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_48 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_2 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_4 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_decap_4 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_152 ();
 sg13g2_decap_4 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_4 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_193 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_378 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_decap_4 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_171 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_290 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_fill_2 FILLER_32_394 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_decap_4 FILLER_34_9 ();
 sg13g2_fill_1 FILLER_34_13 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_decap_4 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_271 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_12 ();
 sg13g2_fill_1 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_decap_4 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_decap_4 FILLER_36_195 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_390 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_12 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
