module tt_um_snake_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire eat;
 wire failure;
 wire \game_inst.apple_inst.apple_x[0] ;
 wire \game_inst.apple_inst.apple_x[1] ;
 wire \game_inst.apple_inst.apple_x[2] ;
 wire \game_inst.apple_inst.apple_x[3] ;
 wire \game_inst.apple_inst.apple_x[4] ;
 wire \game_inst.apple_inst.apple_y[0] ;
 wire \game_inst.apple_inst.apple_y[1] ;
 wire \game_inst.apple_inst.apple_y[2] ;
 wire \game_inst.apple_inst.apple_y[3] ;
 wire \game_inst.apple_inst.i_snake_valid ;
 wire \game_inst.apple_inst.i_snake_x[0] ;
 wire \game_inst.apple_inst.i_snake_x[1] ;
 wire \game_inst.apple_inst.i_snake_x[2] ;
 wire \game_inst.apple_inst.i_snake_x[3] ;
 wire \game_inst.apple_inst.i_snake_x[4] ;
 wire \game_inst.apple_inst.i_snake_y[0] ;
 wire \game_inst.apple_inst.i_snake_y[1] ;
 wire \game_inst.apple_inst.i_snake_y[2] ;
 wire \game_inst.apple_inst.i_snake_y[3] ;
 wire \game_inst.apple_inst.o_ready ;
 wire \game_inst.apple_inst.random_inst.lfsr4[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[4] ;
 wire \game_inst.apple_inst.test ;
 wire \game_inst.control_inst.backwards[1] ;
 wire \game_inst.control_inst.dir[0] ;
 wire \game_inst.control_inst.dir[1] ;
 wire \game_inst.control_inst.i_head_dir[0] ;
 wire \game_inst.control_inst.o_start ;
 wire \game_inst.head_x[0] ;
 wire \game_inst.head_x[1] ;
 wire \game_inst.head_x[2] ;
 wire \game_inst.head_x[3] ;
 wire \game_inst.head_x[4] ;
 wire \game_inst.head_y[0] ;
 wire \game_inst.head_y[1] ;
 wire \game_inst.head_y[2] ;
 wire \game_inst.head_y[3] ;
 wire \game_inst.o_success ;
 wire \game_inst.o_tick ;
 wire \game_inst.o_vga_hsync ;
 wire \game_inst.o_vga_vsync ;
 wire \game_inst.pos_dir[0] ;
 wire \game_inst.pos_dir[1] ;
 wire \game_inst.snake_inst.dir_out[0] ;
 wire \game_inst.snake_inst.dir_out[1] ;
 wire \game_inst.snake_inst.length[0] ;
 wire \game_inst.snake_inst.length[1] ;
 wire \game_inst.snake_inst.length[2] ;
 wire \game_inst.snake_inst.length[3] ;
 wire \game_inst.snake_inst.length[4] ;
 wire \game_inst.snake_inst.length[5] ;
 wire \game_inst.snake_inst.length[6] ;
 wire \game_inst.snake_inst.length[7] ;
 wire \game_inst.snake_inst.pos[0] ;
 wire \game_inst.snake_inst.pos[1] ;
 wire \game_inst.snake_inst.pos[2] ;
 wire \game_inst.snake_inst.pos[3] ;
 wire \game_inst.snake_inst.pos[4] ;
 wire \game_inst.snake_inst.pos[5] ;
 wire \game_inst.snake_inst.pos[6] ;
 wire \game_inst.snake_inst.pos[7] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[100][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[100][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[101][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[101][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[102][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[102][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[103][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[103][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[104][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[104][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[105][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[105][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[106][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[106][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[107][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[107][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[108][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[108][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[109][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[109][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[10][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[10][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[110][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[110][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[111][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[111][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[112][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[112][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[113][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[113][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[114][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[114][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[115][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[115][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[116][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[116][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[117][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[117][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[118][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[118][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[119][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[119][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[11][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[11][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[120][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[120][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[121][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[121][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[122][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[122][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[123][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[123][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[124][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[124][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[125][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[125][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[126][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[126][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[127][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[127][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[128][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[128][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[129][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[129][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[12][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[12][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[130][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[130][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[131][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[131][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[132][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[132][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[133][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[133][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[134][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[134][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[135][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[135][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[136][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[136][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[137][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[137][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[138][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[138][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[139][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[139][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[13][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[13][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[140][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[140][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[141][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[141][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[142][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[142][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[143][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[143][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[144][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[144][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[145][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[145][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[146][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[146][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[147][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[147][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[148][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[148][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[149][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[149][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[14][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[14][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[150][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[150][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[151][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[151][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[152][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[152][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[153][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[153][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[154][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[154][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[155][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[155][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[156][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[156][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[157][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[157][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[158][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[158][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[159][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[159][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[15][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[15][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[160][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[160][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[161][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[161][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[162][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[162][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[163][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[163][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[164][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[164][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[165][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[165][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[166][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[166][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[167][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[167][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[168][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[168][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[169][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[169][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[16][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[16][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[170][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[170][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[171][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[171][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[172][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[172][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[173][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[173][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[174][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[174][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[175][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[175][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[176][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[176][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[177][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[177][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[178][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[178][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[179][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[179][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[17][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[17][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[180][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[180][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[181][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[181][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[182][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[182][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[183][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[183][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[184][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[184][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[185][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[185][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[186][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[186][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[187][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[187][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[188][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[188][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[189][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[189][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[18][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[18][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[190][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[190][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[191][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[191][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[192][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[192][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[193][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[193][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[194][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[194][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[195][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[195][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[196][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[196][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[197][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[197][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[198][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[198][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[199][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[199][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[19][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[19][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[1][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[1][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[200][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[200][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[201][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[201][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[202][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[202][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[203][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[203][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[204][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[204][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[205][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[205][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[206][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[206][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[207][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[207][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[208][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[208][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[209][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[209][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[20][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[20][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[210][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[210][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[211][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[211][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[212][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[212][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[213][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[213][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[214][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[214][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[215][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[215][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[216][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[216][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[217][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[217][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[218][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[218][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[219][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[219][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[21][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[21][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[220][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[220][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[221][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[221][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[222][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[222][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[223][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[223][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[224][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[224][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[225][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[225][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[226][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[226][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[227][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[227][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[228][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[228][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[229][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[229][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[22][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[22][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[230][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[230][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[231][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[231][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[232][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[232][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[23][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[23][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[24][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[24][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[25][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[25][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[26][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[26][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[27][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[27][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[28][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[28][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[29][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[29][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[2][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[2][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[30][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[30][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[31][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[31][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[32][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[32][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[33][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[33][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[34][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[34][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[35][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[35][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[36][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[36][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[37][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[37][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[38][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[38][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[39][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[39][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[3][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[3][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[40][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[40][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[41][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[41][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[42][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[42][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[43][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[43][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[44][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[44][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[45][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[45][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[46][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[46][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[47][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[47][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[48][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[48][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[49][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[49][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[4][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[4][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[50][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[50][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[51][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[51][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[52][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[52][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[53][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[53][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[54][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[54][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[55][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[55][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[56][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[56][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[57][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[57][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[58][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[58][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[59][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[59][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[5][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[5][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[60][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[60][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[61][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[61][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[62][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[62][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[63][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[63][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[64][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[64][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[65][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[65][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[66][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[66][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[67][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[67][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[68][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[68][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[69][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[69][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[6][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[6][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[70][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[70][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[71][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[71][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[72][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[72][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[73][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[73][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[74][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[74][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[75][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[75][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[76][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[76][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[77][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[77][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[78][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[78][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[79][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[79][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[7][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[7][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[80][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[80][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[81][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[81][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[82][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[82][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[83][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[83][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[84][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[84][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[85][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[85][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[86][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[86][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[87][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[87][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[88][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[88][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[89][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[89][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[8][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[8][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[90][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[90][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[91][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[91][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[92][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[92][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[93][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[93][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[94][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[94][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[95][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[95][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[96][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[96][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[97][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[97][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[98][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[98][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[99][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[99][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[9][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[9][1] ;
 wire \game_inst.tick ;
 wire \game_inst.tickgen_inst.counter[0] ;
 wire \game_inst.tickgen_inst.counter[1] ;
 wire \game_inst.tickgen_inst.counter[2] ;
 wire \game_inst.tickgen_inst.counter[3] ;
 wire \game_inst.tickgen_inst.counter_max[1] ;
 wire \game_inst.tickgen_inst.counter_max[2] ;
 wire \game_inst.tickgen_inst.counter_max[3] ;
 wire \game_inst.tickgen_inst.prev_user_input ;
 wire \game_inst.vga_inst.color[1] ;
 wire \game_inst.vga_inst.color[2] ;
 wire \game_inst.vga_inst.color[3] ;
 wire \game_inst.vga_inst.prev_dir[0] ;
 wire \game_inst.vga_inst.px[0] ;
 wire \game_inst.vga_inst.px[1] ;
 wire \game_inst.vga_inst.px[2] ;
 wire \game_inst.vga_inst.px[3] ;
 wire \game_inst.vga_inst.px[4] ;
 wire \game_inst.vga_inst.px[5] ;
 wire \game_inst.vga_inst.px[6] ;
 wire \game_inst.vga_inst.px[7] ;
 wire \game_inst.vga_inst.px[8] ;
 wire \game_inst.vga_inst.px[9] ;
 wire \game_inst.vga_inst.py[0] ;
 wire \game_inst.vga_inst.py[1] ;
 wire \game_inst.vga_inst.py[2] ;
 wire \game_inst.vga_inst.py[3] ;
 wire \game_inst.vga_inst.py[4] ;
 wire \game_inst.vga_inst.py[5] ;
 wire \game_inst.vga_inst.py[6] ;
 wire \game_inst.vga_inst.py[7] ;
 wire \game_inst.vga_inst.py[8] ;
 wire \game_inst.vga_inst.py[9] ;
 wire \game_inst.vga_inst.row_buffer[0][0] ;
 wire \game_inst.vga_inst.row_buffer[0][1] ;
 wire \game_inst.vga_inst.row_buffer[0][2] ;
 wire \game_inst.vga_inst.row_buffer[0][3] ;
 wire \game_inst.vga_inst.row_buffer[1][0] ;
 wire \game_inst.vga_inst.row_buffer[1][1] ;
 wire \game_inst.vga_inst.row_buffer[1][2] ;
 wire \game_inst.vga_inst.row_buffer[1][3] ;
 wire \game_inst.vga_inst.row_buffer[2][0] ;
 wire \game_inst.vga_inst.row_buffer[2][1] ;
 wire \game_inst.vga_inst.row_buffer[2][2] ;
 wire \game_inst.vga_inst.row_buffer[2][3] ;
 wire \game_inst.vga_inst.row_buffer[3][0] ;
 wire \game_inst.vga_inst.row_buffer[3][1] ;
 wire \game_inst.vga_inst.row_buffer[3][2] ;
 wire \game_inst.vga_inst.row_buffer[3][3] ;
 wire \game_inst.vga_inst.row_buffer[4][0] ;
 wire \game_inst.vga_inst.row_buffer[4][1] ;
 wire \game_inst.vga_inst.row_buffer[4][2] ;
 wire \game_inst.vga_inst.row_buffer[4][3] ;
 wire \game_inst.vga_inst.row_buffer[5][0] ;
 wire \game_inst.vga_inst.row_buffer[5][1] ;
 wire \game_inst.vga_inst.row_buffer[5][2] ;
 wire \game_inst.vga_inst.row_buffer[5][3] ;
 wire \game_inst.vga_inst.row_buffer[6][0] ;
 wire \game_inst.vga_inst.row_buffer[6][1] ;
 wire \game_inst.vga_inst.row_buffer[6][2] ;
 wire \game_inst.vga_inst.row_buffer[6][3] ;
 wire \game_inst.vga_inst.row_buffer[7][0] ;
 wire \game_inst.vga_inst.row_buffer[7][1] ;
 wire \game_inst.vga_inst.row_buffer[7][2] ;
 wire \game_inst.vga_inst.row_buffer[7][3] ;
 wire \game_inst.vga_inst.row_buffer[8][0] ;
 wire \game_inst.vga_inst.row_buffer[8][1] ;
 wire \game_inst.vga_inst.row_buffer[8][2] ;
 wire \game_inst.vga_inst.row_buffer[8][3] ;
 wire \game_inst.vga_inst.s_hsync ;
 wire \game_inst.vga_inst.s_vsync ;
 wire net662;
 wire net663;
 wire net664;
 wire clknet_leaf_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;

 sg13g2_inv_1 _1291_ (.Y(_0135_),
    .A(net1342));
 sg13g2_inv_2 _1292_ (.Y(_0136_),
    .A(net1248));
 sg13g2_inv_1 _1293_ (.Y(_0137_),
    .A(\game_inst.head_x[3] ));
 sg13g2_inv_1 _1294_ (.Y(_0138_),
    .A(net1249));
 sg13g2_inv_2 _1295_ (.Y(_0139_),
    .A(net1202));
 sg13g2_inv_2 _1296_ (.Y(_0140_),
    .A(\game_inst.control_inst.dir[0] ));
 sg13g2_inv_1 _1297_ (.Y(_0141_),
    .A(net1198));
 sg13g2_inv_1 _1298_ (.Y(_0142_),
    .A(net1169));
 sg13g2_inv_1 _1299_ (.Y(_0143_),
    .A(net1167));
 sg13g2_inv_1 _1300_ (.Y(_0144_),
    .A(net1188));
 sg13g2_inv_1 _1301_ (.Y(_0145_),
    .A(net1195));
 sg13g2_inv_1 _1302_ (.Y(_0146_),
    .A(net1172));
 sg13g2_inv_2 _1303_ (.Y(_0147_),
    .A(net1241));
 sg13g2_inv_1 _1304_ (.Y(_0148_),
    .A(\game_inst.vga_inst.py[6] ));
 sg13g2_inv_1 _1305_ (.Y(_0149_),
    .A(\game_inst.vga_inst.py[5] ));
 sg13g2_inv_2 _1306_ (.Y(_0150_),
    .A(net1311));
 sg13g2_inv_1 _1307_ (.Y(_0151_),
    .A(net1233));
 sg13g2_inv_1 _1308_ (.Y(_0152_),
    .A(net1221));
 sg13g2_inv_1 _1309_ (.Y(_0153_),
    .A(\game_inst.o_tick ));
 sg13g2_inv_1 _1310_ (.Y(_0154_),
    .A(net1146));
 sg13g2_inv_1 _1311_ (.Y(_0155_),
    .A(\game_inst.snake_inst.pos[4] ));
 sg13g2_inv_1 _1312_ (.Y(_0156_),
    .A(net134));
 sg13g2_inv_2 _1313_ (.Y(_0038_),
    .A(net1131));
 sg13g2_inv_1 _1314_ (.Y(_0157_),
    .A(net122));
 sg13g2_inv_2 _1315_ (.Y(_0158_),
    .A(net1250));
 sg13g2_inv_2 _1316_ (.Y(_0159_),
    .A(net1315));
 sg13g2_inv_2 _1317_ (.Y(_0160_),
    .A(net1197));
 sg13g2_inv_1 _1318_ (.Y(_0161_),
    .A(net1273));
 sg13g2_inv_1 _1319_ (.Y(_0162_),
    .A(net1196));
 sg13g2_inv_1 _1320_ (.Y(_0163_),
    .A(\game_inst.apple_inst.i_snake_y[0] ));
 sg13g2_inv_1 _1321_ (.Y(_0164_),
    .A(\game_inst.apple_inst.i_snake_y[1] ));
 sg13g2_inv_1 _1322_ (.Y(_0165_),
    .A(\game_inst.apple_inst.apple_y[1] ));
 sg13g2_inv_2 _1323_ (.Y(_0166_),
    .A(net129));
 sg13g2_inv_2 _1324_ (.Y(_0167_),
    .A(net125));
 sg13g2_inv_1 _1325_ (.Y(_0168_),
    .A(net2));
 sg13g2_inv_1 _1326_ (.Y(_0169_),
    .A(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ));
 sg13g2_nand4_1 _1327_ (.B(\game_inst.snake_inst.length[5] ),
    .C(\game_inst.snake_inst.length[6] ),
    .A(_0152_),
    .Y(_0170_),
    .D(\game_inst.snake_inst.length[7] ));
 sg13g2_nand2b_1 _1328_ (.Y(_0171_),
    .B(\game_inst.snake_inst.length[3] ),
    .A_N(\game_inst.snake_inst.length[2] ));
 sg13g2_nor4_1 _1329_ (.A(_0150_),
    .B(\game_inst.snake_inst.length[1] ),
    .C(_0170_),
    .D(_0171_),
    .Y(\game_inst.o_success ));
 sg13g2_nor2_1 _1330_ (.A(net2),
    .B(net1),
    .Y(_0172_));
 sg13g2_inv_1 _1331_ (.Y(_0003_),
    .A(_0172_));
 sg13g2_nor3_1 _1332_ (.A(\game_inst.vga_inst.py[8] ),
    .B(\game_inst.vga_inst.py[7] ),
    .C(\game_inst.vga_inst.py[6] ),
    .Y(_0173_));
 sg13g2_nand3_1 _1333_ (.B(\game_inst.vga_inst.py[7] ),
    .C(\game_inst.vga_inst.py[6] ),
    .A(\game_inst.vga_inst.py[8] ),
    .Y(_0174_));
 sg13g2_nand2b_1 _1334_ (.Y(_0175_),
    .B(_0174_),
    .A_N(_0173_));
 sg13g2_and2_1 _1335_ (.A(_0149_),
    .B(_0175_),
    .X(_0176_));
 sg13g2_nor2_1 _1336_ (.A(net129),
    .B(net128),
    .Y(_0177_));
 sg13g2_and2_1 _1337_ (.A(net129),
    .B(\game_inst.vga_inst.px[6] ),
    .X(_0178_));
 sg13g2_nor3_1 _1338_ (.A(net129),
    .B(net124),
    .C(\game_inst.vga_inst.px[6] ),
    .Y(_0179_));
 sg13g2_a21oi_1 _1339_ (.A1(net124),
    .A2(_0178_),
    .Y(_0180_),
    .B1(_0179_));
 sg13g2_nor3_1 _1340_ (.A(net125),
    .B(net127),
    .C(_0180_),
    .Y(_0181_));
 sg13g2_nor2_1 _1341_ (.A(_0176_),
    .B(_0181_),
    .Y(_0182_));
 sg13g2_or2_1 _1342_ (.X(_0183_),
    .B(_0174_),
    .A(_0149_));
 sg13g2_o21ai_1 _1343_ (.B1(net124),
    .Y(_0184_),
    .A1(net1336),
    .A2(net127));
 sg13g2_nand3b_1 _1344_ (.B(_0183_),
    .C(_0184_),
    .Y(_0185_),
    .A_N(net1200));
 sg13g2_nor2_1 _1345_ (.A(_0182_),
    .B(_0185_),
    .Y(_0186_));
 sg13g2_or3_1 _1346_ (.A(_0176_),
    .B(_0181_),
    .C(_0185_),
    .X(_0187_));
 sg13g2_nand3_1 _1347_ (.B(net1209),
    .C(net1213),
    .A(net1157),
    .Y(_0188_));
 sg13g2_or3_1 _1348_ (.A(\game_inst.vga_inst.py[4] ),
    .B(\game_inst.vga_inst.py[3] ),
    .C(\game_inst.vga_inst.py[2] ),
    .X(_0189_));
 sg13g2_and2_1 _1349_ (.A(_0188_),
    .B(_0189_),
    .X(_0190_));
 sg13g2_nand3_1 _1350_ (.B(net1159),
    .C(net1255),
    .A(net1285),
    .Y(_0191_));
 sg13g2_or3_1 _1351_ (.A(net1345),
    .B(net1159),
    .C(net1255),
    .X(_0192_));
 sg13g2_nand3_1 _1352_ (.B(_0191_),
    .C(_0192_),
    .A(_0190_),
    .Y(_0193_));
 sg13g2_nor4_1 _1353_ (.A(net1231),
    .B(net1207),
    .C(net1228),
    .D(net1226),
    .Y(_0194_));
 sg13g2_nand2b_1 _1354_ (.Y(_0195_),
    .B(net1241),
    .A_N(net1217));
 sg13g2_xnor2_1 _1355_ (.Y(_0196_),
    .A(\game_inst.vga_inst.py[5] ),
    .B(net1196));
 sg13g2_xnor2_1 _1356_ (.Y(_0197_),
    .A(net1214),
    .B(net1181));
 sg13g2_o21ai_1 _1357_ (.B1(net121),
    .Y(_0198_),
    .A1(\game_inst.apple_inst.apple_x[0] ),
    .A2(_0166_));
 sg13g2_xnor2_1 _1358_ (.Y(_0199_),
    .A(\game_inst.vga_inst.py[6] ),
    .B(\game_inst.apple_inst.apple_y[1] ));
 sg13g2_a22oi_1 _1359_ (.Y(_0200_),
    .B1(_0166_),
    .B2(net1245),
    .A2(net1217),
    .A1(_0147_));
 sg13g2_xnor2_1 _1360_ (.Y(_0201_),
    .A(net1197),
    .B(net125));
 sg13g2_xor2_1 _1361_ (.B(net128),
    .A(\game_inst.apple_inst.apple_x[1] ),
    .X(_0202_));
 sg13g2_xor2_1 _1362_ (.B(net127),
    .A(\game_inst.apple_inst.apple_x[2] ),
    .X(_0203_));
 sg13g2_xor2_1 _1363_ (.B(net124),
    .A(\game_inst.apple_inst.apple_x[4] ),
    .X(_0204_));
 sg13g2_nor4_1 _1364_ (.A(_0198_),
    .B(_0202_),
    .C(_0203_),
    .D(_0204_),
    .Y(_0205_));
 sg13g2_nand4_1 _1365_ (.B(_0197_),
    .C(_0199_),
    .A(_0194_),
    .Y(_0206_),
    .D(_0205_));
 sg13g2_nand4_1 _1366_ (.B(_0196_),
    .C(_0200_),
    .A(_0195_),
    .Y(_0207_),
    .D(_0201_));
 sg13g2_nor4_1 _1367_ (.A(_0187_),
    .B(_0193_),
    .C(_0206_),
    .D(net1246),
    .Y(_0208_));
 sg13g2_a21o_1 _1368_ (.A2(_0186_),
    .A1(net1134),
    .B1(net1247),
    .X(_0000_));
 sg13g2_nor3_1 _1369_ (.A(net1134),
    .B(_0182_),
    .C(_0185_),
    .Y(_0002_));
 sg13g2_mux2_1 _1370_ (.A0(net1228),
    .A1(net1226),
    .S(net1285),
    .X(_0209_));
 sg13g2_nand2_1 _1371_ (.Y(_0210_),
    .A(_0190_),
    .B(_0209_));
 sg13g2_nor2_1 _1372_ (.A(net1231),
    .B(_0189_),
    .Y(_0211_));
 sg13g2_o21ai_1 _1373_ (.B1(_0188_),
    .Y(_0212_),
    .A1(_0194_),
    .A2(_0211_));
 sg13g2_or2_1 _1374_ (.X(_0213_),
    .B(_0188_),
    .A(net1207));
 sg13g2_nand4_1 _1375_ (.B(_0192_),
    .C(_0212_),
    .A(_0191_),
    .Y(_0214_),
    .D(_0213_));
 sg13g2_a21oi_1 _1376_ (.A1(_0210_),
    .A2(_0214_),
    .Y(_0001_),
    .B1(_0187_));
 sg13g2_nand3b_1 _1377_ (.B(\game_inst.vga_inst.py[3] ),
    .C(\game_inst.vga_inst.py[1] ),
    .Y(_0215_),
    .A_N(\game_inst.vga_inst.py[9] ));
 sg13g2_nor4_1 _1378_ (.A(net1157),
    .B(\game_inst.vga_inst.py[2] ),
    .C(_0183_),
    .D(_0215_),
    .Y(_0037_));
 sg13g2_nor3_1 _1379_ (.A(net1238),
    .B(\game_inst.vga_inst.px[6] ),
    .C(net1285),
    .Y(_0216_));
 sg13g2_a21oi_1 _1380_ (.A1(net1285),
    .A2(_0178_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_and4_1 _1381_ (.A(net124),
    .B(_0167_),
    .C(net127),
    .D(_0217_),
    .X(_0036_));
 sg13g2_nor2b_1 _1382_ (.A(net121),
    .B_N(\game_inst.control_inst.o_start ),
    .Y(eat));
 sg13g2_and3_1 _1383_ (.X(_0218_),
    .A(net1132),
    .B(net1133),
    .C(net1159));
 sg13g2_and2_1 _1384_ (.A(net1255),
    .B(_0218_),
    .X(_0219_));
 sg13g2_and2_1 _1385_ (.A(\game_inst.vga_inst.px[4] ),
    .B(_0219_),
    .X(_0220_));
 sg13g2_nand2_1 _1386_ (.Y(_0221_),
    .A(net1285),
    .B(_0219_));
 sg13g2_xor2_1 _1387_ (.B(\game_inst.snake_inst.pos[0] ),
    .A(\game_inst.snake_inst.length[0] ),
    .X(_0222_));
 sg13g2_xor2_1 _1388_ (.B(\game_inst.snake_inst.pos[7] ),
    .A(\game_inst.snake_inst.length[7] ),
    .X(_0223_));
 sg13g2_xnor2_1 _1389_ (.Y(_0224_),
    .A(\game_inst.snake_inst.length[4] ),
    .B(\game_inst.snake_inst.pos[4] ));
 sg13g2_xor2_1 _1390_ (.B(\game_inst.snake_inst.pos[5] ),
    .A(\game_inst.snake_inst.length[5] ),
    .X(_0225_));
 sg13g2_xor2_1 _1391_ (.B(\game_inst.snake_inst.pos[2] ),
    .A(\game_inst.snake_inst.length[2] ),
    .X(_0226_));
 sg13g2_xor2_1 _1392_ (.B(\game_inst.snake_inst.pos[1] ),
    .A(\game_inst.snake_inst.length[1] ),
    .X(_0227_));
 sg13g2_xor2_1 _1393_ (.B(\game_inst.snake_inst.pos[6] ),
    .A(\game_inst.snake_inst.length[6] ),
    .X(_0228_));
 sg13g2_xor2_1 _1394_ (.B(\game_inst.snake_inst.pos[3] ),
    .A(\game_inst.snake_inst.length[3] ),
    .X(_0229_));
 sg13g2_nor3_1 _1395_ (.A(_0225_),
    .B(_0226_),
    .C(_0228_),
    .Y(_0230_));
 sg13g2_nor4_1 _1396_ (.A(_0222_),
    .B(_0223_),
    .C(_0227_),
    .D(_0229_),
    .Y(_0231_));
 sg13g2_nand3_1 _1397_ (.B(_0230_),
    .C(_0231_),
    .A(_0224_),
    .Y(_0232_));
 sg13g2_and2_1 _1398_ (.A(_0038_),
    .B(_0232_),
    .X(_0233_));
 sg13g2_nand2_1 _1399_ (.Y(_0234_),
    .A(_0157_),
    .B(_0233_));
 sg13g2_nor4_1 _1400_ (.A(\game_inst.snake_inst.pos[3] ),
    .B(\game_inst.snake_inst.pos[4] ),
    .C(\game_inst.snake_inst.pos[5] ),
    .D(\game_inst.snake_inst.pos[6] ),
    .Y(_0235_));
 sg13g2_nor2_1 _1401_ (.A(net1303),
    .B(net1162),
    .Y(_0236_));
 sg13g2_nor4_1 _1402_ (.A(\game_inst.snake_inst.pos[7] ),
    .B(\game_inst.snake_inst.pos[1] ),
    .C(\game_inst.snake_inst.pos[0] ),
    .D(\game_inst.snake_inst.pos[2] ),
    .Y(_0237_));
 sg13g2_and2_1 _1403_ (.A(_0235_),
    .B(_0237_),
    .X(_0238_));
 sg13g2_or2_1 _1404_ (.X(_0239_),
    .B(_0238_),
    .A(\game_inst.vga_inst.prev_dir[0] ));
 sg13g2_o21ai_1 _1405_ (.B1(_0234_),
    .Y(_0240_),
    .A1(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .A2(_0239_));
 sg13g2_nand2b_1 _1406_ (.Y(_0241_),
    .B(net116),
    .A_N(net126));
 sg13g2_nor2b_1 _1407_ (.A(net128),
    .B_N(net117),
    .Y(_0242_));
 sg13g2_nand2b_1 _1408_ (.Y(_0243_),
    .B(net129),
    .A_N(net118));
 sg13g2_nor2b_1 _1409_ (.A(net117),
    .B_N(net128),
    .Y(_0244_));
 sg13g2_xnor2_1 _1410_ (.Y(_0245_),
    .A(net117),
    .B(net128));
 sg13g2_a21oi_1 _1411_ (.A1(_0243_),
    .A2(_0245_),
    .Y(_0246_),
    .B1(_0242_));
 sg13g2_nor2b_1 _1412_ (.A(net116),
    .B_N(net126),
    .Y(_0247_));
 sg13g2_xnor2_1 _1413_ (.Y(_0248_),
    .A(net116),
    .B(net126));
 sg13g2_o21ai_1 _1414_ (.B1(_0241_),
    .Y(_0249_),
    .A1(_0246_),
    .A2(_0247_));
 sg13g2_xnor2_1 _1415_ (.Y(_0250_),
    .A(\game_inst.apple_inst.i_snake_x[3] ),
    .B(net125));
 sg13g2_xnor2_1 _1416_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_inv_1 _1417_ (.Y(_0252_),
    .A(_0251_));
 sg13g2_nand2_1 _1418_ (.Y(_0253_),
    .A(net1174),
    .B(net1160));
 sg13g2_and4_1 _1419_ (.A(net1209),
    .B(\game_inst.vga_inst.py[2] ),
    .C(net1174),
    .D(net1160),
    .X(_0254_));
 sg13g2_nand3_1 _1420_ (.B(net1157),
    .C(_0254_),
    .A(net1266),
    .Y(_0255_));
 sg13g2_nand4_1 _1421_ (.B(\game_inst.vga_inst.py[5] ),
    .C(\game_inst.vga_inst.py[4] ),
    .A(\game_inst.vga_inst.py[6] ),
    .Y(_0256_),
    .D(_0254_));
 sg13g2_xnor2_1 _1422_ (.Y(_0257_),
    .A(\game_inst.vga_inst.py[7] ),
    .B(\game_inst.apple_inst.i_snake_y[2] ));
 sg13g2_nand2_1 _1423_ (.Y(_0258_),
    .A(net1157),
    .B(_0254_));
 sg13g2_xnor2_1 _1424_ (.Y(_0259_),
    .A(\game_inst.vga_inst.py[5] ),
    .B(\game_inst.apple_inst.i_snake_y[0] ));
 sg13g2_xnor2_1 _1425_ (.Y(_0260_),
    .A(_0258_),
    .B(_0259_));
 sg13g2_nor3_2 _1426_ (.A(_0147_),
    .B(_0148_),
    .C(_0255_),
    .Y(_0261_));
 sg13g2_xnor2_1 _1427_ (.Y(_0262_),
    .A(\game_inst.vga_inst.py[8] ),
    .B(\game_inst.apple_inst.i_snake_y[3] ));
 sg13g2_xnor2_1 _1428_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_xnor2_1 _1429_ (.Y(_0264_),
    .A(\game_inst.vga_inst.py[6] ),
    .B(\game_inst.apple_inst.i_snake_y[1] ));
 sg13g2_nand2_1 _1430_ (.Y(_0265_),
    .A(_0161_),
    .B(net124));
 sg13g2_a21oi_1 _1431_ (.A1(\game_inst.apple_inst.i_snake_x[3] ),
    .A2(_0167_),
    .Y(_0266_),
    .B1(_0265_));
 sg13g2_xnor2_1 _1432_ (.Y(_0267_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_xor2_1 _1433_ (.B(_0264_),
    .A(_0255_),
    .X(_0268_));
 sg13g2_nand3_1 _1434_ (.B(_0266_),
    .C(_0267_),
    .A(_0260_),
    .Y(_0269_));
 sg13g2_nor4_2 _1435_ (.A(_0251_),
    .B(_0263_),
    .C(_0268_),
    .Y(_0270_),
    .D(_0269_));
 sg13g2_or4_1 _1436_ (.A(_0251_),
    .B(_0263_),
    .C(_0268_),
    .D(_0269_),
    .X(_0271_));
 sg13g2_nand2_2 _1437_ (.Y(_0272_),
    .A(\game_inst.apple_inst.i_snake_valid ),
    .B(_0270_));
 sg13g2_nand2b_2 _1438_ (.Y(_0273_),
    .B(\game_inst.apple_inst.i_snake_x[4] ),
    .A_N(\game_inst.vga_inst.px[9] ));
 sg13g2_o21ai_1 _1439_ (.B1(_0273_),
    .Y(_0274_),
    .A1(_0159_),
    .A2(net125));
 sg13g2_a21oi_1 _1440_ (.A1(_0249_),
    .A2(_0250_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_nor2b_1 _1441_ (.A(net129),
    .B_N(net118),
    .Y(_0276_));
 sg13g2_nand2b_1 _1442_ (.Y(_0277_),
    .B(net118),
    .A_N(net129));
 sg13g2_and2_1 _1443_ (.A(_0243_),
    .B(_0277_),
    .X(_0278_));
 sg13g2_and2_1 _1444_ (.A(_0248_),
    .B(_0250_),
    .X(_0279_));
 sg13g2_nand4_1 _1445_ (.B(_0273_),
    .C(_0278_),
    .A(_0245_),
    .Y(_0280_),
    .D(_0279_));
 sg13g2_nand3_1 _1446_ (.B(net126),
    .C(net128),
    .A(net129),
    .Y(_0281_));
 sg13g2_nand3b_1 _1447_ (.B(_0281_),
    .C(_0167_),
    .Y(_0282_),
    .A_N(_0273_));
 sg13g2_nand4_1 _1448_ (.B(_0262_),
    .C(_0265_),
    .A(\game_inst.apple_inst.i_snake_valid ),
    .Y(_0283_),
    .D(_0282_));
 sg13g2_nand4_1 _1449_ (.B(_0259_),
    .C(_0264_),
    .A(_0257_),
    .Y(_0284_),
    .D(_0280_));
 sg13g2_nand2b_1 _1450_ (.Y(_0285_),
    .B(_0277_),
    .A_N(_0242_));
 sg13g2_nor3_1 _1451_ (.A(_0178_),
    .B(_0244_),
    .C(_0247_),
    .Y(_0286_));
 sg13g2_nand2_1 _1452_ (.Y(_0287_),
    .A(\game_inst.apple_inst.i_snake_x[3] ),
    .B(net125));
 sg13g2_nand3_1 _1453_ (.B(_0281_),
    .C(_0287_),
    .A(_0241_),
    .Y(_0288_));
 sg13g2_a21oi_1 _1454_ (.A1(_0285_),
    .A2(_0286_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_a21oi_1 _1455_ (.A1(_0159_),
    .A2(net125),
    .Y(_0290_),
    .B1(_0273_));
 sg13g2_a21oi_1 _1456_ (.A1(_0274_),
    .A2(_0281_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_nor2_1 _1457_ (.A(_0289_),
    .B(_0291_),
    .Y(_0292_));
 sg13g2_or4_1 _1458_ (.A(_0275_),
    .B(_0283_),
    .C(_0284_),
    .D(_0292_),
    .X(_0293_));
 sg13g2_o21ai_1 _1459_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0136_),
    .A2(_0271_));
 sg13g2_and3_2 _1460_ (.X(_0295_),
    .A(net118),
    .B(net117),
    .C(net116));
 sg13g2_a21oi_1 _1461_ (.A1(net118),
    .A2(net117),
    .Y(_0296_),
    .B1(net116));
 sg13g2_nor3_1 _1462_ (.A(net126),
    .B(_0295_),
    .C(_0296_),
    .Y(_0297_));
 sg13g2_o21ai_1 _1463_ (.B1(net126),
    .Y(_0298_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_nor2b_1 _1464_ (.A(_0297_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_a22oi_1 _1465_ (.Y(_0300_),
    .B1(_0244_),
    .B2(_0277_),
    .A2(net117),
    .A1(net118));
 sg13g2_or2_1 _1466_ (.X(_0301_),
    .B(_0300_),
    .A(_0177_));
 sg13g2_a21oi_1 _1467_ (.A1(_0298_),
    .A2(_0301_),
    .Y(_0302_),
    .B1(_0297_));
 sg13g2_xnor2_1 _1468_ (.Y(_0303_),
    .A(_0250_),
    .B(_0295_));
 sg13g2_xnor2_1 _1469_ (.Y(_0304_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_o21ai_1 _1470_ (.B1(_0252_),
    .Y(_0305_),
    .A1(_0271_),
    .A2(_0304_));
 sg13g2_nor2b_2 _1471_ (.A(_0305_),
    .B_N(_0294_),
    .Y(_0306_));
 sg13g2_a21oi_1 _1472_ (.A1(_0240_),
    .A2(_0306_),
    .Y(_0307_),
    .B1(net1142));
 sg13g2_nor2_1 _1473_ (.A(net111),
    .B(_0307_),
    .Y(_0032_));
 sg13g2_nor2b_1 _1474_ (.A(_0238_),
    .B_N(\game_inst.vga_inst.prev_dir[0] ),
    .Y(_0308_));
 sg13g2_nand2_1 _1475_ (.Y(_0309_),
    .A(_0169_),
    .B(_0308_));
 sg13g2_nand2_1 _1476_ (.Y(_0310_),
    .A(\game_inst.pos_dir[0] ),
    .B(_0232_));
 sg13g2_o21ai_1 _1477_ (.B1(_0309_),
    .Y(_0311_),
    .A1(net122),
    .A2(_0310_));
 sg13g2_a21oi_1 _1478_ (.A1(_0306_),
    .A2(_0311_),
    .Y(_0312_),
    .B1(net1148));
 sg13g2_nor2_1 _1479_ (.A(net111),
    .B(_0312_),
    .Y(_0033_));
 sg13g2_nand2_1 _1480_ (.Y(_0313_),
    .A(net122),
    .B(_0233_));
 sg13g2_o21ai_1 _1481_ (.B1(_0313_),
    .Y(_0314_),
    .A1(_0169_),
    .A2(_0239_));
 sg13g2_a21oi_1 _1482_ (.A1(_0306_),
    .A2(_0314_),
    .Y(_0315_),
    .B1(net1136));
 sg13g2_nor2_1 _1483_ (.A(net111),
    .B(_0315_),
    .Y(_0034_));
 sg13g2_nand2_1 _1484_ (.Y(_0316_),
    .A(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .B(_0308_));
 sg13g2_o21ai_1 _1485_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0157_),
    .A2(_0310_));
 sg13g2_a21oi_1 _1486_ (.A1(_0306_),
    .A2(_0317_),
    .Y(_0318_),
    .B1(net1144));
 sg13g2_nor2_1 _1487_ (.A(net111),
    .B(_0318_),
    .Y(_0035_));
 sg13g2_nor3_1 _1488_ (.A(_0136_),
    .B(_0271_),
    .C(_0304_),
    .Y(_0319_));
 sg13g2_nand3b_1 _1489_ (.B(_0270_),
    .C(\game_inst.apple_inst.i_snake_valid ),
    .Y(_0320_),
    .A_N(_0304_));
 sg13g2_xor2_1 _1490_ (.B(_0301_),
    .A(_0299_),
    .X(_0321_));
 sg13g2_xnor2_1 _1491_ (.Y(_0322_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_mux2_1 _1492_ (.A0(_0321_),
    .A1(_0322_),
    .S(_0271_),
    .X(_0323_));
 sg13g2_o21ai_1 _1493_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_0251_),
    .A2(_0319_));
 sg13g2_xor2_1 _1494_ (.B(_0245_),
    .A(_0243_),
    .X(_0325_));
 sg13g2_xnor2_1 _1495_ (.Y(_0326_),
    .A(_0245_),
    .B(_0276_));
 sg13g2_mux2_1 _1496_ (.A0(_0325_),
    .A1(_0326_),
    .S(_0270_),
    .X(_0327_));
 sg13g2_nand2_2 _1497_ (.Y(_0328_),
    .A(_0294_),
    .B(_0327_));
 sg13g2_xnor2_1 _1498_ (.Y(_0329_),
    .A(_0272_),
    .B(_0278_));
 sg13g2_xor2_1 _1499_ (.B(_0278_),
    .A(_0272_),
    .X(_0330_));
 sg13g2_nor3_2 _1500_ (.A(_0324_),
    .B(_0328_),
    .C(_0329_),
    .Y(_0331_));
 sg13g2_a21o_1 _1501_ (.A2(_0331_),
    .A1(_0240_),
    .B1(net1277),
    .X(_0332_));
 sg13g2_nor2_1 _1502_ (.A(net108),
    .B(_0307_),
    .Y(_0333_));
 sg13g2_a21o_1 _1503_ (.A2(_0332_),
    .A1(net109),
    .B1(_0333_),
    .X(_0028_));
 sg13g2_a21o_1 _1504_ (.A2(_0331_),
    .A1(_0311_),
    .B1(net1284),
    .X(_0334_));
 sg13g2_nor2_1 _1505_ (.A(net108),
    .B(_0312_),
    .Y(_0335_));
 sg13g2_a21o_1 _1506_ (.A2(_0334_),
    .A1(net108),
    .B1(_0335_),
    .X(_0029_));
 sg13g2_a21o_1 _1507_ (.A2(_0331_),
    .A1(_0314_),
    .B1(net1274),
    .X(_0336_));
 sg13g2_nor2_1 _1508_ (.A(net108),
    .B(_0315_),
    .Y(_0337_));
 sg13g2_a21o_1 _1509_ (.A2(_0336_),
    .A1(net108),
    .B1(_0337_),
    .X(_0030_));
 sg13g2_a21o_1 _1510_ (.A2(_0331_),
    .A1(_0317_),
    .B1(net1283),
    .X(_0338_));
 sg13g2_nor2_1 _1511_ (.A(net108),
    .B(_0318_),
    .Y(_0339_));
 sg13g2_a21o_1 _1512_ (.A2(_0338_),
    .A1(net108),
    .B1(_0339_),
    .X(_0031_));
 sg13g2_nor3_2 _1513_ (.A(_0324_),
    .B(_0328_),
    .C(_0330_),
    .Y(_0340_));
 sg13g2_a21o_1 _1514_ (.A2(_0340_),
    .A1(_0240_),
    .B1(net1293),
    .X(_0341_));
 sg13g2_mux2_1 _1515_ (.A0(_0332_),
    .A1(_0341_),
    .S(net108),
    .X(_0024_));
 sg13g2_a21o_1 _1516_ (.A2(_0340_),
    .A1(_0311_),
    .B1(net1319),
    .X(_0342_));
 sg13g2_mux2_1 _1517_ (.A0(_0334_),
    .A1(_0342_),
    .S(net105),
    .X(_0025_));
 sg13g2_a21o_1 _1518_ (.A2(_0340_),
    .A1(_0314_),
    .B1(net1291),
    .X(_0343_));
 sg13g2_mux2_1 _1519_ (.A0(_0336_),
    .A1(_0343_),
    .S(net106),
    .X(_0026_));
 sg13g2_a21o_1 _1520_ (.A2(_0340_),
    .A1(_0317_),
    .B1(net1289),
    .X(_0344_));
 sg13g2_mux2_1 _1521_ (.A0(_0338_),
    .A1(_0344_),
    .S(net106),
    .X(_0027_));
 sg13g2_a21o_2 _1522_ (.A2(_0293_),
    .A1(_0272_),
    .B1(_0327_),
    .X(_0345_));
 sg13g2_nor3_2 _1523_ (.A(_0324_),
    .B(_0329_),
    .C(_0345_),
    .Y(_0346_));
 sg13g2_a21o_1 _1524_ (.A2(_0346_),
    .A1(_0240_),
    .B1(\game_inst.vga_inst.row_buffer[5][0] ),
    .X(_0347_));
 sg13g2_mux2_1 _1525_ (.A0(_0341_),
    .A1(_0347_),
    .S(net106),
    .X(_0020_));
 sg13g2_a21o_1 _1526_ (.A2(_0346_),
    .A1(_0311_),
    .B1(net1312),
    .X(_0348_));
 sg13g2_mux2_1 _1527_ (.A0(_0342_),
    .A1(_0348_),
    .S(net105),
    .X(_0021_));
 sg13g2_a21o_1 _1528_ (.A2(_0346_),
    .A1(_0314_),
    .B1(net1302),
    .X(_0349_));
 sg13g2_mux2_1 _1529_ (.A0(_0343_),
    .A1(_0349_),
    .S(net105),
    .X(_0022_));
 sg13g2_a21o_1 _1530_ (.A2(_0346_),
    .A1(_0317_),
    .B1(net1301),
    .X(_0350_));
 sg13g2_mux2_1 _1531_ (.A0(_0344_),
    .A1(_0350_),
    .S(net105),
    .X(_0023_));
 sg13g2_nor3_2 _1532_ (.A(_0324_),
    .B(_0330_),
    .C(_0345_),
    .Y(_0351_));
 sg13g2_a21o_1 _1533_ (.A2(_0351_),
    .A1(_0240_),
    .B1(net1307),
    .X(_0352_));
 sg13g2_mux2_1 _1534_ (.A0(_0347_),
    .A1(_0352_),
    .S(net106),
    .X(_0016_));
 sg13g2_a21o_1 _1535_ (.A2(_0351_),
    .A1(_0311_),
    .B1(net1309),
    .X(_0353_));
 sg13g2_mux2_1 _1536_ (.A0(_0348_),
    .A1(_0353_),
    .S(net105),
    .X(_0017_));
 sg13g2_a21o_1 _1537_ (.A2(_0351_),
    .A1(_0314_),
    .B1(net1295),
    .X(_0354_));
 sg13g2_mux2_1 _1538_ (.A0(_0349_),
    .A1(_0354_),
    .S(net105),
    .X(_0018_));
 sg13g2_a21o_1 _1539_ (.A2(_0351_),
    .A1(_0317_),
    .B1(net1297),
    .X(_0355_));
 sg13g2_mux2_1 _1540_ (.A0(_0350_),
    .A1(_0355_),
    .S(net105),
    .X(_0019_));
 sg13g2_a21o_2 _1541_ (.A2(_0320_),
    .A1(_0252_),
    .B1(_0323_),
    .X(_0356_));
 sg13g2_nor3_2 _1542_ (.A(_0328_),
    .B(_0329_),
    .C(_0356_),
    .Y(_0357_));
 sg13g2_a21o_1 _1543_ (.A2(_0357_),
    .A1(_0240_),
    .B1(net1304),
    .X(_0358_));
 sg13g2_mux2_1 _1544_ (.A0(_0352_),
    .A1(_0358_),
    .S(net105),
    .X(_0012_));
 sg13g2_a21o_1 _1545_ (.A2(_0357_),
    .A1(_0311_),
    .B1(net1327),
    .X(_0359_));
 sg13g2_mux2_1 _1546_ (.A0(_0353_),
    .A1(_0359_),
    .S(net107),
    .X(_0013_));
 sg13g2_a21o_1 _1547_ (.A2(_0357_),
    .A1(_0314_),
    .B1(net1313),
    .X(_0360_));
 sg13g2_mux2_1 _1548_ (.A0(_0354_),
    .A1(_0360_),
    .S(net107),
    .X(_0014_));
 sg13g2_a21o_1 _1549_ (.A2(_0357_),
    .A1(_0317_),
    .B1(net1299),
    .X(_0361_));
 sg13g2_mux2_1 _1550_ (.A0(_0355_),
    .A1(_0361_),
    .S(net107),
    .X(_0015_));
 sg13g2_nor3_2 _1551_ (.A(_0328_),
    .B(_0330_),
    .C(_0356_),
    .Y(_0362_));
 sg13g2_a21o_1 _1552_ (.A2(_0362_),
    .A1(_0240_),
    .B1(net1317),
    .X(_0363_));
 sg13g2_mux2_1 _1553_ (.A0(_0358_),
    .A1(_0363_),
    .S(net109),
    .X(_0008_));
 sg13g2_a21o_1 _1554_ (.A2(_0362_),
    .A1(_0311_),
    .B1(\game_inst.vga_inst.row_buffer[2][1] ),
    .X(_0364_));
 sg13g2_mux2_1 _1555_ (.A0(_0359_),
    .A1(_0364_),
    .S(net107),
    .X(_0009_));
 sg13g2_a21o_1 _1556_ (.A2(_0362_),
    .A1(_0314_),
    .B1(\game_inst.vga_inst.row_buffer[2][2] ),
    .X(_0365_));
 sg13g2_mux2_1 _1557_ (.A0(_0360_),
    .A1(_0365_),
    .S(net107),
    .X(_0010_));
 sg13g2_a21o_1 _1558_ (.A2(_0362_),
    .A1(_0317_),
    .B1(\game_inst.vga_inst.row_buffer[2][3] ),
    .X(_0366_));
 sg13g2_mux2_1 _1559_ (.A0(_0361_),
    .A1(_0366_),
    .S(net107),
    .X(_0011_));
 sg13g2_nor3_1 _1560_ (.A(_0329_),
    .B(_0345_),
    .C(_0356_),
    .Y(_0367_));
 sg13g2_a21o_1 _1561_ (.A2(_0367_),
    .A1(_0240_),
    .B1(\game_inst.vga_inst.row_buffer[1][0] ),
    .X(_0368_));
 sg13g2_mux2_1 _1562_ (.A0(_0363_),
    .A1(_0368_),
    .S(net109),
    .X(_0004_));
 sg13g2_a21o_1 _1563_ (.A2(_0367_),
    .A1(_0311_),
    .B1(net1325),
    .X(_0369_));
 sg13g2_mux2_1 _1564_ (.A0(_0364_),
    .A1(_0369_),
    .S(net109),
    .X(_0005_));
 sg13g2_a21o_1 _1565_ (.A2(_0367_),
    .A1(_0314_),
    .B1(net1323),
    .X(_0370_));
 sg13g2_mux2_1 _1566_ (.A0(_0365_),
    .A1(_0370_),
    .S(net109),
    .X(_0006_));
 sg13g2_a21o_1 _1567_ (.A2(_0367_),
    .A1(_0317_),
    .B1(net1320),
    .X(_0371_));
 sg13g2_mux2_1 _1568_ (.A0(_0366_),
    .A1(_0371_),
    .S(net109),
    .X(_0007_));
 sg13g2_or2_1 _1569_ (.X(uo_out[5]),
    .B(\game_inst.vga_inst.color[2] ),
    .A(\game_inst.vga_inst.color[3] ));
 sg13g2_or2_1 _1570_ (.X(uo_out[4]),
    .B(\game_inst.vga_inst.color[3] ),
    .A(\game_inst.vga_inst.color[1] ));
 sg13g2_nor2b_1 _1571_ (.A(net127),
    .B_N(net124),
    .Y(_0372_));
 sg13g2_and4_1 _1572_ (.A(\game_inst.vga_inst.px[8] ),
    .B(_0177_),
    .C(net111),
    .D(_0372_),
    .X(_0373_));
 sg13g2_nand4_1 _1573_ (.B(_0177_),
    .C(net112),
    .A(net1338),
    .Y(_0374_),
    .D(_0372_));
 sg13g2_nor2_2 _1574_ (.A(net132),
    .B(_0373_),
    .Y(_0375_));
 sg13g2_nand2_2 _1575_ (.Y(_0376_),
    .A(net134),
    .B(_0374_));
 sg13g2_nor2_1 _1576_ (.A(net1132),
    .B(net132),
    .Y(_0039_));
 sg13g2_o21ai_1 _1577_ (.B1(_0375_),
    .Y(_0377_),
    .A1(net1132),
    .A2(net1133));
 sg13g2_a21oi_1 _1578_ (.A1(net1132),
    .A2(net1133),
    .Y(_0040_),
    .B1(_0377_));
 sg13g2_a21oi_1 _1579_ (.A1(net1132),
    .A2(net1133),
    .Y(_0378_),
    .B1(net1159));
 sg13g2_nor3_1 _1580_ (.A(net132),
    .B(_0218_),
    .C(_0378_),
    .Y(_0041_));
 sg13g2_o21ai_1 _1581_ (.B1(net134),
    .Y(_0379_),
    .A1(net1255),
    .A2(_0218_));
 sg13g2_nor2_1 _1582_ (.A(_0219_),
    .B(_0379_),
    .Y(_0042_));
 sg13g2_o21ai_1 _1583_ (.B1(net134),
    .Y(_0380_),
    .A1(net1285),
    .A2(_0219_));
 sg13g2_nor2_1 _1584_ (.A(net112),
    .B(_0380_),
    .Y(_0043_));
 sg13g2_o21ai_1 _1585_ (.B1(_0375_),
    .Y(_0381_),
    .A1(_0166_),
    .A2(net110));
 sg13g2_a21oi_1 _1586_ (.A1(_0166_),
    .A2(net110),
    .Y(_0044_),
    .B1(_0381_));
 sg13g2_a21oi_1 _1587_ (.A1(net1238),
    .A2(net112),
    .Y(_0382_),
    .B1(net128));
 sg13g2_and2_1 _1588_ (.A(_0178_),
    .B(net112),
    .X(_0383_));
 sg13g2_nor3_1 _1589_ (.A(_0376_),
    .B(net1239),
    .C(_0383_),
    .Y(_0045_));
 sg13g2_nor2_1 _1590_ (.A(net126),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_and4_1 _1591_ (.A(net1238),
    .B(net126),
    .C(net128),
    .D(net112),
    .X(_0385_));
 sg13g2_nor3_1 _1592_ (.A(_0376_),
    .B(net1333),
    .C(_0385_),
    .Y(_0046_));
 sg13g2_o21ai_1 _1593_ (.B1(_0167_),
    .Y(_0386_),
    .A1(net110),
    .A2(_0281_));
 sg13g2_nand2_1 _1594_ (.Y(_0387_),
    .A(net125),
    .B(_0385_));
 sg13g2_and3_1 _1595_ (.X(_0047_),
    .A(_0375_),
    .B(_0386_),
    .C(_0387_));
 sg13g2_xor2_1 _1596_ (.B(_0387_),
    .A(net124),
    .X(_0388_));
 sg13g2_nor2_1 _1597_ (.A(_0376_),
    .B(_0388_),
    .Y(_0048_));
 sg13g2_nor2_2 _1598_ (.A(net132),
    .B(net6),
    .Y(_0389_));
 sg13g2_nand2b_1 _1599_ (.Y(_0390_),
    .B(net136),
    .A_N(net6));
 sg13g2_nand4_1 _1600_ (.B(_0155_),
    .C(\game_inst.snake_inst.pos[5] ),
    .A(net1146),
    .Y(_0391_),
    .D(\game_inst.snake_inst.pos[6] ));
 sg13g2_nor2b_1 _1601_ (.A(\game_inst.snake_inst.pos[2] ),
    .B_N(\game_inst.snake_inst.pos[3] ),
    .Y(_0392_));
 sg13g2_nand4_1 _1602_ (.B(net121),
    .C(_0236_),
    .A(\game_inst.tick ),
    .Y(_0393_),
    .D(_0392_));
 sg13g2_nor2_2 _1603_ (.A(_0391_),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_or2_1 _1604_ (.X(_0395_),
    .B(_0393_),
    .A(_0391_));
 sg13g2_nand2_1 _1605_ (.Y(_0396_),
    .A(\game_inst.tick ),
    .B(_0236_));
 sg13g2_nand2_1 _1606_ (.Y(_0397_),
    .A(net121),
    .B(_0392_));
 sg13g2_nor3_1 _1607_ (.A(_0391_),
    .B(_0396_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_o21ai_1 _1608_ (.B1(net113),
    .Y(_0049_),
    .A1(net1162),
    .A2(_0394_));
 sg13g2_nand3b_1 _1609_ (.B(\game_inst.snake_inst.pos[0] ),
    .C(_0392_),
    .Y(_0399_),
    .A_N(\game_inst.snake_inst.pos[1] ));
 sg13g2_or2_1 _1610_ (.X(_0400_),
    .B(_0399_),
    .A(_0391_));
 sg13g2_and2_1 _1611_ (.A(net104),
    .B(net101),
    .X(_0401_));
 sg13g2_nand2_2 _1612_ (.Y(_0402_),
    .A(_0395_),
    .B(net101));
 sg13g2_and2_1 _1613_ (.A(net1303),
    .B(net1162),
    .X(_0403_));
 sg13g2_and2_1 _1614_ (.A(net1218),
    .B(_0403_),
    .X(_0404_));
 sg13g2_xnor2_1 _1615_ (.Y(_0405_),
    .A(net1282),
    .B(_0404_));
 sg13g2_o21ai_1 _1616_ (.B1(net113),
    .Y(_0050_),
    .A1(_0402_),
    .A2(_0405_));
 sg13g2_and3_2 _1617_ (.X(_0406_),
    .A(net1282),
    .B(net1190),
    .C(_0404_));
 sg13g2_a21oi_1 _1618_ (.A1(net1306),
    .A2(_0406_),
    .Y(_0407_),
    .B1(_0402_));
 sg13g2_o21ai_1 _1619_ (.B1(_0407_),
    .Y(_0408_),
    .A1(net1306),
    .A2(_0406_));
 sg13g2_nand2_1 _1620_ (.Y(_0051_),
    .A(_0389_),
    .B(_0408_));
 sg13g2_nand3_1 _1621_ (.B(net1252),
    .C(_0406_),
    .A(net1306),
    .Y(_0409_));
 sg13g2_a21oi_1 _1622_ (.A1(\game_inst.snake_inst.pos[5] ),
    .A2(_0406_),
    .Y(_0410_),
    .B1(net1252));
 sg13g2_nand2_1 _1623_ (.Y(_0411_),
    .A(_0401_),
    .B(_0409_));
 sg13g2_o21ai_1 _1624_ (.B1(net114),
    .Y(_0052_),
    .A1(net1253),
    .A2(_0411_));
 sg13g2_xnor2_1 _1625_ (.Y(_0412_),
    .A(_0154_),
    .B(_0409_));
 sg13g2_o21ai_1 _1626_ (.B1(net113),
    .Y(_0053_),
    .A1(net99),
    .A2(_0412_));
 sg13g2_o21ai_1 _1627_ (.B1(net115),
    .Y(_0413_),
    .A1(_0140_),
    .A2(net104));
 sg13g2_a21o_1 _1628_ (.A2(net104),
    .A1(net1155),
    .B1(_0413_),
    .X(_0054_));
 sg13g2_nor2_1 _1629_ (.A(_0139_),
    .B(net103),
    .Y(_0414_));
 sg13g2_nand2_1 _1630_ (.Y(_0415_),
    .A(net119),
    .B(_0394_));
 sg13g2_and2_1 _1631_ (.A(net119),
    .B(_0398_),
    .X(_0416_));
 sg13g2_nand2_1 _1632_ (.Y(_0417_),
    .A(net115),
    .B(_0415_));
 sg13g2_a21o_1 _1633_ (.A2(net104),
    .A1(net1177),
    .B1(_0417_),
    .X(_0055_));
 sg13g2_mux2_1 _1634_ (.A0(net1207),
    .A1(_0368_),
    .S(net112),
    .X(_0056_));
 sg13g2_mux2_1 _1635_ (.A0(net1231),
    .A1(_0369_),
    .S(net111),
    .X(_0057_));
 sg13g2_mux2_1 _1636_ (.A0(net1226),
    .A1(_0370_),
    .S(net111),
    .X(_0058_));
 sg13g2_mux2_1 _1637_ (.A0(net1228),
    .A1(_0371_),
    .S(net111),
    .X(_0059_));
 sg13g2_nand4_1 _1638_ (.B(_0149_),
    .C(\game_inst.vga_inst.py[3] ),
    .A(\game_inst.vga_inst.py[9] ),
    .Y(_0418_),
    .D(\game_inst.vga_inst.py[2] ));
 sg13g2_nor4_1 _1639_ (.A(\game_inst.vga_inst.py[4] ),
    .B(\game_inst.vga_inst.py[1] ),
    .C(\game_inst.vga_inst.py[0] ),
    .D(_0418_),
    .Y(_0419_));
 sg13g2_a21oi_1 _1640_ (.A1(_0173_),
    .A2(_0419_),
    .Y(_0420_),
    .B1(_0374_));
 sg13g2_o21ai_1 _1641_ (.B1(net134),
    .Y(_0421_),
    .A1(net1160),
    .A2(_0420_));
 sg13g2_a21oi_1 _1642_ (.A1(net1160),
    .A2(_0373_),
    .Y(_0060_),
    .B1(_0421_));
 sg13g2_a21oi_1 _1643_ (.A1(net1160),
    .A2(_0373_),
    .Y(_0422_),
    .B1(net1174));
 sg13g2_o21ai_1 _1644_ (.B1(net134),
    .Y(_0423_),
    .A1(_0253_),
    .A2(_0374_));
 sg13g2_nor2_1 _1645_ (.A(net1175),
    .B(_0423_),
    .Y(_0061_));
 sg13g2_nand2_1 _1646_ (.Y(_0424_),
    .A(net1213),
    .B(_0375_));
 sg13g2_nand2_2 _1647_ (.Y(_0425_),
    .A(net134),
    .B(_0420_));
 sg13g2_nand3_1 _1648_ (.B(net1174),
    .C(net1160),
    .A(net1213),
    .Y(_0426_));
 sg13g2_xor2_1 _1649_ (.B(_0253_),
    .A(net1213),
    .X(_0427_));
 sg13g2_o21ai_1 _1650_ (.B1(_0424_),
    .Y(_0062_),
    .A1(_0425_),
    .A2(_0427_));
 sg13g2_nor2b_1 _1651_ (.A(net1209),
    .B_N(_0426_),
    .Y(_0428_));
 sg13g2_nor3_1 _1652_ (.A(_0254_),
    .B(_0425_),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_a21o_1 _1653_ (.A2(_0375_),
    .A1(net1209),
    .B1(_0429_),
    .X(_0063_));
 sg13g2_a21oi_1 _1654_ (.A1(net1210),
    .A2(_0373_),
    .Y(_0430_),
    .B1(net1157));
 sg13g2_nor2_1 _1655_ (.A(_0258_),
    .B(_0374_),
    .Y(_0431_));
 sg13g2_nor3_1 _1656_ (.A(net132),
    .B(net1211),
    .C(_0431_),
    .Y(_0064_));
 sg13g2_nor2_1 _1657_ (.A(net1266),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_nor2_1 _1658_ (.A(_0255_),
    .B(_0374_),
    .Y(_0433_));
 sg13g2_nor3_1 _1659_ (.A(net132),
    .B(net1267),
    .C(_0433_),
    .Y(_0065_));
 sg13g2_or2_1 _1660_ (.X(_0434_),
    .B(_0433_),
    .A(net1337));
 sg13g2_nand2_1 _1661_ (.Y(_0435_),
    .A(net1337),
    .B(_0433_));
 sg13g2_and3_1 _1662_ (.X(_0066_),
    .A(net134),
    .B(_0434_),
    .C(_0435_));
 sg13g2_a221oi_1 _1663_ (.B2(_0147_),
    .C1(net132),
    .B1(_0435_),
    .A1(_0261_),
    .Y(_0067_),
    .A2(_0373_));
 sg13g2_a21oi_1 _1664_ (.A1(_0261_),
    .A2(_0373_),
    .Y(_0436_),
    .B1(net1214));
 sg13g2_nand2_1 _1665_ (.Y(_0437_),
    .A(net1214),
    .B(_0261_));
 sg13g2_inv_1 _1666_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nor2_1 _1667_ (.A(_0374_),
    .B(_0437_),
    .Y(_0439_));
 sg13g2_nor3_1 _1668_ (.A(net132),
    .B(net1215),
    .C(_0439_),
    .Y(_0068_));
 sg13g2_o21ai_1 _1669_ (.B1(_0376_),
    .Y(_0440_),
    .A1(_0425_),
    .A2(_0438_));
 sg13g2_nor3_1 _1670_ (.A(net1200),
    .B(_0425_),
    .C(_0437_),
    .Y(_0441_));
 sg13g2_a21o_1 _1671_ (.A2(_0440_),
    .A1(net1200),
    .B1(_0441_),
    .X(_0069_));
 sg13g2_xor2_1 _1672_ (.B(\game_inst.apple_inst.i_snake_x[3] ),
    .A(\game_inst.head_x[3] ),
    .X(_0442_));
 sg13g2_xor2_1 _1673_ (.B(\game_inst.apple_inst.i_snake_y[0] ),
    .A(net120),
    .X(_0443_));
 sg13g2_xor2_1 _1674_ (.B(\game_inst.apple_inst.i_snake_x[0] ),
    .A(\game_inst.head_x[0] ),
    .X(_0444_));
 sg13g2_xnor2_1 _1675_ (.Y(_0445_),
    .A(\game_inst.head_y[2] ),
    .B(\game_inst.apple_inst.i_snake_y[2] ));
 sg13g2_xnor2_1 _1676_ (.Y(_0446_),
    .A(\game_inst.head_y[1] ),
    .B(\game_inst.apple_inst.i_snake_y[1] ));
 sg13g2_xor2_1 _1677_ (.B(\game_inst.apple_inst.i_snake_y[3] ),
    .A(\game_inst.head_y[3] ),
    .X(_0447_));
 sg13g2_xor2_1 _1678_ (.B(net117),
    .A(\game_inst.head_x[1] ),
    .X(_0448_));
 sg13g2_xor2_1 _1679_ (.B(\game_inst.apple_inst.i_snake_x[4] ),
    .A(\game_inst.head_x[4] ),
    .X(_0449_));
 sg13g2_xor2_1 _1680_ (.B(net116),
    .A(\game_inst.head_x[2] ),
    .X(_0450_));
 sg13g2_nor4_1 _1681_ (.A(_0447_),
    .B(_0448_),
    .C(_0449_),
    .D(_0450_),
    .Y(_0451_));
 sg13g2_nand3_1 _1682_ (.B(_0446_),
    .C(_0451_),
    .A(_0445_),
    .Y(_0452_));
 sg13g2_nor4_1 _1683_ (.A(_0442_),
    .B(_0443_),
    .C(_0444_),
    .D(_0452_),
    .Y(_0453_));
 sg13g2_a21oi_1 _1684_ (.A1(\game_inst.head_x[4] ),
    .A2(\game_inst.head_x[1] ),
    .Y(_0454_),
    .B1(_0138_));
 sg13g2_nor2_1 _1685_ (.A(\game_inst.head_x[4] ),
    .B(\game_inst.head_x[1] ),
    .Y(_0455_));
 sg13g2_nor2_1 _1686_ (.A(\game_inst.head_x[0] ),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nor4_1 _1687_ (.A(\game_inst.head_x[3] ),
    .B(\game_inst.head_x[2] ),
    .C(_0454_),
    .D(_0456_),
    .Y(_0457_));
 sg13g2_nand3_1 _1688_ (.B(\game_inst.head_y[2] ),
    .C(\game_inst.head_y[1] ),
    .A(\game_inst.head_y[3] ),
    .Y(_0458_));
 sg13g2_or3_1 _1689_ (.A(\game_inst.head_y[3] ),
    .B(\game_inst.head_y[2] ),
    .C(\game_inst.head_y[1] ),
    .X(_0459_));
 sg13g2_a21oi_1 _1690_ (.A1(_0458_),
    .A2(_0459_),
    .Y(_0460_),
    .B1(net120));
 sg13g2_nor3_1 _1691_ (.A(_0453_),
    .B(_0457_),
    .C(_0460_),
    .Y(_0461_));
 sg13g2_nor3_1 _1692_ (.A(_0136_),
    .B(_0238_),
    .C(_0461_),
    .Y(_0462_));
 sg13g2_o21ai_1 _1693_ (.B1(net113),
    .Y(_0463_),
    .A1(net1134),
    .A2(_0462_));
 sg13g2_inv_1 _1694_ (.Y(_0070_),
    .A(_0463_));
 sg13g2_nand3_1 _1695_ (.B(\game_inst.apple_inst.apple_y[2] ),
    .C(\game_inst.apple_inst.apple_y[3] ),
    .A(\game_inst.apple_inst.apple_y[1] ),
    .Y(_0464_));
 sg13g2_nand2_1 _1696_ (.Y(_0465_),
    .A(\game_inst.apple_inst.apple_x[0] ),
    .B(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_nand3b_1 _1697_ (.B(_0160_),
    .C(_0465_),
    .Y(_0466_),
    .A_N(\game_inst.apple_inst.apple_x[2] ));
 sg13g2_xor2_1 _1698_ (.B(\game_inst.apple_inst.i_snake_x[4] ),
    .A(\game_inst.apple_inst.apple_x[4] ),
    .X(_0467_));
 sg13g2_xor2_1 _1699_ (.B(\game_inst.apple_inst.apple_y[3] ),
    .A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(_0468_));
 sg13g2_xor2_1 _1700_ (.B(\game_inst.apple_inst.apple_x[2] ),
    .A(net116),
    .X(_0469_));
 sg13g2_xor2_1 _1701_ (.B(net118),
    .A(\game_inst.apple_inst.apple_x[0] ),
    .X(_0470_));
 sg13g2_nand2b_1 _1702_ (.Y(_0471_),
    .B(net117),
    .A_N(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_a221oi_1 _1703_ (.B2(_0160_),
    .C1(_0469_),
    .B1(\game_inst.apple_inst.i_snake_x[3] ),
    .A1(_0158_),
    .Y(_0472_),
    .A2(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_a221oi_1 _1704_ (.B2(_0165_),
    .C1(_0467_),
    .B1(\game_inst.apple_inst.i_snake_y[1] ),
    .A1(_0162_),
    .Y(_0473_),
    .A2(\game_inst.apple_inst.i_snake_y[0] ));
 sg13g2_a221oi_1 _1705_ (.B2(\game_inst.apple_inst.apple_y[1] ),
    .C1(_0470_),
    .B1(_0164_),
    .A1(\game_inst.apple_inst.apple_y[0] ),
    .Y(_0474_),
    .A2(_0163_));
 sg13g2_xor2_1 _1706_ (.B(\game_inst.apple_inst.apple_y[2] ),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .X(_0475_));
 sg13g2_o21ai_1 _1707_ (.B1(_0471_),
    .Y(_0476_),
    .A1(\game_inst.apple_inst.i_snake_x[3] ),
    .A2(_0160_));
 sg13g2_nor3_1 _1708_ (.A(_0468_),
    .B(_0475_),
    .C(_0476_),
    .Y(_0477_));
 sg13g2_and4_1 _1709_ (.A(_0472_),
    .B(_0473_),
    .C(_0474_),
    .D(_0477_),
    .X(_0478_));
 sg13g2_a22oi_1 _1710_ (.Y(_0479_),
    .B1(_0478_),
    .B2(\game_inst.apple_inst.i_snake_valid ),
    .A2(_0466_),
    .A1(\game_inst.apple_inst.apple_x[4] ));
 sg13g2_nand3_1 _1711_ (.B(_0238_),
    .C(_0478_),
    .A(net121),
    .Y(_0480_));
 sg13g2_and4_1 _1712_ (.A(net113),
    .B(_0464_),
    .C(_0479_),
    .D(_0480_),
    .X(_0481_));
 sg13g2_nand2_1 _1713_ (.Y(_0482_),
    .A(\game_inst.apple_inst.apple_x[0] ),
    .B(net96));
 sg13g2_o21ai_1 _1714_ (.B1(_0482_),
    .Y(_0071_),
    .A1(_0146_),
    .A2(net96));
 sg13g2_nand2_1 _1715_ (.Y(_0483_),
    .A(net1183),
    .B(net97));
 sg13g2_o21ai_1 _1716_ (.B1(_0483_),
    .Y(_0072_),
    .A1(_0145_),
    .A2(net96));
 sg13g2_nand2_1 _1717_ (.Y(_0484_),
    .A(net1193),
    .B(net97));
 sg13g2_o21ai_1 _1718_ (.B1(_0484_),
    .Y(_0073_),
    .A1(_0144_),
    .A2(net96));
 sg13g2_nor2_1 _1719_ (.A(net1167),
    .B(net96),
    .Y(_0485_));
 sg13g2_a21oi_1 _1720_ (.A1(_0160_),
    .A2(net97),
    .Y(_0074_),
    .B1(_0485_));
 sg13g2_mux2_1 _1721_ (.A0(net1205),
    .A1(\game_inst.apple_inst.apple_x[4] ),
    .S(net97),
    .X(_0075_));
 sg13g2_a21oi_1 _1722_ (.A1(net1152),
    .A2(_0238_),
    .Y(_0486_),
    .B1(net121));
 sg13g2_nor2b_1 _1723_ (.A(net1153),
    .B_N(net98),
    .Y(_0076_));
 sg13g2_o21ai_1 _1724_ (.B1(net98),
    .Y(_0487_),
    .A1(net1152),
    .A2(_0238_));
 sg13g2_inv_1 _1725_ (.Y(_0077_),
    .A(_0487_));
 sg13g2_o21ai_1 _1726_ (.B1(net1230),
    .Y(_0488_),
    .A1(net2),
    .A2(net1));
 sg13g2_nand2b_1 _1727_ (.Y(_0489_),
    .B(net1230),
    .A_N(net1203));
 sg13g2_nand3_1 _1728_ (.B(_0488_),
    .C(_0489_),
    .A(net4),
    .Y(_0490_));
 sg13g2_nand2_1 _1729_ (.Y(_0491_),
    .A(\game_inst.control_inst.backwards[1] ),
    .B(\game_inst.control_inst.i_head_dir[0] ));
 sg13g2_and3_1 _1730_ (.X(_0492_),
    .A(net3),
    .B(_0488_),
    .C(_0491_));
 sg13g2_nor2_1 _1731_ (.A(net119),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nand2_1 _1732_ (.Y(_0494_),
    .A(_0490_),
    .B(_0493_));
 sg13g2_nor2_1 _1733_ (.A(net4),
    .B(net3),
    .Y(_0495_));
 sg13g2_nor3_1 _1734_ (.A(net1341),
    .B(net4),
    .C(net3),
    .Y(_0496_));
 sg13g2_o21ai_1 _1735_ (.B1(net1),
    .Y(_0497_),
    .A1(net1230),
    .A2(_0496_));
 sg13g2_a21oi_1 _1736_ (.A1(net1341),
    .A2(_0495_),
    .Y(_0498_),
    .B1(net1230));
 sg13g2_nor2_1 _1737_ (.A(_0168_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_o21ai_1 _1738_ (.B1(_0497_),
    .Y(_0500_),
    .A1(_0168_),
    .A2(_0498_));
 sg13g2_o21ai_1 _1739_ (.B1(_0494_),
    .Y(_0501_),
    .A1(_0139_),
    .A2(_0500_));
 sg13g2_a21oi_1 _1740_ (.A1(_0140_),
    .A2(_0490_),
    .Y(_0502_),
    .B1(_0492_));
 sg13g2_o21ai_1 _1741_ (.B1(_0497_),
    .Y(_0503_),
    .A1(_0499_),
    .A2(_0502_));
 sg13g2_xnor2_1 _1742_ (.Y(_0504_),
    .A(_0140_),
    .B(_0503_));
 sg13g2_a21o_1 _1743_ (.A2(_0504_),
    .A1(_0501_),
    .B1(net121),
    .X(_0505_));
 sg13g2_nand3_1 _1744_ (.B(_0501_),
    .C(_0504_),
    .A(net121),
    .Y(_0506_));
 sg13g2_nand3_1 _1745_ (.B(_0505_),
    .C(_0506_),
    .A(net98),
    .Y(_0507_));
 sg13g2_xor2_1 _1746_ (.B(net1188),
    .A(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .X(_0508_));
 sg13g2_a21oi_1 _1747_ (.A1(net94),
    .A2(net1189),
    .Y(_0509_),
    .B1(net133));
 sg13g2_o21ai_1 _1748_ (.B1(_0509_),
    .Y(_0078_),
    .A1(_0146_),
    .A2(net94));
 sg13g2_a21oi_1 _1749_ (.A1(net1172),
    .A2(net95),
    .Y(_0510_),
    .B1(net133));
 sg13g2_o21ai_1 _1750_ (.B1(_0510_),
    .Y(_0079_),
    .A1(_0145_),
    .A2(net94));
 sg13g2_a21oi_1 _1751_ (.A1(net1195),
    .A2(net95),
    .Y(_0511_),
    .B1(net133));
 sg13g2_o21ai_1 _1752_ (.B1(_0511_),
    .Y(_0080_),
    .A1(_0144_),
    .A2(net94));
 sg13g2_o21ai_1 _1753_ (.B1(net135),
    .Y(_0512_),
    .A1(net1167),
    .A2(net94));
 sg13g2_a21oi_1 _1754_ (.A1(_0144_),
    .A2(net94),
    .Y(_0081_),
    .B1(_0512_));
 sg13g2_o21ai_1 _1755_ (.B1(net135),
    .Y(_0513_),
    .A1(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .A2(net94));
 sg13g2_a21oi_1 _1756_ (.A1(_0143_),
    .A2(net94),
    .Y(_0082_),
    .B1(_0513_));
 sg13g2_nand2_1 _1757_ (.Y(_0514_),
    .A(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .B(_0507_));
 sg13g2_a21oi_1 _1758_ (.A1(net1140),
    .A2(_0514_),
    .Y(_0515_),
    .B1(net133));
 sg13g2_o21ai_1 _1759_ (.B1(_0515_),
    .Y(_0083_),
    .A1(net1140),
    .A2(_0514_));
 sg13g2_o21ai_1 _1760_ (.B1(net135),
    .Y(_0516_),
    .A1(_0142_),
    .A2(net95));
 sg13g2_a21o_1 _1761_ (.A2(_0507_),
    .A1(net1140),
    .B1(_0516_),
    .X(_0084_));
 sg13g2_o21ai_1 _1762_ (.B1(net135),
    .Y(_0517_),
    .A1(net1194),
    .A2(net95));
 sg13g2_a21oi_1 _1763_ (.A1(_0142_),
    .A2(net95),
    .Y(_0085_),
    .B1(_0517_));
 sg13g2_a21oi_1 _1764_ (.A1(net1194),
    .A2(net95),
    .Y(_0518_),
    .B1(net133));
 sg13g2_o21ai_1 _1765_ (.B1(_0518_),
    .Y(_0086_),
    .A1(_0141_),
    .A2(net95));
 sg13g2_a21o_1 _1766_ (.A2(net104),
    .A1(net1203),
    .B1(_0413_),
    .X(_0087_));
 sg13g2_a21o_1 _1767_ (.A2(net104),
    .A1(net1230),
    .B1(_0417_),
    .X(_0088_));
 sg13g2_nand2_1 _1768_ (.Y(_0519_),
    .A(net1249),
    .B(net102));
 sg13g2_nor2_2 _1769_ (.A(net119),
    .B(net102),
    .Y(_0520_));
 sg13g2_o21ai_1 _1770_ (.B1(net1249),
    .Y(_0521_),
    .A1(net119),
    .A2(net102));
 sg13g2_nand2_1 _1771_ (.Y(_0522_),
    .A(_0138_),
    .B(_0415_));
 sg13g2_nand2_1 _1772_ (.Y(_0523_),
    .A(_0521_),
    .B(_0522_));
 sg13g2_and2_1 _1773_ (.A(_0139_),
    .B(_0398_),
    .X(_0524_));
 sg13g2_a21oi_1 _1774_ (.A1(_0519_),
    .A2(_0523_),
    .Y(_0089_),
    .B1(net130));
 sg13g2_nand2_2 _1775_ (.Y(_0525_),
    .A(net119),
    .B(\game_inst.control_inst.dir[0] ));
 sg13g2_and2_1 _1776_ (.A(\game_inst.head_x[1] ),
    .B(_0525_),
    .X(_0526_));
 sg13g2_xor2_1 _1777_ (.B(_0525_),
    .A(\game_inst.head_x[1] ),
    .X(_0527_));
 sg13g2_and2_1 _1778_ (.A(\game_inst.head_x[0] ),
    .B(_0527_),
    .X(_0528_));
 sg13g2_xnor2_1 _1779_ (.Y(_0529_),
    .A(_0138_),
    .B(_0527_));
 sg13g2_a22oi_1 _1780_ (.Y(_0530_),
    .B1(_0529_),
    .B2(_0414_),
    .A2(_0520_),
    .A1(net1322));
 sg13g2_nand2_1 _1781_ (.Y(_0531_),
    .A(net1322),
    .B(net102));
 sg13g2_nand3_1 _1782_ (.B(_0530_),
    .C(_0531_),
    .A(net115),
    .Y(_0090_));
 sg13g2_nand2_1 _1783_ (.Y(_0532_),
    .A(net1265),
    .B(net102));
 sg13g2_nand2_1 _1784_ (.Y(_0533_),
    .A(\game_inst.head_x[2] ),
    .B(_0525_));
 sg13g2_xor2_1 _1785_ (.B(_0525_),
    .A(\game_inst.head_x[2] ),
    .X(_0534_));
 sg13g2_nor3_1 _1786_ (.A(_0526_),
    .B(_0528_),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_o21ai_1 _1787_ (.B1(_0534_),
    .Y(_0536_),
    .A1(_0526_),
    .A2(_0528_));
 sg13g2_nor2b_1 _1788_ (.A(_0535_),
    .B_N(_0536_),
    .Y(_0537_));
 sg13g2_a22oi_1 _1789_ (.Y(_0538_),
    .B1(_0537_),
    .B2(_0416_),
    .A2(_0524_),
    .A1(net1265));
 sg13g2_a21oi_1 _1790_ (.A1(_0532_),
    .A2(_0538_),
    .Y(_0091_),
    .B1(net130));
 sg13g2_and2_1 _1791_ (.A(_0533_),
    .B(_0536_),
    .X(_0539_));
 sg13g2_xnor2_1 _1792_ (.Y(_0540_),
    .A(\game_inst.head_x[3] ),
    .B(_0539_));
 sg13g2_xnor2_1 _1793_ (.Y(_0541_),
    .A(\game_inst.control_inst.dir[0] ),
    .B(_0540_));
 sg13g2_a22oi_1 _1794_ (.Y(_0542_),
    .B1(_0541_),
    .B2(_0414_),
    .A2(_0520_),
    .A1(net1280));
 sg13g2_nand2_1 _1795_ (.Y(_0543_),
    .A(net1280),
    .B(net102));
 sg13g2_nand3_1 _1796_ (.B(_0542_),
    .C(_0543_),
    .A(net115),
    .Y(_0092_));
 sg13g2_nand2_1 _1797_ (.Y(_0544_),
    .A(net1261),
    .B(net102));
 sg13g2_and4_1 _1798_ (.A(_0137_),
    .B(net119),
    .C(_0140_),
    .D(_0539_),
    .X(_0545_));
 sg13g2_nor3_1 _1799_ (.A(_0137_),
    .B(_0525_),
    .C(_0536_),
    .Y(_0546_));
 sg13g2_o21ai_1 _1800_ (.B1(net1261),
    .Y(_0547_),
    .A1(_0545_),
    .A2(_0546_));
 sg13g2_nor3_1 _1801_ (.A(net1261),
    .B(_0545_),
    .C(_0546_),
    .Y(_0548_));
 sg13g2_nor2_1 _1802_ (.A(net102),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_nand2_1 _1803_ (.Y(_0550_),
    .A(_0547_),
    .B(_0549_));
 sg13g2_a21oi_1 _1804_ (.A1(_0544_),
    .A2(_0550_),
    .Y(_0093_),
    .B1(net130));
 sg13g2_nand2_1 _1805_ (.Y(_0551_),
    .A(net120),
    .B(_0415_));
 sg13g2_o21ai_1 _1806_ (.B1(_0551_),
    .Y(_0552_),
    .A1(net120),
    .A2(_0520_));
 sg13g2_a21oi_1 _1807_ (.A1(net1257),
    .A2(net103),
    .Y(_0553_),
    .B1(net130));
 sg13g2_nand2_1 _1808_ (.Y(_0094_),
    .A(_0552_),
    .B(_0553_));
 sg13g2_nand2_1 _1809_ (.Y(_0554_),
    .A(_0139_),
    .B(\game_inst.control_inst.dir[0] ));
 sg13g2_and2_1 _1810_ (.A(\game_inst.head_y[1] ),
    .B(_0554_),
    .X(_0555_));
 sg13g2_xor2_1 _1811_ (.B(_0554_),
    .A(\game_inst.head_y[1] ),
    .X(_0556_));
 sg13g2_xor2_1 _1812_ (.B(_0556_),
    .A(net1257),
    .X(_0557_));
 sg13g2_a22oi_1 _1813_ (.Y(_0558_),
    .B1(_0520_),
    .B2(_0557_),
    .A2(_0414_),
    .A1(net1287));
 sg13g2_nand2_1 _1814_ (.Y(_0559_),
    .A(net1287),
    .B(net103));
 sg13g2_nand3_1 _1815_ (.B(_0558_),
    .C(_0559_),
    .A(net115),
    .Y(_0095_));
 sg13g2_nand2_1 _1816_ (.Y(_0560_),
    .A(net1288),
    .B(net103));
 sg13g2_a21oi_1 _1817_ (.A1(net120),
    .A2(_0556_),
    .Y(_0561_),
    .B1(_0555_));
 sg13g2_xor2_1 _1818_ (.B(_0554_),
    .A(\game_inst.head_y[2] ),
    .X(_0562_));
 sg13g2_xnor2_1 _1819_ (.Y(_0563_),
    .A(_0561_),
    .B(_0562_));
 sg13g2_a22oi_1 _1820_ (.Y(_0564_),
    .B1(_0524_),
    .B2(_0563_),
    .A2(_0416_),
    .A1(net1288));
 sg13g2_nand3_1 _1821_ (.B(_0560_),
    .C(_0564_),
    .A(net115),
    .Y(_0096_));
 sg13g2_nand2b_1 _1822_ (.Y(_0565_),
    .B(\game_inst.control_inst.dir[0] ),
    .A_N(net120));
 sg13g2_a21oi_1 _1823_ (.A1(net120),
    .A2(_0140_),
    .Y(_0566_),
    .B1(net119));
 sg13g2_and4_1 _1824_ (.A(_0556_),
    .B(_0562_),
    .C(_0565_),
    .D(_0566_),
    .X(_0567_));
 sg13g2_nor2_1 _1825_ (.A(net1339),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_a21oi_1 _1826_ (.A1(\game_inst.head_y[3] ),
    .A2(_0567_),
    .Y(_0569_),
    .B1(net103));
 sg13g2_nor2b_1 _1827_ (.A(_0568_),
    .B_N(_0569_),
    .Y(_0570_));
 sg13g2_a21o_1 _1828_ (.A2(net103),
    .A1(net1339),
    .B1(_0570_),
    .X(_0571_));
 sg13g2_and2_1 _1829_ (.A(net115),
    .B(_0571_),
    .X(_0097_));
 sg13g2_nor2_1 _1830_ (.A(net130),
    .B(_0503_),
    .Y(_0098_));
 sg13g2_a21oi_1 _1831_ (.A1(_0490_),
    .A2(_0493_),
    .Y(_0572_),
    .B1(_0500_));
 sg13g2_nand2b_1 _1832_ (.Y(_0099_),
    .B(net115),
    .A_N(_0572_));
 sg13g2_nor2_2 _1833_ (.A(net122),
    .B(net99),
    .Y(_0573_));
 sg13g2_a22oi_1 _1834_ (.Y(_0574_),
    .B1(net99),
    .B2(_0519_),
    .A2(net100),
    .A1(net1335));
 sg13g2_a21oi_1 _1835_ (.A1(_0521_),
    .A2(_0522_),
    .Y(_0575_),
    .B1(_0574_));
 sg13g2_xnor2_1 _1836_ (.Y(_0100_),
    .A(_0573_),
    .B(_0575_));
 sg13g2_nor2_1 _1837_ (.A(net100),
    .B(_0531_),
    .Y(_0576_));
 sg13g2_nand2_2 _1838_ (.Y(_0577_),
    .A(\game_inst.pos_dir[0] ),
    .B(net123));
 sg13g2_nor2_1 _1839_ (.A(_0158_),
    .B(_0577_),
    .Y(_0578_));
 sg13g2_xnor2_1 _1840_ (.Y(_0579_),
    .A(\game_inst.apple_inst.i_snake_x[1] ),
    .B(_0577_));
 sg13g2_xnor2_1 _1841_ (.Y(_0580_),
    .A(net118),
    .B(_0579_));
 sg13g2_a21oi_1 _1842_ (.A1(net122),
    .A2(_0580_),
    .Y(_0581_),
    .B1(net99));
 sg13g2_nor2_1 _1843_ (.A(_0576_),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_o21ai_1 _1844_ (.B1(net100),
    .Y(_0583_),
    .A1(net122),
    .A2(_0394_));
 sg13g2_a22oi_1 _1845_ (.Y(_0101_),
    .B1(_0582_),
    .B2(_0530_),
    .A2(_0573_),
    .A1(_0158_));
 sg13g2_nand3_1 _1846_ (.B(net123),
    .C(\game_inst.apple_inst.i_snake_x[2] ),
    .A(\game_inst.pos_dir[0] ),
    .Y(_0584_));
 sg13g2_xor2_1 _1847_ (.B(_0577_),
    .A(\game_inst.apple_inst.i_snake_x[2] ),
    .X(_0585_));
 sg13g2_a21o_1 _1848_ (.A2(_0579_),
    .A1(\game_inst.apple_inst.i_snake_x[0] ),
    .B1(_0578_),
    .X(_0586_));
 sg13g2_nand2b_1 _1849_ (.Y(_0587_),
    .B(_0586_),
    .A_N(_0585_));
 sg13g2_xor2_1 _1850_ (.B(_0586_),
    .A(_0585_),
    .X(_0588_));
 sg13g2_a22oi_1 _1851_ (.Y(_0589_),
    .B1(_0588_),
    .B2(net100),
    .A2(_0532_),
    .A1(net99));
 sg13g2_nand2_1 _1852_ (.Y(_0590_),
    .A(net116),
    .B(_0573_));
 sg13g2_nor2b_1 _1853_ (.A(_0589_),
    .B_N(_0538_),
    .Y(_0591_));
 sg13g2_o21ai_1 _1854_ (.B1(_0590_),
    .Y(_0102_),
    .A1(_0573_),
    .A2(_0591_));
 sg13g2_nand2_1 _1855_ (.Y(_0592_),
    .A(net99),
    .B(_0543_));
 sg13g2_nand2_1 _1856_ (.Y(_0593_),
    .A(_0584_),
    .B(_0587_));
 sg13g2_xnor2_1 _1857_ (.Y(_0594_),
    .A(_0159_),
    .B(_0577_));
 sg13g2_xnor2_1 _1858_ (.Y(_0595_),
    .A(_0593_),
    .B(_0594_));
 sg13g2_o21ai_1 _1859_ (.B1(_0592_),
    .Y(_0596_),
    .A1(_0583_),
    .A2(_0595_));
 sg13g2_a22oi_1 _1860_ (.Y(_0103_),
    .B1(_0596_),
    .B2(_0542_),
    .A2(_0573_),
    .A1(_0159_));
 sg13g2_a21oi_1 _1861_ (.A1(_0584_),
    .A2(_0587_),
    .Y(_0597_),
    .B1(\game_inst.apple_inst.i_snake_x[3] ));
 sg13g2_mux2_1 _1862_ (.A0(_0159_),
    .A1(_0295_),
    .S(_0577_),
    .X(_0598_));
 sg13g2_nor2b_1 _1863_ (.A(_0597_),
    .B_N(_0598_),
    .Y(_0599_));
 sg13g2_xnor2_1 _1864_ (.Y(_0600_),
    .A(net1273),
    .B(_0599_));
 sg13g2_a22oi_1 _1865_ (.Y(_0601_),
    .B1(_0600_),
    .B2(net100),
    .A2(_0544_),
    .A1(net99));
 sg13g2_a221oi_1 _1866_ (.B2(_0549_),
    .C1(_0601_),
    .B1(_0547_),
    .A1(_0157_),
    .Y(_0602_),
    .A2(_0401_));
 sg13g2_a21oi_1 _1867_ (.A1(_0161_),
    .A2(_0573_),
    .Y(_0104_),
    .B1(_0602_));
 sg13g2_nand2_1 _1868_ (.Y(_0603_),
    .A(net1248),
    .B(_0232_));
 sg13g2_a21oi_1 _1869_ (.A1(_0401_),
    .A2(_0603_),
    .Y(_0105_),
    .B1(net130));
 sg13g2_nand2_2 _1870_ (.Y(_0604_),
    .A(net122),
    .B(_0401_));
 sg13g2_o21ai_1 _1871_ (.B1(net103),
    .Y(_0605_),
    .A1(net120),
    .A2(net100));
 sg13g2_a21o_1 _1872_ (.A2(net100),
    .A1(net1340),
    .B1(_0605_),
    .X(_0606_));
 sg13g2_and2_1 _1873_ (.A(_0552_),
    .B(_0606_),
    .X(_0607_));
 sg13g2_xor2_1 _1874_ (.B(_0607_),
    .A(_0604_),
    .X(_0106_));
 sg13g2_nor2_2 _1875_ (.A(_0038_),
    .B(net123),
    .Y(_0608_));
 sg13g2_nand2_1 _1876_ (.Y(_0609_),
    .A(\game_inst.apple_inst.i_snake_y[1] ),
    .B(_0608_));
 sg13g2_xnor2_1 _1877_ (.Y(_0610_),
    .A(_0164_),
    .B(_0608_));
 sg13g2_nand2_1 _1878_ (.Y(_0611_),
    .A(\game_inst.apple_inst.i_snake_y[0] ),
    .B(_0610_));
 sg13g2_xnor2_1 _1879_ (.Y(_0612_),
    .A(_0163_),
    .B(_0610_));
 sg13g2_o21ai_1 _1880_ (.B1(_0401_),
    .Y(_0613_),
    .A1(net123),
    .A2(_0612_));
 sg13g2_o21ai_1 _1881_ (.B1(_0613_),
    .Y(_0614_),
    .A1(net100),
    .A2(_0559_));
 sg13g2_inv_1 _1882_ (.Y(_0615_),
    .A(_0614_));
 sg13g2_nand2_1 _1883_ (.Y(_0616_),
    .A(net101),
    .B(_0604_));
 sg13g2_nor2_1 _1884_ (.A(net1236),
    .B(_0604_),
    .Y(_0617_));
 sg13g2_a21oi_1 _1885_ (.A1(_0558_),
    .A2(_0615_),
    .Y(_0107_),
    .B1(_0617_));
 sg13g2_xnor2_1 _1886_ (.Y(_0618_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(_0608_));
 sg13g2_a21oi_1 _1887_ (.A1(_0609_),
    .A2(_0611_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nand3_1 _1888_ (.B(_0611_),
    .C(_0618_),
    .A(_0609_),
    .Y(_0620_));
 sg13g2_nand2b_1 _1889_ (.Y(_0621_),
    .B(_0620_),
    .A_N(_0619_));
 sg13g2_a22oi_1 _1890_ (.Y(_0622_),
    .B1(_0621_),
    .B2(net101),
    .A2(_0560_),
    .A1(net99));
 sg13g2_nand2b_1 _1891_ (.Y(_0623_),
    .B(_0564_),
    .A_N(_0622_));
 sg13g2_mux2_1 _1892_ (.A0(net1278),
    .A1(_0623_),
    .S(_0604_),
    .X(_0108_));
 sg13g2_a21oi_1 _1893_ (.A1(\game_inst.apple_inst.i_snake_y[2] ),
    .A2(_0608_),
    .Y(_0624_),
    .B1(_0619_));
 sg13g2_xor2_1 _1894_ (.B(_0608_),
    .A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(_0625_));
 sg13g2_xnor2_1 _1895_ (.Y(_0626_),
    .A(_0624_),
    .B(_0625_));
 sg13g2_nor3_1 _1896_ (.A(_0570_),
    .B(_0616_),
    .C(_0626_),
    .Y(_0627_));
 sg13g2_nor2_1 _1897_ (.A(net1275),
    .B(_0604_),
    .Y(_0628_));
 sg13g2_nor2_1 _1898_ (.A(_0401_),
    .B(_0571_),
    .Y(_0629_));
 sg13g2_nor3_1 _1899_ (.A(_0627_),
    .B(_0628_),
    .C(_0629_),
    .Y(_0109_));
 sg13g2_and4_1 _1900_ (.A(net1199),
    .B(\game_inst.snake_inst.length[0] ),
    .C(_0238_),
    .D(_0478_),
    .X(_0630_));
 sg13g2_xnor2_1 _1901_ (.Y(_0631_),
    .A(_0150_),
    .B(_0480_));
 sg13g2_nand2_1 _1902_ (.Y(_0110_),
    .A(net114),
    .B(_0631_));
 sg13g2_nor2_1 _1903_ (.A(net1233),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_nor3_1 _1904_ (.A(_0150_),
    .B(_0151_),
    .C(_0480_),
    .Y(_0633_));
 sg13g2_nor3_1 _1905_ (.A(net130),
    .B(net1234),
    .C(_0633_),
    .Y(_0111_));
 sg13g2_and2_1 _1906_ (.A(net1270),
    .B(_0633_),
    .X(_0634_));
 sg13g2_o21ai_1 _1907_ (.B1(net113),
    .Y(_0635_),
    .A1(net1270),
    .A2(_0633_));
 sg13g2_nor2_1 _1908_ (.A(_0634_),
    .B(net1271),
    .Y(_0112_));
 sg13g2_nor2_1 _1909_ (.A(net1262),
    .B(_0634_),
    .Y(_0636_));
 sg13g2_and4_1 _1910_ (.A(net1233),
    .B(\game_inst.snake_inst.length[2] ),
    .C(net1262),
    .D(_0630_),
    .X(_0637_));
 sg13g2_nand3_1 _1911_ (.B(\game_inst.snake_inst.length[3] ),
    .C(_0633_),
    .A(\game_inst.snake_inst.length[2] ),
    .Y(_0638_));
 sg13g2_nor3_1 _1912_ (.A(net130),
    .B(net1263),
    .C(_0637_),
    .Y(_0113_));
 sg13g2_nor2_1 _1913_ (.A(net1221),
    .B(_0637_),
    .Y(_0639_));
 sg13g2_nor2_1 _1914_ (.A(_0152_),
    .B(_0638_),
    .Y(_0640_));
 sg13g2_nor3_1 _1915_ (.A(net131),
    .B(net1222),
    .C(_0640_),
    .Y(_0114_));
 sg13g2_nor2_1 _1916_ (.A(net1243),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_a21oi_1 _1917_ (.A1(net1243),
    .A2(_0640_),
    .Y(_0642_),
    .B1(net131));
 sg13g2_nor2b_1 _1918_ (.A(net1244),
    .B_N(_0642_),
    .Y(_0115_));
 sg13g2_a21oi_1 _1919_ (.A1(\game_inst.snake_inst.length[5] ),
    .A2(_0640_),
    .Y(_0643_),
    .B1(net1164));
 sg13g2_and4_1 _1920_ (.A(\game_inst.snake_inst.length[4] ),
    .B(\game_inst.snake_inst.length[5] ),
    .C(net1164),
    .D(_0637_),
    .X(_0644_));
 sg13g2_nor3_1 _1921_ (.A(net131),
    .B(net1165),
    .C(_0644_),
    .Y(_0116_));
 sg13g2_o21ai_1 _1922_ (.B1(net113),
    .Y(_0645_),
    .A1(net1138),
    .A2(_0644_));
 sg13g2_a21oi_1 _1923_ (.A1(net1138),
    .A2(_0644_),
    .Y(_0117_),
    .B1(_0645_));
 sg13g2_nand2_1 _1924_ (.Y(_0646_),
    .A(net113),
    .B(_0401_));
 sg13g2_nor3_1 _1925_ (.A(_0236_),
    .B(_0403_),
    .C(_0646_),
    .Y(_0118_));
 sg13g2_nor2_1 _1926_ (.A(net1218),
    .B(_0403_),
    .Y(_0647_));
 sg13g2_nor3_1 _1927_ (.A(_0404_),
    .B(_0646_),
    .C(net1219),
    .Y(_0119_));
 sg13g2_a21oi_1 _1928_ (.A1(\game_inst.snake_inst.pos[3] ),
    .A2(_0404_),
    .Y(_0648_),
    .B1(net1190));
 sg13g2_nor3_1 _1929_ (.A(_0406_),
    .B(_0646_),
    .C(net1191),
    .Y(_0120_));
 sg13g2_o21ai_1 _1930_ (.B1(_0395_),
    .Y(_0121_),
    .A1(_0153_),
    .A2(net1146));
 sg13g2_nor2_1 _1931_ (.A(net1140),
    .B(net96),
    .Y(_0649_));
 sg13g2_a21oi_1 _1932_ (.A1(_0162_),
    .A2(net97),
    .Y(_0122_),
    .B1(_0649_));
 sg13g2_nor2_1 _1933_ (.A(net1169),
    .B(net98),
    .Y(_0650_));
 sg13g2_a21oi_1 _1934_ (.A1(_0165_),
    .A2(net97),
    .Y(_0123_),
    .B1(_0650_));
 sg13g2_mux2_1 _1935_ (.A0(net1194),
    .A1(net1217),
    .S(net96),
    .X(_0124_));
 sg13g2_nand2_1 _1936_ (.Y(_0651_),
    .A(net1181),
    .B(net96));
 sg13g2_o21ai_1 _1937_ (.B1(_0651_),
    .Y(_0125_),
    .A1(_0141_),
    .A2(net97));
 sg13g2_nor3_1 _1938_ (.A(_0139_),
    .B(\game_inst.control_inst.dir[0] ),
    .C(net1224),
    .Y(_0652_));
 sg13g2_nor2_1 _1939_ (.A(net131),
    .B(net1225),
    .Y(_0126_));
 sg13g2_nor3_2 _1940_ (.A(\game_inst.tickgen_inst.prev_user_input ),
    .B(_0172_),
    .C(net114),
    .Y(_0653_));
 sg13g2_xnor2_1 _1941_ (.Y(_0654_),
    .A(net1268),
    .B(_0653_));
 sg13g2_nand2_1 _1942_ (.Y(_0127_),
    .A(net136),
    .B(net1269));
 sg13g2_xnor2_1 _1943_ (.Y(_0655_),
    .A(\game_inst.tickgen_inst.counter_max[2] ),
    .B(net1));
 sg13g2_nand2_1 _1944_ (.Y(_0656_),
    .A(net1268),
    .B(_0655_));
 sg13g2_o21ai_1 _1945_ (.B1(_0653_),
    .Y(_0657_),
    .A1(net1268),
    .A2(_0655_));
 sg13g2_nor2b_1 _1946_ (.A(_0657_),
    .B_N(_0656_),
    .Y(_0658_));
 sg13g2_o21ai_1 _1947_ (.B1(net136),
    .Y(_0659_),
    .A1(_0135_),
    .A2(_0653_));
 sg13g2_or2_1 _1948_ (.X(_0128_),
    .B(net1343),
    .A(_0658_));
 sg13g2_o21ai_1 _1949_ (.B1(_0656_),
    .Y(_0660_),
    .A1(_0135_),
    .A2(net1));
 sg13g2_xor2_1 _1950_ (.B(net1),
    .A(net1258),
    .X(_0661_));
 sg13g2_xnor2_1 _1951_ (.Y(_0662_),
    .A(_0660_),
    .B(_0661_));
 sg13g2_nand2_1 _1952_ (.Y(_0663_),
    .A(_0653_),
    .B(_0662_));
 sg13g2_nand2b_1 _1953_ (.Y(_0664_),
    .B(net1258),
    .A_N(_0653_));
 sg13g2_nand3_1 _1954_ (.B(_0663_),
    .C(net1259),
    .A(net136),
    .Y(_0129_));
 sg13g2_nor2b_1 _1955_ (.A(\game_inst.tickgen_inst.counter[3] ),
    .B_N(\game_inst.tickgen_inst.counter_max[3] ),
    .Y(_0665_));
 sg13g2_nor2b_1 _1956_ (.A(\game_inst.tickgen_inst.counter_max[3] ),
    .B_N(\game_inst.tickgen_inst.counter[3] ),
    .Y(_0666_));
 sg13g2_xor2_1 _1957_ (.B(\game_inst.tickgen_inst.counter_max[2] ),
    .A(\game_inst.tickgen_inst.counter[2] ),
    .X(_0667_));
 sg13g2_nor4_1 _1958_ (.A(net1154),
    .B(_0665_),
    .C(_0666_),
    .D(_0667_),
    .Y(_0668_));
 sg13g2_xnor2_1 _1959_ (.Y(_0669_),
    .A(\game_inst.tickgen_inst.counter[1] ),
    .B(\game_inst.tickgen_inst.counter_max[1] ));
 sg13g2_and2_1 _1960_ (.A(_0668_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_o21ai_1 _1961_ (.B1(net1185),
    .Y(_0671_),
    .A1(_0153_),
    .A2(_0154_));
 sg13g2_nand2b_1 _1962_ (.Y(_0672_),
    .B(net1125),
    .A_N(\game_inst.o_vga_vsync ));
 sg13g2_nand2b_1 _1963_ (.Y(_0673_),
    .B(\game_inst.control_inst.o_start ),
    .A_N(failure));
 sg13g2_or4_1 _1964_ (.A(net5),
    .B(\game_inst.o_success ),
    .C(_0672_),
    .D(_0673_),
    .X(_0674_));
 sg13g2_inv_1 _1965_ (.Y(_0675_),
    .A(_0674_));
 sg13g2_o21ai_1 _1966_ (.B1(net114),
    .Y(_0676_),
    .A1(net1185),
    .A2(_0670_));
 sg13g2_a21oi_1 _1967_ (.A1(net1186),
    .A2(_0674_),
    .Y(_0130_),
    .B1(_0676_));
 sg13g2_nor2_2 _1968_ (.A(_0670_),
    .B(_0674_),
    .Y(_0677_));
 sg13g2_o21ai_1 _1969_ (.B1(net114),
    .Y(_0678_),
    .A1(net1154),
    .A2(_0677_));
 sg13g2_a21oi_1 _1970_ (.A1(net1154),
    .A2(_0675_),
    .Y(_0131_),
    .B1(_0678_));
 sg13g2_and2_1 _1971_ (.A(\game_inst.tickgen_inst.counter[1] ),
    .B(net1154),
    .X(_0679_));
 sg13g2_nand2_1 _1972_ (.Y(_0680_),
    .A(net1256),
    .B(net1154));
 sg13g2_a22oi_1 _1973_ (.Y(_0681_),
    .B1(_0677_),
    .B2(_0680_),
    .A2(_0674_),
    .A1(net1256));
 sg13g2_o21ai_1 _1974_ (.B1(net114),
    .Y(_0682_),
    .A1(net1256),
    .A2(net1154));
 sg13g2_nor2_1 _1975_ (.A(_0681_),
    .B(_0682_),
    .Y(_0132_));
 sg13g2_a21oi_1 _1976_ (.A1(_0677_),
    .A2(_0679_),
    .Y(_0683_),
    .B1(net1179));
 sg13g2_nand2_1 _1977_ (.Y(_0684_),
    .A(net1179),
    .B(_0679_));
 sg13g2_a21oi_1 _1978_ (.A1(_0677_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(_0674_));
 sg13g2_nor3_1 _1979_ (.A(net131),
    .B(net1180),
    .C(_0685_),
    .Y(_0133_));
 sg13g2_nor3_1 _1980_ (.A(_0670_),
    .B(_0674_),
    .C(_0684_),
    .Y(_0686_));
 sg13g2_o21ai_1 _1981_ (.B1(net114),
    .Y(_0687_),
    .A1(net1150),
    .A2(_0686_));
 sg13g2_a21oi_1 _1982_ (.A1(net1150),
    .A2(_0685_),
    .Y(_0134_),
    .B1(_0687_));
 sg13g2_buf_1 _1983_ (.A(\game_inst.vga_inst.color[3] ),
    .X(uo_out[6]));
 sg13g2_dfrbpq_2 _1984_ (.RESET_B(net25),
    .D(_0039_),
    .Q(\game_inst.vga_inst.px[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1985_ (.RESET_B(net93),
    .D(_0040_),
    .Q(\game_inst.vga_inst.px[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1986_ (.RESET_B(net92),
    .D(_0041_),
    .Q(\game_inst.vga_inst.px[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1987_ (.RESET_B(net91),
    .D(_0042_),
    .Q(\game_inst.vga_inst.px[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _1988_ (.RESET_B(net90),
    .D(net1286),
    .Q(\game_inst.vga_inst.px[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _1989_ (.RESET_B(net89),
    .D(_0044_),
    .Q(\game_inst.vga_inst.px[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _1990_ (.RESET_B(net88),
    .D(net1240),
    .Q(\game_inst.vga_inst.px[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1991_ (.RESET_B(net87),
    .D(net1334),
    .Q(\game_inst.vga_inst.px[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _1992_ (.RESET_B(net86),
    .D(_0047_),
    .Q(\game_inst.vga_inst.px[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1993_ (.RESET_B(net26),
    .D(_0048_),
    .Q(\game_inst.vga_inst.px[9] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1994_ (.RESET_B(net27),
    .D(_0000_),
    .Q(\game_inst.vga_inst.color[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1995_ (.RESET_B(net33),
    .D(_0001_),
    .Q(\game_inst.vga_inst.color[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1996_ (.RESET_B(net84),
    .D(net1135),
    .Q(\game_inst.vga_inst.color[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1997_ (.RESET_B(net83),
    .D(net1163),
    .Q(\game_inst.snake_inst.pos[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1998_ (.RESET_B(net82),
    .D(_0050_),
    .Q(\game_inst.snake_inst.pos[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1999_ (.RESET_B(net81),
    .D(_0051_),
    .Q(\game_inst.snake_inst.pos[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2000_ (.RESET_B(net80),
    .D(net1254),
    .Q(\game_inst.snake_inst.pos[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2001_ (.RESET_B(net34),
    .D(_0053_),
    .Q(\game_inst.snake_inst.pos[7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2002_ (.RESET_B(net35),
    .D(net718),
    .Q(\game_inst.o_vga_hsync ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2003_ (.RESET_B(net36),
    .D(net1125),
    .Q(\game_inst.o_vga_vsync ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2004_ (.RESET_B(net37),
    .D(_0038_),
    .Q(\game_inst.vga_inst.prev_dir[0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2005_ (.RESET_B(net38),
    .D(net1143),
    .Q(\game_inst.vga_inst.row_buffer[8][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2006_ (.RESET_B(net39),
    .D(net1149),
    .Q(\game_inst.vga_inst.row_buffer[8][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2007_ (.RESET_B(net42),
    .D(net1137),
    .Q(\game_inst.vga_inst.row_buffer[8][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2008_ (.RESET_B(net79),
    .D(net1145),
    .Q(\game_inst.vga_inst.row_buffer[8][3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2009_ (.RESET_B(net78),
    .D(net1156),
    .Q(\game_inst.pos_dir[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _2010_ (.RESET_B(net43),
    .D(net1178),
    .Q(\game_inst.pos_dir[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2011_ (.RESET_B(net44),
    .D(net1318),
    .Q(\game_inst.vga_inst.row_buffer[1][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2012_ (.RESET_B(net45),
    .D(net1326),
    .Q(\game_inst.vga_inst.row_buffer[1][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2013_ (.RESET_B(net46),
    .D(net1324),
    .Q(\game_inst.vga_inst.row_buffer[1][2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2014_ (.RESET_B(net47),
    .D(net1321),
    .Q(\game_inst.vga_inst.row_buffer[1][3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2015_ (.RESET_B(net48),
    .D(net1305),
    .Q(\game_inst.vga_inst.row_buffer[2][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2016_ (.RESET_B(net49),
    .D(net1328),
    .Q(\game_inst.vga_inst.row_buffer[2][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2017_ (.RESET_B(net50),
    .D(net1314),
    .Q(\game_inst.vga_inst.row_buffer[2][2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2018_ (.RESET_B(net51),
    .D(net1300),
    .Q(\game_inst.vga_inst.row_buffer[2][3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2019_ (.RESET_B(net52),
    .D(_0012_),
    .Q(\game_inst.vga_inst.row_buffer[3][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2020_ (.RESET_B(net53),
    .D(net1310),
    .Q(\game_inst.vga_inst.row_buffer[3][1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2021_ (.RESET_B(net54),
    .D(net1296),
    .Q(\game_inst.vga_inst.row_buffer[3][2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2022_ (.RESET_B(net55),
    .D(net1298),
    .Q(\game_inst.vga_inst.row_buffer[3][3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2023_ (.RESET_B(net56),
    .D(net1308),
    .Q(\game_inst.vga_inst.row_buffer[4][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2024_ (.RESET_B(net57),
    .D(_0017_),
    .Q(\game_inst.vga_inst.row_buffer[4][1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2025_ (.RESET_B(net58),
    .D(_0018_),
    .Q(\game_inst.vga_inst.row_buffer[4][2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2026_ (.RESET_B(net59),
    .D(_0019_),
    .Q(\game_inst.vga_inst.row_buffer[4][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2027_ (.RESET_B(net60),
    .D(net1294),
    .Q(\game_inst.vga_inst.row_buffer[5][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2028_ (.RESET_B(net61),
    .D(_0021_),
    .Q(\game_inst.vga_inst.row_buffer[5][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2029_ (.RESET_B(net62),
    .D(net1292),
    .Q(\game_inst.vga_inst.row_buffer[5][2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2030_ (.RESET_B(net63),
    .D(net1290),
    .Q(\game_inst.vga_inst.row_buffer[5][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2031_ (.RESET_B(net64),
    .D(_0024_),
    .Q(\game_inst.vga_inst.row_buffer[6][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2032_ (.RESET_B(net65),
    .D(_0025_),
    .Q(\game_inst.vga_inst.row_buffer[6][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2033_ (.RESET_B(net66),
    .D(_0026_),
    .Q(\game_inst.vga_inst.row_buffer[6][2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2034_ (.RESET_B(net67),
    .D(_0027_),
    .Q(\game_inst.vga_inst.row_buffer[6][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2035_ (.RESET_B(net68),
    .D(_0028_),
    .Q(\game_inst.vga_inst.row_buffer[7][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2036_ (.RESET_B(net69),
    .D(_0029_),
    .Q(\game_inst.vga_inst.row_buffer[7][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2037_ (.RESET_B(net74),
    .D(_0030_),
    .Q(\game_inst.vga_inst.row_buffer[7][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2038_ (.RESET_B(net77),
    .D(_0031_),
    .Q(\game_inst.vga_inst.row_buffer[7][3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2039_ (.RESET_B(net76),
    .D(net1208),
    .Q(\game_inst.vga_inst.row_buffer[0][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2040_ (.RESET_B(net75),
    .D(net1232),
    .Q(\game_inst.vga_inst.row_buffer[0][1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2041_ (.RESET_B(net73),
    .D(net1227),
    .Q(\game_inst.vga_inst.row_buffer[0][2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2042_ (.RESET_B(net85),
    .D(net1229),
    .Q(\game_inst.vga_inst.row_buffer[0][3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2043_ (.RESET_B(net72),
    .D(net1330),
    .Q(\game_inst.vga_inst.s_hsync ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _2044_ (.RESET_B(net71),
    .D(net1161),
    .Q(\game_inst.vga_inst.py[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2045_ (.RESET_B(net41),
    .D(net1176),
    .Q(\game_inst.vga_inst.py[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2046_ (.RESET_B(net32),
    .D(_0062_),
    .Q(\game_inst.vga_inst.py[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2047_ (.RESET_B(net30),
    .D(_0063_),
    .Q(\game_inst.vga_inst.py[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2048_ (.RESET_B(net28),
    .D(net1212),
    .Q(\game_inst.vga_inst.py[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2049_ (.RESET_B(net23),
    .D(_0065_),
    .Q(\game_inst.vga_inst.py[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2050_ (.RESET_B(net21),
    .D(_0066_),
    .Q(\game_inst.vga_inst.py[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2051_ (.RESET_B(net19),
    .D(net1242),
    .Q(\game_inst.vga_inst.py[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2052_ (.RESET_B(net17),
    .D(net1216),
    .Q(\game_inst.vga_inst.py[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _2053_ (.RESET_B(net180),
    .D(net1201),
    .Q(\game_inst.vga_inst.py[9] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2054_ (.RESET_B(net15),
    .D(net1158),
    .Q(\game_inst.vga_inst.s_vsync ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2055_ (.RESET_B(net659),
    .D(_0070_),
    .Q(failure),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2056_ (.RESET_B(net658),
    .D(net1173),
    .Q(\game_inst.apple_inst.apple_x[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2057_ (.RESET_B(net657),
    .D(net1184),
    .Q(\game_inst.apple_inst.apple_x[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _2058_ (.RESET_B(net655),
    .D(_0073_),
    .Q(\game_inst.apple_inst.apple_x[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2059_ (.RESET_B(net654),
    .D(_0074_),
    .Q(\game_inst.apple_inst.apple_x[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2060_ (.RESET_B(net653),
    .D(net1206),
    .Q(\game_inst.apple_inst.apple_x[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2061_ (.RESET_B(net652),
    .D(_0076_),
    .Q(\game_inst.apple_inst.o_ready ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2062_ (.RESET_B(net650),
    .D(_0077_),
    .Q(\game_inst.apple_inst.test ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2063_ (.RESET_B(net648),
    .D(_0078_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2064_ (.RESET_B(net646),
    .D(_0079_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2065_ (.RESET_B(net178),
    .D(_0080_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2066_ (.RESET_B(net176),
    .D(_0081_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _2067_ (.RESET_B(net174),
    .D(net1168),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _2068_ (.RESET_B(net172),
    .D(net1141),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2069_ (.RESET_B(net170),
    .D(_0084_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2070_ (.RESET_B(net168),
    .D(_0085_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2071_ (.RESET_B(net166),
    .D(_0086_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _2072_ (.RESET_B(net164),
    .D(net1204),
    .Q(\game_inst.control_inst.i_head_dir[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _2073_ (.RESET_B(net162),
    .D(_0088_),
    .Q(\game_inst.control_inst.backwards[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _2074_ (.RESET_B(net160),
    .D(_0089_),
    .Q(\game_inst.head_x[0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2075_ (.RESET_B(net158),
    .D(_0090_),
    .Q(\game_inst.head_x[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2076_ (.RESET_B(net156),
    .D(_0091_),
    .Q(\game_inst.head_x[2] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _2077_ (.RESET_B(net154),
    .D(net1281),
    .Q(\game_inst.head_x[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2078_ (.RESET_B(net152),
    .D(_0093_),
    .Q(\game_inst.head_x[4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _2079_ (.RESET_B(net150),
    .D(_0094_),
    .Q(\game_inst.head_y[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _2080_ (.RESET_B(net148),
    .D(_0095_),
    .Q(\game_inst.head_y[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2081_ (.RESET_B(net146),
    .D(_0096_),
    .Q(\game_inst.head_y[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2082_ (.RESET_B(net144),
    .D(_0097_),
    .Q(\game_inst.head_y[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2083_ (.RESET_B(net142),
    .D(_0098_),
    .Q(\game_inst.control_inst.dir[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2084_ (.RESET_B(net141),
    .D(_0099_),
    .Q(\game_inst.control_inst.dir[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _2085_ (.RESET_B(net140),
    .D(_0100_),
    .Q(\game_inst.apple_inst.i_snake_x[0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2086_ (.RESET_B(net139),
    .D(net1251),
    .Q(\game_inst.apple_inst.i_snake_x[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2087_ (.RESET_B(net138),
    .D(_0102_),
    .Q(\game_inst.apple_inst.i_snake_x[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2088_ (.RESET_B(net137),
    .D(net1316),
    .Q(\game_inst.apple_inst.i_snake_x[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2089_ (.RESET_B(net70),
    .D(_0104_),
    .Q(\game_inst.apple_inst.i_snake_x[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2090_ (.RESET_B(net40),
    .D(_0105_),
    .Q(\game_inst.apple_inst.i_snake_valid ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2091_ (.RESET_B(net29),
    .D(_0106_),
    .Q(\game_inst.apple_inst.i_snake_y[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2092_ (.RESET_B(net24),
    .D(net1237),
    .Q(\game_inst.apple_inst.i_snake_y[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2093_ (.RESET_B(net22),
    .D(net1279),
    .Q(\game_inst.apple_inst.i_snake_y[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2094_ (.RESET_B(net20),
    .D(net1276),
    .Q(\game_inst.apple_inst.i_snake_y[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _2095_ (.RESET_B(net18),
    .D(_0110_),
    .Q(\game_inst.snake_inst.length[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2096_ (.RESET_B(net16),
    .D(net1235),
    .Q(\game_inst.snake_inst.length[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2097_ (.RESET_B(net660),
    .D(net1272),
    .Q(\game_inst.snake_inst.length[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2098_ (.RESET_B(net651),
    .D(net1264),
    .Q(\game_inst.snake_inst.length[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2099_ (.RESET_B(net649),
    .D(net1223),
    .Q(\game_inst.snake_inst.length[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2100_ (.RESET_B(net647),
    .D(_0115_),
    .Q(\game_inst.snake_inst.length[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2101_ (.RESET_B(net179),
    .D(net1166),
    .Q(\game_inst.snake_inst.length[6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2102_ (.RESET_B(net177),
    .D(net1139),
    .Q(\game_inst.snake_inst.length[7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2103_ (.RESET_B(net175),
    .D(_0118_),
    .Q(\game_inst.snake_inst.pos[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2104_ (.RESET_B(net173),
    .D(net1220),
    .Q(\game_inst.snake_inst.pos[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2105_ (.RESET_B(net181),
    .D(net1192),
    .Q(\game_inst.snake_inst.pos[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2106_ (.RESET_B(net182),
    .D(net958),
    .Q(\game_inst.snake_inst.dir_out[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2107_ (.RESET_B(net183),
    .D(net715),
    .Q(\game_inst.snake_inst.dir_out[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2108_ (.RESET_B(net184),
    .D(net881),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[232][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2109_ (.RESET_B(net185),
    .D(net879),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[232][1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2110_ (.RESET_B(net186),
    .D(net1112),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[231][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2111_ (.RESET_B(net187),
    .D(net973),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[231][1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2112_ (.RESET_B(net188),
    .D(net818),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[230][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2113_ (.RESET_B(net189),
    .D(net703),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[230][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2114_ (.RESET_B(net190),
    .D(net908),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[229][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2115_ (.RESET_B(net191),
    .D(net1011),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[229][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2116_ (.RESET_B(net192),
    .D(net762),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[228][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2117_ (.RESET_B(net193),
    .D(net1072),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[228][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2118_ (.RESET_B(net194),
    .D(net777),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[227][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2119_ (.RESET_B(net195),
    .D(net1108),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[227][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2120_ (.RESET_B(net196),
    .D(net945),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[226][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2121_ (.RESET_B(net197),
    .D(net890),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[226][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2122_ (.RESET_B(net198),
    .D(net871),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[225][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2123_ (.RESET_B(net199),
    .D(net1062),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[225][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2124_ (.RESET_B(net200),
    .D(net759),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[224][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2125_ (.RESET_B(net201),
    .D(net1036),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[224][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2126_ (.RESET_B(net202),
    .D(net1078),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[223][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2127_ (.RESET_B(net203),
    .D(net1035),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[223][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2128_ (.RESET_B(net204),
    .D(net894),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[222][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2129_ (.RESET_B(net205),
    .D(net983),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[222][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2130_ (.RESET_B(net206),
    .D(net803),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[221][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2131_ (.RESET_B(net207),
    .D(net1071),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[221][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2132_ (.RESET_B(net208),
    .D(net860),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[220][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2133_ (.RESET_B(net209),
    .D(net749),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[220][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2134_ (.RESET_B(net210),
    .D(net977),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[219][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2135_ (.RESET_B(net211),
    .D(net705),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[219][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2136_ (.RESET_B(net212),
    .D(net723),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[218][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2137_ (.RESET_B(net213),
    .D(net972),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[218][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2138_ (.RESET_B(net214),
    .D(net1033),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[217][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2139_ (.RESET_B(net215),
    .D(net895),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[217][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2140_ (.RESET_B(net216),
    .D(net934),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[216][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2141_ (.RESET_B(net217),
    .D(net1016),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[216][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2142_ (.RESET_B(net218),
    .D(net940),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[215][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2143_ (.RESET_B(net219),
    .D(net982),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[215][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2144_ (.RESET_B(net220),
    .D(net784),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[214][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2145_ (.RESET_B(net221),
    .D(net1101),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[214][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2146_ (.RESET_B(net222),
    .D(net1114),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[213][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2147_ (.RESET_B(net223),
    .D(net781),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[213][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2148_ (.RESET_B(net224),
    .D(net764),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[212][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2149_ (.RESET_B(net225),
    .D(net965),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[212][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2150_ (.RESET_B(net226),
    .D(net800),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[211][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2151_ (.RESET_B(net227),
    .D(net920),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[211][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2152_ (.RESET_B(net228),
    .D(net848),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[210][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2153_ (.RESET_B(net229),
    .D(net914),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[210][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2154_ (.RESET_B(net230),
    .D(net756),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[209][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2155_ (.RESET_B(net231),
    .D(net1094),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[209][1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2156_ (.RESET_B(net232),
    .D(net702),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[208][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2157_ (.RESET_B(net233),
    .D(net722),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[208][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2158_ (.RESET_B(net234),
    .D(net753),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[207][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2159_ (.RESET_B(net235),
    .D(net875),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[207][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2160_ (.RESET_B(net236),
    .D(net1077),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[206][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2161_ (.RESET_B(net237),
    .D(net953),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[206][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2162_ (.RESET_B(net238),
    .D(net775),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[205][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2163_ (.RESET_B(net239),
    .D(net935),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[205][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2164_ (.RESET_B(net240),
    .D(net1084),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[204][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2165_ (.RESET_B(net241),
    .D(net929),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[204][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2166_ (.RESET_B(net242),
    .D(net995),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[203][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2167_ (.RESET_B(net243),
    .D(net867),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[203][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2168_ (.RESET_B(net244),
    .D(net1106),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[202][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2169_ (.RESET_B(net245),
    .D(net809),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[202][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2170_ (.RESET_B(net246),
    .D(net687),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[201][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2171_ (.RESET_B(net247),
    .D(net1099),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[201][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2172_ (.RESET_B(net248),
    .D(net891),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[200][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2173_ (.RESET_B(net249),
    .D(net1075),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[200][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2174_ (.RESET_B(net250),
    .D(net868),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[199][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2175_ (.RESET_B(net251),
    .D(net1083),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[199][1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2176_ (.RESET_B(net252),
    .D(net837),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[198][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2177_ (.RESET_B(net253),
    .D(net1028),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[198][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2178_ (.RESET_B(net254),
    .D(net1050),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[197][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2179_ (.RESET_B(net255),
    .D(net880),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[197][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2180_ (.RESET_B(net256),
    .D(net951),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[196][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2181_ (.RESET_B(net257),
    .D(net993),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[196][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2182_ (.RESET_B(net258),
    .D(net832),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[195][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2183_ (.RESET_B(net259),
    .D(net1089),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[195][1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2184_ (.RESET_B(net260),
    .D(net672),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[194][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2185_ (.RESET_B(net261),
    .D(net1105),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[194][1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2186_ (.RESET_B(net262),
    .D(net980),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[193][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2187_ (.RESET_B(net263),
    .D(net693),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[193][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2188_ (.RESET_B(net264),
    .D(net727),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[192][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2189_ (.RESET_B(net265),
    .D(net696),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[192][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2190_ (.RESET_B(net266),
    .D(net985),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[191][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2191_ (.RESET_B(net267),
    .D(net824),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[191][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2192_ (.RESET_B(net268),
    .D(net1118),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[190][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2193_ (.RESET_B(net269),
    .D(net947),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[190][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2194_ (.RESET_B(net270),
    .D(net968),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[189][0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2195_ (.RESET_B(net271),
    .D(net834),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[189][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2196_ (.RESET_B(net272),
    .D(net767),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[188][0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2197_ (.RESET_B(net273),
    .D(net769),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[188][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2198_ (.RESET_B(net274),
    .D(net1044),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[187][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2199_ (.RESET_B(net275),
    .D(net898),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[187][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2200_ (.RESET_B(net276),
    .D(net694),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[186][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2201_ (.RESET_B(net277),
    .D(net975),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[186][1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2202_ (.RESET_B(net278),
    .D(net1023),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[185][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2203_ (.RESET_B(net279),
    .D(net1102),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[185][1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2204_ (.RESET_B(net280),
    .D(net745),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[184][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2205_ (.RESET_B(net281),
    .D(net872),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[184][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2206_ (.RESET_B(net282),
    .D(net799),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[183][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2207_ (.RESET_B(net283),
    .D(net1041),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[183][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2208_ (.RESET_B(net284),
    .D(net950),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[182][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2209_ (.RESET_B(net285),
    .D(net941),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[182][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2210_ (.RESET_B(net286),
    .D(net1013),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[181][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2211_ (.RESET_B(net287),
    .D(net1070),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[181][1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2212_ (.RESET_B(net288),
    .D(net1004),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[180][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2213_ (.RESET_B(net289),
    .D(net689),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[180][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2214_ (.RESET_B(net290),
    .D(net778),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[179][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2215_ (.RESET_B(net291),
    .D(net1047),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[179][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2216_ (.RESET_B(net292),
    .D(net674),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[178][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2217_ (.RESET_B(net293),
    .D(net1097),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[178][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2218_ (.RESET_B(net294),
    .D(net1080),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[177][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2219_ (.RESET_B(net295),
    .D(net698),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[177][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2220_ (.RESET_B(net296),
    .D(net1065),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[176][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2221_ (.RESET_B(net297),
    .D(net685),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[176][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2222_ (.RESET_B(net298),
    .D(net692),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[175][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2223_ (.RESET_B(net299),
    .D(net918),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[175][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2224_ (.RESET_B(net300),
    .D(net997),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[174][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2225_ (.RESET_B(net301),
    .D(net683),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[174][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2226_ (.RESET_B(net302),
    .D(net971),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[173][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2227_ (.RESET_B(net303),
    .D(net1079),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[173][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2228_ (.RESET_B(net304),
    .D(net1055),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[172][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2229_ (.RESET_B(net305),
    .D(net896),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[172][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2230_ (.RESET_B(net306),
    .D(net1085),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[171][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2231_ (.RESET_B(net307),
    .D(net864),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[171][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2232_ (.RESET_B(net308),
    .D(net724),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[170][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2233_ (.RESET_B(net309),
    .D(net719),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[170][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2234_ (.RESET_B(net310),
    .D(net961),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[169][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2235_ (.RESET_B(net311),
    .D(net998),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[169][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2236_ (.RESET_B(net312),
    .D(net852),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[168][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2237_ (.RESET_B(net313),
    .D(net668),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[168][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2238_ (.RESET_B(net314),
    .D(net675),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[167][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2239_ (.RESET_B(net315),
    .D(net1038),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[167][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2240_ (.RESET_B(net316),
    .D(net1119),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[166][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2241_ (.RESET_B(net317),
    .D(net747),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[166][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2242_ (.RESET_B(net318),
    .D(net1109),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[165][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2243_ (.RESET_B(net319),
    .D(net932),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[165][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2244_ (.RESET_B(net320),
    .D(net967),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[164][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2245_ (.RESET_B(net321),
    .D(net905),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[164][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2246_ (.RESET_B(net322),
    .D(net688),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[163][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2247_ (.RESET_B(net323),
    .D(net960),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[163][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2248_ (.RESET_B(net324),
    .D(net970),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[162][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2249_ (.RESET_B(net325),
    .D(net828),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[162][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2250_ (.RESET_B(net326),
    .D(net1042),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[161][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2251_ (.RESET_B(net327),
    .D(net1063),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[161][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2252_ (.RESET_B(net328),
    .D(net899),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[160][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2253_ (.RESET_B(net329),
    .D(net1081),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[160][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2254_ (.RESET_B(net330),
    .D(net812),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[159][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2255_ (.RESET_B(net331),
    .D(net835),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[159][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2256_ (.RESET_B(net332),
    .D(net816),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[158][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2257_ (.RESET_B(net333),
    .D(net728),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[158][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2258_ (.RESET_B(net334),
    .D(net863),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[157][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2259_ (.RESET_B(net335),
    .D(net819),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[157][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2260_ (.RESET_B(net336),
    .D(net1056),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[156][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2261_ (.RESET_B(net337),
    .D(net900),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[156][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2262_ (.RESET_B(net338),
    .D(net974),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[155][0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2263_ (.RESET_B(net339),
    .D(net732),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[155][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2264_ (.RESET_B(net340),
    .D(net733),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[154][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _2265_ (.RESET_B(net341),
    .D(net912),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[154][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2266_ (.RESET_B(net342),
    .D(net949),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[153][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2267_ (.RESET_B(net343),
    .D(net1018),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[153][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2268_ (.RESET_B(net344),
    .D(net1017),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[152][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2269_ (.RESET_B(net345),
    .D(net886),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[152][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2270_ (.RESET_B(net346),
    .D(net931),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[151][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2271_ (.RESET_B(net347),
    .D(net859),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[151][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2272_ (.RESET_B(net348),
    .D(net810),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[150][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2273_ (.RESET_B(net349),
    .D(net806),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[150][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2274_ (.RESET_B(net350),
    .D(net1121),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[149][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2275_ (.RESET_B(net351),
    .D(net794),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[149][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2276_ (.RESET_B(net352),
    .D(net673),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[148][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2277_ (.RESET_B(net353),
    .D(net746),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[148][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2278_ (.RESET_B(net354),
    .D(net937),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[147][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2279_ (.RESET_B(net355),
    .D(net855),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[147][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2280_ (.RESET_B(net356),
    .D(net776),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[146][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2281_ (.RESET_B(net357),
    .D(net956),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[146][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2282_ (.RESET_B(net358),
    .D(net979),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[145][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2283_ (.RESET_B(net359),
    .D(net869),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[145][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2284_ (.RESET_B(net360),
    .D(net1110),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[144][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2285_ (.RESET_B(net361),
    .D(net1066),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[144][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2286_ (.RESET_B(net362),
    .D(net944),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[143][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2287_ (.RESET_B(net363),
    .D(net1053),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[143][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2288_ (.RESET_B(net364),
    .D(net1069),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[142][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2289_ (.RESET_B(net365),
    .D(net821),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[142][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2290_ (.RESET_B(net366),
    .D(net1032),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[141][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2291_ (.RESET_B(net367),
    .D(net988),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[141][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2292_ (.RESET_B(net368),
    .D(net792),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[140][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2293_ (.RESET_B(net369),
    .D(net1127),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[140][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2294_ (.RESET_B(net370),
    .D(net671),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[139][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2295_ (.RESET_B(net371),
    .D(net962),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[139][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2296_ (.RESET_B(net372),
    .D(net874),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[138][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2297_ (.RESET_B(net373),
    .D(net954),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[138][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2298_ (.RESET_B(net374),
    .D(net670),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[137][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2299_ (.RESET_B(net375),
    .D(net813),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[137][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2300_ (.RESET_B(net376),
    .D(net1123),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[136][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2301_ (.RESET_B(net377),
    .D(net922),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[136][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2302_ (.RESET_B(net378),
    .D(net830),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[135][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2303_ (.RESET_B(net379),
    .D(net815),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[135][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2304_ (.RESET_B(net380),
    .D(net976),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[134][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2305_ (.RESET_B(net381),
    .D(net865),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[134][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2306_ (.RESET_B(net382),
    .D(net797),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[133][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2307_ (.RESET_B(net383),
    .D(net763),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[133][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2308_ (.RESET_B(net384),
    .D(net866),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[132][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2309_ (.RESET_B(net385),
    .D(net933),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[132][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2310_ (.RESET_B(net386),
    .D(net903),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[131][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2311_ (.RESET_B(net387),
    .D(net755),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[131][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2312_ (.RESET_B(net388),
    .D(net957),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[130][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2313_ (.RESET_B(net389),
    .D(net730),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[130][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2314_ (.RESET_B(net390),
    .D(net907),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[129][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net391),
    .D(net770),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[129][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net392),
    .D(net720),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[128][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net393),
    .D(net758),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[128][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net394),
    .D(net1045),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[127][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2319_ (.RESET_B(net395),
    .D(net786),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[127][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net396),
    .D(net854),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[126][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net397),
    .D(net909),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[126][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net398),
    .D(net911),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[125][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2323_ (.RESET_B(net399),
    .D(net858),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[125][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2324_ (.RESET_B(net400),
    .D(net748),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[124][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2325_ (.RESET_B(net401),
    .D(net916),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[124][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2326_ (.RESET_B(net402),
    .D(net772),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[123][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2327_ (.RESET_B(net403),
    .D(net885),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[123][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net404),
    .D(net1026),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[122][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2329_ (.RESET_B(net405),
    .D(net1010),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[122][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2330_ (.RESET_B(net406),
    .D(net740),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[121][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2331_ (.RESET_B(net407),
    .D(net1098),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[121][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2332_ (.RESET_B(net408),
    .D(net987),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[120][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net409),
    .D(net1090),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[120][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net410),
    .D(net990),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[119][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net411),
    .D(net1092),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[119][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2336_ (.RESET_B(net412),
    .D(net739),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[118][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2337_ (.RESET_B(net413),
    .D(net955),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[118][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2338_ (.RESET_B(net414),
    .D(net709),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[117][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2339_ (.RESET_B(net415),
    .D(net1091),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[117][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2340_ (.RESET_B(net416),
    .D(net1122),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[116][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2341_ (.RESET_B(net417),
    .D(net1008),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[116][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2342_ (.RESET_B(net418),
    .D(net846),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[115][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2343_ (.RESET_B(net419),
    .D(net845),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[115][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net420),
    .D(net851),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[114][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net421),
    .D(net793),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[114][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2346_ (.RESET_B(net422),
    .D(net1030),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[113][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2347_ (.RESET_B(net423),
    .D(net805),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[113][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net424),
    .D(net906),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[112][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net425),
    .D(net919),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[112][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net426),
    .D(net1126),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[111][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2351_ (.RESET_B(net427),
    .D(net742),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[111][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2352_ (.RESET_B(net428),
    .D(net744),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[110][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2353_ (.RESET_B(net429),
    .D(net986),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[110][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2354_ (.RESET_B(net430),
    .D(net731),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[109][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2355_ (.RESET_B(net431),
    .D(net699),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[109][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2356_ (.RESET_B(net432),
    .D(net1037),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[108][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2357_ (.RESET_B(net433),
    .D(net774),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[108][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2358_ (.RESET_B(net434),
    .D(net1052),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[107][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2359_ (.RESET_B(net435),
    .D(net817),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[107][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2360_ (.RESET_B(net436),
    .D(net917),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[106][0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2361_ (.RESET_B(net437),
    .D(net928),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[106][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2362_ (.RESET_B(net438),
    .D(net948),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[105][0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2363_ (.RESET_B(net439),
    .D(net936),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[105][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2364_ (.RESET_B(net440),
    .D(net766),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[104][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2365_ (.RESET_B(net441),
    .D(net991),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[104][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2366_ (.RESET_B(net442),
    .D(net676),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[103][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2367_ (.RESET_B(net443),
    .D(net796),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[103][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2368_ (.RESET_B(net444),
    .D(net887),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[102][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2369_ (.RESET_B(net445),
    .D(net771),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[102][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2370_ (.RESET_B(net446),
    .D(net711),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[101][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2371_ (.RESET_B(net447),
    .D(net704),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[101][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2372_ (.RESET_B(net448),
    .D(net757),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[100][0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2373_ (.RESET_B(net449),
    .D(net984),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[100][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2374_ (.RESET_B(net450),
    .D(net888),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[99][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2375_ (.RESET_B(net451),
    .D(net826),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[99][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2376_ (.RESET_B(net452),
    .D(net1124),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[98][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2377_ (.RESET_B(net453),
    .D(net681),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[98][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2378_ (.RESET_B(net454),
    .D(net925),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[97][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2379_ (.RESET_B(net455),
    .D(net710),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[97][1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _2380_ (.RESET_B(net456),
    .D(net1003),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[96][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2381_ (.RESET_B(net457),
    .D(net1005),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[96][1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _2382_ (.RESET_B(net458),
    .D(net969),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[95][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2383_ (.RESET_B(net459),
    .D(net691),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[95][1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _2384_ (.RESET_B(net460),
    .D(net808),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[94][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2385_ (.RESET_B(net461),
    .D(net1001),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[94][1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _2386_ (.RESET_B(net462),
    .D(net849),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[93][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2387_ (.RESET_B(net463),
    .D(net716),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[93][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2388_ (.RESET_B(net464),
    .D(net829),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[92][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2389_ (.RESET_B(net465),
    .D(net897),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[92][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2390_ (.RESET_B(net466),
    .D(net1061),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[91][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2391_ (.RESET_B(net467),
    .D(net892),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[91][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2392_ (.RESET_B(net468),
    .D(net783),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[90][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2393_ (.RESET_B(net469),
    .D(net1115),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[90][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2394_ (.RESET_B(net470),
    .D(net836),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[89][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2395_ (.RESET_B(net471),
    .D(net938),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[89][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2396_ (.RESET_B(net472),
    .D(net737),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[88][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2397_ (.RESET_B(net473),
    .D(net1012),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[88][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2398_ (.RESET_B(net474),
    .D(net996),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[87][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2399_ (.RESET_B(net475),
    .D(net999),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[87][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2400_ (.RESET_B(net476),
    .D(net1051),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[86][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2401_ (.RESET_B(net477),
    .D(net1074),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[86][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2402_ (.RESET_B(net478),
    .D(net1029),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[85][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2403_ (.RESET_B(net479),
    .D(net1015),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[85][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2404_ (.RESET_B(net480),
    .D(net754),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[84][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2405_ (.RESET_B(net481),
    .D(net1002),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[84][1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2406_ (.RESET_B(net482),
    .D(net677),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[83][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2407_ (.RESET_B(net483),
    .D(net743),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[83][1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2408_ (.RESET_B(net484),
    .D(net1060),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[82][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2409_ (.RESET_B(net485),
    .D(net790),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[82][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2410_ (.RESET_B(net486),
    .D(net1113),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[81][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2411_ (.RESET_B(net487),
    .D(net780),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[81][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2412_ (.RESET_B(net488),
    .D(net989),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[80][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2413_ (.RESET_B(net489),
    .D(net1039),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[80][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2414_ (.RESET_B(net490),
    .D(net721),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[79][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2415_ (.RESET_B(net491),
    .D(net802),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[79][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2416_ (.RESET_B(net492),
    .D(net678),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[78][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2417_ (.RESET_B(net493),
    .D(net736),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[78][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2418_ (.RESET_B(net494),
    .D(net798),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[77][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2419_ (.RESET_B(net495),
    .D(net915),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[77][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2420_ (.RESET_B(net496),
    .D(net1020),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[76][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2421_ (.RESET_B(net497),
    .D(net923),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[76][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2422_ (.RESET_B(net498),
    .D(net734),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[75][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2423_ (.RESET_B(net499),
    .D(net825),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[75][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2424_ (.RESET_B(net500),
    .D(net686),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[74][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2425_ (.RESET_B(net501),
    .D(net697),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[74][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2426_ (.RESET_B(net502),
    .D(net1058),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[73][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2427_ (.RESET_B(net503),
    .D(net1027),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[73][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2428_ (.RESET_B(net504),
    .D(net667),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[72][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2429_ (.RESET_B(net505),
    .D(net840),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[72][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2430_ (.RESET_B(net506),
    .D(net714),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[71][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2431_ (.RESET_B(net507),
    .D(net1117),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[71][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2432_ (.RESET_B(net508),
    .D(net889),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[70][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2433_ (.RESET_B(net509),
    .D(net712),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[70][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2434_ (.RESET_B(net510),
    .D(net1034),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[69][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2435_ (.RESET_B(net511),
    .D(net1009),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[69][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2436_ (.RESET_B(net512),
    .D(net785),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[68][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2437_ (.RESET_B(net513),
    .D(net1043),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[68][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2438_ (.RESET_B(net514),
    .D(net1064),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[67][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2439_ (.RESET_B(net515),
    .D(net690),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[67][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2440_ (.RESET_B(net516),
    .D(net1019),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[66][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2441_ (.RESET_B(net517),
    .D(net706),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[66][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2442_ (.RESET_B(net518),
    .D(net1059),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[65][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2443_ (.RESET_B(net519),
    .D(net700),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[65][1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2444_ (.RESET_B(net520),
    .D(net1088),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[64][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2445_ (.RESET_B(net521),
    .D(net901),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[64][1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2446_ (.RESET_B(net522),
    .D(net877),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[63][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2447_ (.RESET_B(net523),
    .D(net1073),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[63][1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2448_ (.RESET_B(net524),
    .D(net952),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[62][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2449_ (.RESET_B(net525),
    .D(net1111),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[62][1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2450_ (.RESET_B(net526),
    .D(net669),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[61][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2451_ (.RESET_B(net527),
    .D(net707),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[61][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2452_ (.RESET_B(net528),
    .D(net788),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[60][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2453_ (.RESET_B(net529),
    .D(net1031),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[60][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2454_ (.RESET_B(net530),
    .D(net921),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[59][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2455_ (.RESET_B(net531),
    .D(net1024),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[59][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2456_ (.RESET_B(net532),
    .D(net811),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[58][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2457_ (.RESET_B(net533),
    .D(net1068),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[58][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2458_ (.RESET_B(net534),
    .D(net814),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[57][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2459_ (.RESET_B(net535),
    .D(net789),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[57][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2460_ (.RESET_B(net536),
    .D(net1022),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[56][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2461_ (.RESET_B(net537),
    .D(net820),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[56][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2462_ (.RESET_B(net538),
    .D(net1093),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[55][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2463_ (.RESET_B(net539),
    .D(net1087),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[55][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2464_ (.RESET_B(net540),
    .D(net943),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[54][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2465_ (.RESET_B(net541),
    .D(net913),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[54][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2466_ (.RESET_B(net542),
    .D(net1104),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[53][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2467_ (.RESET_B(net543),
    .D(net876),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[53][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2468_ (.RESET_B(net544),
    .D(net666),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[52][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2469_ (.RESET_B(net545),
    .D(net822),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[52][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2470_ (.RESET_B(net546),
    .D(net1049),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[51][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2471_ (.RESET_B(net547),
    .D(net878),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[51][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2472_ (.RESET_B(net548),
    .D(net930),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[50][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2473_ (.RESET_B(net549),
    .D(net942),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[50][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2474_ (.RESET_B(net550),
    .D(net1116),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[49][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2475_ (.RESET_B(net551),
    .D(net684),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[49][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2476_ (.RESET_B(net552),
    .D(net847),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[48][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2477_ (.RESET_B(net553),
    .D(net680),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[48][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2478_ (.RESET_B(net554),
    .D(net751),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[47][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2479_ (.RESET_B(net555),
    .D(net861),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[47][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2480_ (.RESET_B(net556),
    .D(net939),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[46][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2481_ (.RESET_B(net557),
    .D(net883),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[46][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2482_ (.RESET_B(net558),
    .D(net838),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[45][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2483_ (.RESET_B(net559),
    .D(net862),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[45][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2484_ (.RESET_B(net560),
    .D(net787),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[44][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2485_ (.RESET_B(net561),
    .D(net804),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[44][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2486_ (.RESET_B(net562),
    .D(net1006),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[43][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2487_ (.RESET_B(net563),
    .D(net752),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[43][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2488_ (.RESET_B(net564),
    .D(net850),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[42][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2489_ (.RESET_B(net565),
    .D(net779),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[42][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2490_ (.RESET_B(net566),
    .D(net801),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[41][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2491_ (.RESET_B(net567),
    .D(net827),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[41][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2492_ (.RESET_B(net568),
    .D(net665),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[40][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2493_ (.RESET_B(net569),
    .D(net717),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[40][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2494_ (.RESET_B(net570),
    .D(net1095),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[39][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2495_ (.RESET_B(net571),
    .D(net1103),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[39][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2496_ (.RESET_B(net572),
    .D(net765),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[38][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2497_ (.RESET_B(net573),
    .D(net926),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[38][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2498_ (.RESET_B(net574),
    .D(net959),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[37][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2499_ (.RESET_B(net575),
    .D(net963),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[37][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2500_ (.RESET_B(net576),
    .D(net1120),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[36][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2501_ (.RESET_B(net577),
    .D(net1076),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[36][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2502_ (.RESET_B(net578),
    .D(net1057),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[35][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2503_ (.RESET_B(net579),
    .D(net964),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[35][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2504_ (.RESET_B(net580),
    .D(net682),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[34][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2505_ (.RESET_B(net581),
    .D(net841),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[34][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2506_ (.RESET_B(net582),
    .D(net1021),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[33][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2507_ (.RESET_B(net583),
    .D(net893),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[33][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2508_ (.RESET_B(net584),
    .D(net738),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[32][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2509_ (.RESET_B(net585),
    .D(net1000),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[32][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2510_ (.RESET_B(net586),
    .D(net1054),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[31][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2511_ (.RESET_B(net587),
    .D(net695),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[31][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2512_ (.RESET_B(net588),
    .D(net1128),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[30][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2513_ (.RESET_B(net589),
    .D(net856),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[30][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2514_ (.RESET_B(net590),
    .D(net1046),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[29][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2515_ (.RESET_B(net591),
    .D(net741),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[29][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2516_ (.RESET_B(net592),
    .D(net833),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[28][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2517_ (.RESET_B(net593),
    .D(net1096),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[28][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2518_ (.RESET_B(net594),
    .D(net844),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[27][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2519_ (.RESET_B(net595),
    .D(net853),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[27][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2520_ (.RESET_B(net596),
    .D(net708),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[26][0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2521_ (.RESET_B(net597),
    .D(net884),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[26][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2522_ (.RESET_B(net598),
    .D(net701),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[25][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2523_ (.RESET_B(net599),
    .D(net994),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[25][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2524_ (.RESET_B(net600),
    .D(net713),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[24][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2525_ (.RESET_B(net601),
    .D(net1086),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[24][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2526_ (.RESET_B(net602),
    .D(net857),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[23][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2527_ (.RESET_B(net603),
    .D(net1082),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[23][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2528_ (.RESET_B(net604),
    .D(net1007),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[22][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2529_ (.RESET_B(net605),
    .D(net1067),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[22][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2530_ (.RESET_B(net606),
    .D(net726),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[21][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2531_ (.RESET_B(net607),
    .D(net831),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[21][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2532_ (.RESET_B(net608),
    .D(net1025),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[20][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2533_ (.RESET_B(net609),
    .D(net842),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[20][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2534_ (.RESET_B(net610),
    .D(net773),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[19][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2535_ (.RESET_B(net611),
    .D(net924),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[19][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2536_ (.RESET_B(net612),
    .D(net1129),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[18][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2537_ (.RESET_B(net613),
    .D(net1040),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[18][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2538_ (.RESET_B(net614),
    .D(net679),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[17][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2539_ (.RESET_B(net615),
    .D(net843),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[17][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2540_ (.RESET_B(net616),
    .D(net725),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[16][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2541_ (.RESET_B(net617),
    .D(net927),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[16][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2542_ (.RESET_B(net618),
    .D(net904),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[15][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2543_ (.RESET_B(net619),
    .D(net1107),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[15][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2544_ (.RESET_B(net620),
    .D(net760),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[14][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2545_ (.RESET_B(net621),
    .D(net966),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[14][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2546_ (.RESET_B(net622),
    .D(net1014),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[13][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2547_ (.RESET_B(net623),
    .D(net768),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[13][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2548_ (.RESET_B(net624),
    .D(net823),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[12][0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2549_ (.RESET_B(net625),
    .D(net750),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[12][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2550_ (.RESET_B(net626),
    .D(net807),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[11][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2551_ (.RESET_B(net627),
    .D(net870),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[11][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2552_ (.RESET_B(net628),
    .D(net882),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[10][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2553_ (.RESET_B(net629),
    .D(net981),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[10][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2554_ (.RESET_B(net630),
    .D(net1100),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[9][0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2555_ (.RESET_B(net631),
    .D(net839),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[9][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2556_ (.RESET_B(net632),
    .D(net992),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[8][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2557_ (.RESET_B(net633),
    .D(net1048),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[8][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2558_ (.RESET_B(net634),
    .D(net978),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[7][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2559_ (.RESET_B(net635),
    .D(net735),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[7][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2560_ (.RESET_B(net636),
    .D(net946),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[6][0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2561_ (.RESET_B(net637),
    .D(net873),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[6][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2562_ (.RESET_B(net638),
    .D(net729),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[5][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2563_ (.RESET_B(net639),
    .D(net902),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[5][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2564_ (.RESET_B(net640),
    .D(net795),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[4][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2565_ (.RESET_B(net641),
    .D(net910),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[4][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2566_ (.RESET_B(net642),
    .D(net782),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[3][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2567_ (.RESET_B(net643),
    .D(net791),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[3][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2568_ (.RESET_B(net644),
    .D(net761),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[2][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2569_ (.RESET_B(net645),
    .D(net1130),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[2][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2570_ (.RESET_B(net656),
    .D(net1131),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[1][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2571_ (.RESET_B(net171),
    .D(net122),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2572_ (.RESET_B(net169),
    .D(net1147),
    .Q(\game_inst.o_tick ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2573_ (.RESET_B(net167),
    .D(_0122_),
    .Q(\game_inst.apple_inst.apple_y[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2574_ (.RESET_B(net165),
    .D(net1170),
    .Q(\game_inst.apple_inst.apple_y[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2575_ (.RESET_B(net163),
    .D(_0124_),
    .Q(\game_inst.apple_inst.apple_y[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _2576_ (.RESET_B(net161),
    .D(net1182),
    .Q(\game_inst.apple_inst.apple_y[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2577_ (.RESET_B(net159),
    .D(_0126_),
    .Q(\game_inst.control_inst.o_start ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2578_ (.RESET_B(net157),
    .D(_0127_),
    .Q(\game_inst.tickgen_inst.counter_max[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2579_ (.RESET_B(net153),
    .D(net1344),
    .Q(\game_inst.tickgen_inst.counter_max[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2580_ (.RESET_B(net149),
    .D(net1260),
    .Q(\game_inst.tickgen_inst.counter_max[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2581_ (.RESET_B(net155),
    .D(net1187),
    .Q(\game_inst.tick ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2582_ (.RESET_B(net145),
    .D(_0003_),
    .Q(\game_inst.tickgen_inst.prev_user_input ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2583_ (.RESET_B(net31),
    .D(_0131_),
    .Q(\game_inst.tickgen_inst.counter[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2584_ (.RESET_B(net151),
    .D(_0132_),
    .Q(\game_inst.tickgen_inst.counter[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2585_ (.RESET_B(net143),
    .D(_0133_),
    .Q(\game_inst.tickgen_inst.counter[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2586_ (.RESET_B(net147),
    .D(net1151),
    .Q(\game_inst.tickgen_inst.counter[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_tiehi _2096__16 (.L_HI(net16));
 sg13g2_tiehi _2052__17 (.L_HI(net17));
 sg13g2_tiehi _2095__18 (.L_HI(net18));
 sg13g2_tiehi _2051__19 (.L_HI(net19));
 sg13g2_tiehi _2094__20 (.L_HI(net20));
 sg13g2_tiehi _2050__21 (.L_HI(net21));
 sg13g2_tiehi _2093__22 (.L_HI(net22));
 sg13g2_tiehi _2049__23 (.L_HI(net23));
 sg13g2_tiehi _2092__24 (.L_HI(net24));
 sg13g2_tiehi _1984__25 (.L_HI(net25));
 sg13g2_tiehi _1993__26 (.L_HI(net26));
 sg13g2_tiehi _1994__27 (.L_HI(net27));
 sg13g2_tiehi _2048__28 (.L_HI(net28));
 sg13g2_tiehi _2091__29 (.L_HI(net29));
 sg13g2_tiehi _2047__30 (.L_HI(net30));
 sg13g2_tiehi _2583__31 (.L_HI(net31));
 sg13g2_tiehi _2046__32 (.L_HI(net32));
 sg13g2_tiehi _1995__33 (.L_HI(net33));
 sg13g2_tiehi _2001__34 (.L_HI(net34));
 sg13g2_tiehi _2002__35 (.L_HI(net35));
 sg13g2_tiehi _2003__36 (.L_HI(net36));
 sg13g2_tiehi _2004__37 (.L_HI(net37));
 sg13g2_tiehi _2005__38 (.L_HI(net38));
 sg13g2_tiehi _2006__39 (.L_HI(net39));
 sg13g2_tiehi _2090__40 (.L_HI(net40));
 sg13g2_tiehi _2045__41 (.L_HI(net41));
 sg13g2_tiehi _2007__42 (.L_HI(net42));
 sg13g2_tiehi _2010__43 (.L_HI(net43));
 sg13g2_tiehi _2011__44 (.L_HI(net44));
 sg13g2_tiehi _2012__45 (.L_HI(net45));
 sg13g2_tiehi _2013__46 (.L_HI(net46));
 sg13g2_tiehi _2014__47 (.L_HI(net47));
 sg13g2_tiehi _2015__48 (.L_HI(net48));
 sg13g2_tiehi _2016__49 (.L_HI(net49));
 sg13g2_tiehi _2017__50 (.L_HI(net50));
 sg13g2_tiehi _2018__51 (.L_HI(net51));
 sg13g2_tiehi _2019__52 (.L_HI(net52));
 sg13g2_tiehi _2020__53 (.L_HI(net53));
 sg13g2_tiehi _2021__54 (.L_HI(net54));
 sg13g2_tiehi _2022__55 (.L_HI(net55));
 sg13g2_tiehi _2023__56 (.L_HI(net56));
 sg13g2_tiehi _2024__57 (.L_HI(net57));
 sg13g2_tiehi _2025__58 (.L_HI(net58));
 sg13g2_tiehi _2026__59 (.L_HI(net59));
 sg13g2_tiehi _2027__60 (.L_HI(net60));
 sg13g2_tiehi _2028__61 (.L_HI(net61));
 sg13g2_tiehi _2029__62 (.L_HI(net62));
 sg13g2_tiehi _2030__63 (.L_HI(net63));
 sg13g2_tiehi _2031__64 (.L_HI(net64));
 sg13g2_tiehi _2032__65 (.L_HI(net65));
 sg13g2_tiehi _2033__66 (.L_HI(net66));
 sg13g2_tiehi _2034__67 (.L_HI(net67));
 sg13g2_tiehi _2035__68 (.L_HI(net68));
 sg13g2_tiehi _2036__69 (.L_HI(net69));
 sg13g2_tiehi _2089__70 (.L_HI(net70));
 sg13g2_tiehi _2044__71 (.L_HI(net71));
 sg13g2_tiehi _2043__72 (.L_HI(net72));
 sg13g2_tiehi _2041__73 (.L_HI(net73));
 sg13g2_tiehi _2037__74 (.L_HI(net74));
 sg13g2_tiehi _2040__75 (.L_HI(net75));
 sg13g2_tiehi _2039__76 (.L_HI(net76));
 sg13g2_tiehi _2038__77 (.L_HI(net77));
 sg13g2_tiehi _2009__78 (.L_HI(net78));
 sg13g2_tiehi _2008__79 (.L_HI(net79));
 sg13g2_tiehi _2000__80 (.L_HI(net80));
 sg13g2_tiehi _1999__81 (.L_HI(net81));
 sg13g2_tiehi _1998__82 (.L_HI(net82));
 sg13g2_tiehi _1997__83 (.L_HI(net83));
 sg13g2_tiehi _1996__84 (.L_HI(net84));
 sg13g2_tiehi _2042__85 (.L_HI(net85));
 sg13g2_tiehi _1992__86 (.L_HI(net86));
 sg13g2_tiehi _1991__87 (.L_HI(net87));
 sg13g2_tiehi _1990__88 (.L_HI(net88));
 sg13g2_tiehi _1989__89 (.L_HI(net89));
 sg13g2_tiehi _1988__90 (.L_HI(net90));
 sg13g2_tiehi _1987__91 (.L_HI(net91));
 sg13g2_tiehi _1986__92 (.L_HI(net92));
 sg13g2_tiehi _1985__93 (.L_HI(net93));
 sg13g2_tiehi _2088__94 (.L_HI(net137));
 sg13g2_tiehi _2087__95 (.L_HI(net138));
 sg13g2_tiehi _2086__96 (.L_HI(net139));
 sg13g2_tiehi _2085__97 (.L_HI(net140));
 sg13g2_tiehi _2084__98 (.L_HI(net141));
 sg13g2_tiehi _2083__99 (.L_HI(net142));
 sg13g2_tiehi _2585__100 (.L_HI(net143));
 sg13g2_tiehi _2082__101 (.L_HI(net144));
 sg13g2_tiehi _2582__102 (.L_HI(net145));
 sg13g2_tiehi _2081__103 (.L_HI(net146));
 sg13g2_tiehi _2586__104 (.L_HI(net147));
 sg13g2_tiehi _2080__105 (.L_HI(net148));
 sg13g2_tiehi _2580__106 (.L_HI(net149));
 sg13g2_tiehi _2079__107 (.L_HI(net150));
 sg13g2_tiehi _2584__108 (.L_HI(net151));
 sg13g2_tiehi _2078__109 (.L_HI(net152));
 sg13g2_tiehi _2579__110 (.L_HI(net153));
 sg13g2_tiehi _2077__111 (.L_HI(net154));
 sg13g2_tiehi _2581__112 (.L_HI(net155));
 sg13g2_tiehi _2076__113 (.L_HI(net156));
 sg13g2_tiehi _2578__114 (.L_HI(net157));
 sg13g2_tiehi _2075__115 (.L_HI(net158));
 sg13g2_tiehi _2577__116 (.L_HI(net159));
 sg13g2_tiehi _2074__117 (.L_HI(net160));
 sg13g2_tiehi _2576__118 (.L_HI(net161));
 sg13g2_tiehi _2073__119 (.L_HI(net162));
 sg13g2_tiehi _2575__120 (.L_HI(net163));
 sg13g2_tiehi _2072__121 (.L_HI(net164));
 sg13g2_tiehi _2574__122 (.L_HI(net165));
 sg13g2_tiehi _2071__123 (.L_HI(net166));
 sg13g2_tiehi _2573__124 (.L_HI(net167));
 sg13g2_tiehi _2070__125 (.L_HI(net168));
 sg13g2_tiehi _2572__126 (.L_HI(net169));
 sg13g2_tiehi _2069__127 (.L_HI(net170));
 sg13g2_tiehi _2571__128 (.L_HI(net171));
 sg13g2_tiehi _2068__129 (.L_HI(net172));
 sg13g2_tiehi _2104__130 (.L_HI(net173));
 sg13g2_tiehi _2067__131 (.L_HI(net174));
 sg13g2_tiehi _2103__132 (.L_HI(net175));
 sg13g2_tiehi _2066__133 (.L_HI(net176));
 sg13g2_tiehi _2102__134 (.L_HI(net177));
 sg13g2_tiehi _2065__135 (.L_HI(net178));
 sg13g2_tiehi _2101__136 (.L_HI(net179));
 sg13g2_tiehi _2053__137 (.L_HI(net180));
 sg13g2_tiehi _2105__138 (.L_HI(net181));
 sg13g2_tiehi _2106__139 (.L_HI(net182));
 sg13g2_tiehi _2107__140 (.L_HI(net183));
 sg13g2_tiehi _2108__141 (.L_HI(net184));
 sg13g2_tiehi _2109__142 (.L_HI(net185));
 sg13g2_tiehi _2110__143 (.L_HI(net186));
 sg13g2_tiehi _2111__144 (.L_HI(net187));
 sg13g2_tiehi _2112__145 (.L_HI(net188));
 sg13g2_tiehi _2113__146 (.L_HI(net189));
 sg13g2_tiehi _2114__147 (.L_HI(net190));
 sg13g2_tiehi _2115__148 (.L_HI(net191));
 sg13g2_tiehi _2116__149 (.L_HI(net192));
 sg13g2_tiehi _2117__150 (.L_HI(net193));
 sg13g2_tiehi _2118__151 (.L_HI(net194));
 sg13g2_tiehi _2119__152 (.L_HI(net195));
 sg13g2_tiehi _2120__153 (.L_HI(net196));
 sg13g2_tiehi _2121__154 (.L_HI(net197));
 sg13g2_tiehi _2122__155 (.L_HI(net198));
 sg13g2_tiehi _2123__156 (.L_HI(net199));
 sg13g2_tiehi _2124__157 (.L_HI(net200));
 sg13g2_tiehi _2125__158 (.L_HI(net201));
 sg13g2_tiehi _2126__159 (.L_HI(net202));
 sg13g2_tiehi _2127__160 (.L_HI(net203));
 sg13g2_tiehi _2128__161 (.L_HI(net204));
 sg13g2_tiehi _2129__162 (.L_HI(net205));
 sg13g2_tiehi _2130__163 (.L_HI(net206));
 sg13g2_tiehi _2131__164 (.L_HI(net207));
 sg13g2_tiehi _2132__165 (.L_HI(net208));
 sg13g2_tiehi _2133__166 (.L_HI(net209));
 sg13g2_tiehi _2134__167 (.L_HI(net210));
 sg13g2_tiehi _2135__168 (.L_HI(net211));
 sg13g2_tiehi _2136__169 (.L_HI(net212));
 sg13g2_tiehi _2137__170 (.L_HI(net213));
 sg13g2_tiehi _2138__171 (.L_HI(net214));
 sg13g2_tiehi _2139__172 (.L_HI(net215));
 sg13g2_tiehi _2140__173 (.L_HI(net216));
 sg13g2_tiehi _2141__174 (.L_HI(net217));
 sg13g2_tiehi _2142__175 (.L_HI(net218));
 sg13g2_tiehi _2143__176 (.L_HI(net219));
 sg13g2_tiehi _2144__177 (.L_HI(net220));
 sg13g2_tiehi _2145__178 (.L_HI(net221));
 sg13g2_tiehi _2146__179 (.L_HI(net222));
 sg13g2_tiehi _2147__180 (.L_HI(net223));
 sg13g2_tiehi _2148__181 (.L_HI(net224));
 sg13g2_tiehi _2149__182 (.L_HI(net225));
 sg13g2_tiehi _2150__183 (.L_HI(net226));
 sg13g2_tiehi _2151__184 (.L_HI(net227));
 sg13g2_tiehi _2152__185 (.L_HI(net228));
 sg13g2_tiehi _2153__186 (.L_HI(net229));
 sg13g2_tiehi _2154__187 (.L_HI(net230));
 sg13g2_tiehi _2155__188 (.L_HI(net231));
 sg13g2_tiehi _2156__189 (.L_HI(net232));
 sg13g2_tiehi _2157__190 (.L_HI(net233));
 sg13g2_tiehi _2158__191 (.L_HI(net234));
 sg13g2_tiehi _2159__192 (.L_HI(net235));
 sg13g2_tiehi _2160__193 (.L_HI(net236));
 sg13g2_tiehi _2161__194 (.L_HI(net237));
 sg13g2_tiehi _2162__195 (.L_HI(net238));
 sg13g2_tiehi _2163__196 (.L_HI(net239));
 sg13g2_tiehi _2164__197 (.L_HI(net240));
 sg13g2_tiehi _2165__198 (.L_HI(net241));
 sg13g2_tiehi _2166__199 (.L_HI(net242));
 sg13g2_tiehi _2167__200 (.L_HI(net243));
 sg13g2_tiehi _2168__201 (.L_HI(net244));
 sg13g2_tiehi _2169__202 (.L_HI(net245));
 sg13g2_tiehi _2170__203 (.L_HI(net246));
 sg13g2_tiehi _2171__204 (.L_HI(net247));
 sg13g2_tiehi _2172__205 (.L_HI(net248));
 sg13g2_tiehi _2173__206 (.L_HI(net249));
 sg13g2_tiehi _2174__207 (.L_HI(net250));
 sg13g2_tiehi _2175__208 (.L_HI(net251));
 sg13g2_tiehi _2176__209 (.L_HI(net252));
 sg13g2_tiehi _2177__210 (.L_HI(net253));
 sg13g2_tiehi _2178__211 (.L_HI(net254));
 sg13g2_tiehi _2179__212 (.L_HI(net255));
 sg13g2_tiehi _2180__213 (.L_HI(net256));
 sg13g2_tiehi _2181__214 (.L_HI(net257));
 sg13g2_tiehi _2182__215 (.L_HI(net258));
 sg13g2_tiehi _2183__216 (.L_HI(net259));
 sg13g2_tiehi _2184__217 (.L_HI(net260));
 sg13g2_tiehi _2185__218 (.L_HI(net261));
 sg13g2_tiehi _2186__219 (.L_HI(net262));
 sg13g2_tiehi _2187__220 (.L_HI(net263));
 sg13g2_tiehi _2188__221 (.L_HI(net264));
 sg13g2_tiehi _2189__222 (.L_HI(net265));
 sg13g2_tiehi _2190__223 (.L_HI(net266));
 sg13g2_tiehi _2191__224 (.L_HI(net267));
 sg13g2_tiehi _2192__225 (.L_HI(net268));
 sg13g2_tiehi _2193__226 (.L_HI(net269));
 sg13g2_tiehi _2194__227 (.L_HI(net270));
 sg13g2_tiehi _2195__228 (.L_HI(net271));
 sg13g2_tiehi _2196__229 (.L_HI(net272));
 sg13g2_tiehi _2197__230 (.L_HI(net273));
 sg13g2_tiehi _2198__231 (.L_HI(net274));
 sg13g2_tiehi _2199__232 (.L_HI(net275));
 sg13g2_tiehi _2200__233 (.L_HI(net276));
 sg13g2_tiehi _2201__234 (.L_HI(net277));
 sg13g2_tiehi _2202__235 (.L_HI(net278));
 sg13g2_tiehi _2203__236 (.L_HI(net279));
 sg13g2_tiehi _2204__237 (.L_HI(net280));
 sg13g2_tiehi _2205__238 (.L_HI(net281));
 sg13g2_tiehi _2206__239 (.L_HI(net282));
 sg13g2_tiehi _2207__240 (.L_HI(net283));
 sg13g2_tiehi _2208__241 (.L_HI(net284));
 sg13g2_tiehi _2209__242 (.L_HI(net285));
 sg13g2_tiehi _2210__243 (.L_HI(net286));
 sg13g2_tiehi _2211__244 (.L_HI(net287));
 sg13g2_tiehi _2212__245 (.L_HI(net288));
 sg13g2_tiehi _2213__246 (.L_HI(net289));
 sg13g2_tiehi _2214__247 (.L_HI(net290));
 sg13g2_tiehi _2215__248 (.L_HI(net291));
 sg13g2_tiehi _2216__249 (.L_HI(net292));
 sg13g2_tiehi _2217__250 (.L_HI(net293));
 sg13g2_tiehi _2218__251 (.L_HI(net294));
 sg13g2_tiehi _2219__252 (.L_HI(net295));
 sg13g2_tiehi _2220__253 (.L_HI(net296));
 sg13g2_tiehi _2221__254 (.L_HI(net297));
 sg13g2_tiehi _2222__255 (.L_HI(net298));
 sg13g2_tiehi _2223__256 (.L_HI(net299));
 sg13g2_tiehi _2224__257 (.L_HI(net300));
 sg13g2_tiehi _2225__258 (.L_HI(net301));
 sg13g2_tiehi _2226__259 (.L_HI(net302));
 sg13g2_tiehi _2227__260 (.L_HI(net303));
 sg13g2_tiehi _2228__261 (.L_HI(net304));
 sg13g2_tiehi _2229__262 (.L_HI(net305));
 sg13g2_tiehi _2230__263 (.L_HI(net306));
 sg13g2_tiehi _2231__264 (.L_HI(net307));
 sg13g2_tiehi _2232__265 (.L_HI(net308));
 sg13g2_tiehi _2233__266 (.L_HI(net309));
 sg13g2_tiehi _2234__267 (.L_HI(net310));
 sg13g2_tiehi _2235__268 (.L_HI(net311));
 sg13g2_tiehi _2236__269 (.L_HI(net312));
 sg13g2_tiehi _2237__270 (.L_HI(net313));
 sg13g2_tiehi _2238__271 (.L_HI(net314));
 sg13g2_tiehi _2239__272 (.L_HI(net315));
 sg13g2_tiehi _2240__273 (.L_HI(net316));
 sg13g2_tiehi _2241__274 (.L_HI(net317));
 sg13g2_tiehi _2242__275 (.L_HI(net318));
 sg13g2_tiehi _2243__276 (.L_HI(net319));
 sg13g2_tiehi _2244__277 (.L_HI(net320));
 sg13g2_tiehi _2245__278 (.L_HI(net321));
 sg13g2_tiehi _2246__279 (.L_HI(net322));
 sg13g2_tiehi _2247__280 (.L_HI(net323));
 sg13g2_tiehi _2248__281 (.L_HI(net324));
 sg13g2_tiehi _2249__282 (.L_HI(net325));
 sg13g2_tiehi _2250__283 (.L_HI(net326));
 sg13g2_tiehi _2251__284 (.L_HI(net327));
 sg13g2_tiehi _2252__285 (.L_HI(net328));
 sg13g2_tiehi _2253__286 (.L_HI(net329));
 sg13g2_tiehi _2254__287 (.L_HI(net330));
 sg13g2_tiehi _2255__288 (.L_HI(net331));
 sg13g2_tiehi _2256__289 (.L_HI(net332));
 sg13g2_tiehi _2257__290 (.L_HI(net333));
 sg13g2_tiehi _2258__291 (.L_HI(net334));
 sg13g2_tiehi _2259__292 (.L_HI(net335));
 sg13g2_tiehi _2260__293 (.L_HI(net336));
 sg13g2_tiehi _2261__294 (.L_HI(net337));
 sg13g2_tiehi _2262__295 (.L_HI(net338));
 sg13g2_tiehi _2263__296 (.L_HI(net339));
 sg13g2_tiehi _2264__297 (.L_HI(net340));
 sg13g2_tiehi _2265__298 (.L_HI(net341));
 sg13g2_tiehi _2266__299 (.L_HI(net342));
 sg13g2_tiehi _2267__300 (.L_HI(net343));
 sg13g2_tiehi _2268__301 (.L_HI(net344));
 sg13g2_tiehi _2269__302 (.L_HI(net345));
 sg13g2_tiehi _2270__303 (.L_HI(net346));
 sg13g2_tiehi _2271__304 (.L_HI(net347));
 sg13g2_tiehi _2272__305 (.L_HI(net348));
 sg13g2_tiehi _2273__306 (.L_HI(net349));
 sg13g2_tiehi _2274__307 (.L_HI(net350));
 sg13g2_tiehi _2275__308 (.L_HI(net351));
 sg13g2_tiehi _2276__309 (.L_HI(net352));
 sg13g2_tiehi _2277__310 (.L_HI(net353));
 sg13g2_tiehi _2278__311 (.L_HI(net354));
 sg13g2_tiehi _2279__312 (.L_HI(net355));
 sg13g2_tiehi _2280__313 (.L_HI(net356));
 sg13g2_tiehi _2281__314 (.L_HI(net357));
 sg13g2_tiehi _2282__315 (.L_HI(net358));
 sg13g2_tiehi _2283__316 (.L_HI(net359));
 sg13g2_tiehi _2284__317 (.L_HI(net360));
 sg13g2_tiehi _2285__318 (.L_HI(net361));
 sg13g2_tiehi _2286__319 (.L_HI(net362));
 sg13g2_tiehi _2287__320 (.L_HI(net363));
 sg13g2_tiehi _2288__321 (.L_HI(net364));
 sg13g2_tiehi _2289__322 (.L_HI(net365));
 sg13g2_tiehi _2290__323 (.L_HI(net366));
 sg13g2_tiehi _2291__324 (.L_HI(net367));
 sg13g2_tiehi _2292__325 (.L_HI(net368));
 sg13g2_tiehi _2293__326 (.L_HI(net369));
 sg13g2_tiehi _2294__327 (.L_HI(net370));
 sg13g2_tiehi _2295__328 (.L_HI(net371));
 sg13g2_tiehi _2296__329 (.L_HI(net372));
 sg13g2_tiehi _2297__330 (.L_HI(net373));
 sg13g2_tiehi _2298__331 (.L_HI(net374));
 sg13g2_tiehi _2299__332 (.L_HI(net375));
 sg13g2_tiehi _2300__333 (.L_HI(net376));
 sg13g2_tiehi _2301__334 (.L_HI(net377));
 sg13g2_tiehi _2302__335 (.L_HI(net378));
 sg13g2_tiehi _2303__336 (.L_HI(net379));
 sg13g2_tiehi _2304__337 (.L_HI(net380));
 sg13g2_tiehi _2305__338 (.L_HI(net381));
 sg13g2_tiehi _2306__339 (.L_HI(net382));
 sg13g2_tiehi _2307__340 (.L_HI(net383));
 sg13g2_tiehi _2308__341 (.L_HI(net384));
 sg13g2_tiehi _2309__342 (.L_HI(net385));
 sg13g2_tiehi _2310__343 (.L_HI(net386));
 sg13g2_tiehi _2311__344 (.L_HI(net387));
 sg13g2_tiehi _2312__345 (.L_HI(net388));
 sg13g2_tiehi _2313__346 (.L_HI(net389));
 sg13g2_tiehi _2314__347 (.L_HI(net390));
 sg13g2_tiehi _2315__348 (.L_HI(net391));
 sg13g2_tiehi _2316__349 (.L_HI(net392));
 sg13g2_tiehi _2317__350 (.L_HI(net393));
 sg13g2_tiehi _2318__351 (.L_HI(net394));
 sg13g2_tiehi _2319__352 (.L_HI(net395));
 sg13g2_tiehi _2320__353 (.L_HI(net396));
 sg13g2_tiehi _2321__354 (.L_HI(net397));
 sg13g2_tiehi _2322__355 (.L_HI(net398));
 sg13g2_tiehi _2323__356 (.L_HI(net399));
 sg13g2_tiehi _2324__357 (.L_HI(net400));
 sg13g2_tiehi _2325__358 (.L_HI(net401));
 sg13g2_tiehi _2326__359 (.L_HI(net402));
 sg13g2_tiehi _2327__360 (.L_HI(net403));
 sg13g2_tiehi _2328__361 (.L_HI(net404));
 sg13g2_tiehi _2329__362 (.L_HI(net405));
 sg13g2_tiehi _2330__363 (.L_HI(net406));
 sg13g2_tiehi _2331__364 (.L_HI(net407));
 sg13g2_tiehi _2332__365 (.L_HI(net408));
 sg13g2_tiehi _2333__366 (.L_HI(net409));
 sg13g2_tiehi _2334__367 (.L_HI(net410));
 sg13g2_tiehi _2335__368 (.L_HI(net411));
 sg13g2_tiehi _2336__369 (.L_HI(net412));
 sg13g2_tiehi _2337__370 (.L_HI(net413));
 sg13g2_tiehi _2338__371 (.L_HI(net414));
 sg13g2_tiehi _2339__372 (.L_HI(net415));
 sg13g2_tiehi _2340__373 (.L_HI(net416));
 sg13g2_tiehi _2341__374 (.L_HI(net417));
 sg13g2_tiehi _2342__375 (.L_HI(net418));
 sg13g2_tiehi _2343__376 (.L_HI(net419));
 sg13g2_tiehi _2344__377 (.L_HI(net420));
 sg13g2_tiehi _2345__378 (.L_HI(net421));
 sg13g2_tiehi _2346__379 (.L_HI(net422));
 sg13g2_tiehi _2347__380 (.L_HI(net423));
 sg13g2_tiehi _2348__381 (.L_HI(net424));
 sg13g2_tiehi _2349__382 (.L_HI(net425));
 sg13g2_tiehi _2350__383 (.L_HI(net426));
 sg13g2_tiehi _2351__384 (.L_HI(net427));
 sg13g2_tiehi _2352__385 (.L_HI(net428));
 sg13g2_tiehi _2353__386 (.L_HI(net429));
 sg13g2_tiehi _2354__387 (.L_HI(net430));
 sg13g2_tiehi _2355__388 (.L_HI(net431));
 sg13g2_tiehi _2356__389 (.L_HI(net432));
 sg13g2_tiehi _2357__390 (.L_HI(net433));
 sg13g2_tiehi _2358__391 (.L_HI(net434));
 sg13g2_tiehi _2359__392 (.L_HI(net435));
 sg13g2_tiehi _2360__393 (.L_HI(net436));
 sg13g2_tiehi _2361__394 (.L_HI(net437));
 sg13g2_tiehi _2362__395 (.L_HI(net438));
 sg13g2_tiehi _2363__396 (.L_HI(net439));
 sg13g2_tiehi _2364__397 (.L_HI(net440));
 sg13g2_tiehi _2365__398 (.L_HI(net441));
 sg13g2_tiehi _2366__399 (.L_HI(net442));
 sg13g2_tiehi _2367__400 (.L_HI(net443));
 sg13g2_tiehi _2368__401 (.L_HI(net444));
 sg13g2_tiehi _2369__402 (.L_HI(net445));
 sg13g2_tiehi _2370__403 (.L_HI(net446));
 sg13g2_tiehi _2371__404 (.L_HI(net447));
 sg13g2_tiehi _2372__405 (.L_HI(net448));
 sg13g2_tiehi _2373__406 (.L_HI(net449));
 sg13g2_tiehi _2374__407 (.L_HI(net450));
 sg13g2_tiehi _2375__408 (.L_HI(net451));
 sg13g2_tiehi _2376__409 (.L_HI(net452));
 sg13g2_tiehi _2377__410 (.L_HI(net453));
 sg13g2_tiehi _2378__411 (.L_HI(net454));
 sg13g2_tiehi _2379__412 (.L_HI(net455));
 sg13g2_tiehi _2380__413 (.L_HI(net456));
 sg13g2_tiehi _2381__414 (.L_HI(net457));
 sg13g2_tiehi _2382__415 (.L_HI(net458));
 sg13g2_tiehi _2383__416 (.L_HI(net459));
 sg13g2_tiehi _2384__417 (.L_HI(net460));
 sg13g2_tiehi _2385__418 (.L_HI(net461));
 sg13g2_tiehi _2386__419 (.L_HI(net462));
 sg13g2_tiehi _2387__420 (.L_HI(net463));
 sg13g2_tiehi _2388__421 (.L_HI(net464));
 sg13g2_tiehi _2389__422 (.L_HI(net465));
 sg13g2_tiehi _2390__423 (.L_HI(net466));
 sg13g2_tiehi _2391__424 (.L_HI(net467));
 sg13g2_tiehi _2392__425 (.L_HI(net468));
 sg13g2_tiehi _2393__426 (.L_HI(net469));
 sg13g2_tiehi _2394__427 (.L_HI(net470));
 sg13g2_tiehi _2395__428 (.L_HI(net471));
 sg13g2_tiehi _2396__429 (.L_HI(net472));
 sg13g2_tiehi _2397__430 (.L_HI(net473));
 sg13g2_tiehi _2398__431 (.L_HI(net474));
 sg13g2_tiehi _2399__432 (.L_HI(net475));
 sg13g2_tiehi _2400__433 (.L_HI(net476));
 sg13g2_tiehi _2401__434 (.L_HI(net477));
 sg13g2_tiehi _2402__435 (.L_HI(net478));
 sg13g2_tiehi _2403__436 (.L_HI(net479));
 sg13g2_tiehi _2404__437 (.L_HI(net480));
 sg13g2_tiehi _2405__438 (.L_HI(net481));
 sg13g2_tiehi _2406__439 (.L_HI(net482));
 sg13g2_tiehi _2407__440 (.L_HI(net483));
 sg13g2_tiehi _2408__441 (.L_HI(net484));
 sg13g2_tiehi _2409__442 (.L_HI(net485));
 sg13g2_tiehi _2410__443 (.L_HI(net486));
 sg13g2_tiehi _2411__444 (.L_HI(net487));
 sg13g2_tiehi _2412__445 (.L_HI(net488));
 sg13g2_tiehi _2413__446 (.L_HI(net489));
 sg13g2_tiehi _2414__447 (.L_HI(net490));
 sg13g2_tiehi _2415__448 (.L_HI(net491));
 sg13g2_tiehi _2416__449 (.L_HI(net492));
 sg13g2_tiehi _2417__450 (.L_HI(net493));
 sg13g2_tiehi _2418__451 (.L_HI(net494));
 sg13g2_tiehi _2419__452 (.L_HI(net495));
 sg13g2_tiehi _2420__453 (.L_HI(net496));
 sg13g2_tiehi _2421__454 (.L_HI(net497));
 sg13g2_tiehi _2422__455 (.L_HI(net498));
 sg13g2_tiehi _2423__456 (.L_HI(net499));
 sg13g2_tiehi _2424__457 (.L_HI(net500));
 sg13g2_tiehi _2425__458 (.L_HI(net501));
 sg13g2_tiehi _2426__459 (.L_HI(net502));
 sg13g2_tiehi _2427__460 (.L_HI(net503));
 sg13g2_tiehi _2428__461 (.L_HI(net504));
 sg13g2_tiehi _2429__462 (.L_HI(net505));
 sg13g2_tiehi _2430__463 (.L_HI(net506));
 sg13g2_tiehi _2431__464 (.L_HI(net507));
 sg13g2_tiehi _2432__465 (.L_HI(net508));
 sg13g2_tiehi _2433__466 (.L_HI(net509));
 sg13g2_tiehi _2434__467 (.L_HI(net510));
 sg13g2_tiehi _2435__468 (.L_HI(net511));
 sg13g2_tiehi _2436__469 (.L_HI(net512));
 sg13g2_tiehi _2437__470 (.L_HI(net513));
 sg13g2_tiehi _2438__471 (.L_HI(net514));
 sg13g2_tiehi _2439__472 (.L_HI(net515));
 sg13g2_tiehi _2440__473 (.L_HI(net516));
 sg13g2_tiehi _2441__474 (.L_HI(net517));
 sg13g2_tiehi _2442__475 (.L_HI(net518));
 sg13g2_tiehi _2443__476 (.L_HI(net519));
 sg13g2_tiehi _2444__477 (.L_HI(net520));
 sg13g2_tiehi _2445__478 (.L_HI(net521));
 sg13g2_tiehi _2446__479 (.L_HI(net522));
 sg13g2_tiehi _2447__480 (.L_HI(net523));
 sg13g2_tiehi _2448__481 (.L_HI(net524));
 sg13g2_tiehi _2449__482 (.L_HI(net525));
 sg13g2_tiehi _2450__483 (.L_HI(net526));
 sg13g2_tiehi _2451__484 (.L_HI(net527));
 sg13g2_tiehi _2452__485 (.L_HI(net528));
 sg13g2_tiehi _2453__486 (.L_HI(net529));
 sg13g2_tiehi _2454__487 (.L_HI(net530));
 sg13g2_tiehi _2455__488 (.L_HI(net531));
 sg13g2_tiehi _2456__489 (.L_HI(net532));
 sg13g2_tiehi _2457__490 (.L_HI(net533));
 sg13g2_tiehi _2458__491 (.L_HI(net534));
 sg13g2_tiehi _2459__492 (.L_HI(net535));
 sg13g2_tiehi _2460__493 (.L_HI(net536));
 sg13g2_tiehi _2461__494 (.L_HI(net537));
 sg13g2_tiehi _2462__495 (.L_HI(net538));
 sg13g2_tiehi _2463__496 (.L_HI(net539));
 sg13g2_tiehi _2464__497 (.L_HI(net540));
 sg13g2_tiehi _2465__498 (.L_HI(net541));
 sg13g2_tiehi _2466__499 (.L_HI(net542));
 sg13g2_tiehi _2467__500 (.L_HI(net543));
 sg13g2_tiehi _2468__501 (.L_HI(net544));
 sg13g2_tiehi _2469__502 (.L_HI(net545));
 sg13g2_tiehi _2470__503 (.L_HI(net546));
 sg13g2_tiehi _2471__504 (.L_HI(net547));
 sg13g2_tiehi _2472__505 (.L_HI(net548));
 sg13g2_tiehi _2473__506 (.L_HI(net549));
 sg13g2_tiehi _2474__507 (.L_HI(net550));
 sg13g2_tiehi _2475__508 (.L_HI(net551));
 sg13g2_tiehi _2476__509 (.L_HI(net552));
 sg13g2_tiehi _2477__510 (.L_HI(net553));
 sg13g2_tiehi _2478__511 (.L_HI(net554));
 sg13g2_tiehi _2479__512 (.L_HI(net555));
 sg13g2_tiehi _2480__513 (.L_HI(net556));
 sg13g2_tiehi _2481__514 (.L_HI(net557));
 sg13g2_tiehi _2482__515 (.L_HI(net558));
 sg13g2_tiehi _2483__516 (.L_HI(net559));
 sg13g2_tiehi _2484__517 (.L_HI(net560));
 sg13g2_tiehi _2485__518 (.L_HI(net561));
 sg13g2_tiehi _2486__519 (.L_HI(net562));
 sg13g2_tiehi _2487__520 (.L_HI(net563));
 sg13g2_tiehi _2488__521 (.L_HI(net564));
 sg13g2_tiehi _2489__522 (.L_HI(net565));
 sg13g2_tiehi _2490__523 (.L_HI(net566));
 sg13g2_tiehi _2491__524 (.L_HI(net567));
 sg13g2_tiehi _2492__525 (.L_HI(net568));
 sg13g2_tiehi _2493__526 (.L_HI(net569));
 sg13g2_tiehi _2494__527 (.L_HI(net570));
 sg13g2_tiehi _2495__528 (.L_HI(net571));
 sg13g2_tiehi _2496__529 (.L_HI(net572));
 sg13g2_tiehi _2497__530 (.L_HI(net573));
 sg13g2_tiehi _2498__531 (.L_HI(net574));
 sg13g2_tiehi _2499__532 (.L_HI(net575));
 sg13g2_tiehi _2500__533 (.L_HI(net576));
 sg13g2_tiehi _2501__534 (.L_HI(net577));
 sg13g2_tiehi _2502__535 (.L_HI(net578));
 sg13g2_tiehi _2503__536 (.L_HI(net579));
 sg13g2_tiehi _2504__537 (.L_HI(net580));
 sg13g2_tiehi _2505__538 (.L_HI(net581));
 sg13g2_tiehi _2506__539 (.L_HI(net582));
 sg13g2_tiehi _2507__540 (.L_HI(net583));
 sg13g2_tiehi _2508__541 (.L_HI(net584));
 sg13g2_tiehi _2509__542 (.L_HI(net585));
 sg13g2_tiehi _2510__543 (.L_HI(net586));
 sg13g2_tiehi _2511__544 (.L_HI(net587));
 sg13g2_tiehi _2512__545 (.L_HI(net588));
 sg13g2_tiehi _2513__546 (.L_HI(net589));
 sg13g2_tiehi _2514__547 (.L_HI(net590));
 sg13g2_tiehi _2515__548 (.L_HI(net591));
 sg13g2_tiehi _2516__549 (.L_HI(net592));
 sg13g2_tiehi _2517__550 (.L_HI(net593));
 sg13g2_tiehi _2518__551 (.L_HI(net594));
 sg13g2_tiehi _2519__552 (.L_HI(net595));
 sg13g2_tiehi _2520__553 (.L_HI(net596));
 sg13g2_tiehi _2521__554 (.L_HI(net597));
 sg13g2_tiehi _2522__555 (.L_HI(net598));
 sg13g2_tiehi _2523__556 (.L_HI(net599));
 sg13g2_tiehi _2524__557 (.L_HI(net600));
 sg13g2_tiehi _2525__558 (.L_HI(net601));
 sg13g2_tiehi _2526__559 (.L_HI(net602));
 sg13g2_tiehi _2527__560 (.L_HI(net603));
 sg13g2_tiehi _2528__561 (.L_HI(net604));
 sg13g2_tiehi _2529__562 (.L_HI(net605));
 sg13g2_tiehi _2530__563 (.L_HI(net606));
 sg13g2_tiehi _2531__564 (.L_HI(net607));
 sg13g2_tiehi _2532__565 (.L_HI(net608));
 sg13g2_tiehi _2533__566 (.L_HI(net609));
 sg13g2_tiehi _2534__567 (.L_HI(net610));
 sg13g2_tiehi _2535__568 (.L_HI(net611));
 sg13g2_tiehi _2536__569 (.L_HI(net612));
 sg13g2_tiehi _2537__570 (.L_HI(net613));
 sg13g2_tiehi _2538__571 (.L_HI(net614));
 sg13g2_tiehi _2539__572 (.L_HI(net615));
 sg13g2_tiehi _2540__573 (.L_HI(net616));
 sg13g2_tiehi _2541__574 (.L_HI(net617));
 sg13g2_tiehi _2542__575 (.L_HI(net618));
 sg13g2_tiehi _2543__576 (.L_HI(net619));
 sg13g2_tiehi _2544__577 (.L_HI(net620));
 sg13g2_tiehi _2545__578 (.L_HI(net621));
 sg13g2_tiehi _2546__579 (.L_HI(net622));
 sg13g2_tiehi _2547__580 (.L_HI(net623));
 sg13g2_tiehi _2548__581 (.L_HI(net624));
 sg13g2_tiehi _2549__582 (.L_HI(net625));
 sg13g2_tiehi _2550__583 (.L_HI(net626));
 sg13g2_tiehi _2551__584 (.L_HI(net627));
 sg13g2_tiehi _2552__585 (.L_HI(net628));
 sg13g2_tiehi _2553__586 (.L_HI(net629));
 sg13g2_tiehi _2554__587 (.L_HI(net630));
 sg13g2_tiehi _2555__588 (.L_HI(net631));
 sg13g2_tiehi _2556__589 (.L_HI(net632));
 sg13g2_tiehi _2557__590 (.L_HI(net633));
 sg13g2_tiehi _2558__591 (.L_HI(net634));
 sg13g2_tiehi _2559__592 (.L_HI(net635));
 sg13g2_tiehi _2560__593 (.L_HI(net636));
 sg13g2_tiehi _2561__594 (.L_HI(net637));
 sg13g2_tiehi _2562__595 (.L_HI(net638));
 sg13g2_tiehi _2563__596 (.L_HI(net639));
 sg13g2_tiehi _2564__597 (.L_HI(net640));
 sg13g2_tiehi _2565__598 (.L_HI(net641));
 sg13g2_tiehi _2566__599 (.L_HI(net642));
 sg13g2_tiehi _2567__600 (.L_HI(net643));
 sg13g2_tiehi _2568__601 (.L_HI(net644));
 sg13g2_tiehi _2569__602 (.L_HI(net645));
 sg13g2_tiehi _2064__603 (.L_HI(net646));
 sg13g2_tiehi _2100__604 (.L_HI(net647));
 sg13g2_tiehi _2063__605 (.L_HI(net648));
 sg13g2_tiehi _2099__606 (.L_HI(net649));
 sg13g2_tiehi _2062__607 (.L_HI(net650));
 sg13g2_tiehi _2098__608 (.L_HI(net651));
 sg13g2_tiehi _2061__609 (.L_HI(net652));
 sg13g2_tiehi _2060__610 (.L_HI(net653));
 sg13g2_tiehi _2059__611 (.L_HI(net654));
 sg13g2_tiehi _2058__612 (.L_HI(net655));
 sg13g2_tiehi _2570__613 (.L_HI(net656));
 sg13g2_tiehi _2057__614 (.L_HI(net657));
 sg13g2_tiehi _2056__615 (.L_HI(net658));
 sg13g2_tiehi _2055__616 (.L_HI(net659));
 sg13g2_tiehi _2097__617 (.L_HI(net660));
 sg13g2_tiehi tt_um_snake_game_618 (.L_HI(net661));
 sg13g2_tiehi tt_um_snake_game_619 (.L_HI(net662));
 sg13g2_tiehi tt_um_snake_game_620 (.L_HI(net663));
 sg13g2_tiehi tt_um_snake_game_621 (.L_HI(net664));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_snake_game_8 (.L_LO(net8));
 sg13g2_tielo tt_um_snake_game_9 (.L_LO(net9));
 sg13g2_tielo tt_um_snake_game_10 (.L_LO(net10));
 sg13g2_tielo tt_um_snake_game_11 (.L_LO(net11));
 sg13g2_tielo tt_um_snake_game_12 (.L_LO(net12));
 sg13g2_tielo tt_um_snake_game_13 (.L_LO(net13));
 sg13g2_tielo tt_um_snake_game_14 (.L_LO(net14));
 sg13g2_tiehi _2054__15 (.L_HI(net15));
 sg13g2_buf_1 _3202_ (.A(failure),
    .X(uio_out[0]));
 sg13g2_buf_1 _3203_ (.A(\game_inst.o_success ),
    .X(uio_out[1]));
 sg13g2_buf_1 _3204_ (.A(eat),
    .X(uio_out[2]));
 sg13g2_buf_1 _3205_ (.A(\game_inst.o_tick ),
    .X(uio_out[3]));
 sg13g2_buf_1 _3206_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _3207_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _3208_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _3209_ (.A(\game_inst.o_vga_vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _3210_ (.A(\game_inst.o_vga_hsync ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(_0507_),
    .X(net95));
 sg13g2_buf_8 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(_0481_),
    .X(net98));
 sg13g2_buf_8 fanout99 (.A(_0402_),
    .X(net99));
 sg13g2_buf_8 fanout100 (.A(_0400_),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(_0400_),
    .X(net101));
 sg13g2_buf_8 fanout102 (.A(net104),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_8 fanout104 (.A(_0395_),
    .X(net104));
 sg13g2_buf_8 fanout105 (.A(net107),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_8 fanout107 (.A(net110),
    .X(net107));
 sg13g2_buf_8 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_8 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_8 fanout110 (.A(_0221_),
    .X(net110));
 sg13g2_buf_8 fanout111 (.A(_0220_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0220_),
    .X(net112));
 sg13g2_buf_8 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_8 fanout114 (.A(_0389_),
    .X(net114));
 sg13g2_buf_8 fanout115 (.A(_0389_),
    .X(net115));
 sg13g2_buf_8 fanout116 (.A(net1331),
    .X(net116));
 sg13g2_buf_8 fanout117 (.A(\game_inst.apple_inst.i_snake_x[1] ),
    .X(net117));
 sg13g2_buf_8 fanout118 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(net1202),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(net1257),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net1199),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(net1171),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(\game_inst.pos_dir[1] ),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(net1329),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net1336),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net1332),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(\game_inst.vga_inst.px[7] ),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(\game_inst.vga_inst.px[6] ),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net1238),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0390_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0390_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0156_),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(_0156_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(rst_n),
    .X(net136));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_tielo tt_um_snake_game_7 (.L_LO(net7));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_76_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_9_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_28_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\game_inst.snake_inst.shiftreg_inst.memory[39][0] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold2 (.A(\game_inst.snake_inst.shiftreg_inst.memory[51][0] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold3 (.A(\game_inst.snake_inst.shiftreg_inst.memory[71][0] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold4 (.A(\game_inst.snake_inst.shiftreg_inst.memory[167][1] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold5 (.A(\game_inst.snake_inst.shiftreg_inst.memory[60][0] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold6 (.A(\game_inst.snake_inst.shiftreg_inst.memory[136][0] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold7 (.A(\game_inst.snake_inst.shiftreg_inst.memory[138][0] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold8 (.A(\game_inst.snake_inst.shiftreg_inst.memory[193][0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold9 (.A(\game_inst.snake_inst.shiftreg_inst.memory[147][0] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold10 (.A(\game_inst.snake_inst.shiftreg_inst.memory[177][0] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold11 (.A(\game_inst.snake_inst.shiftreg_inst.memory[166][0] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold12 (.A(\game_inst.snake_inst.shiftreg_inst.memory[102][0] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold13 (.A(\game_inst.snake_inst.shiftreg_inst.memory[82][0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold14 (.A(\game_inst.snake_inst.shiftreg_inst.memory[77][0] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold15 (.A(\game_inst.snake_inst.shiftreg_inst.memory[16][0] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold16 (.A(\game_inst.snake_inst.shiftreg_inst.memory[47][1] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold17 (.A(\game_inst.snake_inst.shiftreg_inst.memory[97][1] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold18 (.A(\game_inst.snake_inst.shiftreg_inst.memory[33][0] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold19 (.A(\game_inst.snake_inst.shiftreg_inst.memory[173][1] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold20 (.A(\game_inst.snake_inst.shiftreg_inst.memory[48][1] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold21 (.A(\game_inst.snake_inst.shiftreg_inst.memory[175][1] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game_inst.snake_inst.shiftreg_inst.memory[73][0] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold23 (.A(\game_inst.snake_inst.shiftreg_inst.memory[200][0] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold24 (.A(\game_inst.snake_inst.shiftreg_inst.memory[162][0] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold25 (.A(\game_inst.snake_inst.shiftreg_inst.memory[179][1] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold26 (.A(\game_inst.snake_inst.shiftreg_inst.memory[66][1] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold27 (.A(\game_inst.snake_inst.shiftreg_inst.memory[94][1] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold28 (.A(\game_inst.snake_inst.shiftreg_inst.memory[174][0] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold29 (.A(\game_inst.snake_inst.shiftreg_inst.memory[192][1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold30 (.A(\game_inst.snake_inst.shiftreg_inst.memory[185][0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold31 (.A(\game_inst.snake_inst.shiftreg_inst.memory[30][1] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold32 (.A(\game_inst.snake_inst.shiftreg_inst.memory[191][1] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold33 (.A(\game_inst.snake_inst.shiftreg_inst.memory[73][1] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold34 (.A(\game_inst.snake_inst.shiftreg_inst.memory[176][1] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold35 (.A(\game_inst.snake_inst.shiftreg_inst.memory[108][1] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold36 (.A(\game_inst.snake_inst.shiftreg_inst.memory[64][1] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold37 (.A(\game_inst.snake_inst.shiftreg_inst.memory[24][0] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold38 (.A(\game_inst.snake_inst.shiftreg_inst.memory[207][0] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold39 (.A(\game_inst.snake_inst.shiftreg_inst.memory[229][1] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game_inst.snake_inst.shiftreg_inst.memory[100][1] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold41 (.A(\game_inst.snake_inst.shiftreg_inst.memory[218][1] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold42 (.A(\game_inst.snake_inst.shiftreg_inst.memory[65][1] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold43 (.A(\game_inst.snake_inst.shiftreg_inst.memory[60][1] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold44 (.A(\game_inst.snake_inst.shiftreg_inst.memory[25][0] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold45 (.A(\game_inst.snake_inst.shiftreg_inst.memory[116][0] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold46 (.A(\game_inst.snake_inst.shiftreg_inst.memory[96][1] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game_inst.snake_inst.shiftreg_inst.memory[100][0] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold48 (.A(\game_inst.snake_inst.shiftreg_inst.memory[69][1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold49 (.A(\game_inst.snake_inst.shiftreg_inst.memory[23][0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold50 (.A(\game_inst.snake_inst.shiftreg_inst.memory[70][0] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold51 (.A(\game_inst.snake_inst.shiftreg_inst.memory[232][1] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold52 (.A(\game_inst.snake_inst.shiftreg_inst.memory[92][1] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold53 (.A(\game_inst.snake_inst.shiftreg_inst.memory[39][1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold54 (.A(\game_inst.vga_inst.s_hsync ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold55 (.A(\game_inst.snake_inst.shiftreg_inst.memory[169][1] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold56 (.A(\game_inst.snake_inst.shiftreg_inst.memory[127][0] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold57 (.A(\game_inst.snake_inst.shiftreg_inst.memory[78][0] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold58 (.A(\game_inst.snake_inst.shiftreg_inst.memory[207][1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold59 (.A(\game_inst.snake_inst.shiftreg_inst.memory[217][0] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold60 (.A(\game_inst.snake_inst.shiftreg_inst.memory[169][0] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game_inst.snake_inst.shiftreg_inst.memory[15][0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold62 (.A(\game_inst.snake_inst.shiftreg_inst.memory[20][0] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold63 (.A(\game_inst.snake_inst.shiftreg_inst.memory[191][0] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold64 (.A(\game_inst.snake_inst.shiftreg_inst.memory[157][1] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold65 (.A(\game_inst.snake_inst.shiftreg_inst.memory[4][0] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold66 (.A(\game_inst.snake_inst.shiftreg_inst.memory[129][1] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold67 (.A(\game_inst.snake_inst.shiftreg_inst.memory[108][0] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game_inst.snake_inst.shiftreg_inst.memory[154][1] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold69 (.A(\game_inst.snake_inst.shiftreg_inst.memory[153][0] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold70 (.A(\game_inst.snake_inst.shiftreg_inst.memory[74][0] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold71 (.A(\game_inst.snake_inst.shiftreg_inst.memory[6][1] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold72 (.A(\game_inst.snake_inst.shiftreg_inst.memory[77][1] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold73 (.A(\game_inst.snake_inst.shiftreg_inst.memory[87][0] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold74 (.A(\game_inst.snake_inst.shiftreg_inst.memory[31][0] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold75 (.A(\game_inst.snake_inst.shiftreg_inst.memory[117][0] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold76 (.A(\game_inst.snake_inst.shiftreg_inst.memory[120][0] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold77 (.A(\game_inst.snake_inst.shiftreg_inst.memory[28][1] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold78 (.A(\game_inst.snake_inst.shiftreg_inst.memory[110][1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold79 (.A(\game_inst.snake_inst.shiftreg_inst.memory[82][1] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold80 (.A(\game_inst.snake_inst.shiftreg_inst.memory[109][0] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold81 (.A(\game_inst.snake_inst.shiftreg_inst.memory[183][0] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold82 (.A(\game_inst.snake_inst.shiftreg_inst.memory[147][1] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold83 (.A(\game_inst.snake_inst.shiftreg_inst.memory[165][1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game_inst.snake_inst.shiftreg_inst.memory[123][0] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold85 (.A(\game_inst.snake_inst.shiftreg_inst.memory[219][1] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold86 (.A(\game_inst.snake_inst.shiftreg_inst.memory[11][1] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold87 (.A(\game_inst.snake_inst.shiftreg_inst.memory[46][0] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold88 (.A(\game_inst.snake_inst.shiftreg_inst.memory[42][1] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold89 (.A(\game_inst.snake_inst.shiftreg_inst.memory[206][0] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold90 (.A(\game_inst.snake_inst.shiftreg_inst.memory[83][0] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold91 (.A(\game_inst.snake_inst.shiftreg_inst.memory[130][1] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold92 (.A(\game_inst.snake_inst.shiftreg_inst.memory[208][0] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold93 (.A(\game_inst.snake_inst.shiftreg_inst.memory[99][0] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold94 (.A(\game_inst.snake_inst.shiftreg_inst.memory[127][1] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold95 (.A(\game_inst.snake_inst.shiftreg_inst.memory[223][0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold96 (.A(\game_inst.snake_inst.shiftreg_inst.memory[13][0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold97 (.A(\game_inst.snake_inst.shiftreg_inst.memory[1][0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold98 (.A(\game_inst.snake_inst.shiftreg_inst.memory[227][0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold99 (.A(\game_inst.snake_inst.shiftreg_inst.memory[132][1] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold100 (.A(\game_inst.snake_inst.shiftreg_inst.memory[211][0] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game_inst.snake_inst.shiftreg_inst.memory[37][0] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold102 (.A(\game_inst.snake_inst.shiftreg_inst.memory[103][0] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold103 (.A(\game_inst.snake_inst.shiftreg_inst.memory[187][0] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold104 (.A(\game_inst.snake_inst.shiftreg_inst.memory[12][1] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold105 (.A(\game_inst.snake_inst.shiftreg_inst.memory[187][1] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold106 (.A(\game_inst.snake_inst.shiftreg_inst.memory[128][1] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold107 (.A(\game_inst.snake_inst.shiftreg_inst.memory[101][1] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold108 (.A(\game_inst.snake_inst.shiftreg_inst.memory[122][0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold109 (.A(\game_inst.snake_inst.shiftreg_inst.memory[18][0] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold110 (.A(\game_inst.snake_inst.shiftreg_inst.memory[107][1] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold111 (.A(\game_inst.snake_inst.shiftreg_inst.memory[204][0] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold112 (.A(\game_inst.snake_inst.shiftreg_inst.memory[145][0] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold113 (.A(\game_inst.snake_inst.shiftreg_inst.memory[226][0] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold114 (.A(\game_inst.snake_inst.shiftreg_inst.memory[178][0] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold115 (.A(\game_inst.snake_inst.shiftreg_inst.memory[41][1] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold116 (.A(\game_inst.snake_inst.shiftreg_inst.memory[80][1] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold117 (.A(\game_inst.snake_inst.shiftreg_inst.memory[212][1] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold118 (.A(\game_inst.snake_inst.shiftreg_inst.memory[2][0] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold119 (.A(\game_inst.snake_inst.shiftreg_inst.memory[89][0] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold120 (.A(\game_inst.snake_inst.shiftreg_inst.memory[213][0] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold121 (.A(\game_inst.snake_inst.shiftreg_inst.memory[67][0] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold122 (.A(\game_inst.snake_inst.shiftreg_inst.memory[126][1] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold123 (.A(\game_inst.snake_inst.shiftreg_inst.memory[43][0] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold124 (.A(\game_inst.snake_inst.shiftreg_inst.memory[59][0] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold125 (.A(\game_inst.snake_inst.shiftreg_inst.memory[56][1] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold126 (.A(\game_inst.snake_inst.shiftreg_inst.memory[81][1] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold127 (.A(\game_inst.snake_inst.shiftreg_inst.memory[2][1] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold128 (.A(\game_inst.snake_inst.shiftreg_inst.memory[139][0] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold129 (.A(\game_inst.snake_inst.shiftreg_inst.memory[113][1] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold130 (.A(\game_inst.snake_inst.shiftreg_inst.memory[148][1] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold131 (.A(\game_inst.snake_inst.shiftreg_inst.memory[3][0] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game_inst.snake_inst.shiftreg_inst.memory[102][1] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold133 (.A(\game_inst.snake_inst.shiftreg_inst.memory[132][0] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold134 (.A(\game_inst.snake_inst.shiftreg_inst.memory[76][0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold135 (.A(\game_inst.snake_inst.shiftreg_inst.memory[182][0] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold136 (.A(\game_inst.snake_inst.shiftreg_inst.memory[210][0] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold137 (.A(\game_inst.snake_inst.shiftreg_inst.memory[40][0] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold138 (.A(\game_inst.snake_inst.shiftreg_inst.memory[78][1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold139 (.A(\game_inst.snake_inst.shiftreg_inst.memory[220][0] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold140 (.A(\game_inst.snake_inst.shiftreg_inst.memory[43][1] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold141 (.A(\game_inst.snake_inst.shiftreg_inst.memory[112][1] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold142 (.A(\game_inst.snake_inst.shiftreg_inst.memory[149][1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold143 (.A(\game_inst.snake_inst.shiftreg_inst.memory[10][0] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold144 (.A(\game_inst.snake_inst.shiftreg_inst.memory[93][0] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold145 (.A(\game_inst.snake_inst.shiftreg_inst.memory[201][1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold146 (.A(\game_inst.snake_inst.shiftreg_inst.memory[149][0] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold147 (.A(\game_inst.snake_inst.shiftreg_inst.memory[57][0] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold148 (.A(\game_inst.snake_inst.shiftreg_inst.memory[158][0] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold149 (.A(\game_inst.snake_inst.shiftreg_inst.memory[136][1] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold150 (.A(\game_inst.snake_inst.shiftreg_inst.memory[56][0] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold151 (.A(\game_inst.snake_inst.shiftreg_inst.memory[134][1] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold152 (.A(\game_inst.snake_inst.shiftreg_inst.memory[157][0] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold153 (.A(\game_inst.snake_inst.shiftreg_inst.memory[106][1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold154 (.A(\game_inst.snake_inst.shiftreg_inst.memory[229][0] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold155 (.A(\game_inst.snake_inst.shiftreg_inst.memory[156][1] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold156 (.A(\game_inst.snake_inst.shiftreg_inst.memory[55][1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold157 (.A(\game_inst.snake_inst.shiftreg_inst.memory[141][1] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold158 (.A(\game_inst.snake_inst.shiftreg_inst.memory[51][1] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold159 (.A(\game_inst.snake_inst.shiftreg_inst.memory[11][0] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold160 (.A(\game_inst.snake_inst.shiftreg_inst.memory[190][1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold161 (.A(\game_inst.snake_inst.shiftreg_inst.memory[74][1] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game_inst.snake_inst.shiftreg_inst.memory[98][1] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold163 (.A(\game_inst.snake_inst.shiftreg_inst.memory[40][1] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold164 (.A(\game_inst.snake_inst.shiftreg_inst.memory[161][1] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold165 (.A(\game_inst.snake_inst.shiftreg_inst.memory[91][0] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold166 (.A(\game_inst.snake_inst.shiftreg_inst.memory[134][0] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold167 (.A(\game_inst.snake_inst.shiftreg_inst.memory[20][1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold168 (.A(\game_inst.snake_inst.shiftreg_inst.memory[194][0] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold169 (.A(\game_inst.snake_inst.shiftreg_inst.memory[27][0] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold170 (.A(\game_inst.snake_inst.shiftreg_inst.memory[188][1] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold171 (.A(\game_inst.snake_inst.shiftreg_inst.memory[158][1] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold172 (.A(\game_inst.snake_inst.shiftreg_inst.memory[88][0] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold173 (.A(\game_inst.snake_inst.shiftreg_inst.memory[197][0] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold174 (.A(\game_inst.snake_inst.shiftreg_inst.memory[44][0] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold175 (.A(\game_inst.snake_inst.shiftreg_inst.memory[8][1] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold176 (.A(\game_inst.snake_inst.shiftreg_inst.memory[71][1] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold177 (.A(\game_inst.snake_inst.shiftreg_inst.memory[33][1] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold178 (.A(\game_inst.snake_inst.shiftreg_inst.memory[19][1] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold179 (.A(\game_inst.snake_inst.shiftreg_inst.memory[16][1] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold180 (.A(\game_inst.snake_inst.shiftreg_inst.memory[26][0] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold181 (.A(\game_inst.snake_inst.shiftreg_inst.memory[114][1] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold182 (.A(\game_inst.snake_inst.shiftreg_inst.memory[114][0] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold183 (.A(\game_inst.snake_inst.shiftreg_inst.memory[47][0] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold184 (.A(\game_inst.snake_inst.shiftreg_inst.memory[209][0] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold185 (.A(\game_inst.snake_inst.shiftreg_inst.memory[92][0] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold186 (.A(\game_inst.snake_inst.shiftreg_inst.memory[41][0] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold187 (.A(\game_inst.snake_inst.shiftreg_inst.memory[113][0] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold188 (.A(\game_inst.snake_inst.shiftreg_inst.memory[167][0] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold189 (.A(\game_inst.snake_inst.shiftreg_inst.memory[26][1] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold190 (.A(\game_inst.snake_inst.shiftreg_inst.memory[125][0] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold191 (.A(\game_inst.snake_inst.shiftreg_inst.memory[146][1] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold192 (.A(\game_inst.snake_inst.shiftreg_inst.memory[29][1] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold193 (.A(\game_inst.snake_inst.shiftreg_inst.memory[22][0] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold194 (.A(\game_inst.snake_inst.shiftreg_inst.memory[124][1] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold195 (.A(\game_inst.snake_inst.shiftreg_inst.memory[150][1] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold196 (.A(\game_inst.snake_inst.shiftreg_inst.memory[219][0] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold197 (.A(\game_inst.snake_inst.shiftreg_inst.memory[46][1] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold198 (.A(\game_inst.snake_inst.shiftreg_inst.memory[44][1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold199 (.A(\game_inst.snake_inst.shiftreg_inst.memory[156][0] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold200 (.A(\game_inst.snake_inst.shiftreg_inst.memory[170][1] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold201 (.A(\game_inst.snake_inst.shiftreg_inst.memory[133][1] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold202 (.A(\game_inst.snake_inst.shiftreg_inst.memory[131][0] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold203 (.A(\game_inst.snake_inst.shiftreg_inst.memory[202][1] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold204 (.A(\game_inst.snake_inst.shiftreg_inst.memory[198][0] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold205 (.A(\game_inst.snake_inst.shiftreg_inst.memory[144][1] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold206 (.A(\game_inst.snake_inst.shiftreg_inst.memory[10][1] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold207 (.A(\game_inst.snake_inst.shiftreg_inst.memory[224][0] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold208 (.A(\game_inst.snake_inst.shiftreg_inst.memory[183][1] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold209 (.A(\game_inst.snake_inst.shiftreg_inst.memory[5][1] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold210 (.A(\game_inst.snake_inst.shiftreg_inst.memory[137][0] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold211 (.A(\game_inst.snake_inst.shiftreg_inst.memory[206][1] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold212 (.A(\game_inst.snake_inst.shiftreg_inst.memory[52][1] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold213 (.A(\game_inst.snake_inst.shiftreg_inst.memory[62][0] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold214 (.A(\game_inst.snake_inst.shiftreg_inst.memory[50][1] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold215 (.A(\game_inst.snake_inst.shiftreg_inst.memory[231][1] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold216 (.A(\game_inst.snake_inst.shiftreg_inst.memory[196][1] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold217 (.A(\game_inst.snake_inst.shiftreg_inst.memory[231][0] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold218 (.A(\game_inst.snake_inst.shiftreg_inst.memory[9][0] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold219 (.A(\game_inst.snake_inst.shiftreg_inst.memory[45][1] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold220 (.A(\game_inst.snake_inst.shiftreg_inst.memory[25][1] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold221 (.A(\game_inst.snake_inst.shiftreg_inst.memory[122][1] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold222 (.A(\game_inst.snake_inst.shiftreg_inst.memory[151][1] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold223 (.A(\game_inst.snake_inst.shiftreg_inst.memory[101][0] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold224 (.A(\game_inst.snake_inst.shiftreg_inst.memory[98][0] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold225 (.A(\game_inst.snake_inst.shiftreg_inst.memory[69][0] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold226 (.A(\game_inst.snake_inst.shiftreg_inst.memory[225][1] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold227 (.A(\game_inst.snake_inst.shiftreg_inst.memory[199][0] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold228 (.A(\game_inst.snake_inst.shiftreg_inst.memory[90][1] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold229 (.A(\game_inst.snake_inst.shiftreg_inst.memory[32][1] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold230 (.A(\game_inst.snake_inst.shiftreg_inst.memory[221][0] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold231 (.A(\game_inst.snake_inst.shiftreg_inst.memory[216][1] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold232 (.A(\game_inst.snake_inst.shiftreg_inst.memory[171][1] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold233 (.A(\game_inst.snake_inst.shiftreg_inst.memory[91][1] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold234 (.A(\game_inst.snake_inst.shiftreg_inst.memory[186][1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold235 (.A(\game_inst.snake_inst.shiftreg_inst.memory[159][0] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold236 (.A(\game_inst.snake_inst.shiftreg_inst.memory[155][1] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold237 (.A(\game_inst.snake_inst.shiftreg_inst.memory[63][1] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold238 (.A(\game_inst.snake_inst.shiftreg_inst.memory[4][1] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold239 (.A(\game_inst.snake_inst.shiftreg_inst.memory[130][0] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold240 (.A(\game_inst.snake_inst.shiftreg_inst.memory[14][0] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold241 (.A(\game_inst.snake_inst.shiftreg_inst.memory[163][1] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold242 (.A(\game_inst.snake_inst.shiftreg_inst.memory[111][0] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold243 (.A(\game_inst.snake_inst.shiftreg_inst.memory[128][0] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold244 (.A(\game_inst.snake_inst.shiftreg_inst.memory[228][0] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold245 (.A(\game_inst.snake_inst.shiftreg_inst.memory[125][1] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold246 (.A(\game_inst.snake_inst.shiftreg_inst.memory[3][1] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold247 (.A(\game_inst.snake_inst.shiftreg_inst.memory[124][0] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold248 (.A(\game_inst.snake_inst.shiftreg_inst.memory[153][1] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold249 (.A(\game_inst.snake_inst.shiftreg_inst.memory[53][1] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold250 (.A(\game_inst.snake_inst.shiftreg_inst.memory[209][1] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold251 (.A(\game_inst.snake_inst.shiftreg_inst.memory[76][1] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold252 (.A(\game_inst.snake_inst.shiftreg_inst.memory[123][1] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold253 (.A(\game_inst.snake_inst.shiftreg_inst.memory[105][0] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold254 (.A(\game_inst.snake_inst.shiftreg_inst.memory[174][1] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold255 (.A(\game_inst.snake_inst.shiftreg_inst.memory[111][1] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold256 (.A(\game_inst.snake_inst.shiftreg_inst.memory[210][1] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold257 (.A(\game_inst.snake_inst.shiftreg_inst.memory[58][0] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold258 (.A(\game_inst.snake_inst.shiftreg_inst.memory[135][1] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold259 (.A(\game_inst.snake_inst.shiftreg_inst.memory[75][1] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold260 (.A(\game_inst.snake_inst.shiftreg_inst.memory[18][1] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold261 (.A(\game_inst.snake_inst.shiftreg_inst.memory[96][0] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold262 (.A(\game_inst.snake_inst.shiftreg_inst.memory[37][1] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold263 (.A(\game_inst.snake_inst.shiftreg_inst.memory[15][1] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold264 (.A(\game_inst.snake_inst.shiftreg_inst.memory[105][1] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold265 (.A(\game_inst.snake_inst.shiftreg_inst.memory[203][1] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold266 (.A(\game_inst.snake_inst.shiftreg_inst.memory[49][0] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold267 (.A(\game_inst.snake_inst.shiftreg_inst.memory[150][0] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold268 (.A(\game_inst.snake_inst.shiftreg_inst.memory[164][1] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold269 (.A(\game_inst.snake_inst.shiftreg_inst.memory[131][1] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold270 (.A(\game_inst.snake_inst.shiftreg_inst.memory[215][0] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold271 (.A(\game_inst.snake_inst.shiftreg_inst.memory[204][1] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold272 (.A(\game_inst.snake_inst.shiftreg_inst.memory[104][1] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold273 (.A(\game_inst.snake_inst.shiftreg_inst.memory[146][0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold274 (.A(\game_inst.snake_inst.shiftreg_inst.memory[88][1] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold275 (.A(\game_inst.snake_inst.shiftreg_inst.memory[45][0] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold276 (.A(\game_inst.snake_inst.shiftreg_inst.memory[214][0] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold277 (.A(\game_inst.snake_inst.shiftreg_inst.memory[181][1] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold278 (.A(\game_inst.snake_inst.shiftreg_inst.memory[49][1] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold279 (.A(\game_inst.snake_inst.shiftreg_inst.memory[53][0] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold280 (.A(\game_inst.snake_inst.shiftreg_inst.memory[142][0] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold281 (.A(\game_inst.snake_inst.shiftreg_inst.memory[225][0] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold282 (.A(\game_inst.snake_inst.shiftreg_inst.memory[5][0] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold283 (.A(\game_inst.snake_inst.shiftreg_inst.memory[189][1] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold284 (.A(\game_inst.snake_inst.shiftreg_inst.memory[104][0] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold285 (.A(\game_inst.snake_inst.shiftreg_inst.memory[152][0] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold286 (.A(\game_inst.snake_inst.shiftreg_inst.memory[181][0] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold287 (.A(\game_inst.snake_inst.shiftreg_inst.memory[195][0] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold288 (.A(\game_inst.snake_inst.shiftreg_inst.memory[61][0] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold289 (.A(\game_inst.snake_inst.shiftreg_inst.memory[205][1] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold290 (.A(\game_inst.snake_inst.shiftreg_inst.memory[137][1] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold291 (.A(\game_inst.snake_inst.shiftreg_inst.memory[117][1] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold292 (.A(\game_inst.snake_inst.shiftreg_inst.memory[145][1] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold293 (.A(\game_inst.snake_inst.shiftreg_inst.memory[129][0] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold294 (.A(\game_inst.snake_inst.shiftreg_inst.memory[232][0] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold295 (.A(\game_inst.snake_inst.shiftreg_inst.memory[36][0] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold296 (.A(\game_inst.snake_inst.shiftreg_inst.memory[162][1] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold297 (.A(\game_inst.snake_inst.shiftreg_inst.memory[168][0] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold298 (.A(\game_inst.snake_inst.shiftreg_inst.memory[138][1] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold299 (.A(\game_inst.snake_inst.shiftreg_inst.memory[36][1] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold300 (.A(\game_inst.snake_inst.shiftreg_inst.memory[34][1] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold301 (.A(\game_inst.snake_inst.shiftreg_inst.memory[211][1] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold302 (.A(\game_inst.snake_inst.shiftreg_inst.memory[13][1] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold303 (.A(\game_inst.snake_inst.shiftreg_inst.memory[163][0] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold304 (.A(\game_inst.snake_inst.shiftreg_inst.memory[188][0] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold305 (.A(\game_inst.snake_inst.shiftreg_inst.memory[94][0] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold306 (.A(\game_inst.snake_inst.shiftreg_inst.memory[161][0] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold307 (.A(\game_inst.snake_inst.shiftreg_inst.memory[172][0] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold308 (.A(\game_inst.snake_inst.shiftreg_inst.memory[217][1] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold309 (.A(\game_inst.snake_inst.shiftreg_inst.memory[230][1] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold310 (.A(\game_inst.snake_inst.shiftreg_inst.memory[154][0] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold311 (.A(\game_inst.snake_inst.shiftreg_inst.memory[185][1] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold312 (.A(\game_inst.snake_inst.shiftreg_inst.memory[133][0] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold313 (.A(\game_inst.snake_inst.shiftreg_inst.memory[218][0] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold314 (.A(\game_inst.snake_inst.shiftreg_inst.memory[6][0] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold315 (.A(\game_inst.snake_inst.shiftreg_inst.memory[144][0] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold316 (.A(\game_inst.snake_inst.shiftreg_inst.memory[192][0] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold317 (.A(\game_inst.snake_inst.shiftreg_inst.memory[9][1] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold318 (.A(\game_inst.snake_inst.shiftreg_inst.memory[214][1] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold319 (.A(\game_inst.snake_inst.shiftreg_inst.memory[221][1] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold320 (.A(\game_inst.snake_inst.shiftreg_inst.memory[99][1] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold321 (.A(\game_inst.snake_inst.shiftreg_inst.memory[190][0] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold322 (.A(\game_inst.snake_inst.shiftreg_inst.memory[109][1] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold323 (.A(\game_inst.snake_inst.shiftreg_inst.memory[119][0] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold324 (.A(\game_inst.snake_inst.shiftreg_inst.memory[140][1] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold325 (.A(\game_inst.snake_inst.shiftreg_inst.memory[79][0] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold326 (.A(\game_inst.snake_inst.shiftreg_inst.memory[118][0] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold327 (.A(\game_inst.snake_inst.shiftreg_inst.memory[103][1] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold328 (.A(\game_inst.snake_inst.shiftreg_inst.memory[7][0] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold329 (.A(\game_inst.snake_inst.shiftreg_inst.memory[195][1] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold330 (.A(\game_inst.snake_inst.shiftreg_inst.memory[24][1] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold331 (.A(\game_inst.snake_inst.shiftreg_inst.memory[202][0] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold332 (.A(\game_inst.snake_inst.shiftreg_inst.memory[86][0] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold333 (.A(\game_inst.snake_inst.shiftreg_inst.memory[173][0] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold334 (.A(\game_inst.snake_inst.shiftreg_inst.memory[168][1] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold335 (.A(\game_inst.snake_inst.shiftreg_inst.memory[86][1] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold336 (.A(\game_inst.snake_inst.shiftreg_inst.memory[31][1] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold337 (.A(\game_inst.snake_inst.shiftreg_inst.memory[93][1] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold338 (.A(\game_inst.snake_inst.shiftreg_inst.memory[83][1] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold339 (.A(\game_inst.snake_inst.shiftreg_inst.memory[95][0] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold340 (.A(\game_inst.snake_inst.shiftreg_inst.memory[179][0] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold341 (.A(\game_inst.snake_inst.shiftreg_inst.memory[95][1] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold342 (.A(\game_inst.snake_inst.shiftreg_inst.memory[42][0] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold343 (.A(\game_inst.snake_inst.shiftreg_inst.memory[21][0] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold344 (.A(\game_inst.snake_inst.shiftreg_inst.memory[115][1] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold345 (.A(\game_inst.snake_inst.shiftreg_inst.memory[68][1] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold346 (.A(\game_inst.snake_inst.shiftreg_inst.memory[121][1] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold347 (.A(\game_inst.snake_inst.shiftreg_inst.memory[228][1] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold348 (.A(\game_inst.snake_inst.shiftreg_inst.memory[87][1] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold349 (.A(\game_inst.snake_inst.shiftreg_inst.memory[180][0] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold350 (.A(\game_inst.snake_inst.shiftreg_inst.memory[12][0] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold351 (.A(\game_inst.snake_inst.shiftreg_inst.memory[84][1] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold352 (.A(\game_inst.snake_inst.shiftreg_inst.memory[215][1] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold353 (.A(\game_inst.snake_inst.shiftreg_inst.memory[151][0] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold354 (.A(\game_inst.snake_inst.shiftreg_inst.memory[152][1] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold355 (.A(\game_inst.snake_inst.shiftreg_inst.memory[65][0] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold356 (.A(\game_inst.snake_inst.shiftreg_inst.memory[75][0] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold357 (.A(\game_inst.snake_inst.shiftreg_inst.memory[32][0] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold358 (.A(\game_inst.snake_inst.shiftreg_inst.memory[55][0] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold359 (.A(\game_inst.snake_inst.shiftreg_inst.memory[184][0] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold360 (.A(\game_inst.snake_inst.shiftreg_inst.memory[58][1] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold361 (.A(\game_inst.snake_inst.shiftreg_inst.memory[19][0] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold362 (.A(\game_inst.snake_inst.shiftreg_inst.memory[121][0] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold363 (.A(\game_inst.snake_inst.shiftreg_inst.memory[72][1] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold364 (.A(\game_inst.snake_inst.shiftreg_inst.memory[197][1] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold365 (.A(\game_inst.snake_inst.shiftreg_inst.memory[84][0] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold366 (.A(\game_inst.snake_inst.shiftreg_inst.memory[112][0] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold367 (.A(\game_inst.snake_inst.shiftreg_inst.memory[59][1] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold368 (.A(\game_inst.snake_inst.shiftreg_inst.memory[140][0] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold369 (.A(\game_inst.snake_inst.shiftreg_inst.memory[216][0] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold370 (.A(\game_inst.snake_inst.shiftreg_inst.memory[68][0] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold371 (.A(\game_inst.snake_inst.shiftreg_inst.memory[222][1] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold372 (.A(\game_inst.snake_inst.shiftreg_inst.memory[223][1] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold373 (.A(\game_inst.snake_inst.shiftreg_inst.memory[107][0] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold374 (.A(\game_inst.snake_inst.shiftreg_inst.memory[166][1] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold375 (.A(\game_inst.snake_inst.shiftreg_inst.memory[79][1] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold376 (.A(\game_inst.snake_inst.shiftreg_inst.memory[17][1] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold377 (.A(\game_inst.snake_inst.shiftreg_inst.memory[182][1] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold378 (.A(\game_inst.snake_inst.shiftreg_inst.memory[160][0] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold379 (.A(\game_inst.snake_inst.shiftreg_inst.memory[67][1] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold380 (.A(\game_inst.snake_inst.shiftreg_inst.memory[186][0] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold381 (.A(\game_inst.snake_inst.shiftreg_inst.memory[126][0] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold382 (.A(\game_inst.snake_inst.shiftreg_inst.memory[28][0] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold383 (.A(\game_inst.snake_inst.shiftreg_inst.memory[178][1] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold384 (.A(\game_inst.snake_inst.shiftreg_inst.memory[7][1] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold385 (.A(\game_inst.snake_inst.shiftreg_inst.memory[50][0] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold386 (.A(\game_inst.snake_inst.shiftreg_inst.memory[196][0] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold387 (.A(\game_inst.snake_inst.shiftreg_inst.memory[85][0] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold388 (.A(\game_inst.snake_inst.shiftreg_inst.memory[106][0] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold389 (.A(\game_inst.snake_inst.shiftreg_inst.memory[142][1] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold390 (.A(\game_inst.snake_inst.shiftreg_inst.memory[30][0] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold391 (.A(\game_inst.snake_inst.shiftreg_inst.memory[171][0] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold392 (.A(\game_inst.snake_inst.shiftreg_inst.memory[155][0] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold393 (.A(\game_inst.snake_inst.shiftreg_inst.memory[34][0] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold394 (.A(\game_inst.snake_inst.shiftreg_inst.memory[72][0] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold395 (.A(\game_inst.snake_inst.shiftreg_inst.memory[64][0] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold396 (.A(\game_inst.snake_inst.shiftreg_inst.memory[81][0] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold397 (.A(\game_inst.snake_inst.shiftreg_inst.memory[90][0] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold398 (.A(\game_inst.snake_inst.shiftreg_inst.memory[224][1] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold399 (.A(\game_inst.snake_inst.shiftreg_inst.memory[160][1] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold400 (.A(\game_inst.snake_inst.shiftreg_inst.memory[66][0] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold401 (.A(\game_inst.snake_inst.shiftreg_inst.memory[175][0] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold402 (.A(\game_inst.snake_inst.shiftreg_inst.memory[143][1] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold403 (.A(\game_inst.snake_inst.shiftreg_inst.memory[21][1] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold404 (.A(\game_inst.snake_inst.shiftreg_inst.memory[57][1] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold405 (.A(\game_inst.snake_inst.shiftreg_inst.memory[141][0] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold406 (.A(\game_inst.snake_inst.shiftreg_inst.memory[180][1] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold407 (.A(\game_inst.snake_inst.shiftreg_inst.memory[220][1] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold408 (.A(\game_inst.snake_inst.shiftreg_inst.memory[227][1] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold409 (.A(\game_inst.snake_inst.shiftreg_inst.memory[62][1] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold410 (.A(\game_inst.snake_inst.shiftreg_inst.memory[85][1] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold411 (.A(\game_inst.snake_inst.shiftreg_inst.memory[199][1] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold412 (.A(\game_inst.snake_inst.shiftreg_inst.memory[35][1] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold413 (.A(\game_inst.snake_inst.shiftreg_inst.memory[205][0] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold414 (.A(\game_inst.snake_inst.shiftreg_inst.memory[222][0] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold415 (.A(\game_inst.snake_inst.shiftreg_inst.memory[172][1] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold416 (.A(\game_inst.snake_inst.shiftreg_inst.memory[176][0] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold417 (.A(\game_inst.snake_inst.shiftreg_inst.memory[159][1] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold418 (.A(\game_inst.snake_inst.shiftreg_inst.memory[22][1] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold419 (.A(\game_inst.snake_inst.shiftreg_inst.memory[198][1] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold420 (.A(\game_inst.snake_inst.shiftreg_inst.memory[203][0] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold421 (.A(\game_inst.snake_inst.shiftreg_inst.memory[170][0] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold422 (.A(\game_inst.snake_inst.shiftreg_inst.memory[23][1] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold423 (.A(\game_inst.snake_inst.shiftreg_inst.memory[54][1] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold424 (.A(\game_inst.snake_inst.shiftreg_inst.memory[63][0] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold425 (.A(\game_inst.snake_inst.shiftreg_inst.memory[194][1] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold426 (.A(\game_inst.snake_inst.shiftreg_inst.memory[119][1] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold427 (.A(\game_inst.snake_inst.shiftreg_inst.memory[116][1] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold428 (.A(\game_inst.snake_inst.shiftreg_inst.memory[118][1] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold429 (.A(\game_inst.snake_inst.shiftreg_inst.memory[54][0] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold430 (.A(\game_inst.snake_inst.shiftreg_inst.memory[208][1] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold431 (.A(\game_inst.snake_inst.shiftreg_inst.memory[38][0] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold432 (.A(\game_inst.snake_inst.shiftreg_inst.memory[27][1] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold433 (.A(\game_inst.snake_inst.shiftreg_inst.memory[177][1] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold434 (.A(\game_inst.snake_inst.shiftreg_inst.memory[120][1] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold435 (.A(\game_inst.snake_inst.shiftreg_inst.memory[200][1] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold436 (.A(\game_inst.snake_inst.shiftreg_inst.memory[8][0] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold437 (.A(\game_inst.snake_inst.shiftreg_inst.memory[213][1] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold438 (.A(\game_inst.snake_inst.shiftreg_inst.memory[184][1] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold439 (.A(\game_inst.snake_inst.shiftreg_inst.memory[38][1] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold440 (.A(\game_inst.snake_inst.shiftreg_inst.memory[52][0] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold441 (.A(\game_inst.snake_inst.shiftreg_inst.memory[193][1] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold442 (.A(\game_inst.snake_inst.shiftreg_inst.memory[201][0] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold443 (.A(\game_inst.snake_inst.shiftreg_inst.memory[14][1] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold444 (.A(\game_inst.snake_inst.shiftreg_inst.memory[226][1] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold445 (.A(\game_inst.snake_inst.shiftreg_inst.memory[164][0] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold446 (.A(\game_inst.snake_inst.shiftreg_inst.memory[143][0] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold447 (.A(\game_inst.snake_inst.shiftreg_inst.memory[61][1] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold448 (.A(\game_inst.snake_inst.shiftreg_inst.memory[230][0] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold449 (.A(\game_inst.snake_inst.shiftreg_inst.memory[80][0] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold450 (.A(\game_inst.snake_inst.shiftreg_inst.memory[212][0] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold451 (.A(\game_inst.snake_inst.shiftreg_inst.memory[89][1] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold452 (.A(\game_inst.snake_inst.shiftreg_inst.memory[48][0] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold453 (.A(\game_inst.snake_inst.shiftreg_inst.memory[70][1] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold454 (.A(\game_inst.snake_inst.shiftreg_inst.memory[189][0] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold455 (.A(\game_inst.snake_inst.shiftreg_inst.memory[165][0] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold456 (.A(\game_inst.snake_inst.shiftreg_inst.memory[35][0] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold457 (.A(\game_inst.snake_inst.shiftreg_inst.memory[148][0] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold458 (.A(\game_inst.snake_inst.shiftreg_inst.memory[115][0] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold459 (.A(\game_inst.snake_inst.shiftreg_inst.memory[135][0] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold460 (.A(\game_inst.snake_inst.shiftreg_inst.memory[97][0] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold461 (.A(\game_inst.vga_inst.s_vsync ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold462 (.A(\game_inst.snake_inst.shiftreg_inst.memory[110][0] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold463 (.A(\game_inst.snake_inst.shiftreg_inst.memory[139][1] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold464 (.A(\game_inst.snake_inst.shiftreg_inst.memory[29][0] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold465 (.A(\game_inst.snake_inst.shiftreg_inst.memory[17][0] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold466 (.A(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold467 (.A(\game_inst.pos_dir[0] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold468 (.A(\game_inst.vga_inst.px[0] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold469 (.A(\game_inst.vga_inst.px[1] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold470 (.A(failure),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0002_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold472 (.A(\game_inst.vga_inst.row_buffer[8][2] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0034_),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold474 (.A(\game_inst.snake_inst.length[7] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0117_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold476 (.A(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0083_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold478 (.A(\game_inst.vga_inst.row_buffer[8][0] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0032_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold480 (.A(\game_inst.vga_inst.row_buffer[8][3] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0035_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold482 (.A(\game_inst.snake_inst.pos[7] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0121_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold484 (.A(\game_inst.vga_inst.row_buffer[8][1] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0033_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold486 (.A(\game_inst.tickgen_inst.counter[3] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0134_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold488 (.A(\game_inst.apple_inst.test ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0486_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold490 (.A(\game_inst.tickgen_inst.counter[0] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold491 (.A(\game_inst.snake_inst.dir_out[0] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0054_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold493 (.A(\game_inst.vga_inst.py[4] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0037_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold495 (.A(\game_inst.vga_inst.px[2] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold496 (.A(\game_inst.vga_inst.py[0] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0060_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold498 (.A(\game_inst.snake_inst.pos[0] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0049_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold500 (.A(\game_inst.snake_inst.length[6] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0643_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0116_),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold503 (.A(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0082_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold505 (.A(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0123_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold507 (.A(\game_inst.pos_dir[1] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold508 (.A(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0071_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold510 (.A(\game_inst.vga_inst.py[1] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0422_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0061_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold513 (.A(\game_inst.snake_inst.dir_out[1] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0055_),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold515 (.A(\game_inst.tickgen_inst.counter[2] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0683_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold517 (.A(\game_inst.apple_inst.apple_y[3] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0125_),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold519 (.A(\game_inst.apple_inst.apple_x[1] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0072_),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold521 (.A(\game_inst.tick ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0671_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0130_),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold524 (.A(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold525 (.A(_0508_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold526 (.A(\game_inst.snake_inst.pos[4] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0648_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0120_),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold529 (.A(\game_inst.apple_inst.apple_x[2] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold530 (.A(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold531 (.A(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold532 (.A(\game_inst.apple_inst.apple_y[0] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold533 (.A(\game_inst.apple_inst.apple_x[3] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold534 (.A(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold535 (.A(\game_inst.apple_inst.o_ready ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold536 (.A(\game_inst.vga_inst.py[9] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0069_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold538 (.A(\game_inst.control_inst.dir[1] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold539 (.A(\game_inst.control_inst.i_head_dir[0] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0087_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold541 (.A(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0075_),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold543 (.A(\game_inst.vga_inst.row_buffer[0][0] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0056_),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold545 (.A(\game_inst.vga_inst.py[3] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0254_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0430_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0064_),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold549 (.A(\game_inst.vga_inst.py[2] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold550 (.A(\game_inst.vga_inst.py[8] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0436_),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0068_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold553 (.A(\game_inst.apple_inst.apple_y[2] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold554 (.A(\game_inst.snake_inst.pos[2] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0647_),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0119_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold557 (.A(\game_inst.snake_inst.length[4] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0639_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0114_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold560 (.A(\game_inst.control_inst.o_start ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0652_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold562 (.A(\game_inst.vga_inst.row_buffer[0][2] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold563 (.A(_0058_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold564 (.A(\game_inst.vga_inst.row_buffer[0][3] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0059_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold566 (.A(\game_inst.control_inst.backwards[1] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold567 (.A(\game_inst.vga_inst.row_buffer[0][1] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0057_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold569 (.A(\game_inst.snake_inst.length[1] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0632_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0111_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold572 (.A(\game_inst.apple_inst.i_snake_y[1] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0107_),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold574 (.A(\game_inst.vga_inst.px[5] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0382_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0045_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold577 (.A(\game_inst.vga_inst.py[7] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold578 (.A(_0067_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold579 (.A(\game_inst.snake_inst.length[5] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0641_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold581 (.A(\game_inst.apple_inst.apple_x[0] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0207_),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold583 (.A(_0208_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold584 (.A(\game_inst.apple_inst.i_snake_valid ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold585 (.A(\game_inst.head_x[0] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold586 (.A(\game_inst.apple_inst.i_snake_x[1] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0101_),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold588 (.A(\game_inst.snake_inst.pos[6] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0410_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0052_),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold591 (.A(\game_inst.vga_inst.px[3] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold592 (.A(\game_inst.tickgen_inst.counter[1] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold593 (.A(\game_inst.head_y[0] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold594 (.A(\game_inst.tickgen_inst.counter_max[3] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0664_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0129_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold597 (.A(\game_inst.head_x[4] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold598 (.A(\game_inst.snake_inst.length[3] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0636_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0113_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold601 (.A(\game_inst.head_x[2] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold602 (.A(\game_inst.vga_inst.py[5] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0432_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold604 (.A(\game_inst.tickgen_inst.counter_max[1] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0654_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold606 (.A(\game_inst.snake_inst.length[2] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0635_),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0112_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold609 (.A(\game_inst.apple_inst.i_snake_x[4] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold610 (.A(\game_inst.vga_inst.row_buffer[7][2] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold611 (.A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0109_),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold613 (.A(\game_inst.vga_inst.row_buffer[7][0] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold614 (.A(\game_inst.apple_inst.i_snake_y[2] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0108_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold616 (.A(\game_inst.head_x[3] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0092_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold618 (.A(\game_inst.snake_inst.pos[3] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold619 (.A(\game_inst.vga_inst.row_buffer[7][3] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold620 (.A(\game_inst.vga_inst.row_buffer[7][1] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold621 (.A(\game_inst.vga_inst.px[4] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0043_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold623 (.A(\game_inst.head_y[1] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold624 (.A(\game_inst.head_y[2] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold625 (.A(\game_inst.vga_inst.row_buffer[6][3] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold626 (.A(_0023_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold627 (.A(\game_inst.vga_inst.row_buffer[6][2] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0022_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold629 (.A(\game_inst.vga_inst.row_buffer[6][0] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0020_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold631 (.A(\game_inst.vga_inst.row_buffer[4][2] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0014_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold633 (.A(\game_inst.vga_inst.row_buffer[4][3] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0015_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold635 (.A(\game_inst.vga_inst.row_buffer[3][3] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold636 (.A(_0011_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold637 (.A(\game_inst.vga_inst.row_buffer[5][3] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold638 (.A(\game_inst.vga_inst.row_buffer[5][2] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold639 (.A(\game_inst.snake_inst.pos[1] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold640 (.A(\game_inst.vga_inst.row_buffer[3][0] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0008_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold642 (.A(\game_inst.snake_inst.pos[5] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold643 (.A(\game_inst.vga_inst.row_buffer[4][0] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold644 (.A(_0016_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold645 (.A(\game_inst.vga_inst.row_buffer[4][1] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold646 (.A(_0013_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold647 (.A(\game_inst.snake_inst.length[0] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold648 (.A(\game_inst.vga_inst.row_buffer[5][1] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold649 (.A(\game_inst.vga_inst.row_buffer[3][2] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0010_),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold651 (.A(\game_inst.apple_inst.i_snake_x[3] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold652 (.A(_0103_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold653 (.A(\game_inst.vga_inst.row_buffer[2][0] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold654 (.A(_0004_),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold655 (.A(\game_inst.vga_inst.row_buffer[6][1] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold656 (.A(\game_inst.vga_inst.row_buffer[1][3] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold657 (.A(_0007_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold658 (.A(\game_inst.head_x[1] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold659 (.A(\game_inst.vga_inst.row_buffer[1][2] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0006_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold661 (.A(\game_inst.vga_inst.row_buffer[1][1] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0005_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold663 (.A(\game_inst.vga_inst.row_buffer[3][1] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0009_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold665 (.A(\game_inst.vga_inst.px[9] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0036_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold667 (.A(\game_inst.apple_inst.i_snake_x[2] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold668 (.A(\game_inst.vga_inst.px[7] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0384_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold670 (.A(_0046_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold671 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold672 (.A(\game_inst.vga_inst.px[8] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold673 (.A(\game_inst.vga_inst.py[6] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold674 (.A(\game_inst.vga_inst.px[8] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold675 (.A(\game_inst.head_y[3] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold676 (.A(\game_inst.apple_inst.i_snake_y[0] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold677 (.A(\game_inst.control_inst.i_head_dir[0] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold678 (.A(\game_inst.tickgen_inst.counter_max[2] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold679 (.A(_0659_),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0128_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold681 (.A(\game_inst.vga_inst.px[4] ),
    .X(net1345));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_fill_2 FILLER_0_84 ();
 sg13g2_fill_1 FILLER_0_86 ();
 sg13g2_fill_2 FILLER_0_139 ();
 sg13g2_fill_1 FILLER_0_141 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_fill_2 FILLER_0_207 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_215 ();
 sg13g2_fill_2 FILLER_0_261 ();
 sg13g2_fill_2 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_fill_1 FILLER_1_81 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_2 FILLER_1_177 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_fill_2 FILLER_1_216 ();
 sg13g2_fill_1 FILLER_1_218 ();
 sg13g2_fill_1 FILLER_1_282 ();
 sg13g2_fill_1 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_32 ();
 sg13g2_decap_4 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_46 ();
 sg13g2_fill_1 FILLER_2_51 ();
 sg13g2_decap_4 FILLER_2_61 ();
 sg13g2_fill_2 FILLER_2_73 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_4 ();
 sg13g2_fill_2 FILLER_3_13 ();
 sg13g2_fill_1 FILLER_3_15 ();
 sg13g2_fill_2 FILLER_3_20 ();
 sg13g2_fill_2 FILLER_3_76 ();
 sg13g2_fill_1 FILLER_3_78 ();
 sg13g2_fill_1 FILLER_3_115 ();
 sg13g2_fill_2 FILLER_3_129 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_250 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_fill_2 FILLER_4_31 ();
 sg13g2_fill_1 FILLER_4_33 ();
 sg13g2_fill_2 FILLER_4_88 ();
 sg13g2_fill_1 FILLER_4_90 ();
 sg13g2_fill_2 FILLER_4_122 ();
 sg13g2_fill_1 FILLER_4_124 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_fill_2 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_297 ();
 sg13g2_fill_1 FILLER_4_299 ();
 sg13g2_fill_2 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_47 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_320 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_fill_2 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_1 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_229 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_2 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_334 ();
 sg13g2_fill_1 FILLER_6_336 ();
 sg13g2_fill_2 FILLER_6_364 ();
 sg13g2_fill_2 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_2 FILLER_6_386 ();
 sg13g2_fill_1 FILLER_6_388 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_1 FILLER_7_37 ();
 sg13g2_fill_1 FILLER_7_65 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_2 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_2 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_fill_2 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_325 ();
 sg13g2_fill_2 FILLER_7_370 ();
 sg13g2_fill_1 FILLER_7_372 ();
 sg13g2_fill_2 FILLER_7_382 ();
 sg13g2_fill_1 FILLER_7_393 ();
 sg13g2_fill_2 FILLER_7_403 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_2 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_8_382 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_32 ();
 sg13g2_fill_1 FILLER_9_51 ();
 sg13g2_fill_1 FILLER_9_115 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_238 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_fill_2 FILLER_9_327 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_393 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_2 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_11_31 ();
 sg13g2_fill_1 FILLER_11_33 ();
 sg13g2_fill_1 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_317 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_fill_1 FILLER_12_16 ();
 sg13g2_fill_1 FILLER_12_177 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_4 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_23 ();
 sg13g2_fill_1 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_fill_2 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_351 ();
 sg13g2_fill_2 FILLER_14_379 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_51 ();
 sg13g2_fill_2 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_11 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_365 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_17_8 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_13 ();
 sg13g2_fill_1 FILLER_18_15 ();
 sg13g2_fill_1 FILLER_18_51 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_fill_2 FILLER_19_103 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_fill_2 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_100 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_19 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_29 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_5 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_43 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_decap_4 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_fill_2 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_decap_4 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_decap_4 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_decap_4 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_decap_4 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_213 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_106 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_fill_2 FILLER_39_82 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_154 ();
 sg13g2_fill_1 FILLER_39_185 ();
 sg13g2_fill_2 FILLER_39_202 ();
 sg13g2_fill_1 FILLER_39_204 ();
 sg13g2_fill_1 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_fill_1 FILLER_39_285 ();
 sg13g2_fill_2 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_fill_2 FILLER_40_58 ();
 sg13g2_fill_1 FILLER_40_95 ();
 sg13g2_fill_2 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_fill_1 FILLER_40_148 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_184 ();
 sg13g2_decap_8 FILLER_40_191 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_fill_1 FILLER_41_39 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_decap_8 FILLER_41_152 ();
 sg13g2_decap_4 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_47 ();
 sg13g2_fill_2 FILLER_42_92 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_fill_2 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_166 ();
 sg13g2_fill_2 FILLER_42_216 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_fill_2 FILLER_42_317 ();
 sg13g2_fill_1 FILLER_42_319 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_2 FILLER_42_380 ();
 sg13g2_fill_2 FILLER_43_80 ();
 sg13g2_fill_2 FILLER_43_136 ();
 sg13g2_fill_1 FILLER_43_138 ();
 sg13g2_decap_4 FILLER_43_160 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_238 ();
 sg13g2_fill_2 FILLER_43_292 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_182 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_55 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_118 ();
 sg13g2_fill_1 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_130 ();
 sg13g2_fill_2 FILLER_45_145 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_decap_4 FILLER_45_164 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_fill_2 FILLER_45_310 ();
 sg13g2_fill_1 FILLER_45_348 ();
 sg13g2_fill_2 FILLER_45_380 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_2 FILLER_46_30 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_fill_2 FILLER_46_73 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_decap_4 FILLER_46_174 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_274 ();
 sg13g2_fill_2 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_47 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_2 FILLER_47_292 ();
 sg13g2_fill_2 FILLER_47_307 ();
 sg13g2_fill_2 FILLER_47_318 ();
 sg13g2_fill_1 FILLER_47_320 ();
 sg13g2_fill_2 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_48_27 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_143 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_fill_2 FILLER_48_229 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_305 ();
 sg13g2_fill_2 FILLER_48_343 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_96 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_184 ();
 sg13g2_decap_4 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_2 FILLER_49_276 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_355 ();
 sg13g2_fill_1 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_398 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_fill_1 FILLER_50_48 ();
 sg13g2_fill_2 FILLER_50_85 ();
 sg13g2_fill_1 FILLER_50_87 ();
 sg13g2_fill_2 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_207 ();
 sg13g2_fill_1 FILLER_50_225 ();
 sg13g2_fill_2 FILLER_50_250 ();
 sg13g2_fill_2 FILLER_50_284 ();
 sg13g2_fill_1 FILLER_50_335 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_29 ();
 sg13g2_fill_1 FILLER_51_66 ();
 sg13g2_fill_2 FILLER_51_76 ();
 sg13g2_fill_2 FILLER_51_97 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_fill_2 FILLER_51_249 ();
 sg13g2_fill_1 FILLER_51_372 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_1 FILLER_52_126 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_decap_4 FILLER_52_181 ();
 sg13g2_fill_1 FILLER_52_185 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_fill_2 FILLER_53_149 ();
 sg13g2_fill_1 FILLER_53_151 ();
 sg13g2_fill_1 FILLER_53_177 ();
 sg13g2_fill_2 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_53_215 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_fill_2 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_336 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_108 ();
 sg13g2_fill_1 FILLER_54_133 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_251 ();
 sg13g2_fill_1 FILLER_54_253 ();
 sg13g2_fill_2 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_2 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_62 ();
 sg13g2_fill_2 FILLER_55_103 ();
 sg13g2_fill_1 FILLER_55_134 ();
 sg13g2_fill_1 FILLER_55_150 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_220 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_fill_1 FILLER_55_284 ();
 sg13g2_fill_1 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_1 FILLER_56_40 ();
 sg13g2_fill_2 FILLER_56_81 ();
 sg13g2_fill_1 FILLER_56_83 ();
 sg13g2_fill_2 FILLER_56_117 ();
 sg13g2_fill_1 FILLER_56_119 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_fill_2 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_331 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_2 FILLER_56_397 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_45 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_208 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_fill_1 FILLER_57_296 ();
 sg13g2_fill_1 FILLER_57_301 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_51 ();
 sg13g2_fill_1 FILLER_58_53 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_127 ();
 sg13g2_fill_1 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_200 ();
 sg13g2_fill_2 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_316 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_29 ();
 sg13g2_fill_1 FILLER_59_31 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_fill_2 FILLER_59_97 ();
 sg13g2_fill_2 FILLER_59_159 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_37 ();
 sg13g2_fill_1 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_131 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_2 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_263 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_82 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_fill_2 FILLER_61_136 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_197 ();
 sg13g2_fill_2 FILLER_61_216 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_2 FILLER_61_284 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_fill_2 FILLER_62_13 ();
 sg13g2_fill_1 FILLER_62_64 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_341 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_15 ();
 sg13g2_fill_2 FILLER_63_79 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_fill_2 FILLER_63_192 ();
 sg13g2_fill_1 FILLER_63_208 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_359 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_2 FILLER_64_38 ();
 sg13g2_fill_1 FILLER_64_40 ();
 sg13g2_fill_2 FILLER_64_50 ();
 sg13g2_fill_1 FILLER_64_52 ();
 sg13g2_fill_2 FILLER_64_67 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_83 ();
 sg13g2_fill_2 FILLER_64_113 ();
 sg13g2_fill_1 FILLER_64_115 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_fill_1 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_decap_4 FILLER_64_394 ();
 sg13g2_fill_1 FILLER_64_398 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_55 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_2 FILLER_65_72 ();
 sg13g2_fill_2 FILLER_65_139 ();
 sg13g2_fill_2 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_fill_1 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_57 ();
 sg13g2_fill_1 FILLER_66_59 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_2 FILLER_66_158 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_310 ();
 sg13g2_fill_2 FILLER_66_334 ();
 sg13g2_decap_8 FILLER_66_398 ();
 sg13g2_decap_4 FILLER_66_405 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_fill_1 FILLER_67_16 ();
 sg13g2_fill_2 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_142 ();
 sg13g2_fill_1 FILLER_67_282 ();
 sg13g2_fill_1 FILLER_67_302 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_11 ();
 sg13g2_fill_2 FILLER_68_84 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_fill_1 FILLER_68_185 ();
 sg13g2_fill_1 FILLER_68_203 ();
 sg13g2_fill_2 FILLER_68_222 ();
 sg13g2_fill_1 FILLER_68_224 ();
 sg13g2_fill_1 FILLER_68_246 ();
 sg13g2_fill_2 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_fill_2 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_167 ();
 sg13g2_fill_2 FILLER_69_205 ();
 sg13g2_fill_2 FILLER_69_212 ();
 sg13g2_fill_2 FILLER_69_218 ();
 sg13g2_fill_2 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_fill_1 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_399 ();
 sg13g2_fill_1 FILLER_70_53 ();
 sg13g2_fill_1 FILLER_70_230 ();
 sg13g2_fill_1 FILLER_70_239 ();
 sg13g2_fill_2 FILLER_70_293 ();
 sg13g2_fill_2 FILLER_70_361 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_fill_2 FILLER_71_31 ();
 sg13g2_fill_1 FILLER_71_33 ();
 sg13g2_fill_2 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_fill_2 FILLER_71_256 ();
 sg13g2_fill_1 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_265 ();
 sg13g2_fill_1 FILLER_71_381 ();
 sg13g2_fill_2 FILLER_72_4 ();
 sg13g2_fill_1 FILLER_72_6 ();
 sg13g2_fill_2 FILLER_72_38 ();
 sg13g2_fill_1 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_77 ();
 sg13g2_fill_1 FILLER_72_115 ();
 sg13g2_fill_1 FILLER_72_143 ();
 sg13g2_fill_2 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_fill_2 FILLER_72_310 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_fill_1 FILLER_72_372 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_69 ();
 sg13g2_fill_2 FILLER_73_83 ();
 sg13g2_fill_2 FILLER_73_166 ();
 sg13g2_fill_2 FILLER_73_262 ();
 sg13g2_fill_1 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_fill_2 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_379 ();
 sg13g2_fill_2 FILLER_74_397 ();
 sg13g2_fill_1 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_10 ();
 sg13g2_fill_2 FILLER_75_51 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_2 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_2 FILLER_75_318 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_1 FILLER_76_236 ();
 sg13g2_fill_1 FILLER_76_294 ();
 sg13g2_fill_2 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_350 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_381 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_36 ();
 sg13g2_fill_2 FILLER_77_99 ();
 sg13g2_fill_1 FILLER_77_101 ();
 sg13g2_fill_1 FILLER_77_169 ();
 sg13g2_fill_1 FILLER_77_183 ();
 sg13g2_fill_2 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_301 ();
 sg13g2_fill_2 FILLER_77_351 ();
 sg13g2_fill_1 FILLER_77_353 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_fill_1 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_fill_2 FILLER_77_398 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_fill_2 FILLER_78_30 ();
 sg13g2_fill_1 FILLER_78_49 ();
 sg13g2_fill_1 FILLER_78_120 ();
 sg13g2_fill_1 FILLER_78_194 ();
 sg13g2_fill_2 FILLER_78_305 ();
 sg13g2_fill_2 FILLER_78_311 ();
 sg13g2_fill_1 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_78_335 ();
 sg13g2_decap_4 FILLER_78_342 ();
 sg13g2_fill_2 FILLER_78_346 ();
 sg13g2_decap_8 FILLER_78_352 ();
 sg13g2_fill_2 FILLER_78_359 ();
 sg13g2_fill_1 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_366 ();
 sg13g2_decap_4 FILLER_78_373 ();
 sg13g2_fill_1 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_2 FILLER_79_20 ();
 sg13g2_fill_1 FILLER_79_30 ();
 sg13g2_fill_1 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_66 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_fill_1 FILLER_79_78 ();
 sg13g2_fill_1 FILLER_79_109 ();
 sg13g2_fill_1 FILLER_79_159 ();
 sg13g2_fill_1 FILLER_79_186 ();
 sg13g2_fill_1 FILLER_79_192 ();
 sg13g2_fill_1 FILLER_79_207 ();
 sg13g2_fill_2 FILLER_79_234 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_312 ();
 sg13g2_decap_4 FILLER_79_319 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_328 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_decap_8 FILLER_79_342 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_fill_2 FILLER_80_20 ();
 sg13g2_fill_1 FILLER_80_66 ();
 sg13g2_fill_1 FILLER_80_83 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_266 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_315 ();
 sg13g2_decap_4 FILLER_80_322 ();
 sg13g2_fill_2 FILLER_80_326 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net661;
 assign uio_oe[1] = net662;
 assign uio_oe[2] = net663;
 assign uio_oe[3] = net664;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[4] = net11;
 assign uio_out[5] = net12;
 assign uio_out[6] = net13;
 assign uio_out[7] = net14;
endmodule
