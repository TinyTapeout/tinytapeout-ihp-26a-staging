module tt_um_embeddedinn_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire \frame_cnt[0] ;
 wire \frame_cnt[10] ;
 wire \frame_cnt[11] ;
 wire \frame_cnt[12] ;
 wire \frame_cnt[13] ;
 wire \frame_cnt[1] ;
 wire \frame_cnt[2] ;
 wire \frame_cnt[3] ;
 wire \frame_cnt[4] ;
 wire \frame_cnt[5] ;
 wire \frame_cnt[6] ;
 wire \frame_cnt[7] ;
 wire \frame_cnt[8] ;
 wire \frame_cnt[9] ;
 wire hsync;
 wire \hvsync_gen.display_on ;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \tx[0] ;
 wire \tx[1] ;
 wire \tx[3] ;
 wire \tx[4] ;
 wire \tx[7] ;
 wire \tx[8] ;
 wire \ty[0] ;
 wire \ty[1] ;
 wire \ty[3] ;
 wire \ty[4] ;
 wire \ty[7] ;
 wire \ty[8] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire vsync_prev;
 wire x_dir;
 wire y_dir;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;

 sg13g2_inv_1 _426_ (.Y(_063_),
    .A(net84));
 sg13g2_inv_1 _427_ (.Y(_064_),
    .A(_014_));
 sg13g2_inv_1 _428_ (.Y(_065_),
    .A(net114));
 sg13g2_inv_2 _429_ (.Y(_066_),
    .A(net128));
 sg13g2_inv_1 _430_ (.Y(_067_),
    .A(\frame_cnt[0] ));
 sg13g2_inv_1 _431_ (.Y(_068_),
    .A(net139));
 sg13g2_inv_1 _432_ (.Y(_069_),
    .A(\ty[7] ));
 sg13g2_inv_1 _433_ (.Y(_070_),
    .A(\ty[4] ));
 sg13g2_inv_1 _434_ (.Y(_071_),
    .A(\ty[8] ));
 sg13g2_inv_2 _435_ (.Y(_072_),
    .A(net98));
 sg13g2_inv_4 _436_ (.A(net80),
    .Y(_073_));
 sg13g2_inv_1 _437_ (.Y(_074_),
    .A(\hvsync_gen.vpos[4] ));
 sg13g2_inv_1 _438_ (.Y(_075_),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_inv_1 _439_ (.Y(_076_),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_inv_1 _440_ (.Y(_077_),
    .A(\frame_cnt[1] ));
 sg13g2_inv_1 _441_ (.Y(_078_),
    .A(net46));
 sg13g2_inv_1 _442_ (.Y(_079_),
    .A(net4));
 sg13g2_inv_2 _443_ (.Y(_080_),
    .A(net3));
 sg13g2_inv_1 _444_ (.Y(_081_),
    .A(\hvsync_gen.display_on ));
 sg13g2_inv_4 _445_ (.A(net54),
    .Y(_082_));
 sg13g2_inv_2 _446_ (.Y(_083_),
    .A(net57));
 sg13g2_nand2_1 _447_ (.Y(_084_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net95));
 sg13g2_nor3_2 _448_ (.A(_072_),
    .B(_073_),
    .C(_084_),
    .Y(_085_));
 sg13g2_nor3_1 _449_ (.A(_075_),
    .B(\hvsync_gen.vpos[2] ),
    .C(net44),
    .Y(_086_));
 sg13g2_nand4_1 _450_ (.B(_074_),
    .C(net81),
    .A(net86),
    .Y(_012_),
    .D(_086_));
 sg13g2_nor3_1 _451_ (.A(\hvsync_gen.hpos[6] ),
    .B(\hvsync_gen.hpos[4] ),
    .C(net56),
    .Y(_087_));
 sg13g2_nand4_1 _452_ (.B(\hvsync_gen.hpos[6] ),
    .C(\hvsync_gen.hpos[4] ),
    .A(net55),
    .Y(_088_),
    .D(net56));
 sg13g2_nor2_1 _453_ (.A(\hvsync_gen.hpos[8] ),
    .B(_087_),
    .Y(_089_));
 sg13g2_nand4_1 _454_ (.B(net55),
    .C(_088_),
    .A(net91),
    .Y(_011_),
    .D(_089_));
 sg13g2_nand2_2 _455_ (.Y(_090_),
    .A(net91),
    .B(net93));
 sg13g2_o21ai_1 _456_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_091_),
    .A1(\hvsync_gen.hpos[8] ),
    .A2(net55));
 sg13g2_inv_1 _457_ (.Y(_092_),
    .A(_091_));
 sg13g2_nor3_1 _458_ (.A(net44),
    .B(_085_),
    .C(_092_),
    .Y(_000_));
 sg13g2_and3_1 _459_ (.X(_093_),
    .A(net125),
    .B(net77),
    .C(net88));
 sg13g2_and2_1 _460_ (.A(net120),
    .B(_093_),
    .X(_094_));
 sg13g2_and2_1 _461_ (.A(net127),
    .B(_094_),
    .X(_095_));
 sg13g2_nor4_2 _462_ (.A(net55),
    .B(\hvsync_gen.hpos[6] ),
    .C(net56),
    .Y(_096_),
    .D(_095_));
 sg13g2_nor2_1 _463_ (.A(_090_),
    .B(_096_),
    .Y(_097_));
 sg13g2_nor2_1 _464_ (.A(net77),
    .B(net47),
    .Y(_001_));
 sg13g2_xnor2_1 _465_ (.Y(_098_),
    .A(net125),
    .B(net77));
 sg13g2_nor2_1 _466_ (.A(net47),
    .B(_098_),
    .Y(_002_));
 sg13g2_a21oi_1 _467_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(net77),
    .Y(_099_),
    .B1(net88));
 sg13g2_nor3_1 _468_ (.A(_093_),
    .B(net48),
    .C(net89),
    .Y(_003_));
 sg13g2_nor2_1 _469_ (.A(net120),
    .B(_093_),
    .Y(_100_));
 sg13g2_nor3_1 _470_ (.A(_094_),
    .B(net47),
    .C(net121),
    .Y(_004_));
 sg13g2_nor2_1 _471_ (.A(net127),
    .B(_094_),
    .Y(_101_));
 sg13g2_nor3_1 _472_ (.A(_095_),
    .B(net47),
    .C(_101_),
    .Y(_005_));
 sg13g2_and2_1 _473_ (.A(net56),
    .B(_095_),
    .X(_102_));
 sg13g2_o21ai_1 _474_ (.B1(_090_),
    .Y(_103_),
    .A1(net56),
    .A2(_095_));
 sg13g2_nor2_1 _475_ (.A(_102_),
    .B(_103_),
    .Y(_006_));
 sg13g2_nor2_1 _476_ (.A(net119),
    .B(_102_),
    .Y(_104_));
 sg13g2_and2_1 _477_ (.A(net119),
    .B(_102_),
    .X(_105_));
 sg13g2_nor3_1 _478_ (.A(net47),
    .B(_104_),
    .C(_105_),
    .Y(_007_));
 sg13g2_and2_1 _479_ (.A(net55),
    .B(_105_),
    .X(_106_));
 sg13g2_nor2_1 _480_ (.A(net55),
    .B(_105_),
    .Y(_107_));
 sg13g2_nor3_1 _481_ (.A(net47),
    .B(_106_),
    .C(_107_),
    .Y(_008_));
 sg13g2_xnor2_1 _482_ (.Y(_108_),
    .A(net93),
    .B(_106_));
 sg13g2_nor2_1 _483_ (.A(net47),
    .B(_108_),
    .Y(_009_));
 sg13g2_a21oi_1 _484_ (.A1(net93),
    .A2(_106_),
    .Y(_109_),
    .B1(net91));
 sg13g2_nor2_1 _485_ (.A(net47),
    .B(net94),
    .Y(_010_));
 sg13g2_nor2b_1 _486_ (.A(\tx[8] ),
    .B_N(\hvsync_gen.hpos[8] ),
    .Y(_110_));
 sg13g2_xnor2_1 _487_ (.Y(_111_),
    .A(\tx[8] ),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_and2_1 _488_ (.A(_013_),
    .B(\hvsync_gen.hpos[2] ),
    .X(_112_));
 sg13g2_xor2_1 _489_ (.B(\hvsync_gen.hpos[2] ),
    .A(_013_),
    .X(_113_));
 sg13g2_nor2b_1 _490_ (.A(\hvsync_gen.hpos[1] ),
    .B_N(\tx[1] ),
    .Y(_114_));
 sg13g2_nand2b_1 _491_ (.Y(_115_),
    .B(\hvsync_gen.hpos[1] ),
    .A_N(\tx[1] ));
 sg13g2_nor2b_1 _492_ (.A(\hvsync_gen.hpos[0] ),
    .B_N(\tx[0] ),
    .Y(_116_));
 sg13g2_o21ai_1 _493_ (.B1(_115_),
    .Y(_117_),
    .A1(_114_),
    .A2(_116_));
 sg13g2_a221oi_1 _494_ (.B2(_117_),
    .C1(_112_),
    .B1(_113_),
    .A1(_066_),
    .Y(_118_),
    .A2(\hvsync_gen.hpos[3] ));
 sg13g2_a21oi_1 _495_ (.A1(\tx[3] ),
    .A2(_076_),
    .Y(_119_),
    .B1(_118_));
 sg13g2_nor2b_1 _496_ (.A(\tx[4] ),
    .B_N(\hvsync_gen.hpos[4] ),
    .Y(_120_));
 sg13g2_xnor2_1 _497_ (.Y(_121_),
    .A(\tx[4] ),
    .B(\hvsync_gen.hpos[4] ));
 sg13g2_or2_1 _498_ (.X(_122_),
    .B(net56),
    .A(_014_));
 sg13g2_xor2_1 _499_ (.B(net56),
    .A(_014_),
    .X(_123_));
 sg13g2_and2_1 _500_ (.A(_121_),
    .B(_123_),
    .X(_124_));
 sg13g2_a21o_1 _501_ (.A2(\hvsync_gen.hpos[5] ),
    .A1(_014_),
    .B1(_120_),
    .X(_125_));
 sg13g2_a22oi_1 _502_ (.Y(_126_),
    .B1(_125_),
    .B2(_122_),
    .A2(_124_),
    .A1(_119_));
 sg13g2_nor2b_1 _503_ (.A(\tx[7] ),
    .B_N(net55),
    .Y(_127_));
 sg13g2_nand2b_1 _504_ (.Y(_128_),
    .B(net55),
    .A_N(\tx[7] ));
 sg13g2_nand2_1 _505_ (.Y(_129_),
    .A(_015_),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_nor2b_1 _506_ (.A(\hvsync_gen.hpos[7] ),
    .B_N(\tx[7] ),
    .Y(_130_));
 sg13g2_nor2_1 _507_ (.A(_129_),
    .B(_130_),
    .Y(_131_));
 sg13g2_nor2_1 _508_ (.A(_127_),
    .B(_131_),
    .Y(_132_));
 sg13g2_nor2_1 _509_ (.A(_015_),
    .B(\hvsync_gen.hpos[6] ),
    .Y(_133_));
 sg13g2_a221oi_1 _510_ (.B2(_128_),
    .C1(_130_),
    .B1(_133_),
    .A1(_126_),
    .Y(_134_),
    .A2(_132_));
 sg13g2_xor2_1 _511_ (.B(_134_),
    .A(_111_),
    .X(_135_));
 sg13g2_xnor2_1 _512_ (.Y(_136_),
    .A(_111_),
    .B(_134_));
 sg13g2_nor2_1 _513_ (.A(_127_),
    .B(_130_),
    .Y(_137_));
 sg13g2_xnor2_1 _514_ (.Y(_138_),
    .A(_015_),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_o21ai_1 _515_ (.B1(_129_),
    .Y(_139_),
    .A1(_126_),
    .A2(_133_));
 sg13g2_xnor2_1 _516_ (.Y(_140_),
    .A(_137_),
    .B(_139_));
 sg13g2_xor2_1 _517_ (.B(_138_),
    .A(_126_),
    .X(_141_));
 sg13g2_inv_1 _518_ (.Y(_142_),
    .A(_141_));
 sg13g2_a21oi_1 _519_ (.A1(_119_),
    .A2(_121_),
    .Y(_143_),
    .B1(_120_));
 sg13g2_xor2_1 _520_ (.B(_143_),
    .A(_123_),
    .X(_144_));
 sg13g2_and2_1 _521_ (.A(_141_),
    .B(_144_),
    .X(_145_));
 sg13g2_nand2_1 _522_ (.Y(_146_),
    .A(_141_),
    .B(_144_));
 sg13g2_nor2_1 _523_ (.A(_141_),
    .B(_144_),
    .Y(_147_));
 sg13g2_xor2_1 _524_ (.B(_144_),
    .A(_141_),
    .X(_148_));
 sg13g2_nand3b_1 _525_ (.B(_140_),
    .C(_135_),
    .Y(_149_),
    .A_N(_148_));
 sg13g2_nand3_1 _526_ (.B(_140_),
    .C(_147_),
    .A(_136_),
    .Y(_150_));
 sg13g2_nand2_1 _527_ (.Y(_151_),
    .A(_149_),
    .B(_150_));
 sg13g2_and2_1 _528_ (.A(_017_),
    .B(\hvsync_gen.vpos[5] ),
    .X(_152_));
 sg13g2_xor2_1 _529_ (.B(\hvsync_gen.vpos[5] ),
    .A(_017_),
    .X(_153_));
 sg13g2_nand2_1 _530_ (.Y(_154_),
    .A(_070_),
    .B(\hvsync_gen.vpos[4] ));
 sg13g2_xor2_1 _531_ (.B(\hvsync_gen.vpos[4] ),
    .A(\ty[4] ),
    .X(_155_));
 sg13g2_nor2b_1 _532_ (.A(\ty[3] ),
    .B_N(\hvsync_gen.vpos[3] ),
    .Y(_156_));
 sg13g2_nand2_1 _533_ (.Y(_157_),
    .A(_016_),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_xnor2_1 _534_ (.Y(_158_),
    .A(_016_),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_nand2b_1 _535_ (.Y(_159_),
    .B(\ty[1] ),
    .A_N(\hvsync_gen.vpos[1] ));
 sg13g2_nor2b_1 _536_ (.A(\ty[1] ),
    .B_N(\hvsync_gen.vpos[1] ),
    .Y(_160_));
 sg13g2_nand2b_1 _537_ (.Y(_161_),
    .B(\ty[0] ),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_a21oi_1 _538_ (.A1(_159_),
    .A2(_161_),
    .Y(_162_),
    .B1(_160_));
 sg13g2_o21ai_1 _539_ (.B1(_157_),
    .Y(_163_),
    .A1(_158_),
    .A2(_162_));
 sg13g2_xnor2_1 _540_ (.Y(_164_),
    .A(\ty[3] ),
    .B(\hvsync_gen.vpos[3] ));
 sg13g2_a21oi_1 _541_ (.A1(_163_),
    .A2(_164_),
    .Y(_165_),
    .B1(_156_));
 sg13g2_o21ai_1 _542_ (.B1(_154_),
    .Y(_166_),
    .A1(_155_),
    .A2(_165_));
 sg13g2_xor2_1 _543_ (.B(_166_),
    .A(_153_),
    .X(_167_));
 sg13g2_xnor2_1 _544_ (.Y(_168_),
    .A(_153_),
    .B(_166_));
 sg13g2_xor2_1 _545_ (.B(_165_),
    .A(_155_),
    .X(_169_));
 sg13g2_inv_1 _546_ (.Y(_170_),
    .A(_169_));
 sg13g2_xnor2_1 _547_ (.Y(_171_),
    .A(_163_),
    .B(_164_));
 sg13g2_nor2_1 _548_ (.A(_170_),
    .B(_171_),
    .Y(_172_));
 sg13g2_xnor2_1 _549_ (.Y(_173_),
    .A(_113_),
    .B(_117_));
 sg13g2_xnor2_1 _550_ (.Y(_174_),
    .A(\tx[3] ),
    .B(\hvsync_gen.hpos[3] ));
 sg13g2_a21oi_1 _551_ (.A1(_113_),
    .A2(_117_),
    .Y(_175_),
    .B1(_112_));
 sg13g2_xnor2_1 _552_ (.Y(_176_),
    .A(_174_),
    .B(_175_));
 sg13g2_xnor2_1 _553_ (.Y(_177_),
    .A(_119_),
    .B(_121_));
 sg13g2_inv_1 _554_ (.Y(_178_),
    .A(_177_));
 sg13g2_nand3_1 _555_ (.B(_176_),
    .C(_177_),
    .A(_173_),
    .Y(_179_));
 sg13g2_nor3_1 _556_ (.A(_167_),
    .B(_172_),
    .C(_179_),
    .Y(_180_));
 sg13g2_and2_1 _557_ (.A(_149_),
    .B(_180_),
    .X(_181_));
 sg13g2_nand2b_2 _558_ (.Y(_182_),
    .B(_173_),
    .A_N(_176_));
 sg13g2_inv_1 _559_ (.Y(_183_),
    .A(_182_));
 sg13g2_xor2_1 _560_ (.B(_177_),
    .A(_176_),
    .X(_184_));
 sg13g2_xor2_1 _561_ (.B(_162_),
    .A(_158_),
    .X(_185_));
 sg13g2_xnor2_1 _562_ (.Y(_186_),
    .A(_173_),
    .B(_185_));
 sg13g2_nor2b_2 _563_ (.A(_169_),
    .B_N(_171_),
    .Y(_187_));
 sg13g2_nand2b_1 _564_ (.Y(_188_),
    .B(_167_),
    .A_N(_187_));
 sg13g2_xnor2_1 _565_ (.Y(_189_),
    .A(_171_),
    .B(_176_));
 sg13g2_o21ai_1 _566_ (.B1(_189_),
    .Y(_190_),
    .A1(_169_),
    .A2(_184_));
 sg13g2_a221oi_1 _567_ (.B2(_168_),
    .C1(_186_),
    .B1(_187_),
    .A1(_169_),
    .Y(_191_),
    .A2(_184_));
 sg13g2_nand3b_1 _568_ (.B(_191_),
    .C(_188_),
    .Y(_192_),
    .A_N(_190_));
 sg13g2_o21ai_1 _569_ (.B1(_182_),
    .Y(_193_),
    .A1(_149_),
    .A2(_192_));
 sg13g2_o21ai_1 _570_ (.B1(_151_),
    .Y(_194_),
    .A1(_181_),
    .A2(_193_));
 sg13g2_nand3_1 _571_ (.B(_171_),
    .C(_185_),
    .A(_169_),
    .Y(_195_));
 sg13g2_or2_1 _572_ (.X(_196_),
    .B(_195_),
    .A(_167_));
 sg13g2_xnor2_1 _573_ (.Y(_197_),
    .A(_167_),
    .B(_185_));
 sg13g2_a21oi_1 _574_ (.A1(_187_),
    .A2(_197_),
    .Y(_198_),
    .B1(_183_));
 sg13g2_nand3_1 _575_ (.B(_140_),
    .C(_145_),
    .A(_136_),
    .Y(_199_));
 sg13g2_nand2b_1 _576_ (.Y(_200_),
    .B(_177_),
    .A_N(_182_));
 sg13g2_o21ai_1 _577_ (.B1(_200_),
    .Y(_201_),
    .A1(_167_),
    .A2(_195_));
 sg13g2_a21oi_1 _578_ (.A1(_187_),
    .A2(_197_),
    .Y(_202_),
    .B1(_201_));
 sg13g2_a21o_1 _579_ (.A2(_197_),
    .A1(_187_),
    .B1(_201_),
    .X(_203_));
 sg13g2_nor2_1 _580_ (.A(_177_),
    .B(_182_),
    .Y(_204_));
 sg13g2_a221oi_1 _581_ (.B2(_204_),
    .C1(_199_),
    .B1(_203_),
    .A1(_196_),
    .Y(_205_),
    .A2(_198_));
 sg13g2_and3_1 _582_ (.X(_206_),
    .A(_178_),
    .B(_187_),
    .C(_197_));
 sg13g2_or2_1 _583_ (.X(_207_),
    .B(_140_),
    .A(_135_));
 sg13g2_nor4_1 _584_ (.A(_145_),
    .B(_198_),
    .C(_206_),
    .D(_207_),
    .Y(_208_));
 sg13g2_nand4_1 _585_ (.B(_140_),
    .C(_142_),
    .A(_135_),
    .Y(_209_),
    .D(_144_));
 sg13g2_nor2_1 _586_ (.A(_179_),
    .B(_209_),
    .Y(_210_));
 sg13g2_or3_1 _587_ (.A(_135_),
    .B(_140_),
    .C(_146_),
    .X(_211_));
 sg13g2_nand3_1 _588_ (.B(_140_),
    .C(_148_),
    .A(_136_),
    .Y(_212_));
 sg13g2_a21oi_1 _589_ (.A1(_211_),
    .A2(_212_),
    .Y(_213_),
    .B1(_202_));
 sg13g2_nor4_1 _590_ (.A(_205_),
    .B(_208_),
    .C(_210_),
    .D(_213_),
    .Y(_214_));
 sg13g2_nand3_1 _591_ (.B(_149_),
    .C(_209_),
    .A(_135_),
    .Y(_215_));
 sg13g2_a21oi_1 _592_ (.A1(_111_),
    .A2(_134_),
    .Y(_216_),
    .B1(_110_));
 sg13g2_xnor2_1 _593_ (.Y(_217_),
    .A(\hvsync_gen.hpos[9] ),
    .B(_216_));
 sg13g2_nand2_1 _594_ (.Y(_218_),
    .A(_018_),
    .B(\hvsync_gen.vpos[6] ));
 sg13g2_a21oi_1 _595_ (.A1(_153_),
    .A2(_166_),
    .Y(_219_),
    .B1(_152_));
 sg13g2_a21oi_1 _596_ (.A1(_071_),
    .A2(\hvsync_gen.vpos[8] ),
    .Y(_220_),
    .B1(\hvsync_gen.vpos[9] ));
 sg13g2_nor3_1 _597_ (.A(_069_),
    .B(\hvsync_gen.vpos[7] ),
    .C(_220_),
    .Y(_221_));
 sg13g2_nand2_1 _598_ (.Y(_222_),
    .A(\ty[8] ),
    .B(_072_));
 sg13g2_a22oi_1 _599_ (.Y(_223_),
    .B1(_073_),
    .B2(\ty[7] ),
    .A2(\hvsync_gen.vpos[8] ),
    .A1(_071_));
 sg13g2_a21oi_1 _600_ (.A1(_222_),
    .A2(_223_),
    .Y(_224_),
    .B1(_221_));
 sg13g2_a221oi_1 _601_ (.B2(\hvsync_gen.vpos[9] ),
    .C1(_224_),
    .B1(_222_),
    .A1(_178_),
    .Y(_225_),
    .A2(_182_));
 sg13g2_o21ai_1 _602_ (.B1(_225_),
    .Y(_226_),
    .A1(_218_),
    .A2(_219_));
 sg13g2_nor2b_1 _603_ (.A(_226_),
    .B_N(_188_),
    .Y(_227_));
 sg13g2_nor2_1 _604_ (.A(_018_),
    .B(\hvsync_gen.vpos[6] ),
    .Y(_228_));
 sg13g2_o21ai_1 _605_ (.B1(_220_),
    .Y(_229_),
    .A1(\ty[7] ),
    .A2(_073_));
 sg13g2_o21ai_1 _606_ (.B1(_218_),
    .Y(_230_),
    .A1(_219_),
    .A2(_228_));
 sg13g2_nor2_1 _607_ (.A(_229_),
    .B(_230_),
    .Y(_231_));
 sg13g2_nand2_1 _608_ (.Y(_232_),
    .A(_219_),
    .B(_228_));
 sg13g2_a21oi_1 _609_ (.A1(_229_),
    .A2(_232_),
    .Y(_233_),
    .B1(_231_));
 sg13g2_nand4_1 _610_ (.B(_217_),
    .C(_227_),
    .A(_215_),
    .Y(_234_),
    .D(_233_));
 sg13g2_a21o_2 _611_ (.A2(_214_),
    .A1(_194_),
    .B1(_234_),
    .X(_235_));
 sg13g2_xor2_1 _612_ (.B(\frame_cnt[9] ),
    .A(\frame_cnt[3] ),
    .X(_236_));
 sg13g2_xnor2_1 _613_ (.Y(_237_),
    .A(\hvsync_gen.vpos[3] ),
    .B(\hvsync_gen.hpos[3] ));
 sg13g2_xnor2_1 _614_ (.Y(_238_),
    .A(_236_),
    .B(_237_));
 sg13g2_xnor2_1 _615_ (.Y(_239_),
    .A(\frame_cnt[4] ),
    .B(\frame_cnt[10] ));
 sg13g2_xor2_1 _616_ (.B(\hvsync_gen.hpos[4] ),
    .A(\hvsync_gen.vpos[4] ),
    .X(_240_));
 sg13g2_xnor2_1 _617_ (.Y(_241_),
    .A(_239_),
    .B(_240_));
 sg13g2_xor2_1 _618_ (.B(\hvsync_gen.hpos[1] ),
    .A(\hvsync_gen.vpos[1] ),
    .X(_242_));
 sg13g2_xnor2_1 _619_ (.Y(_243_),
    .A(\frame_cnt[1] ),
    .B(\frame_cnt[7] ));
 sg13g2_xnor2_1 _620_ (.Y(_244_),
    .A(_242_),
    .B(_243_));
 sg13g2_xor2_1 _621_ (.B(\frame_cnt[6] ),
    .A(\hvsync_gen.hpos[0] ),
    .X(_245_));
 sg13g2_xor2_1 _622_ (.B(\hvsync_gen.vpos[0] ),
    .A(\frame_cnt[0] ),
    .X(_246_));
 sg13g2_xnor2_1 _623_ (.Y(_247_),
    .A(_245_),
    .B(_246_));
 sg13g2_xnor2_1 _624_ (.Y(_248_),
    .A(\hvsync_gen.vpos[2] ),
    .B(\hvsync_gen.hpos[2] ));
 sg13g2_xnor2_1 _625_ (.Y(_249_),
    .A(\frame_cnt[8] ),
    .B(\frame_cnt[2] ));
 sg13g2_xor2_1 _626_ (.B(_249_),
    .A(_248_),
    .X(_250_));
 sg13g2_xnor2_1 _627_ (.Y(_251_),
    .A(\hvsync_gen.vpos[5] ),
    .B(net56));
 sg13g2_xnor2_1 _628_ (.Y(_252_),
    .A(\frame_cnt[5] ),
    .B(\frame_cnt[11] ));
 sg13g2_xnor2_1 _629_ (.Y(_253_),
    .A(_251_),
    .B(_252_));
 sg13g2_nor4_1 _630_ (.A(_238_),
    .B(_241_),
    .C(_244_),
    .D(_250_),
    .Y(_254_));
 sg13g2_nand3_1 _631_ (.B(_253_),
    .C(_254_),
    .A(_247_),
    .Y(_255_));
 sg13g2_xor2_1 _632_ (.B(\frame_cnt[13] ),
    .A(\frame_cnt[7] ),
    .X(_256_));
 sg13g2_xnor2_1 _633_ (.Y(_257_),
    .A(_251_),
    .B(_256_));
 sg13g2_xnor2_1 _634_ (.Y(_258_),
    .A(_237_),
    .B(_252_));
 sg13g2_xnor2_1 _635_ (.Y(_259_),
    .A(_236_),
    .B(_242_));
 sg13g2_xor2_1 _636_ (.B(\hvsync_gen.hpos[0] ),
    .A(\hvsync_gen.vpos[0] ),
    .X(_260_));
 sg13g2_xnor2_1 _637_ (.Y(_261_),
    .A(_249_),
    .B(_260_));
 sg13g2_xor2_1 _638_ (.B(_248_),
    .A(_239_),
    .X(_262_));
 sg13g2_xnor2_1 _639_ (.Y(_263_),
    .A(\frame_cnt[6] ),
    .B(\frame_cnt[12] ));
 sg13g2_xnor2_1 _640_ (.Y(_264_),
    .A(_240_),
    .B(_263_));
 sg13g2_nor4_1 _641_ (.A(_257_),
    .B(_261_),
    .C(_262_),
    .D(_264_),
    .Y(_265_));
 sg13g2_nand3_1 _642_ (.B(_259_),
    .C(_265_),
    .A(_258_),
    .Y(_266_));
 sg13g2_inv_1 _643_ (.Y(_267_),
    .A(_266_));
 sg13g2_nand2_1 _644_ (.Y(_268_),
    .A(net4),
    .B(_266_));
 sg13g2_a22oi_1 _645_ (.Y(_269_),
    .B1(_255_),
    .B2(_268_),
    .A2(_080_),
    .A1(net4));
 sg13g2_inv_1 _646_ (.Y(_270_),
    .A(_269_));
 sg13g2_o21ai_1 _647_ (.B1(\hvsync_gen.display_on ),
    .Y(_271_),
    .A1(\frame_cnt[8] ),
    .A2(_235_));
 sg13g2_a21oi_1 _648_ (.A1(_235_),
    .A2(_270_),
    .Y(uo_out[4]),
    .B1(_271_));
 sg13g2_nand2_1 _649_ (.Y(_272_),
    .A(_255_),
    .B(_266_));
 sg13g2_o21ai_1 _650_ (.B1(net3),
    .Y(_273_),
    .A1(_079_),
    .A2(_272_));
 sg13g2_a21oi_1 _651_ (.A1(_235_),
    .A2(_273_),
    .Y(uo_out[0]),
    .B1(_081_));
 sg13g2_and3_1 _652_ (.X(_274_),
    .A(net4),
    .B(_255_),
    .C(_267_));
 sg13g2_nor2_1 _653_ (.A(net4),
    .B(_267_),
    .Y(_275_));
 sg13g2_o21ai_1 _654_ (.B1(_235_),
    .Y(_276_),
    .A1(_274_),
    .A2(_275_));
 sg13g2_and2_1 _655_ (.A(\hvsync_gen.display_on ),
    .B(_276_),
    .X(uo_out[5]));
 sg13g2_o21ai_1 _656_ (.B1(_079_),
    .Y(_277_),
    .A1(_080_),
    .A2(_266_));
 sg13g2_nand2_1 _657_ (.Y(_278_),
    .A(_272_),
    .B(_277_));
 sg13g2_o21ai_1 _658_ (.B1(\hvsync_gen.display_on ),
    .Y(_279_),
    .A1(\frame_cnt[9] ),
    .A2(_235_));
 sg13g2_a21oi_1 _659_ (.A1(_235_),
    .A2(_278_),
    .Y(uo_out[1]),
    .B1(_279_));
 sg13g2_nor3_1 _660_ (.A(net4),
    .B(net3),
    .C(_255_),
    .Y(_280_));
 sg13g2_nand2b_1 _661_ (.Y(_281_),
    .B(\hvsync_gen.vpos[0] ),
    .A_N(net5));
 sg13g2_o21ai_1 _662_ (.B1(_080_),
    .Y(_282_),
    .A1(net4),
    .A2(_281_));
 sg13g2_a21oi_1 _663_ (.A1(net3),
    .A2(_274_),
    .Y(_283_),
    .B1(_280_));
 sg13g2_o21ai_1 _664_ (.B1(_283_),
    .Y(_284_),
    .A1(_267_),
    .A2(_282_));
 sg13g2_a21oi_1 _665_ (.A1(_235_),
    .A2(_284_),
    .Y(uo_out[6]),
    .B1(_081_));
 sg13g2_nand4_1 _666_ (.B(_080_),
    .C(\hvsync_gen.display_on ),
    .A(_079_),
    .Y(_285_),
    .D(_272_));
 sg13g2_nand2b_1 _667_ (.Y(uo_out[2]),
    .B(_285_),
    .A_N(uo_out[0]));
 sg13g2_and2_1 _668_ (.A(net106),
    .B(net48),
    .X(_286_));
 sg13g2_nor3_1 _669_ (.A(\hvsync_gen.vpos[5] ),
    .B(net95),
    .C(net141),
    .Y(_287_));
 sg13g2_nand2_1 _670_ (.Y(_288_),
    .A(net86),
    .B(net105));
 sg13g2_nand4_1 _671_ (.B(_073_),
    .C(_287_),
    .A(_072_),
    .Y(_289_),
    .D(_288_));
 sg13g2_nand2_2 _672_ (.Y(_290_),
    .A(net44),
    .B(_289_));
 sg13g2_nor3_2 _673_ (.A(_090_),
    .B(_096_),
    .C(_290_),
    .Y(_291_));
 sg13g2_a21oi_1 _674_ (.A1(net48),
    .A2(_290_),
    .Y(_292_),
    .B1(net106));
 sg13g2_nor2_1 _675_ (.A(_286_),
    .B(_292_),
    .Y(_019_));
 sg13g2_and2_1 _676_ (.A(net102),
    .B(_286_),
    .X(_293_));
 sg13g2_nor2_1 _677_ (.A(net102),
    .B(_286_),
    .Y(_294_));
 sg13g2_nor3_1 _678_ (.A(_291_),
    .B(_293_),
    .C(_294_),
    .Y(_020_));
 sg13g2_xnor2_1 _679_ (.Y(_295_),
    .A(net105),
    .B(_293_));
 sg13g2_nor2_1 _680_ (.A(_291_),
    .B(_295_),
    .Y(_021_));
 sg13g2_a21oi_1 _681_ (.A1(net105),
    .A2(_293_),
    .Y(_296_),
    .B1(net86));
 sg13g2_nor2b_1 _682_ (.A(_288_),
    .B_N(_293_),
    .Y(_297_));
 sg13g2_nor3_1 _683_ (.A(_291_),
    .B(_296_),
    .C(_297_),
    .Y(_022_));
 sg13g2_and2_1 _684_ (.A(net130),
    .B(_297_),
    .X(_298_));
 sg13g2_nor2_1 _685_ (.A(net130),
    .B(_297_),
    .Y(_299_));
 sg13g2_nor3_1 _686_ (.A(_291_),
    .B(_298_),
    .C(_299_),
    .Y(_023_));
 sg13g2_xnor2_1 _687_ (.Y(_300_),
    .A(net133),
    .B(_298_));
 sg13g2_nor2_1 _688_ (.A(_291_),
    .B(_300_),
    .Y(_024_));
 sg13g2_a21oi_1 _689_ (.A1(\hvsync_gen.vpos[5] ),
    .A2(_298_),
    .Y(_301_),
    .B1(net95));
 sg13g2_nand3_1 _690_ (.B(net102),
    .C(\hvsync_gen.vpos[0] ),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_302_));
 sg13g2_nor3_1 _691_ (.A(_084_),
    .B(_288_),
    .C(net103),
    .Y(_303_));
 sg13g2_a21o_1 _692_ (.A2(_303_),
    .A1(net48),
    .B1(_291_),
    .X(_304_));
 sg13g2_nor2_1 _693_ (.A(net96),
    .B(_304_),
    .Y(_025_));
 sg13g2_nand4_1 _694_ (.B(net48),
    .C(_290_),
    .A(_073_),
    .Y(_305_),
    .D(net104));
 sg13g2_o21ai_1 _695_ (.B1(_305_),
    .Y(_026_),
    .A1(_073_),
    .A2(_304_));
 sg13g2_nand4_1 _696_ (.B(\hvsync_gen.vpos[5] ),
    .C(net95),
    .A(net80),
    .Y(_306_),
    .D(_298_));
 sg13g2_a221oi_1 _697_ (.B2(_072_),
    .C1(_291_),
    .B1(_306_),
    .A1(net81),
    .Y(_027_),
    .A2(_298_));
 sg13g2_a21oi_1 _698_ (.A1(net81),
    .A2(_298_),
    .Y(_307_),
    .B1(net44));
 sg13g2_nor2_1 _699_ (.A(_291_),
    .B(net82),
    .Y(_028_));
 sg13g2_nor2b_1 _700_ (.A(net2),
    .B_N(net1),
    .Y(_308_));
 sg13g2_nand2b_2 _701_ (.Y(_309_),
    .B(net1),
    .A_N(net2));
 sg13g2_nor2b_2 _702_ (.A(net137),
    .B_N(net22),
    .Y(_310_));
 sg13g2_nand2_1 _703_ (.Y(_311_),
    .A(_309_),
    .B(_310_));
 sg13g2_xnor2_1 _704_ (.Y(_029_),
    .A(net40),
    .B(_311_));
 sg13g2_o21ai_1 _705_ (.B1(_310_),
    .Y(_312_),
    .A1(net40),
    .A2(_308_));
 sg13g2_nor2_1 _706_ (.A(_077_),
    .B(_312_),
    .Y(_313_));
 sg13g2_xnor2_1 _707_ (.Y(_030_),
    .A(net75),
    .B(_312_));
 sg13g2_and2_1 _708_ (.A(net23),
    .B(_313_),
    .X(_314_));
 sg13g2_xor2_1 _709_ (.B(_313_),
    .A(net23),
    .X(_031_));
 sg13g2_xor2_1 _710_ (.B(_314_),
    .A(net33),
    .X(_032_));
 sg13g2_and3_2 _711_ (.X(_315_),
    .A(net33),
    .B(net70),
    .C(_314_));
 sg13g2_a21oi_1 _712_ (.A1(net33),
    .A2(_314_),
    .Y(_316_),
    .B1(net70));
 sg13g2_nor2_1 _713_ (.A(_315_),
    .B(_316_),
    .Y(_033_));
 sg13g2_xor2_1 _714_ (.B(_315_),
    .A(net29),
    .X(_034_));
 sg13g2_nand3_1 _715_ (.B(net29),
    .C(_315_),
    .A(net140),
    .Y(_317_));
 sg13g2_a21o_1 _716_ (.A2(_315_),
    .A1(net29),
    .B1(net140),
    .X(_318_));
 sg13g2_and2_1 _717_ (.A(_317_),
    .B(_318_),
    .X(_035_));
 sg13g2_nor2_1 _718_ (.A(_078_),
    .B(_317_),
    .Y(_319_));
 sg13g2_xnor2_1 _719_ (.Y(_036_),
    .A(net46),
    .B(_317_));
 sg13g2_and2_1 _720_ (.A(net42),
    .B(_319_),
    .X(_320_));
 sg13g2_xor2_1 _721_ (.B(_319_),
    .A(net42),
    .X(_037_));
 sg13g2_xor2_1 _722_ (.B(_320_),
    .A(net73),
    .X(_038_));
 sg13g2_and3_2 _723_ (.X(_321_),
    .A(\frame_cnt[9] ),
    .B(net37),
    .C(_320_));
 sg13g2_a21oi_1 _724_ (.A1(\frame_cnt[9] ),
    .A2(_320_),
    .Y(_322_),
    .B1(net37));
 sg13g2_nor2_1 _725_ (.A(_321_),
    .B(net38),
    .Y(_039_));
 sg13g2_xor2_1 _726_ (.B(_321_),
    .A(net27),
    .X(_040_));
 sg13g2_nand3_1 _727_ (.B(net134),
    .C(_321_),
    .A(net27),
    .Y(_323_));
 sg13g2_a21o_1 _728_ (.A2(_321_),
    .A1(net27),
    .B1(net134),
    .X(_324_));
 sg13g2_and2_1 _729_ (.A(_323_),
    .B(net135),
    .X(_041_));
 sg13g2_xnor2_1 _730_ (.Y(_042_),
    .A(net25),
    .B(_323_));
 sg13g2_o21ai_1 _731_ (.B1(net2),
    .Y(_325_),
    .A1(net1),
    .A2(_067_));
 sg13g2_and2_1 _732_ (.A(_310_),
    .B(_325_),
    .X(_326_));
 sg13g2_nand2_2 _733_ (.Y(_327_),
    .A(_310_),
    .B(_325_));
 sg13g2_nor2_1 _734_ (.A(net1),
    .B(_327_),
    .Y(_328_));
 sg13g2_xor2_1 _735_ (.B(_328_),
    .A(net71),
    .X(_043_));
 sg13g2_nand2b_1 _736_ (.Y(_329_),
    .B(_309_),
    .A_N(net71));
 sg13g2_and3_1 _737_ (.X(_330_),
    .A(net107),
    .B(net58),
    .C(_309_));
 sg13g2_a21oi_1 _738_ (.A1(net58),
    .A2(_309_),
    .Y(_331_),
    .B1(net107));
 sg13g2_or2_1 _739_ (.X(_332_),
    .B(_331_),
    .A(_330_));
 sg13g2_nor2b_1 _740_ (.A(_332_),
    .B_N(_329_),
    .Y(_333_));
 sg13g2_xnor2_1 _741_ (.Y(_334_),
    .A(_329_),
    .B(_332_));
 sg13g2_mux2_1 _742_ (.A0(net107),
    .A1(_334_),
    .S(net52),
    .X(_044_));
 sg13g2_nand2_1 _743_ (.Y(_335_),
    .A(_065_),
    .B(net58));
 sg13g2_xnor2_1 _744_ (.Y(_336_),
    .A(net114),
    .B(net58));
 sg13g2_o21ai_1 _745_ (.B1(_336_),
    .Y(_337_),
    .A1(_330_),
    .A2(_333_));
 sg13g2_nor3_1 _746_ (.A(_330_),
    .B(_333_),
    .C(_336_),
    .Y(_338_));
 sg13g2_nor2_1 _747_ (.A(net49),
    .B(_338_),
    .Y(_339_));
 sg13g2_a22oi_1 _748_ (.Y(_045_),
    .B1(_337_),
    .B2(_339_),
    .A2(net49),
    .A1(_065_));
 sg13g2_and2_1 _749_ (.A(_335_),
    .B(_337_),
    .X(_340_));
 sg13g2_nand2_1 _750_ (.Y(_341_),
    .A(_066_),
    .B(_083_));
 sg13g2_xnor2_1 _751_ (.Y(_342_),
    .A(net128),
    .B(net58));
 sg13g2_a21oi_1 _752_ (.A1(_340_),
    .A2(_342_),
    .Y(_343_),
    .B1(net49));
 sg13g2_o21ai_1 _753_ (.B1(_343_),
    .Y(_344_),
    .A1(_340_),
    .A2(_342_));
 sg13g2_o21ai_1 _754_ (.B1(_344_),
    .Y(_046_),
    .A1(_066_),
    .A2(net52));
 sg13g2_nand2_1 _755_ (.Y(_345_),
    .A(\tx[4] ),
    .B(net57));
 sg13g2_or2_1 _756_ (.X(_346_),
    .B(net57),
    .A(\tx[4] ));
 sg13g2_o21ai_1 _757_ (.B1(_340_),
    .Y(_347_),
    .A1(_066_),
    .A2(_083_));
 sg13g2_and4_1 _758_ (.A(_341_),
    .B(_345_),
    .C(_346_),
    .D(_347_),
    .X(_348_));
 sg13g2_a22oi_1 _759_ (.Y(_349_),
    .B1(_347_),
    .B2(_341_),
    .A2(_346_),
    .A1(_345_));
 sg13g2_nor3_1 _760_ (.A(net49),
    .B(_348_),
    .C(_349_),
    .Y(_350_));
 sg13g2_a21o_1 _761_ (.A2(net49),
    .A1(net122),
    .B1(_350_),
    .X(_047_));
 sg13g2_xnor2_1 _762_ (.Y(_351_),
    .A(net117),
    .B(net57));
 sg13g2_a21oi_1 _763_ (.A1(\tx[4] ),
    .A2(net57),
    .Y(_352_),
    .B1(_348_));
 sg13g2_xnor2_1 _764_ (.Y(_353_),
    .A(_351_),
    .B(_352_));
 sg13g2_nor2_1 _765_ (.A(net117),
    .B(net52),
    .Y(_354_));
 sg13g2_a21oi_1 _766_ (.A1(net52),
    .A2(_353_),
    .Y(_048_),
    .B1(_354_));
 sg13g2_xnor2_1 _767_ (.Y(_355_),
    .A(net84),
    .B(net57));
 sg13g2_and2_1 _768_ (.A(_348_),
    .B(_351_),
    .X(_356_));
 sg13g2_o21ai_1 _769_ (.B1(_345_),
    .Y(_357_),
    .A1(_014_),
    .A2(_083_));
 sg13g2_or3_1 _770_ (.A(_355_),
    .B(_356_),
    .C(_357_),
    .X(_358_));
 sg13g2_o21ai_1 _771_ (.B1(_355_),
    .Y(_359_),
    .A1(_356_),
    .A2(_357_));
 sg13g2_and2_1 _772_ (.A(net52),
    .B(_359_),
    .X(_360_));
 sg13g2_a22oi_1 _773_ (.Y(_049_),
    .B1(_358_),
    .B2(_360_),
    .A2(net49),
    .A1(_063_));
 sg13g2_xor2_1 _774_ (.B(net57),
    .A(net116),
    .X(_361_));
 sg13g2_o21ai_1 _775_ (.B1(_359_),
    .Y(_362_),
    .A1(net84),
    .A2(_083_));
 sg13g2_xnor2_1 _776_ (.Y(_363_),
    .A(_361_),
    .B(_362_));
 sg13g2_nor2_1 _777_ (.A(net116),
    .B(net52),
    .Y(_364_));
 sg13g2_a21oi_1 _778_ (.A1(net52),
    .A2(_363_),
    .Y(_050_),
    .B1(_364_));
 sg13g2_nor4_1 _779_ (.A(_063_),
    .B(\tx[7] ),
    .C(_083_),
    .D(_357_),
    .Y(_365_));
 sg13g2_and3_1 _780_ (.X(_366_),
    .A(_355_),
    .B(_356_),
    .C(_361_));
 sg13g2_a21oi_1 _781_ (.A1(net57),
    .A2(_366_),
    .Y(_367_),
    .B1(net49));
 sg13g2_o21ai_1 _782_ (.B1(_367_),
    .Y(_368_),
    .A1(_365_),
    .A2(_366_));
 sg13g2_xnor2_1 _783_ (.Y(_051_),
    .A(net78),
    .B(_368_));
 sg13g2_xor2_1 _784_ (.B(_328_),
    .A(net31),
    .X(_052_));
 sg13g2_nor2_1 _785_ (.A(net97),
    .B(net50),
    .Y(_369_));
 sg13g2_nor2_1 _786_ (.A(net31),
    .B(_308_),
    .Y(_370_));
 sg13g2_nand3_1 _787_ (.B(net53),
    .C(_309_),
    .A(net97),
    .Y(_371_));
 sg13g2_a21o_1 _788_ (.A2(_309_),
    .A1(net54),
    .B1(net97),
    .X(_372_));
 sg13g2_nand2_1 _789_ (.Y(_373_),
    .A(_371_),
    .B(_372_));
 sg13g2_xnor2_1 _790_ (.Y(_374_),
    .A(_370_),
    .B(_373_));
 sg13g2_a21oi_1 _791_ (.A1(net50),
    .A2(_374_),
    .Y(_053_),
    .B1(_369_));
 sg13g2_nor2_1 _792_ (.A(net126),
    .B(_082_),
    .Y(_375_));
 sg13g2_nand2_1 _793_ (.Y(_376_),
    .A(_016_),
    .B(_082_));
 sg13g2_nor2b_1 _794_ (.A(_375_),
    .B_N(_376_),
    .Y(_377_));
 sg13g2_o21ai_1 _795_ (.B1(_371_),
    .Y(_378_),
    .A1(_370_),
    .A2(_373_));
 sg13g2_xnor2_1 _796_ (.Y(_379_),
    .A(_377_),
    .B(_378_));
 sg13g2_mux2_1 _797_ (.A0(net126),
    .A1(_379_),
    .S(net51),
    .X(_054_));
 sg13g2_a21oi_1 _798_ (.A1(_376_),
    .A2(_378_),
    .Y(_380_),
    .B1(_375_));
 sg13g2_xnor2_1 _799_ (.Y(_381_),
    .A(net139),
    .B(net53));
 sg13g2_a21oi_1 _800_ (.A1(_380_),
    .A2(_381_),
    .Y(_382_),
    .B1(_327_));
 sg13g2_o21ai_1 _801_ (.B1(_382_),
    .Y(_383_),
    .A1(_380_),
    .A2(_381_));
 sg13g2_o21ai_1 _802_ (.B1(_383_),
    .Y(_055_),
    .A1(_068_),
    .A2(net50));
 sg13g2_nor2_1 _803_ (.A(net110),
    .B(net50),
    .Y(_384_));
 sg13g2_xnor2_1 _804_ (.Y(_385_),
    .A(net110),
    .B(net54));
 sg13g2_o21ai_1 _805_ (.B1(_380_),
    .Y(_386_),
    .A1(_068_),
    .A2(_082_));
 sg13g2_o21ai_1 _806_ (.B1(_386_),
    .Y(_387_),
    .A1(\ty[3] ),
    .A2(net54));
 sg13g2_nor2_1 _807_ (.A(_385_),
    .B(_387_),
    .Y(_388_));
 sg13g2_xnor2_1 _808_ (.Y(_389_),
    .A(_385_),
    .B(_387_));
 sg13g2_a21oi_1 _809_ (.A1(net50),
    .A2(_389_),
    .Y(_056_),
    .B1(_384_));
 sg13g2_xnor2_1 _810_ (.Y(_390_),
    .A(net112),
    .B(net53));
 sg13g2_a21oi_1 _811_ (.A1(net110),
    .A2(net53),
    .Y(_391_),
    .B1(_388_));
 sg13g2_xnor2_1 _812_ (.Y(_392_),
    .A(_390_),
    .B(_391_));
 sg13g2_nor2_1 _813_ (.A(net112),
    .B(net50),
    .Y(_393_));
 sg13g2_a21oi_1 _814_ (.A1(net50),
    .A2(_392_),
    .Y(_057_),
    .B1(_393_));
 sg13g2_nor2_1 _815_ (.A(net108),
    .B(net51),
    .Y(_394_));
 sg13g2_nand2b_1 _816_ (.Y(_395_),
    .B(net53),
    .A_N(net108));
 sg13g2_xor2_1 _817_ (.B(net53),
    .A(net108),
    .X(_396_));
 sg13g2_and2_1 _818_ (.A(_388_),
    .B(_390_),
    .X(_397_));
 sg13g2_a21oi_1 _819_ (.A1(_017_),
    .A2(_070_),
    .Y(_398_),
    .B1(_082_));
 sg13g2_nor2_1 _820_ (.A(_397_),
    .B(net113),
    .Y(_399_));
 sg13g2_xor2_1 _821_ (.B(_399_),
    .A(_396_),
    .X(_400_));
 sg13g2_a21oi_1 _822_ (.A1(net51),
    .A2(_400_),
    .Y(_058_),
    .B1(_394_));
 sg13g2_xor2_1 _823_ (.B(net53),
    .A(net100),
    .X(_401_));
 sg13g2_o21ai_1 _824_ (.B1(_395_),
    .Y(_402_),
    .A1(_396_),
    .A2(_399_));
 sg13g2_xnor2_1 _825_ (.Y(_403_),
    .A(_401_),
    .B(_402_));
 sg13g2_nor2_1 _826_ (.A(net100),
    .B(net51),
    .Y(_404_));
 sg13g2_a21oi_1 _827_ (.A1(net51),
    .A2(net109),
    .Y(_059_),
    .B1(_404_));
 sg13g2_nor2b_1 _828_ (.A(_396_),
    .B_N(_401_),
    .Y(_405_));
 sg13g2_a21oi_1 _829_ (.A1(_018_),
    .A2(_069_),
    .Y(_406_),
    .B1(_082_));
 sg13g2_a21o_1 _830_ (.A2(_405_),
    .A1(_397_),
    .B1(_406_),
    .X(_407_));
 sg13g2_o21ai_1 _831_ (.B1(net53),
    .Y(_408_),
    .A1(_398_),
    .A2(_407_));
 sg13g2_nand2b_1 _832_ (.Y(_409_),
    .B(_082_),
    .A_N(_407_));
 sg13g2_nand3_1 _833_ (.B(_408_),
    .C(_409_),
    .A(net51),
    .Y(_410_));
 sg13g2_xnor2_1 _834_ (.Y(_060_),
    .A(net35),
    .B(_410_));
 sg13g2_nand2_1 _835_ (.Y(_411_),
    .A(net78),
    .B(net52));
 sg13g2_nand2_1 _836_ (.Y(_412_),
    .A(\tx[0] ),
    .B(\tx[1] ));
 sg13g2_a21oi_1 _837_ (.A1(_013_),
    .A2(_412_),
    .Y(_413_),
    .B1(_066_));
 sg13g2_nor4_1 _838_ (.A(\tx[4] ),
    .B(net78),
    .C(net49),
    .D(_413_),
    .Y(_414_));
 sg13g2_nand2_1 _839_ (.Y(_415_),
    .A(_341_),
    .B(_346_));
 sg13g2_nor2_1 _840_ (.A(_414_),
    .B(_415_),
    .Y(_416_));
 sg13g2_nor3_1 _841_ (.A(_064_),
    .B(\tx[7] ),
    .C(_416_),
    .Y(_417_));
 sg13g2_a22oi_1 _842_ (.Y(_061_),
    .B1(_417_),
    .B2(net84),
    .A2(_411_),
    .A1(_083_));
 sg13g2_nand4_1 _843_ (.B(_069_),
    .C(_071_),
    .A(_017_),
    .Y(_418_),
    .D(net50));
 sg13g2_o21ai_1 _844_ (.B1(_418_),
    .Y(_419_),
    .A1(\ty[3] ),
    .A2(_376_));
 sg13g2_nand2_1 _845_ (.Y(_420_),
    .A(\ty[0] ),
    .B(\ty[1] ));
 sg13g2_a21oi_1 _846_ (.A1(_016_),
    .A2(_420_),
    .Y(_421_),
    .B1(_068_));
 sg13g2_nor2_1 _847_ (.A(\ty[4] ),
    .B(_421_),
    .Y(_422_));
 sg13g2_a22oi_1 _848_ (.Y(_423_),
    .B1(_419_),
    .B2(_422_),
    .A2(_082_),
    .A1(_017_));
 sg13g2_nor2b_1 _849_ (.A(_423_),
    .B_N(_018_),
    .Y(_424_));
 sg13g2_nand3_1 _850_ (.B(net35),
    .C(net51),
    .A(net100),
    .Y(_425_));
 sg13g2_a21oi_1 _851_ (.A1(_082_),
    .A2(_425_),
    .Y(_062_),
    .B1(_424_));
 sg13g2_dfrbpq_2 _852_ (.RESET_B(net64),
    .D(_019_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _853_ (.RESET_B(net64),
    .D(_020_),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _854_ (.RESET_B(net64),
    .D(_021_),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _855_ (.RESET_B(net64),
    .D(_022_),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _856_ (.RESET_B(net64),
    .D(_023_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _857_ (.RESET_B(net64),
    .D(_024_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _858_ (.RESET_B(net67),
    .D(_025_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _859_ (.RESET_B(net67),
    .D(_026_),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _860_ (.RESET_B(net67),
    .D(net99),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _861_ (.RESET_B(net64),
    .D(net83),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _862_ (.RESET_B(net65),
    .D(net41),
    .Q(\frame_cnt[0] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _863_ (.RESET_B(net65),
    .D(net76),
    .Q(\frame_cnt[1] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _864_ (.RESET_B(net64),
    .D(net24),
    .Q(\frame_cnt[2] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _865_ (.RESET_B(net63),
    .D(net34),
    .Q(\frame_cnt[3] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _866_ (.RESET_B(net63),
    .D(_033_),
    .Q(\frame_cnt[4] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _867_ (.RESET_B(net62),
    .D(net30),
    .Q(\frame_cnt[5] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _868_ (.RESET_B(net62),
    .D(_035_),
    .Q(\frame_cnt[6] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _869_ (.RESET_B(net63),
    .D(net69),
    .Q(\frame_cnt[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _870_ (.RESET_B(net62),
    .D(net43),
    .Q(\frame_cnt[8] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _871_ (.RESET_B(net62),
    .D(net74),
    .Q(\frame_cnt[9] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _872_ (.RESET_B(net61),
    .D(net39),
    .Q(\frame_cnt[10] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _873_ (.RESET_B(net61),
    .D(net28),
    .Q(\frame_cnt[11] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _874_ (.RESET_B(net62),
    .D(net136),
    .Q(\frame_cnt[12] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _875_ (.RESET_B(net61),
    .D(net26),
    .Q(\frame_cnt[13] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _876_ (.RESET_B(net66),
    .D(net72),
    .Q(\tx[0] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _877_ (.RESET_B(net63),
    .D(_044_),
    .Q(\tx[1] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _878_ (.RESET_B(net60),
    .D(net115),
    .Q(_013_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _879_ (.RESET_B(net60),
    .D(net129),
    .Q(\tx[3] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _880_ (.RESET_B(net59),
    .D(net123),
    .Q(\tx[4] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _881_ (.RESET_B(net60),
    .D(net118),
    .Q(_014_),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _882_ (.RESET_B(net59),
    .D(net138),
    .Q(_015_),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _883_ (.RESET_B(net60),
    .D(_050_),
    .Q(\tx[7] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _884_ (.RESET_B(net59),
    .D(net79),
    .Q(\tx[8] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _885_ (.RESET_B(net65),
    .D(net32),
    .Q(\ty[0] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _886_ (.RESET_B(net65),
    .D(_053_),
    .Q(\ty[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _887_ (.RESET_B(net65),
    .D(_054_),
    .Q(_016_),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _888_ (.RESET_B(net65),
    .D(_055_),
    .Q(\ty[3] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _889_ (.RESET_B(net65),
    .D(net111),
    .Q(\ty[4] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _890_ (.RESET_B(net67),
    .D(_057_),
    .Q(_017_),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _891_ (.RESET_B(net67),
    .D(_058_),
    .Q(_018_),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _892_ (.RESET_B(net67),
    .D(_059_),
    .Q(\ty[7] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _893_ (.RESET_B(net67),
    .D(net36),
    .Q(\ty[8] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _894_ (.RESET_B(net60),
    .D(net85),
    .Q(x_dir),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _895_ (.RESET_B(net65),
    .D(net22),
    .Q(vsync_prev),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _896_ (.RESET_B(net61),
    .D(_001_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _897_ (.RESET_B(net61),
    .D(_002_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _898_ (.RESET_B(net63),
    .D(net90),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _899_ (.RESET_B(net61),
    .D(_004_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _900_ (.RESET_B(net61),
    .D(_005_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _901_ (.RESET_B(net59),
    .D(_006_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _902_ (.RESET_B(net59),
    .D(_007_),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _903_ (.RESET_B(net59),
    .D(_008_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _904_ (.RESET_B(net59),
    .D(_009_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _905_ (.RESET_B(net59),
    .D(_010_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _906_ (.RESET_B(net66),
    .D(net87),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _907_ (.RESET_B(net66),
    .D(net45),
    .Q(\hvsync_gen.display_on ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _908_ (.RESET_B(net61),
    .D(net92),
    .Q(hsync),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _909_ (.RESET_B(net67),
    .D(net101),
    .Q(y_dir),
    .CLK(clknet_4_11_0_clk));
 sg13g2_tielo tt_um_embeddedinn_vga_7 (.L_LO(net7));
 sg13g2_tielo tt_um_embeddedinn_vga_8 (.L_LO(net8));
 sg13g2_tielo tt_um_embeddedinn_vga_9 (.L_LO(net9));
 sg13g2_tielo tt_um_embeddedinn_vga_10 (.L_LO(net10));
 sg13g2_tielo tt_um_embeddedinn_vga_11 (.L_LO(net11));
 sg13g2_tielo tt_um_embeddedinn_vga_12 (.L_LO(net12));
 sg13g2_tielo tt_um_embeddedinn_vga_13 (.L_LO(net13));
 sg13g2_tielo tt_um_embeddedinn_vga_14 (.L_LO(net14));
 sg13g2_tielo tt_um_embeddedinn_vga_15 (.L_LO(net15));
 sg13g2_tielo tt_um_embeddedinn_vga_16 (.L_LO(net16));
 sg13g2_tielo tt_um_embeddedinn_vga_17 (.L_LO(net17));
 sg13g2_tielo tt_um_embeddedinn_vga_18 (.L_LO(net18));
 sg13g2_tielo tt_um_embeddedinn_vga_19 (.L_LO(net19));
 sg13g2_tielo tt_um_embeddedinn_vga_20 (.L_LO(net20));
 sg13g2_tielo tt_um_embeddedinn_vga_21 (.L_LO(net21));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _926_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _927_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_8 fanout48 (.A(_097_),
    .X(net48));
 sg13g2_buf_8 fanout49 (.A(_327_),
    .X(net49));
 sg13g2_buf_8 fanout50 (.A(net51),
    .X(net50));
 sg13g2_buf_8 fanout51 (.A(_326_),
    .X(net51));
 sg13g2_buf_8 fanout52 (.A(_326_),
    .X(net52));
 sg13g2_buf_8 fanout53 (.A(net124),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(y_dir),
    .X(net54));
 sg13g2_buf_8 fanout55 (.A(net132),
    .X(net55));
 sg13g2_buf_8 fanout56 (.A(net131),
    .X(net56));
 sg13g2_buf_8 fanout57 (.A(x_dir),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(x_dir),
    .X(net58));
 sg13g2_buf_8 fanout59 (.A(net68),
    .X(net59));
 sg13g2_buf_8 fanout60 (.A(net68),
    .X(net60));
 sg13g2_buf_8 fanout61 (.A(net63),
    .X(net61));
 sg13g2_buf_8 fanout62 (.A(net63),
    .X(net62));
 sg13g2_buf_8 fanout63 (.A(net68),
    .X(net63));
 sg13g2_buf_8 fanout64 (.A(net66),
    .X(net64));
 sg13g2_buf_8 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_8 fanout66 (.A(net68),
    .X(net66));
 sg13g2_buf_8 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_8 fanout68 (.A(rst_n),
    .X(net68));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_tielo tt_um_embeddedinn_vga_6 (.L_LO(net6));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.vsync ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold2 (.A(\frame_cnt[2] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold3 (.A(_031_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold4 (.A(\frame_cnt[13] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold5 (.A(_042_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold6 (.A(\frame_cnt[11] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold7 (.A(_040_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold8 (.A(\frame_cnt[5] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold9 (.A(_034_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ty[0] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold11 (.A(_052_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold12 (.A(\frame_cnt[3] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold13 (.A(_032_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ty[8] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold15 (.A(_060_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold16 (.A(\frame_cnt[10] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold17 (.A(_322_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold18 (.A(_039_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold19 (.A(\frame_cnt[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold20 (.A(_029_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold21 (.A(\frame_cnt[8] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold22 (.A(_037_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.vpos[9] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold24 (.A(_000_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold25 (.A(\frame_cnt[7] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold26 (.A(_036_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold27 (.A(\frame_cnt[4] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold28 (.A(\tx[0] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold29 (.A(_043_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold30 (.A(\frame_cnt[9] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold31 (.A(_038_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold32 (.A(\frame_cnt[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold33 (.A(_030_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.hpos[0] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold35 (.A(\tx[8] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold36 (.A(_051_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold37 (.A(\hvsync_gen.vpos[7] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold38 (.A(_085_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold39 (.A(_307_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold40 (.A(_028_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold41 (.A(_015_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold42 (.A(_061_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hvsync_gen.vpos[3] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold44 (.A(_012_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hvsync_gen.hpos[2] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold46 (.A(_099_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold47 (.A(_003_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hvsync_gen.hpos[9] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold49 (.A(_011_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hvsync_gen.hpos[8] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold51 (.A(_109_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold52 (.A(\hvsync_gen.vpos[6] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold53 (.A(_301_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ty[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold55 (.A(\hvsync_gen.vpos[8] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold56 (.A(_027_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ty[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold58 (.A(_062_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold59 (.A(\hvsync_gen.vpos[1] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold60 (.A(_302_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold61 (.A(_303_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hvsync_gen.vpos[2] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold63 (.A(\hvsync_gen.vpos[0] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold64 (.A(\tx[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold65 (.A(_018_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold66 (.A(_403_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ty[4] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold68 (.A(_056_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold69 (.A(_017_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold70 (.A(_398_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold71 (.A(_013_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold72 (.A(_045_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold73 (.A(\tx[7] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold74 (.A(_014_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold75 (.A(_048_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold76 (.A(\hvsync_gen.hpos[6] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold77 (.A(\hvsync_gen.hpos[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold78 (.A(_100_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold79 (.A(\tx[4] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold80 (.A(_047_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold81 (.A(y_dir),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold82 (.A(\hvsync_gen.hpos[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold83 (.A(_016_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold84 (.A(\hvsync_gen.hpos[4] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold85 (.A(\tx[3] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold86 (.A(_046_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold87 (.A(\hvsync_gen.vpos[4] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold88 (.A(\hvsync_gen.hpos[5] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold89 (.A(\hvsync_gen.hpos[7] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold90 (.A(\hvsync_gen.vpos[5] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold91 (.A(\frame_cnt[12] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold92 (.A(_324_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold93 (.A(_041_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold94 (.A(vsync_prev),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold95 (.A(_049_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ty[3] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold97 (.A(\frame_cnt[6] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold98 (.A(\hvsync_gen.vpos[4] ),
    .X(net141));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_170 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_166 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_114 ();
 sg13g2_decap_4 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_95 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_decap_4 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_4 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_decap_4 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_4 FILLER_21_245 ();
 sg13g2_fill_2 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_4 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_decap_4 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_4 FILLER_22_293 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_decap_4 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_117 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_decap_4 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_209 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_386 ();
 sg13g2_fill_1 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_378 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_227 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_4 FILLER_26_305 ();
 sg13g2_decap_4 FILLER_26_322 ();
 sg13g2_decap_4 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_167 ();
 sg13g2_decap_4 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_4 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_2 FILLER_28_291 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_192 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_decap_4 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_157 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_decap_4 FILLER_31_189 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_decap_4 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_381 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_decap_4 FILLER_32_393 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_decap_4 FILLER_33_66 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_decap_4 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_decap_4 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_decap_4 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_decap_4 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_4 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_decap_4 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_2 FILLER_37_73 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_decap_4 FILLER_37_238 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_82 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_decap_4 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_366 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
