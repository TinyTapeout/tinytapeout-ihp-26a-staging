module tt_um_herald (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire clknet_leaf_0_clk;
 wire \byte_counter[0] ;
 wire \byte_counter[1] ;
 wire \byte_counter[2] ;
 wire \cmd_reg[0] ;
 wire \cmd_reg[1] ;
 wire \cmd_reg[2] ;
 wire \cmd_reg[3] ;
 wire \cmd_reg[4] ;
 wire \cmd_reg[5] ;
 wire \cmd_reg[6] ;
 wire \cmd_reg[7] ;
 wire \cordic_atan2_result[0] ;
 wire \cordic_atan2_result[10] ;
 wire \cordic_atan2_result[11] ;
 wire \cordic_atan2_result[12] ;
 wire \cordic_atan2_result[13] ;
 wire \cordic_atan2_result[14] ;
 wire \cordic_atan2_result[15] ;
 wire \cordic_atan2_result[16] ;
 wire \cordic_atan2_result[17] ;
 wire \cordic_atan2_result[18] ;
 wire \cordic_atan2_result[19] ;
 wire \cordic_atan2_result[1] ;
 wire \cordic_atan2_result[20] ;
 wire \cordic_atan2_result[21] ;
 wire \cordic_atan2_result[22] ;
 wire \cordic_atan2_result[23] ;
 wire \cordic_atan2_result[2] ;
 wire \cordic_atan2_result[3] ;
 wire \cordic_atan2_result[4] ;
 wire \cordic_atan2_result[5] ;
 wire \cordic_atan2_result[6] ;
 wire \cordic_atan2_result[7] ;
 wire \cordic_atan2_result[8] ;
 wire \cordic_atan2_result[9] ;
 wire cordic_busy;
 wire cordic_en_atan2;
 wire cordic_en_get_atan2;
 wire cordic_en_get_sin_cos;
 wire cordic_en_get_sqrt;
 wire cordic_en_sin_cos;
 wire cordic_en_sqrt;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ;
 wire \cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ;
 wire \cordic_inst.cordic_state[0] ;
 wire \cordic_inst.cordic_state[32] ;
 wire \cordic_inst.cordic_state[33] ;
 wire \cordic_inst.cordic_state[34] ;
 wire \cordic_inst.cordic_state[35] ;
 wire \cordic_inst.cordic_state[36] ;
 wire \cordic_inst.cordic_state[37] ;
 wire \cordic_inst.cordic_state[38] ;
 wire \cordic_inst.cordic_state[39] ;
 wire \cordic_inst.cordic_state[3] ;
 wire \cordic_inst.cordic_state[40] ;
 wire \cordic_inst.cordic_state[41] ;
 wire \cordic_inst.cordic_state[42] ;
 wire \cordic_inst.cordic_state[43] ;
 wire \cordic_inst.cordic_state[44] ;
 wire \cordic_inst.cordic_state[45] ;
 wire \cordic_inst.cordic_state[46] ;
 wire \cordic_inst.cordic_state[47] ;
 wire \cordic_inst.cordic_state[48] ;
 wire \cordic_inst.cordic_state[49] ;
 wire \cordic_inst.cordic_state[4] ;
 wire \cordic_inst.cordic_state[50] ;
 wire \cordic_inst.cordic_state[51] ;
 wire \cordic_inst.cordic_state[52] ;
 wire \cordic_inst.cordic_state[53] ;
 wire \cordic_inst.cordic_state[54] ;
 wire \cordic_inst.cordic_state[55] ;
 wire \cordic_inst.cordic_state[56] ;
 wire \cordic_inst.cordic_state[57] ;
 wire \cordic_inst.cordic_state[58] ;
 wire \cordic_inst.cordic_state[59] ;
 wire \cordic_inst.cordic_state[5] ;
 wire \cordic_inst.cordic_state[60] ;
 wire \cordic_inst.cordic_state[61] ;
 wire \cordic_inst.cordic_state[62] ;
 wire \cordic_inst.cordic_state[63] ;
 wire \cordic_inst.cordic_state[64] ;
 wire \cordic_inst.cordic_state[65] ;
 wire \cordic_inst.cordic_state[66] ;
 wire \cordic_inst.cordic_state[67] ;
 wire \cordic_inst.cordic_state[68] ;
 wire \cordic_inst.cordic_state[69] ;
 wire \cordic_inst.cordic_state[6] ;
 wire \cordic_inst.cordic_state[70] ;
 wire \cordic_inst.cordic_state[71] ;
 wire \cordic_inst.cordic_state[72] ;
 wire \cordic_inst.cordic_state[73] ;
 wire \cordic_inst.cordic_state[74] ;
 wire \cordic_inst.cordic_state[75] ;
 wire \cordic_inst.cordic_state[76] ;
 wire \cordic_inst.cordic_state[77] ;
 wire \cordic_inst.cordic_state[78] ;
 wire \cordic_inst.cordic_state[79] ;
 wire \cordic_inst.cordic_state[7] ;
 wire \cordic_inst.current_op[0] ;
 wire \cordic_inst.current_op[1] ;
 wire \cordic_inst.current_op[2] ;
 wire \cordic_inst.operation_pending ;
 wire \cordic_inst.result_ready ;
 wire \exec_phase[1] ;
 wire \exec_phase[2] ;
 wire mac_en_clear;
 wire mac_en_get_mac;
 wire mac_en_get_multiply;
 wire mac_en_mac;
 wire mac_en_multiply;
 wire \mac_inst.RDY_get_mac ;
 wire \mac_inst.RDY_get_multiply ;
 wire \mac_inst.accumulator[0] ;
 wire \mac_inst.accumulator[10] ;
 wire \mac_inst.accumulator[11] ;
 wire \mac_inst.accumulator[12] ;
 wire \mac_inst.accumulator[13] ;
 wire \mac_inst.accumulator[14] ;
 wire \mac_inst.accumulator[15] ;
 wire \mac_inst.accumulator[16] ;
 wire \mac_inst.accumulator[17] ;
 wire \mac_inst.accumulator[18] ;
 wire \mac_inst.accumulator[19] ;
 wire \mac_inst.accumulator[1] ;
 wire \mac_inst.accumulator[20] ;
 wire \mac_inst.accumulator[21] ;
 wire \mac_inst.accumulator[22] ;
 wire \mac_inst.accumulator[23] ;
 wire \mac_inst.accumulator[2] ;
 wire \mac_inst.accumulator[3] ;
 wire \mac_inst.accumulator[4] ;
 wire \mac_inst.accumulator[5] ;
 wire \mac_inst.accumulator[6] ;
 wire \mac_inst.accumulator[7] ;
 wire \mac_inst.accumulator[8] ;
 wire \mac_inst.accumulator[9] ;
 wire \mac_inst.get_multiply[0] ;
 wire \mac_inst.get_multiply[10] ;
 wire \mac_inst.get_multiply[11] ;
 wire \mac_inst.get_multiply[12] ;
 wire \mac_inst.get_multiply[13] ;
 wire \mac_inst.get_multiply[14] ;
 wire \mac_inst.get_multiply[15] ;
 wire \mac_inst.get_multiply[16] ;
 wire \mac_inst.get_multiply[17] ;
 wire \mac_inst.get_multiply[18] ;
 wire \mac_inst.get_multiply[19] ;
 wire \mac_inst.get_multiply[1] ;
 wire \mac_inst.get_multiply[20] ;
 wire \mac_inst.get_multiply[21] ;
 wire \mac_inst.get_multiply[22] ;
 wire \mac_inst.get_multiply[23] ;
 wire \mac_inst.get_multiply[2] ;
 wire \mac_inst.get_multiply[3] ;
 wire \mac_inst.get_multiply[4] ;
 wire \mac_inst.get_multiply[5] ;
 wire \mac_inst.get_multiply[6] ;
 wire \mac_inst.get_multiply[7] ;
 wire \mac_inst.get_multiply[8] ;
 wire \mac_inst.get_multiply[9] ;
 wire rd_prev;
 wire \result_reg[0] ;
 wire \result_reg[10] ;
 wire \result_reg[11] ;
 wire \result_reg[12] ;
 wire \result_reg[13] ;
 wire \result_reg[14] ;
 wire \result_reg[15] ;
 wire \result_reg[16] ;
 wire \result_reg[17] ;
 wire \result_reg[18] ;
 wire \result_reg[19] ;
 wire \result_reg[1] ;
 wire \result_reg[20] ;
 wire \result_reg[21] ;
 wire \result_reg[22] ;
 wire \result_reg[23] ;
 wire \result_reg[24] ;
 wire \result_reg[25] ;
 wire \result_reg[26] ;
 wire \result_reg[27] ;
 wire \result_reg[28] ;
 wire \result_reg[29] ;
 wire \result_reg[2] ;
 wire \result_reg[30] ;
 wire \result_reg[31] ;
 wire \result_reg[32] ;
 wire \result_reg[33] ;
 wire \result_reg[34] ;
 wire \result_reg[35] ;
 wire \result_reg[36] ;
 wire \result_reg[37] ;
 wire \result_reg[38] ;
 wire \result_reg[39] ;
 wire \result_reg[3] ;
 wire \result_reg[40] ;
 wire \result_reg[41] ;
 wire \result_reg[42] ;
 wire \result_reg[43] ;
 wire \result_reg[44] ;
 wire \result_reg[45] ;
 wire \result_reg[46] ;
 wire \result_reg[47] ;
 wire \result_reg[4] ;
 wire \result_reg[5] ;
 wire \result_reg[6] ;
 wire \result_reg[7] ;
 wire \result_reg[8] ;
 wire \result_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire wr_prev;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;

 sg13g2_inv_1 _05215_ (.Y(_04762_),
    .A(\mac_inst.RDY_get_mac ));
 sg13g2_inv_1 _05216_ (.Y(_04763_),
    .A(\mac_inst.accumulator[22] ));
 sg13g2_inv_1 _05217_ (.Y(_04764_),
    .A(\mac_inst.accumulator[20] ));
 sg13g2_inv_1 _05218_ (.Y(_04765_),
    .A(\mac_inst.accumulator[16] ));
 sg13g2_inv_1 _05219_ (.Y(_04766_),
    .A(\mac_inst.accumulator[11] ));
 sg13g2_inv_1 _05220_ (.Y(_04767_),
    .A(\mac_inst.accumulator[8] ));
 sg13g2_inv_1 _05221_ (.Y(_04768_),
    .A(\mac_inst.accumulator[2] ));
 sg13g2_inv_1 _05222_ (.Y(_04769_),
    .A(net190));
 sg13g2_inv_1 _05223_ (.Y(_04770_),
    .A(net1297));
 sg13g2_inv_1 _05224_ (.Y(_04771_),
    .A(net196));
 sg13g2_inv_1 _05225_ (.Y(_04772_),
    .A(net185));
 sg13g2_inv_1 _05226_ (.Y(_04773_),
    .A(net181));
 sg13g2_inv_1 _05227_ (.Y(_04774_),
    .A(net183));
 sg13g2_inv_1 _05228_ (.Y(_04775_),
    .A(net186));
 sg13g2_inv_1 _05229_ (.Y(_04776_),
    .A(net187));
 sg13g2_inv_1 _05230_ (.Y(_04777_),
    .A(net193));
 sg13g2_inv_1 _05231_ (.Y(_04778_),
    .A(net188));
 sg13g2_inv_1 _05232_ (.Y(_04779_),
    .A(net182));
 sg13g2_inv_1 _05233_ (.Y(_04780_),
    .A(net184));
 sg13g2_inv_1 _05234_ (.Y(_04781_),
    .A(net189));
 sg13g2_inv_2 _05235_ (.Y(_04782_),
    .A(\cordic_inst.result_ready ));
 sg13g2_inv_2 _05236_ (.Y(_04783_),
    .A(net1230));
 sg13g2_inv_1 _05237_ (.Y(_04784_),
    .A(net436));
 sg13g2_inv_1 _05238_ (.Y(_04785_),
    .A(net1235));
 sg13g2_inv_1 _05239_ (.Y(_04786_),
    .A(net471));
 sg13g2_inv_1 _05240_ (.Y(_04787_),
    .A(net464));
 sg13g2_inv_1 _05241_ (.Y(_04788_),
    .A(net469));
 sg13g2_inv_1 _05242_ (.Y(_04789_),
    .A(net465));
 sg13g2_inv_2 _05243_ (.Y(_04790_),
    .A(net428));
 sg13g2_inv_1 _05244_ (.Y(_04791_),
    .A(net179));
 sg13g2_inv_2 _05245_ (.Y(_04792_),
    .A(net1256));
 sg13g2_inv_1 _05246_ (.Y(_04793_),
    .A(net1266));
 sg13g2_inv_2 _05247_ (.Y(_04794_),
    .A(net1269));
 sg13g2_inv_1 _05248_ (.Y(_04795_),
    .A(net1274));
 sg13g2_inv_2 _05249_ (.Y(_04796_),
    .A(net492));
 sg13g2_inv_2 _05250_ (.Y(_04797_),
    .A(net432));
 sg13g2_inv_2 _05251_ (.Y(_04798_),
    .A(net450));
 sg13g2_inv_1 _05252_ (.Y(_04799_),
    .A(\byte_counter[0] ));
 sg13g2_inv_1 _05253_ (.Y(_04800_),
    .A(net1519));
 sg13g2_inv_2 _05254_ (.Y(_04801_),
    .A(net1307));
 sg13g2_inv_1 _05255_ (.Y(_04802_),
    .A(net203));
 sg13g2_inv_8 _05256_ (.Y(_04803_),
    .A(net1295));
 sg13g2_inv_4 _05257_ (.A(net1408),
    .Y(_04804_));
 sg13g2_inv_8 _05258_ (.Y(_04805_),
    .A(net1395));
 sg13g2_inv_4 _05259_ (.A(net1392),
    .Y(_04806_));
 sg13g2_inv_2 _05260_ (.Y(_04807_),
    .A(net1385));
 sg13g2_inv_4 _05261_ (.A(net1378),
    .Y(_04808_));
 sg13g2_inv_4 _05262_ (.A(net1370),
    .Y(_04809_));
 sg13g2_inv_2 _05263_ (.Y(_04810_),
    .A(net1355));
 sg13g2_inv_2 _05264_ (.Y(_04811_),
    .A(net1474));
 sg13g2_inv_2 _05265_ (.Y(_04812_),
    .A(net1469));
 sg13g2_inv_1 _05266_ (.Y(_04813_),
    .A(net1461));
 sg13g2_inv_4 _05267_ (.A(net1458),
    .Y(_04814_));
 sg13g2_inv_1 _05268_ (.Y(_04815_),
    .A(net1452));
 sg13g2_inv_1 _05269_ (.Y(_04816_),
    .A(net1448));
 sg13g2_inv_1 _05270_ (.Y(_04817_),
    .A(net1438));
 sg13g2_inv_1 _05271_ (.Y(_04818_),
    .A(net1430));
 sg13g2_inv_1 _05272_ (.Y(_04819_),
    .A(net1422));
 sg13g2_inv_1 _05273_ (.Y(_04820_),
    .A(net1417));
 sg13g2_inv_4 _05274_ (.A(net1413),
    .Y(_04821_));
 sg13g2_inv_4 _05275_ (.A(net1410),
    .Y(_04822_));
 sg13g2_inv_8 _05276_ (.Y(_04823_),
    .A(net1223));
 sg13g2_inv_4 _05277_ (.A(net406),
    .Y(_04824_));
 sg13g2_inv_4 _05278_ (.A(net1208),
    .Y(_04825_));
 sg13g2_inv_4 _05279_ (.A(net1206),
    .Y(_04826_));
 sg13g2_inv_1 _05280_ (.Y(_04827_),
    .A(net1204));
 sg13g2_inv_1 _05281_ (.Y(_04828_),
    .A(net1195));
 sg13g2_inv_1 _05282_ (.Y(_04829_),
    .A(net1193));
 sg13g2_inv_4 _05283_ (.A(net1184),
    .Y(_04830_));
 sg13g2_inv_1 _05284_ (.Y(_04831_),
    .A(net1177));
 sg13g2_inv_8 _05285_ (.Y(_04832_),
    .A(net1173));
 sg13g2_inv_2 _05286_ (.Y(_04833_),
    .A(net1161));
 sg13g2_inv_1 _05287_ (.Y(_04834_),
    .A(net1151));
 sg13g2_inv_1 _05288_ (.Y(_04835_),
    .A(net1348));
 sg13g2_inv_4 _05289_ (.A(net1342),
    .Y(_04836_));
 sg13g2_inv_1 _05290_ (.Y(_04837_),
    .A(net1327));
 sg13g2_nor2_1 _05291_ (.A(net221),
    .B(net211),
    .Y(_04838_));
 sg13g2_nand3b_1 _05292_ (.B(net340),
    .C(_04838_),
    .Y(_04839_),
    .A_N(net299));
 sg13g2_nor3_1 _05293_ (.A(net419),
    .B(net328),
    .C(net303),
    .Y(_04840_));
 sg13g2_nor2b_2 _05294_ (.A(_04839_),
    .B_N(_04840_),
    .Y(_04841_));
 sg13g2_nand2_1 _05295_ (.Y(_04842_),
    .A(net299),
    .B(_04838_));
 sg13g2_nor2_1 _05296_ (.A(net340),
    .B(_04842_),
    .Y(_04843_));
 sg13g2_nor3_1 _05297_ (.A(net470),
    .B(net328),
    .C(net303),
    .Y(_04844_));
 sg13g2_nand2_1 _05298_ (.Y(_04845_),
    .A(net419),
    .B(_04844_));
 sg13g2_and2_1 _05299_ (.A(_04843_),
    .B(_04844_),
    .X(_04846_));
 sg13g2_nand2_2 _05300_ (.Y(_04847_),
    .A(net419),
    .B(_04846_));
 sg13g2_and3_2 _05301_ (.X(_04848_),
    .A(\cmd_reg[0] ),
    .B(_04840_),
    .C(_04843_));
 sg13g2_nand3_1 _05302_ (.B(_04840_),
    .C(_04843_),
    .A(net329),
    .Y(_04849_));
 sg13g2_nor2_2 _05303_ (.A(_04841_),
    .B(net1061),
    .Y(_04850_));
 sg13g2_nand2_2 _05304_ (.Y(_04851_),
    .A(_04847_),
    .B(net1035));
 sg13g2_nor3_2 _05305_ (.A(_04798_),
    .B(\byte_counter[0] ),
    .C(net1475),
    .Y(_04852_));
 sg13g2_nand3b_1 _05306_ (.B(\byte_counter[1] ),
    .C(_04799_),
    .Y(_04853_),
    .A_N(net1475));
 sg13g2_nor2b_2 _05307_ (.A(net429),
    .B_N(net9),
    .Y(_04854_));
 sg13g2_nand2b_2 _05308_ (.Y(_04855_),
    .B(net9),
    .A_N(wr_prev));
 sg13g2_nor2b_2 _05309_ (.A(net1409),
    .B_N(net447),
    .Y(_04856_));
 sg13g2_nand2b_1 _05310_ (.Y(_04857_),
    .B(net447),
    .A_N(net462));
 sg13g2_nor2_1 _05311_ (.A(\state[0] ),
    .B(_04857_),
    .Y(_04858_));
 sg13g2_nand3_1 _05312_ (.B(_04854_),
    .C(_04858_),
    .A(net1111),
    .Y(_04859_));
 sg13g2_nor2_1 _05313_ (.A(_04851_),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_nor2b_2 _05314_ (.A(net447),
    .B_N(\state[0] ),
    .Y(_04861_));
 sg13g2_nand2b_2 _05315_ (.Y(_04862_),
    .B(_04861_),
    .A_N(net1409));
 sg13g2_or2_1 _05316_ (.X(_04863_),
    .B(_04845_),
    .A(_04839_));
 sg13g2_nor2_1 _05317_ (.A(_04862_),
    .B(_04863_),
    .Y(_04864_));
 sg13g2_nand3_1 _05318_ (.B(_04854_),
    .C(_04856_),
    .A(\state[0] ),
    .Y(_04865_));
 sg13g2_nor2_1 _05319_ (.A(_04853_),
    .B(_04865_),
    .Y(_04866_));
 sg13g2_nor3_1 _05320_ (.A(_04860_),
    .B(_04864_),
    .C(net1100),
    .Y(_04867_));
 sg13g2_nor2_1 _05321_ (.A(\state[0] ),
    .B(\state[1] ),
    .Y(_04868_));
 sg13g2_and2_1 _05322_ (.A(net462),
    .B(_04868_),
    .X(_04869_));
 sg13g2_nand2_1 _05323_ (.Y(_04870_),
    .A(_04841_),
    .B(net1110));
 sg13g2_nor2_1 _05324_ (.A(_04846_),
    .B(net1061),
    .Y(_04871_));
 sg13g2_nor2b_2 _05325_ (.A(_04871_),
    .B_N(net1110),
    .Y(_04872_));
 sg13g2_a21oi_2 _05326_ (.B1(_04872_),
    .Y(_04873_),
    .A2(_04869_),
    .A1(_04841_));
 sg13g2_nand2b_1 _05327_ (.Y(_04874_),
    .B(_04873_),
    .A_N(net1229));
 sg13g2_and2_1 _05328_ (.A(_04867_),
    .B(_04874_),
    .X(_00024_));
 sg13g2_nor2_1 _05329_ (.A(\mac_inst.RDY_get_mac ),
    .B(\mac_inst.RDY_get_multiply ),
    .Y(_04875_));
 sg13g2_a21oi_1 _05330_ (.A1(net1228),
    .A2(_04875_),
    .Y(_04876_),
    .B1(net352));
 sg13g2_or2_1 _05331_ (.X(_04877_),
    .B(_04876_),
    .A(_04870_));
 sg13g2_nand2b_1 _05332_ (.Y(_04878_),
    .B(_04851_),
    .A_N(net456));
 sg13g2_nor2b_1 _05333_ (.A(_04862_),
    .B_N(_04863_),
    .Y(_04879_));
 sg13g2_a21o_1 _05334_ (.A2(_04858_),
    .A1(_04851_),
    .B1(_04879_),
    .X(_04880_));
 sg13g2_o21ai_1 _05335_ (.B1(_04873_),
    .Y(_04881_),
    .A1(net462),
    .A2(_04868_));
 sg13g2_a21oi_1 _05336_ (.A1(_04852_),
    .A2(_04854_),
    .Y(_04882_),
    .B1(_04857_));
 sg13g2_nor2_1 _05337_ (.A(_04880_),
    .B(_04882_),
    .Y(_04883_));
 sg13g2_nand2_1 _05338_ (.Y(_04884_),
    .A(_04881_),
    .B(_04883_));
 sg13g2_a21oi_1 _05339_ (.A1(net352),
    .A2(_04884_),
    .Y(_04885_),
    .B1(_04872_));
 sg13g2_a21oi_1 _05340_ (.A1(_04797_),
    .A2(net1228),
    .Y(_04886_),
    .B1(net352));
 sg13g2_o21ai_1 _05341_ (.B1(_04877_),
    .Y(_00021_),
    .A1(_04885_),
    .A2(net353));
 sg13g2_nor2_2 _05342_ (.A(net1317),
    .B(net1315),
    .Y(_04887_));
 sg13g2_or2_1 _05343_ (.X(_04888_),
    .B(net1315),
    .A(net1318));
 sg13g2_a21oi_1 _05344_ (.A1(net220),
    .A2(_04887_),
    .Y(_04889_),
    .B1(net1309));
 sg13g2_nor2_1 _05345_ (.A(net1479),
    .B(_04889_),
    .Y(_00019_));
 sg13g2_nor2_2 _05346_ (.A(net1309),
    .B(net1316),
    .Y(_04890_));
 sg13g2_o21ai_1 _05347_ (.B1(_04890_),
    .Y(_04891_),
    .A1(net1318),
    .A2(net417));
 sg13g2_nand2_1 _05348_ (.Y(_00018_),
    .A(net1512),
    .B(net418));
 sg13g2_nor2b_1 _05349_ (.A(\cmd_reg[0] ),
    .B_N(_04841_),
    .Y(_04892_));
 sg13g2_nand2b_2 _05350_ (.Y(_04893_),
    .B(_04841_),
    .A_N(net329));
 sg13g2_nand2b_2 _05351_ (.Y(_04894_),
    .B(net1110),
    .A_N(net1229));
 sg13g2_nor2_1 _05352_ (.A(_04893_),
    .B(_04894_),
    .Y(_00017_));
 sg13g2_nor2_1 _05353_ (.A(_04847_),
    .B(_04894_),
    .Y(_00012_));
 sg13g2_nor2_1 _05354_ (.A(_04849_),
    .B(_04894_),
    .Y(_00007_));
 sg13g2_nor2b_2 _05355_ (.A(net419),
    .B_N(_04846_),
    .Y(_04895_));
 sg13g2_inv_1 _05356_ (.Y(_04896_),
    .A(_04895_));
 sg13g2_nor2_1 _05357_ (.A(_04894_),
    .B(_04896_),
    .Y(_00011_));
 sg13g2_and2_1 _05358_ (.A(\cmd_reg[0] ),
    .B(_04841_),
    .X(_04897_));
 sg13g2_nand2_1 _05359_ (.Y(_04898_),
    .A(net329),
    .B(_04841_));
 sg13g2_nor2_1 _05360_ (.A(_04894_),
    .B(net330),
    .Y(_00016_));
 sg13g2_nand2_1 _05361_ (.Y(_04899_),
    .A(net432),
    .B(_04872_));
 sg13g2_o21ai_1 _05362_ (.B1(_04899_),
    .Y(_04900_),
    .A1(_04870_),
    .A2(_04875_));
 sg13g2_o21ai_1 _05363_ (.B1(net1228),
    .Y(_04901_),
    .A1(_04884_),
    .A2(_04900_));
 sg13g2_o21ai_1 _05364_ (.B1(net478),
    .Y(_00022_),
    .A1(net1229),
    .A2(_04873_));
 sg13g2_nor2b_2 _05365_ (.A(net1301),
    .B_N(net1312),
    .Y(_04902_));
 sg13g2_nand2_2 _05366_ (.Y(_04903_),
    .A(net1128),
    .B(net1315));
 sg13g2_nand2_1 _05367_ (.Y(_04904_),
    .A(net1510),
    .B(net1125));
 sg13g2_nor2_2 _05368_ (.A(net1309),
    .B(_04888_),
    .Y(_04905_));
 sg13g2_nand2_2 _05369_ (.Y(_04906_),
    .A(net1127),
    .B(_04887_));
 sg13g2_nand2_1 _05370_ (.Y(_04907_),
    .A(net1510),
    .B(net1108));
 sg13g2_o21ai_1 _05371_ (.B1(_04904_),
    .Y(_00020_),
    .A1(_04802_),
    .A2(_04907_));
 sg13g2_nor2_2 _05372_ (.A(\cordic_inst.cordic_state[0] ),
    .B(_04797_),
    .Y(_04908_));
 sg13g2_nand2_2 _05373_ (.Y(_04909_),
    .A(_04796_),
    .B(cordic_busy));
 sg13g2_nor2_1 _05374_ (.A(net1318),
    .B(_04909_),
    .Y(_04910_));
 sg13g2_nand2b_2 _05375_ (.Y(_04911_),
    .B(net1107),
    .A_N(net1318));
 sg13g2_nor2_1 _05376_ (.A(_04888_),
    .B(_04909_),
    .Y(_04912_));
 sg13g2_nand2_2 _05377_ (.Y(_04913_),
    .A(_04887_),
    .B(net1107));
 sg13g2_nand2_1 _05378_ (.Y(_04914_),
    .A(_04890_),
    .B(net1097));
 sg13g2_and2_1 _05379_ (.A(net1281),
    .B(net1292),
    .X(_04915_));
 sg13g2_nand2_2 _05380_ (.Y(_04916_),
    .A(net1276),
    .B(net1282));
 sg13g2_nand2_2 _05381_ (.Y(_04917_),
    .A(net1273),
    .B(_04915_));
 sg13g2_nand3_1 _05382_ (.B(net1273),
    .C(_04915_),
    .A(net1268),
    .Y(_04918_));
 sg13g2_xnor2_1 _05383_ (.Y(_04919_),
    .A(net1259),
    .B(_04918_));
 sg13g2_nand3_1 _05384_ (.B(net1095),
    .C(_04919_),
    .A(net1127),
    .Y(_04920_));
 sg13g2_nor2_1 _05385_ (.A(_04906_),
    .B(_04908_),
    .Y(_04921_));
 sg13g2_nand2_1 _05386_ (.Y(_04922_),
    .A(net1108),
    .B(_04909_));
 sg13g2_nand2_1 _05387_ (.Y(_04923_),
    .A(net1259),
    .B(net1088));
 sg13g2_and3_2 _05388_ (.X(_04924_),
    .A(net1515),
    .B(_04920_),
    .C(_04923_));
 sg13g2_inv_2 _05389_ (.Y(_00141_),
    .A(_04924_));
 sg13g2_nand2_2 _05390_ (.Y(_04925_),
    .A(net1132),
    .B(_04916_));
 sg13g2_nand2_1 _05391_ (.Y(_04926_),
    .A(_04917_),
    .B(_04925_));
 sg13g2_o21ai_1 _05392_ (.B1(net1513),
    .Y(_04927_),
    .A1(net1049),
    .A2(_04926_));
 sg13g2_a21oi_2 _05393_ (.B1(_04927_),
    .Y(_04928_),
    .A2(net1091),
    .A1(net1273));
 sg13g2_inv_4 _05394_ (.A(_04928_),
    .Y(_00139_));
 sg13g2_nand2_2 _05395_ (.Y(_04929_),
    .A(net1136),
    .B(_04917_));
 sg13g2_nor2b_1 _05396_ (.A(net1049),
    .B_N(_04918_),
    .Y(_04930_));
 sg13g2_a22oi_1 _05397_ (.Y(_04931_),
    .B1(_04929_),
    .B2(_04930_),
    .A2(net1087),
    .A1(net1268));
 sg13g2_nand2b_1 _05398_ (.Y(_04932_),
    .B(net1515),
    .A_N(_04931_));
 sg13g2_inv_2 _05399_ (.Y(_00140_),
    .A(_04932_));
 sg13g2_nor2_1 _05400_ (.A(_00139_),
    .B(_00140_),
    .Y(_04933_));
 sg13g2_o21ai_1 _05401_ (.B1(_00141_),
    .Y(_04934_),
    .A1(_00139_),
    .A2(_00140_));
 sg13g2_inv_1 _05402_ (.Y(_00025_),
    .A(_04934_));
 sg13g2_nand2_1 _05403_ (.Y(_04935_),
    .A(_04924_),
    .B(_04928_));
 sg13g2_nor2_2 _05404_ (.A(net1281),
    .B(net1292),
    .Y(_04936_));
 sg13g2_nor3_1 _05405_ (.A(net1049),
    .B(_04915_),
    .C(_04936_),
    .Y(_04937_));
 sg13g2_a21oi_2 _05406_ (.B1(_04937_),
    .Y(_04938_),
    .A2(net1091),
    .A1(net1281));
 sg13g2_nor2_1 _05407_ (.A(net1484),
    .B(_04938_),
    .Y(_00138_));
 sg13g2_o21ai_1 _05408_ (.B1(net1515),
    .Y(_04939_),
    .A1(net1292),
    .A2(_04914_));
 sg13g2_a21oi_2 _05409_ (.B1(_04939_),
    .Y(_04940_),
    .A2(net1091),
    .A1(net1292));
 sg13g2_inv_2 _05410_ (.Y(_00137_),
    .A(_04940_));
 sg13g2_o21ai_1 _05411_ (.B1(_00138_),
    .Y(_04941_),
    .A1(_04931_),
    .A2(_00137_));
 sg13g2_nand2_1 _05412_ (.Y(_04942_),
    .A(_04924_),
    .B(_04931_));
 sg13g2_nand2_1 _05413_ (.Y(_04943_),
    .A(_04924_),
    .B(_04933_));
 sg13g2_nand2_1 _05414_ (.Y(_04944_),
    .A(_04928_),
    .B(_00137_));
 sg13g2_o21ai_1 _05415_ (.B1(_04934_),
    .Y(_00001_),
    .A1(_04935_),
    .A2(_04941_));
 sg13g2_nand2_1 _05416_ (.Y(_04945_),
    .A(_00140_),
    .B(_04938_));
 sg13g2_o21ai_1 _05417_ (.B1(_04934_),
    .Y(_00006_),
    .A1(_04944_),
    .A2(_04945_));
 sg13g2_nand2_2 _05418_ (.Y(_04946_),
    .A(_04938_),
    .B(_04940_));
 sg13g2_a21oi_1 _05419_ (.A1(_04933_),
    .A2(_04946_),
    .Y(_04947_),
    .B1(_00006_));
 sg13g2_a21oi_1 _05420_ (.A1(_00141_),
    .A2(_04933_),
    .Y(_00002_),
    .B1(_04947_));
 sg13g2_nand3_1 _05421_ (.B(_04933_),
    .C(_04946_),
    .A(_04924_),
    .Y(_04948_));
 sg13g2_nor3_1 _05422_ (.A(net1484),
    .B(_04938_),
    .C(_04940_),
    .Y(_04949_));
 sg13g2_nand2b_1 _05423_ (.Y(_04950_),
    .B(_04949_),
    .A_N(_04942_));
 sg13g2_nand3_1 _05424_ (.B(_04948_),
    .C(_04950_),
    .A(_04934_),
    .Y(_00003_));
 sg13g2_o21ai_1 _05425_ (.B1(_00137_),
    .Y(_04951_),
    .A1(net1484),
    .A2(_04938_));
 sg13g2_xnor2_1 _05426_ (.Y(_04952_),
    .A(_00139_),
    .B(_04951_));
 sg13g2_o21ai_1 _05427_ (.B1(_04934_),
    .Y(_00004_),
    .A1(_04942_),
    .A2(_04952_));
 sg13g2_o21ai_1 _05428_ (.B1(_04934_),
    .Y(_00005_),
    .A1(_04948_),
    .A2(_04949_));
 sg13g2_or2_1 _05429_ (.X(_04953_),
    .B(_04946_),
    .A(_04935_));
 sg13g2_o21ai_1 _05430_ (.B1(_04934_),
    .Y(_00000_),
    .A1(_04943_),
    .A2(_04946_));
 sg13g2_nor2_1 _05431_ (.A(_00138_),
    .B(_04943_),
    .Y(_00050_));
 sg13g2_nor2b_1 _05432_ (.A(net1228),
    .B_N(net352),
    .Y(_04954_));
 sg13g2_nand2_1 _05433_ (.Y(_04955_),
    .A(net1229),
    .B(net1110));
 sg13g2_nand3_1 _05434_ (.B(_04869_),
    .C(_04954_),
    .A(net1229),
    .Y(_04956_));
 sg13g2_nor2_1 _05435_ (.A(net330),
    .B(_04956_),
    .Y(_00014_));
 sg13g2_nor2_1 _05436_ (.A(_04893_),
    .B(net378),
    .Y(_00015_));
 sg13g2_nor2_1 _05437_ (.A(net420),
    .B(net378),
    .Y(_00010_));
 sg13g2_nor2_1 _05438_ (.A(_04849_),
    .B(net378),
    .Y(_00008_));
 sg13g2_nor2_1 _05439_ (.A(_04896_),
    .B(_04956_),
    .Y(_00009_));
 sg13g2_nor2_1 _05440_ (.A(_04863_),
    .B(_04894_),
    .Y(_00013_));
 sg13g2_nand2b_2 _05441_ (.Y(_04957_),
    .B(_04940_),
    .A_N(_04938_));
 sg13g2_nand2b_1 _05442_ (.Y(_04958_),
    .B(_04954_),
    .A_N(\mac_inst.RDY_get_multiply ));
 sg13g2_and2_1 _05443_ (.A(net1229),
    .B(_04958_),
    .X(_04959_));
 sg13g2_a22oi_1 _05444_ (.Y(_04960_),
    .B1(net1052),
    .B2(_04762_),
    .A2(net1061),
    .A1(_04802_));
 sg13g2_o21ai_1 _05445_ (.B1(_04960_),
    .Y(_04961_),
    .A1(\cordic_inst.current_op[1] ),
    .A2(_04847_));
 sg13g2_nor2_1 _05446_ (.A(net1228),
    .B(\exec_phase[1] ),
    .Y(_04962_));
 sg13g2_nor2_1 _05447_ (.A(_04782_),
    .B(_04796_),
    .Y(_04963_));
 sg13g2_a221oi_1 _05448_ (.B2(\exec_phase[1] ),
    .C1(\exec_phase[2] ),
    .B1(_04963_),
    .A1(_04847_),
    .Y(_04964_),
    .A2(_04849_));
 sg13g2_or2_1 _05449_ (.X(_04965_),
    .B(_04895_),
    .A(_04841_));
 sg13g2_a221oi_1 _05450_ (.B2(_04965_),
    .C1(_04964_),
    .B1(_04962_),
    .A1(_04954_),
    .Y(_04966_),
    .A2(_04961_));
 sg13g2_nand2b_1 _05451_ (.Y(_04967_),
    .B(net1229),
    .A_N(_04966_));
 sg13g2_o21ai_1 _05452_ (.B1(_04967_),
    .Y(_04968_),
    .A1(_04893_),
    .A2(_04959_));
 sg13g2_nor3_1 _05453_ (.A(_04846_),
    .B(net1061),
    .C(net1052),
    .Y(_04969_));
 sg13g2_nor2_1 _05454_ (.A(_04894_),
    .B(_04969_),
    .Y(_04970_));
 sg13g2_a21oi_1 _05455_ (.A1(_04855_),
    .A2(_04879_),
    .Y(_04971_),
    .B1(_04970_));
 sg13g2_nand2b_1 _05456_ (.Y(_04972_),
    .B(_04849_),
    .A_N(net1229));
 sg13g2_nand4_1 _05457_ (.B(_04851_),
    .C(net1110),
    .A(net1228),
    .Y(_04973_),
    .D(_04972_));
 sg13g2_nand2_1 _05458_ (.Y(_04974_),
    .A(\cordic_inst.current_op[0] ),
    .B(_04963_));
 sg13g2_nand2_1 _05459_ (.Y(_04975_),
    .A(_00009_),
    .B(_04974_));
 sg13g2_nand4_1 _05460_ (.B(_00023_),
    .C(net1110),
    .A(net1228),
    .Y(_04976_),
    .D(_04895_));
 sg13g2_nand2_1 _05461_ (.Y(_04977_),
    .A(_04975_),
    .B(_04976_));
 sg13g2_nand4_1 _05462_ (.B(_04973_),
    .C(_04975_),
    .A(_04971_),
    .Y(_04978_),
    .D(_04976_));
 sg13g2_a21oi_1 _05463_ (.A1(net1110),
    .A2(_04968_),
    .Y(_04979_),
    .B1(_04978_));
 sg13g2_and2_1 _05464_ (.A(net1409),
    .B(_04861_),
    .X(_04980_));
 sg13g2_nand2_1 _05465_ (.Y(_04981_),
    .A(net1409),
    .B(_04861_));
 sg13g2_nand2b_2 _05466_ (.Y(_04982_),
    .B(net10),
    .A_N(rd_prev));
 sg13g2_nor2_2 _05467_ (.A(_04981_),
    .B(_04982_),
    .Y(_04983_));
 sg13g2_and3_2 _05468_ (.X(_04984_),
    .A(_04798_),
    .B(\byte_counter[0] ),
    .C(net1475));
 sg13g2_nand2_1 _05469_ (.Y(_04985_),
    .A(_04895_),
    .B(net1106));
 sg13g2_o21ai_1 _05470_ (.B1(_04985_),
    .Y(_04986_),
    .A1(_04853_),
    .A2(_04895_));
 sg13g2_nand3b_1 _05471_ (.B(net1035),
    .C(net1110),
    .Y(_04987_),
    .A_N(_04846_));
 sg13g2_o21ai_1 _05472_ (.B1(\state[1] ),
    .Y(_04988_),
    .A1(net1409),
    .A2(_04855_));
 sg13g2_nand2_1 _05473_ (.Y(_04989_),
    .A(_04980_),
    .B(_04982_));
 sg13g2_nand4_1 _05474_ (.B(_04987_),
    .C(_04988_),
    .A(_04867_),
    .Y(_04990_),
    .D(_04989_));
 sg13g2_a21oi_1 _05475_ (.A1(net1072),
    .A2(_04986_),
    .Y(_04991_),
    .B1(_04990_));
 sg13g2_and2_1 _05476_ (.A(_04979_),
    .B(_04991_),
    .X(_04992_));
 sg13g2_a221oi_1 _05477_ (.B2(net1409),
    .C1(_04853_),
    .B1(_04861_),
    .A1(\state[0] ),
    .Y(_04993_),
    .A2(_04856_));
 sg13g2_o21ai_1 _05478_ (.B1(_04862_),
    .Y(_04994_),
    .A1(net452),
    .A2(_04993_));
 sg13g2_o21ai_1 _05479_ (.B1(_04994_),
    .Y(_04995_),
    .A1(_04856_),
    .A2(_04861_));
 sg13g2_nor2_1 _05480_ (.A(net452),
    .B(_04992_),
    .Y(_04996_));
 sg13g2_a21oi_1 _05481_ (.A1(_04992_),
    .A2(_04995_),
    .Y(_00026_),
    .B1(_04996_));
 sg13g2_nor2_1 _05482_ (.A(_04856_),
    .B(_04980_),
    .Y(_04997_));
 sg13g2_nand2_1 _05483_ (.Y(_04998_),
    .A(\byte_counter[1] ),
    .B(\byte_counter[0] ));
 sg13g2_xnor2_1 _05484_ (.Y(_04999_),
    .A(net450),
    .B(\byte_counter[0] ));
 sg13g2_nor3_1 _05485_ (.A(_04993_),
    .B(_04997_),
    .C(_04999_),
    .Y(_05000_));
 sg13g2_nand2_1 _05486_ (.Y(_05001_),
    .A(_04992_),
    .B(_05000_));
 sg13g2_o21ai_1 _05487_ (.B1(_05001_),
    .Y(_00027_),
    .A1(_04798_),
    .A2(_04992_));
 sg13g2_nor2_1 _05488_ (.A(net1475),
    .B(_04998_),
    .Y(_05002_));
 sg13g2_and2_1 _05489_ (.A(net1475),
    .B(_04998_),
    .X(_05003_));
 sg13g2_o21ai_1 _05490_ (.B1(_04992_),
    .Y(_05004_),
    .A1(_05002_),
    .A2(_05003_));
 sg13g2_nand2b_1 _05491_ (.Y(_05005_),
    .B(net201),
    .A_N(_04992_));
 sg13g2_o21ai_1 _05492_ (.B1(_05005_),
    .Y(_00028_),
    .A1(_04997_),
    .A2(_05004_));
 sg13g2_nor3_2 _05493_ (.A(\byte_counter[1] ),
    .B(_04799_),
    .C(net1475),
    .Y(_05006_));
 sg13g2_nand3_1 _05494_ (.B(_04858_),
    .C(_05006_),
    .A(_04854_),
    .Y(_05007_));
 sg13g2_nor2_1 _05495_ (.A(net1),
    .B(net1070),
    .Y(_05008_));
 sg13g2_a21oi_1 _05496_ (.A1(_04811_),
    .A2(net1070),
    .Y(_00029_),
    .B1(_05008_));
 sg13g2_nor2_1 _05497_ (.A(net2),
    .B(net1071),
    .Y(_05009_));
 sg13g2_a21oi_1 _05498_ (.A1(_04812_),
    .A2(net1071),
    .Y(_00030_),
    .B1(_05009_));
 sg13g2_nor2_1 _05499_ (.A(net3),
    .B(net1070),
    .Y(_05010_));
 sg13g2_a21oi_1 _05500_ (.A1(_04813_),
    .A2(net1070),
    .Y(_00031_),
    .B1(_05010_));
 sg13g2_nor2_1 _05501_ (.A(net4),
    .B(net1070),
    .Y(_05011_));
 sg13g2_a21oi_1 _05502_ (.A1(_04814_),
    .A2(net1071),
    .Y(_00032_),
    .B1(_05011_));
 sg13g2_nor2_1 _05503_ (.A(net5),
    .B(net1070),
    .Y(_05012_));
 sg13g2_a21oi_1 _05504_ (.A1(_04815_),
    .A2(net1070),
    .Y(_00033_),
    .B1(_05012_));
 sg13g2_nor2_1 _05505_ (.A(net6),
    .B(net1071),
    .Y(_05013_));
 sg13g2_a21oi_1 _05506_ (.A1(_04816_),
    .A2(net1071),
    .Y(_00034_),
    .B1(_05013_));
 sg13g2_mux2_1 _05507_ (.A0(net7),
    .A1(net1442),
    .S(net1070),
    .X(_00035_));
 sg13g2_nor2_1 _05508_ (.A(net8),
    .B(net1071),
    .Y(_05014_));
 sg13g2_a21oi_1 _05509_ (.A1(_04817_),
    .A2(net1071),
    .Y(_00036_),
    .B1(_05014_));
 sg13g2_mux2_1 _05510_ (.A0(net1),
    .A1(net1433),
    .S(net1101),
    .X(_00037_));
 sg13g2_nor2_1 _05511_ (.A(net2),
    .B(net1101),
    .Y(_05015_));
 sg13g2_a21oi_1 _05512_ (.A1(_04818_),
    .A2(net1101),
    .Y(_00038_),
    .B1(_05015_));
 sg13g2_mux2_1 _05513_ (.A0(net3),
    .A1(net1425),
    .S(net1101),
    .X(_00039_));
 sg13g2_nor2_1 _05514_ (.A(net4),
    .B(net1101),
    .Y(_05016_));
 sg13g2_a21oi_1 _05515_ (.A1(_04819_),
    .A2(net1102),
    .Y(_00040_),
    .B1(_05016_));
 sg13g2_mux2_1 _05516_ (.A0(net5),
    .A1(net1419),
    .S(net1101),
    .X(_00041_));
 sg13g2_nor2_1 _05517_ (.A(net6),
    .B(net1102),
    .Y(_05017_));
 sg13g2_a21oi_1 _05518_ (.A1(_04820_),
    .A2(net1102),
    .Y(_00042_),
    .B1(_05017_));
 sg13g2_nor2_1 _05519_ (.A(net7),
    .B(net1101),
    .Y(_05018_));
 sg13g2_a21oi_1 _05520_ (.A1(_04821_),
    .A2(net1101),
    .Y(_00043_),
    .B1(_05018_));
 sg13g2_nor2_1 _05521_ (.A(net8),
    .B(net1102),
    .Y(_05019_));
 sg13g2_a21oi_1 _05522_ (.A1(_04822_),
    .A2(net1102),
    .Y(_00044_),
    .B1(_05019_));
 sg13g2_and3_1 _05523_ (.X(_05020_),
    .A(_04928_),
    .B(_00140_),
    .C(_04957_));
 sg13g2_a22oi_1 _05524_ (.Y(_05021_),
    .B1(_04957_),
    .B2(_04928_),
    .A2(_04938_),
    .A1(_00140_));
 sg13g2_nor3_1 _05525_ (.A(_00141_),
    .B(_05020_),
    .C(_05021_),
    .Y(_00045_));
 sg13g2_o21ai_1 _05526_ (.B1(_04948_),
    .Y(_00046_),
    .A1(_04935_),
    .A2(_04957_));
 sg13g2_o21ai_1 _05527_ (.B1(_04953_),
    .Y(_00047_),
    .A1(_00139_),
    .A2(_04950_));
 sg13g2_a21oi_1 _05528_ (.A1(_04944_),
    .A2(_04957_),
    .Y(_00048_),
    .B1(_04942_));
 sg13g2_nand2b_1 _05529_ (.Y(_05022_),
    .B(_00139_),
    .A_N(_04946_));
 sg13g2_o21ai_1 _05530_ (.B1(_04948_),
    .Y(_00049_),
    .A1(_04942_),
    .A2(_05022_));
 sg13g2_nand3_1 _05531_ (.B(_00023_),
    .C(_04851_),
    .A(net1228),
    .Y(_05023_));
 sg13g2_o21ai_1 _05532_ (.B1(_05023_),
    .Y(_05024_),
    .A1(_00023_),
    .A2(_04969_));
 sg13g2_nor4_2 _05533_ (.A(_04873_),
    .B(_04968_),
    .C(_04977_),
    .Y(_05025_),
    .D(_05024_));
 sg13g2_a22oi_1 _05534_ (.Y(_05026_),
    .B1(net1053),
    .B2(net397),
    .A2(net1063),
    .A1(net413));
 sg13g2_a22oi_1 _05535_ (.Y(_05027_),
    .B1(net1058),
    .B2(net189),
    .A2(net1037),
    .A1(net415));
 sg13g2_nand2_1 _05536_ (.Y(_05028_),
    .A(_05026_),
    .B(_05027_));
 sg13g2_mux2_1 _05537_ (.A0(net427),
    .A1(_05028_),
    .S(net1025),
    .X(_00051_));
 sg13g2_a22oi_1 _05538_ (.Y(_05029_),
    .B1(net1053),
    .B2(\mac_inst.accumulator[1] ),
    .A2(net1062),
    .A1(\cordic_atan2_result[1] ));
 sg13g2_a22oi_1 _05539_ (.Y(_05030_),
    .B1(net1057),
    .B2(\mac_inst.get_multiply[1] ),
    .A2(net1036),
    .A1(\cordic_inst.cordic_state[57] ));
 sg13g2_nand2_2 _05540_ (.Y(_05031_),
    .A(_05029_),
    .B(_05030_));
 sg13g2_mux2_1 _05541_ (.A0(net243),
    .A1(_05031_),
    .S(net1021),
    .X(_00052_));
 sg13g2_a22oi_1 _05542_ (.Y(_05032_),
    .B1(net1053),
    .B2(net315),
    .A2(net1062),
    .A1(net362));
 sg13g2_a22oi_1 _05543_ (.Y(_05033_),
    .B1(net1057),
    .B2(net310),
    .A2(net1036),
    .A1(\cordic_inst.cordic_state[58] ));
 sg13g2_nand2_1 _05544_ (.Y(_05034_),
    .A(_05032_),
    .B(_05033_));
 sg13g2_mux2_1 _05545_ (.A0(net407),
    .A1(_05034_),
    .S(net1024),
    .X(_00053_));
 sg13g2_a22oi_1 _05546_ (.Y(_05035_),
    .B1(net1053),
    .B2(\mac_inst.accumulator[3] ),
    .A2(net1062),
    .A1(\cordic_atan2_result[3] ));
 sg13g2_a22oi_1 _05547_ (.Y(_05036_),
    .B1(net1057),
    .B2(net300),
    .A2(net1036),
    .A1(\cordic_inst.cordic_state[59] ));
 sg13g2_nand2_1 _05548_ (.Y(_05037_),
    .A(_05035_),
    .B(_05036_));
 sg13g2_mux2_1 _05549_ (.A0(net370),
    .A1(_05037_),
    .S(net1024),
    .X(_00054_));
 sg13g2_nor2_1 _05550_ (.A(net200),
    .B(net1021),
    .Y(_05038_));
 sg13g2_a22oi_1 _05551_ (.Y(_05039_),
    .B1(net1053),
    .B2(net559),
    .A2(net1062),
    .A1(\cordic_atan2_result[4] ));
 sg13g2_inv_1 _05552_ (.Y(_05040_),
    .A(_05039_));
 sg13g2_a221oi_1 _05553_ (.B2(net184),
    .C1(_05040_),
    .B1(net1058),
    .A1(\cordic_inst.cordic_state[60] ),
    .Y(_05041_),
    .A2(net1036));
 sg13g2_a21oi_1 _05554_ (.A1(net1021),
    .A2(_05041_),
    .Y(_00055_),
    .B1(_05038_));
 sg13g2_a22oi_1 _05555_ (.Y(_05042_),
    .B1(net1054),
    .B2(net267),
    .A2(net1062),
    .A1(net398));
 sg13g2_a22oi_1 _05556_ (.Y(_05043_),
    .B1(net1057),
    .B2(net182),
    .A2(net1036),
    .A1(\cordic_inst.cordic_state[61] ));
 sg13g2_nand2_1 _05557_ (.Y(_05044_),
    .A(_05042_),
    .B(_05043_));
 sg13g2_mux2_1 _05558_ (.A0(net445),
    .A1(_05044_),
    .S(net1025),
    .X(_00056_));
 sg13g2_a22oi_1 _05559_ (.Y(_05045_),
    .B1(net1053),
    .B2(net387),
    .A2(net1057),
    .A1(net188));
 sg13g2_a22oi_1 _05560_ (.Y(_05046_),
    .B1(net1037),
    .B2(\cordic_inst.cordic_state[62] ),
    .A2(net1062),
    .A1(net376));
 sg13g2_nand2_1 _05561_ (.Y(_05047_),
    .A(_05045_),
    .B(_05046_));
 sg13g2_mux2_1 _05562_ (.A0(net391),
    .A1(_05047_),
    .S(net1025),
    .X(_00057_));
 sg13g2_a22oi_1 _05563_ (.Y(_05048_),
    .B1(net1054),
    .B2(net347),
    .A2(net1062),
    .A1(net400));
 sg13g2_a22oi_1 _05564_ (.Y(_05049_),
    .B1(net1057),
    .B2(net297),
    .A2(net1036),
    .A1(net561));
 sg13g2_nand2_1 _05565_ (.Y(_05050_),
    .A(_05048_),
    .B(_05049_));
 sg13g2_mux2_1 _05566_ (.A0(net424),
    .A1(_05050_),
    .S(net1025),
    .X(_00058_));
 sg13g2_a22oi_1 _05567_ (.Y(_05051_),
    .B1(net1053),
    .B2(net254),
    .A2(net1057),
    .A1(\mac_inst.get_multiply[8] ));
 sg13g2_a22oi_1 _05568_ (.Y(_05052_),
    .B1(net1036),
    .B2(\cordic_inst.cordic_state[64] ),
    .A2(net1062),
    .A1(\cordic_atan2_result[8] ));
 sg13g2_nand2_2 _05569_ (.Y(_05053_),
    .A(_05051_),
    .B(_05052_));
 sg13g2_mux2_1 _05570_ (.A0(net258),
    .A1(_05053_),
    .S(net1022),
    .X(_00059_));
 sg13g2_a22oi_1 _05571_ (.Y(_05054_),
    .B1(net1054),
    .B2(net411),
    .A2(net1063),
    .A1(net437));
 sg13g2_a22oi_1 _05572_ (.Y(_05055_),
    .B1(net1057),
    .B2(net256),
    .A2(net1036),
    .A1(\cordic_inst.cordic_state[65] ));
 sg13g2_nand2_1 _05573_ (.Y(_05056_),
    .A(_05054_),
    .B(_05055_));
 sg13g2_mux2_1 _05574_ (.A0(net444),
    .A1(_05056_),
    .S(net1025),
    .X(_00060_));
 sg13g2_a22oi_1 _05575_ (.Y(_05057_),
    .B1(net1054),
    .B2(net381),
    .A2(net1063),
    .A1(net380));
 sg13g2_a22oi_1 _05576_ (.Y(_05058_),
    .B1(net1058),
    .B2(net193),
    .A2(net1037),
    .A1(\cordic_inst.cordic_state[66] ));
 sg13g2_nand2_1 _05577_ (.Y(_05059_),
    .A(_05057_),
    .B(_05058_));
 sg13g2_mux2_1 _05578_ (.A0(net399),
    .A1(_05059_),
    .S(net1024),
    .X(_00061_));
 sg13g2_nor2_1 _05579_ (.A(net228),
    .B(net1022),
    .Y(_05060_));
 sg13g2_a22oi_1 _05580_ (.Y(_05061_),
    .B1(net1053),
    .B2(net204),
    .A2(net1063),
    .A1(\cordic_atan2_result[11] ));
 sg13g2_inv_1 _05581_ (.Y(_05062_),
    .A(_05061_));
 sg13g2_a221oi_1 _05582_ (.B2(\mac_inst.get_multiply[11] ),
    .C1(_05062_),
    .B1(net1056),
    .A1(\cordic_inst.cordic_state[67] ),
    .Y(_05063_),
    .A2(net1034));
 sg13g2_a21oi_1 _05583_ (.A1(net1022),
    .A2(_05063_),
    .Y(_00062_),
    .B1(_05060_));
 sg13g2_a22oi_1 _05584_ (.Y(_05064_),
    .B1(net1051),
    .B2(net249),
    .A2(net1060),
    .A1(\cordic_atan2_result[12] ));
 sg13g2_a22oi_1 _05585_ (.Y(_05065_),
    .B1(net1056),
    .B2(net187),
    .A2(net1034),
    .A1(\cordic_inst.cordic_state[68] ));
 sg13g2_nand2_1 _05586_ (.Y(_05066_),
    .A(_05064_),
    .B(_05065_));
 sg13g2_mux2_1 _05587_ (.A0(net345),
    .A1(_05066_),
    .S(net1023),
    .X(_00063_));
 sg13g2_nor2_1 _05588_ (.A(net214),
    .B(net1024),
    .Y(_00282_));
 sg13g2_a22oi_1 _05589_ (.Y(_00283_),
    .B1(net1051),
    .B2(\mac_inst.accumulator[13] ),
    .A2(net1060),
    .A1(\cordic_atan2_result[13] ));
 sg13g2_inv_1 _05590_ (.Y(_00284_),
    .A(_00283_));
 sg13g2_a221oi_1 _05591_ (.B2(net186),
    .C1(_00284_),
    .B1(net1056),
    .A1(\cordic_inst.cordic_state[69] ),
    .Y(_00285_),
    .A2(net1034));
 sg13g2_a21oi_1 _05592_ (.A1(net1024),
    .A2(_00285_),
    .Y(_00064_),
    .B1(_00282_));
 sg13g2_a22oi_1 _05593_ (.Y(_00286_),
    .B1(net1051),
    .B2(net240),
    .A2(net1060),
    .A1(\cordic_atan2_result[14] ));
 sg13g2_a22oi_1 _05594_ (.Y(_00287_),
    .B1(net1056),
    .B2(net183),
    .A2(net1034),
    .A1(\cordic_inst.cordic_state[70] ));
 sg13g2_nand2_1 _05595_ (.Y(_00288_),
    .A(_00286_),
    .B(_00287_));
 sg13g2_mux2_1 _05596_ (.A0(net308),
    .A1(_00288_),
    .S(net1024),
    .X(_00065_));
 sg13g2_a22oi_1 _05597_ (.Y(_00289_),
    .B1(net1051),
    .B2(\mac_inst.accumulator[15] ),
    .A2(net1056),
    .A1(net181));
 sg13g2_a22oi_1 _05598_ (.Y(_00290_),
    .B1(net1034),
    .B2(\cordic_inst.cordic_state[71] ),
    .A2(net1060),
    .A1(\cordic_atan2_result[15] ));
 sg13g2_nand2_2 _05599_ (.Y(_00291_),
    .A(_00289_),
    .B(_00290_));
 sg13g2_mux2_1 _05600_ (.A0(net212),
    .A1(_00291_),
    .S(net1021),
    .X(_00066_));
 sg13g2_nor2_1 _05601_ (.A(net191),
    .B(net1021),
    .Y(_00292_));
 sg13g2_a22oi_1 _05602_ (.Y(_00293_),
    .B1(net1050),
    .B2(\mac_inst.accumulator[16] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[16] ));
 sg13g2_inv_1 _05603_ (.Y(_00294_),
    .A(_00293_));
 sg13g2_a221oi_1 _05604_ (.B2(\mac_inst.get_multiply[16] ),
    .C1(_00294_),
    .B1(net1055),
    .A1(\cordic_inst.cordic_state[72] ),
    .Y(_00295_),
    .A2(net1033));
 sg13g2_a21oi_1 _05605_ (.A1(net1021),
    .A2(_00295_),
    .Y(_00067_),
    .B1(_00292_));
 sg13g2_nor2_1 _05606_ (.A(net247),
    .B(net1022),
    .Y(_00296_));
 sg13g2_a22oi_1 _05607_ (.Y(_00297_),
    .B1(net1050),
    .B2(\mac_inst.accumulator[17] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[17] ));
 sg13g2_inv_1 _05608_ (.Y(_00298_),
    .A(_00297_));
 sg13g2_a221oi_1 _05609_ (.B2(net185),
    .C1(_00298_),
    .B1(net1055),
    .A1(\cordic_inst.cordic_state[73] ),
    .Y(_00299_),
    .A2(net1033));
 sg13g2_a21oi_1 _05610_ (.A1(net1022),
    .A2(_00299_),
    .Y(_00068_),
    .B1(_00296_));
 sg13g2_nor2_1 _05611_ (.A(net209),
    .B(net1021),
    .Y(_00300_));
 sg13g2_a22oi_1 _05612_ (.Y(_00301_),
    .B1(net1050),
    .B2(\mac_inst.accumulator[18] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[18] ));
 sg13g2_inv_1 _05613_ (.Y(_00302_),
    .A(_00301_));
 sg13g2_a221oi_1 _05614_ (.B2(net196),
    .C1(_00302_),
    .B1(net1055),
    .A1(\cordic_inst.cordic_state[74] ),
    .Y(_00303_),
    .A2(net1033));
 sg13g2_a21oi_1 _05615_ (.A1(net1021),
    .A2(_00303_),
    .Y(_00069_),
    .B1(_00300_));
 sg13g2_nor2_1 _05616_ (.A(net207),
    .B(net1024),
    .Y(_00304_));
 sg13g2_a22oi_1 _05617_ (.Y(_00305_),
    .B1(net1050),
    .B2(\mac_inst.accumulator[19] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[19] ));
 sg13g2_inv_1 _05618_ (.Y(_00306_),
    .A(_00305_));
 sg13g2_a221oi_1 _05619_ (.B2(\mac_inst.get_multiply[19] ),
    .C1(_00306_),
    .B1(net1055),
    .A1(\cordic_inst.cordic_state[75] ),
    .Y(_00307_),
    .A2(net1033));
 sg13g2_a21oi_1 _05620_ (.A1(net1024),
    .A2(_00307_),
    .Y(_00070_),
    .B1(_00304_));
 sg13g2_nor2_1 _05621_ (.A(net198),
    .B(net1023),
    .Y(_00308_));
 sg13g2_a22oi_1 _05622_ (.Y(_00309_),
    .B1(net1050),
    .B2(net197),
    .A2(net1059),
    .A1(\cordic_atan2_result[20] ));
 sg13g2_inv_1 _05623_ (.Y(_00310_),
    .A(_00309_));
 sg13g2_a221oi_1 _05624_ (.B2(\mac_inst.get_multiply[20] ),
    .C1(_00310_),
    .B1(net1055),
    .A1(\cordic_inst.cordic_state[76] ),
    .Y(_00311_),
    .A2(net1033));
 sg13g2_a21oi_1 _05625_ (.A1(net1023),
    .A2(_00311_),
    .Y(_00071_),
    .B1(_00308_));
 sg13g2_a22oi_1 _05626_ (.Y(_00312_),
    .B1(net1050),
    .B2(\mac_inst.accumulator[21] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[21] ));
 sg13g2_a22oi_1 _05627_ (.Y(_00313_),
    .B1(net1055),
    .B2(\mac_inst.get_multiply[21] ),
    .A2(net1033),
    .A1(\cordic_inst.cordic_state[77] ));
 sg13g2_nand2_1 _05628_ (.Y(_00314_),
    .A(_00312_),
    .B(_00313_));
 sg13g2_mux2_1 _05629_ (.A0(net230),
    .A1(_00314_),
    .S(net1023),
    .X(_00072_));
 sg13g2_a22oi_1 _05630_ (.Y(_00315_),
    .B1(net1050),
    .B2(net263),
    .A2(net1059),
    .A1(\cordic_atan2_result[22] ));
 sg13g2_a22oi_1 _05631_ (.Y(_00316_),
    .B1(net1055),
    .B2(net260),
    .A2(net1033),
    .A1(\cordic_inst.cordic_state[78] ));
 sg13g2_nand2_1 _05632_ (.Y(_00317_),
    .A(_00315_),
    .B(_00316_));
 sg13g2_mux2_1 _05633_ (.A0(net306),
    .A1(_00317_),
    .S(net1022),
    .X(_00073_));
 sg13g2_a22oi_1 _05634_ (.Y(_00318_),
    .B1(net1050),
    .B2(net242),
    .A2(net1055),
    .A1(net190));
 sg13g2_a22oi_1 _05635_ (.Y(_00319_),
    .B1(net1033),
    .B2(\cordic_inst.cordic_state[79] ),
    .A2(net1059),
    .A1(\cordic_atan2_result[23] ));
 sg13g2_nand2_1 _05636_ (.Y(_00320_),
    .A(_00318_),
    .B(_00319_));
 sg13g2_mux2_1 _05637_ (.A0(net374),
    .A1(_00320_),
    .S(net1023),
    .X(_00074_));
 sg13g2_nor3_2 _05638_ (.A(net1409),
    .B(\state[0] ),
    .C(net447),
    .Y(_00321_));
 sg13g2_nor2_2 _05639_ (.A(_04861_),
    .B(_00321_),
    .Y(_00322_));
 sg13g2_a22oi_1 _05640_ (.Y(_00323_),
    .B1(net1104),
    .B2(net258),
    .A2(_04984_),
    .A1(net359));
 sg13g2_and3_2 _05641_ (.X(_00324_),
    .A(_04798_),
    .B(_04799_),
    .C(net1475));
 sg13g2_nor3_1 _05642_ (.A(\byte_counter[1] ),
    .B(\byte_counter[0] ),
    .C(net1475),
    .Y(_00325_));
 sg13g2_a22oi_1 _05643_ (.Y(_00326_),
    .B1(_00324_),
    .B2(net343),
    .A2(net1111),
    .A1(net191));
 sg13g2_a22oi_1 _05644_ (.Y(_00327_),
    .B1(net1123),
    .B2(\result_reg[0] ),
    .A2(net1105),
    .A1(net218));
 sg13g2_nand3_1 _05645_ (.B(_00326_),
    .C(_00327_),
    .A(_00323_),
    .Y(_00328_));
 sg13g2_a22oi_1 _05646_ (.Y(_00329_),
    .B1(_00328_),
    .B2(_04983_),
    .A2(_00322_),
    .A1(net365));
 sg13g2_inv_1 _05647_ (.Y(_00075_),
    .A(net366));
 sg13g2_a22oi_1 _05648_ (.Y(_00330_),
    .B1(net1104),
    .B2(\result_reg[9] ),
    .A2(net1106),
    .A1(\result_reg[41] ));
 sg13g2_a22oi_1 _05649_ (.Y(_00331_),
    .B1(net1105),
    .B2(net222),
    .A2(net1111),
    .A1(net247));
 sg13g2_a22oi_1 _05650_ (.Y(_00332_),
    .B1(net1123),
    .B2(net243),
    .A2(_00324_),
    .A1(net274));
 sg13g2_nand3_1 _05651_ (.B(_00331_),
    .C(_00332_),
    .A(_00330_),
    .Y(_00333_));
 sg13g2_a22oi_1 _05652_ (.Y(_00334_),
    .B1(_00333_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net319));
 sg13g2_inv_1 _05653_ (.Y(_00076_),
    .A(net320));
 sg13g2_a22oi_1 _05654_ (.Y(_00335_),
    .B1(_00324_),
    .B2(net336),
    .A2(net1111),
    .A1(net209));
 sg13g2_a22oi_1 _05655_ (.Y(_00336_),
    .B1(net1105),
    .B2(\result_reg[26] ),
    .A2(net1106),
    .A1(net295));
 sg13g2_a22oi_1 _05656_ (.Y(_00337_),
    .B1(net1123),
    .B2(\result_reg[2] ),
    .A2(net1104),
    .A1(\result_reg[10] ));
 sg13g2_nand3_1 _05657_ (.B(_00336_),
    .C(_00337_),
    .A(_00335_),
    .Y(_00338_));
 sg13g2_a22oi_1 _05658_ (.Y(_00339_),
    .B1(_00338_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net341));
 sg13g2_inv_1 _05659_ (.Y(_00077_),
    .A(net342));
 sg13g2_a22oi_1 _05660_ (.Y(_00340_),
    .B1(net1123),
    .B2(\result_reg[3] ),
    .A2(net1111),
    .A1(net207));
 sg13g2_a22oi_1 _05661_ (.Y(_00341_),
    .B1(net1104),
    .B2(net228),
    .A2(net1106),
    .A1(\result_reg[43] ));
 sg13g2_a22oi_1 _05662_ (.Y(_00342_),
    .B1(_00324_),
    .B2(\result_reg[35] ),
    .A2(net1105),
    .A1(net226));
 sg13g2_nand3_1 _05663_ (.B(_00341_),
    .C(_00342_),
    .A(_00340_),
    .Y(_00343_));
 sg13g2_a22oi_1 _05664_ (.Y(_00344_),
    .B1(_00343_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net311));
 sg13g2_inv_1 _05665_ (.Y(_00078_),
    .A(net312));
 sg13g2_a22oi_1 _05666_ (.Y(_00345_),
    .B1(net1123),
    .B2(net200),
    .A2(_00324_),
    .A1(\result_reg[36] ));
 sg13g2_a22oi_1 _05667_ (.Y(_00346_),
    .B1(net1104),
    .B2(\result_reg[12] ),
    .A2(net1111),
    .A1(net198));
 sg13g2_a22oi_1 _05668_ (.Y(_00347_),
    .B1(net1105),
    .B2(net232),
    .A2(net1106),
    .A1(net269));
 sg13g2_nand3_1 _05669_ (.B(_00346_),
    .C(_00347_),
    .A(_00345_),
    .Y(_00348_));
 sg13g2_a22oi_1 _05670_ (.Y(_00349_),
    .B1(_00348_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net279));
 sg13g2_inv_1 _05671_ (.Y(_00079_),
    .A(net280));
 sg13g2_a22oi_1 _05672_ (.Y(_00350_),
    .B1(net1123),
    .B2(\result_reg[5] ),
    .A2(net1106),
    .A1(\result_reg[45] ));
 sg13g2_a22oi_1 _05673_ (.Y(_00351_),
    .B1(net1104),
    .B2(net214),
    .A2(net1111),
    .A1(net230));
 sg13g2_a22oi_1 _05674_ (.Y(_00352_),
    .B1(_00324_),
    .B2(net317),
    .A2(net1105),
    .A1(net245));
 sg13g2_nand3_1 _05675_ (.B(_00351_),
    .C(_00352_),
    .A(_00350_),
    .Y(_00353_));
 sg13g2_a22oi_1 _05676_ (.Y(_00354_),
    .B1(_00353_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net332));
 sg13g2_inv_1 _05677_ (.Y(_00080_),
    .A(net333));
 sg13g2_a22oi_1 _05678_ (.Y(_00355_),
    .B1(_00324_),
    .B2(\result_reg[38] ),
    .A2(net1111),
    .A1(net306));
 sg13g2_a22oi_1 _05679_ (.Y(_00356_),
    .B1(net1105),
    .B2(net238),
    .A2(net1106),
    .A1(net265));
 sg13g2_a22oi_1 _05680_ (.Y(_00357_),
    .B1(net1123),
    .B2(\result_reg[6] ),
    .A2(_05006_),
    .A1(net308));
 sg13g2_nand3_1 _05681_ (.B(_00356_),
    .C(_00357_),
    .A(_00355_),
    .Y(_00358_));
 sg13g2_a22oi_1 _05682_ (.Y(_00359_),
    .B1(_00358_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net363));
 sg13g2_inv_1 _05683_ (.Y(_00081_),
    .A(net364));
 sg13g2_a22oi_1 _05684_ (.Y(_00360_),
    .B1(_00325_),
    .B2(net424),
    .A2(_04852_),
    .A1(net374));
 sg13g2_a22oi_1 _05685_ (.Y(_00361_),
    .B1(net1104),
    .B2(net212),
    .A2(net1105),
    .A1(net334));
 sg13g2_a22oi_1 _05686_ (.Y(_00362_),
    .B1(_00324_),
    .B2(net291),
    .A2(net1106),
    .A1(net252));
 sg13g2_nand3_1 _05687_ (.B(_00361_),
    .C(_00362_),
    .A(_00360_),
    .Y(_00363_));
 sg13g2_a22oi_1 _05688_ (.Y(_00364_),
    .B1(_00363_),
    .B2(net1072),
    .A2(_00322_),
    .A1(net442));
 sg13g2_nand2_1 _05689_ (.Y(_00082_),
    .A(_04862_),
    .B(_00364_));
 sg13g2_nor3_1 _05690_ (.A(_04981_),
    .B(_04982_),
    .C(_04986_),
    .Y(_00365_));
 sg13g2_a21oi_1 _05691_ (.A1(_04855_),
    .A2(_00321_),
    .Y(_00366_),
    .B1(_04882_));
 sg13g2_nand2b_1 _05692_ (.Y(_00367_),
    .B(_00013_),
    .A_N(_04875_));
 sg13g2_o21ai_1 _05693_ (.B1(_00367_),
    .Y(_00368_),
    .A1(_04863_),
    .A2(_04955_));
 sg13g2_nor3_1 _05694_ (.A(_00012_),
    .B(_00365_),
    .C(_00368_),
    .Y(_00369_));
 sg13g2_and4_1 _05695_ (.A(_04979_),
    .B(_04989_),
    .C(_00366_),
    .D(_00369_),
    .X(_00370_));
 sg13g2_nor2b_1 _05696_ (.A(_00321_),
    .B_N(_04873_),
    .Y(_00371_));
 sg13g2_o21ai_1 _05697_ (.B1(_00371_),
    .Y(_00372_),
    .A1(_04857_),
    .A2(_04878_));
 sg13g2_mux2_1 _05698_ (.A0(net456),
    .A1(_00372_),
    .S(_00370_),
    .X(_00083_));
 sg13g2_a21o_1 _05699_ (.A2(_00370_),
    .A1(_04880_),
    .B1(_04882_),
    .X(_00084_));
 sg13g2_a21oi_1 _05700_ (.A1(_04856_),
    .A2(_04878_),
    .Y(_00373_),
    .B1(_04864_));
 sg13g2_nand2_1 _05701_ (.Y(_00374_),
    .A(_04873_),
    .B(_00373_));
 sg13g2_mux2_1 _05702_ (.A0(net1409),
    .A1(_00374_),
    .S(_00370_),
    .X(_00085_));
 sg13g2_nand2_2 _05703_ (.Y(_00375_),
    .A(_04854_),
    .B(_00321_));
 sg13g2_mux2_1 _05704_ (.A0(net1),
    .A1(net329),
    .S(_00375_),
    .X(_00086_));
 sg13g2_mux2_1 _05705_ (.A0(net2),
    .A1(net419),
    .S(_00375_),
    .X(_00087_));
 sg13g2_mux2_1 _05706_ (.A0(net3),
    .A1(net303),
    .S(_00375_),
    .X(_00088_));
 sg13g2_mux2_1 _05707_ (.A0(net4),
    .A1(net328),
    .S(_00375_),
    .X(_00089_));
 sg13g2_mux2_1 _05708_ (.A0(net5),
    .A1(net299),
    .S(_00375_),
    .X(_00090_));
 sg13g2_mux2_1 _05709_ (.A0(net6),
    .A1(net340),
    .S(_00375_),
    .X(_00091_));
 sg13g2_mux2_1 _05710_ (.A0(net7),
    .A1(net211),
    .S(_00375_),
    .X(_00092_));
 sg13g2_mux2_1 _05711_ (.A0(net8),
    .A1(net221),
    .S(_00375_),
    .X(_00093_));
 sg13g2_nand2_1 _05712_ (.Y(_00376_),
    .A(_04854_),
    .B(_04879_));
 sg13g2_nor2_1 _05713_ (.A(net1),
    .B(net1031),
    .Y(_00377_));
 sg13g2_a21oi_1 _05714_ (.A1(_04804_),
    .A2(net1031),
    .Y(_00094_),
    .B1(_00377_));
 sg13g2_nor2_1 _05715_ (.A(net2),
    .B(net1032),
    .Y(_00378_));
 sg13g2_a21oi_1 _05716_ (.A1(_04805_),
    .A2(net1032),
    .Y(_00095_),
    .B1(_00378_));
 sg13g2_nor2_1 _05717_ (.A(net3),
    .B(net1031),
    .Y(_00379_));
 sg13g2_a21oi_1 _05718_ (.A1(_04806_),
    .A2(net1031),
    .Y(_00096_),
    .B1(_00379_));
 sg13g2_nor2_1 _05719_ (.A(net4),
    .B(net1031),
    .Y(_00380_));
 sg13g2_a21oi_1 _05720_ (.A1(_04807_),
    .A2(net1031),
    .Y(_00097_),
    .B1(_00380_));
 sg13g2_nor2_1 _05721_ (.A(net5),
    .B(net1031),
    .Y(_00381_));
 sg13g2_a21oi_1 _05722_ (.A1(_04808_),
    .A2(net1032),
    .Y(_00098_),
    .B1(_00381_));
 sg13g2_nor2_1 _05723_ (.A(net6),
    .B(net1032),
    .Y(_00382_));
 sg13g2_a21oi_1 _05724_ (.A1(_04809_),
    .A2(net1032),
    .Y(_00099_),
    .B1(_00382_));
 sg13g2_mux2_1 _05725_ (.A0(net7),
    .A1(net1364),
    .S(net1031),
    .X(_00100_));
 sg13g2_nor2_1 _05726_ (.A(net8),
    .B(net1032),
    .Y(_00383_));
 sg13g2_a21oi_1 _05727_ (.A1(_04810_),
    .A2(net1032),
    .Y(_00101_),
    .B1(_00383_));
 sg13g2_nand2_1 _05728_ (.Y(_00384_),
    .A(net1),
    .B(net1099));
 sg13g2_o21ai_1 _05729_ (.B1(_00384_),
    .Y(_00102_),
    .A1(_04835_),
    .A2(net1099));
 sg13g2_nand2_1 _05730_ (.Y(_00385_),
    .A(net2),
    .B(net1099));
 sg13g2_o21ai_1 _05731_ (.B1(_00385_),
    .Y(_00103_),
    .A1(_04836_),
    .A2(net1099));
 sg13g2_mux2_1 _05732_ (.A0(net1338),
    .A1(net3),
    .S(net1100),
    .X(_00104_));
 sg13g2_mux2_1 _05733_ (.A0(net457),
    .A1(net4),
    .S(net1099),
    .X(_00105_));
 sg13g2_mux2_1 _05734_ (.A0(net1332),
    .A1(net5),
    .S(net1099),
    .X(_00106_));
 sg13g2_mux2_1 _05735_ (.A0(net1330),
    .A1(net6),
    .S(net1100),
    .X(_00107_));
 sg13g2_nand2_1 _05736_ (.Y(_00386_),
    .A(net7),
    .B(net1099));
 sg13g2_o21ai_1 _05737_ (.B1(_00386_),
    .Y(_00108_),
    .A1(_04837_),
    .A2(net1099));
 sg13g2_mux2_1 _05738_ (.A0(net1325),
    .A1(net8),
    .S(net1100),
    .X(_00109_));
 sg13g2_nor3_2 _05739_ (.A(_04896_),
    .B(_04956_),
    .C(_04974_),
    .Y(_00387_));
 sg13g2_mux2_1 _05740_ (.A0(net218),
    .A1(\cordic_inst.cordic_state[32] ),
    .S(net1029),
    .X(_00110_));
 sg13g2_mux2_1 _05741_ (.A0(net222),
    .A1(\cordic_inst.cordic_state[33] ),
    .S(net1029),
    .X(_00111_));
 sg13g2_nor2_1 _05742_ (.A(\result_reg[26] ),
    .B(net1029),
    .Y(_00388_));
 sg13g2_a21oi_1 _05743_ (.A1(_04791_),
    .A2(net1029),
    .Y(_00112_),
    .B1(_00388_));
 sg13g2_mux2_1 _05744_ (.A0(net226),
    .A1(\cordic_inst.cordic_state[35] ),
    .S(net1029),
    .X(_00113_));
 sg13g2_mux2_1 _05745_ (.A0(net232),
    .A1(\cordic_inst.cordic_state[36] ),
    .S(net1028),
    .X(_00114_));
 sg13g2_mux2_1 _05746_ (.A0(net245),
    .A1(\cordic_inst.cordic_state[37] ),
    .S(net1028),
    .X(_00115_));
 sg13g2_mux2_1 _05747_ (.A0(net238),
    .A1(\cordic_inst.cordic_state[38] ),
    .S(net1028),
    .X(_00116_));
 sg13g2_nor2_1 _05748_ (.A(net334),
    .B(net1027),
    .Y(_00389_));
 sg13g2_a21oi_1 _05749_ (.A1(_04790_),
    .A2(net1027),
    .Y(_00117_),
    .B1(_00389_));
 sg13g2_mux2_1 _05750_ (.A0(net343),
    .A1(\cordic_inst.cordic_state[40] ),
    .S(net1026),
    .X(_00118_));
 sg13g2_nor2_1 _05751_ (.A(net274),
    .B(net1026),
    .Y(_00390_));
 sg13g2_a21oi_1 _05752_ (.A1(_04789_),
    .A2(net1026),
    .Y(_00119_),
    .B1(_00390_));
 sg13g2_mux2_1 _05753_ (.A0(net336),
    .A1(\cordic_inst.cordic_state[42] ),
    .S(net1026),
    .X(_00120_));
 sg13g2_mux2_1 _05754_ (.A0(net323),
    .A1(\cordic_inst.cordic_state[43] ),
    .S(net1027),
    .X(_00121_));
 sg13g2_mux2_1 _05755_ (.A0(net383),
    .A1(net1249),
    .S(net1026),
    .X(_00122_));
 sg13g2_mux2_1 _05756_ (.A0(net317),
    .A1(net1248),
    .S(net1027),
    .X(_00123_));
 sg13g2_mux2_1 _05757_ (.A0(\result_reg[38] ),
    .A1(net338),
    .S(net1026),
    .X(_00124_));
 sg13g2_mux2_1 _05758_ (.A0(net291),
    .A1(net1246),
    .S(net1027),
    .X(_00125_));
 sg13g2_mux2_1 _05759_ (.A0(net359),
    .A1(net1245),
    .S(net1026),
    .X(_00126_));
 sg13g2_mux2_1 _05760_ (.A0(net357),
    .A1(net1244),
    .S(net1026),
    .X(_00127_));
 sg13g2_mux2_1 _05761_ (.A0(net295),
    .A1(net1243),
    .S(net1028),
    .X(_00128_));
 sg13g2_mux2_1 _05762_ (.A0(net313),
    .A1(net1242),
    .S(net1027),
    .X(_00129_));
 sg13g2_mux2_1 _05763_ (.A0(net269),
    .A1(net1241),
    .S(net1028),
    .X(_00130_));
 sg13g2_mux2_1 _05764_ (.A0(net355),
    .A1(\cordic_inst.cordic_state[53] ),
    .S(net1027),
    .X(_00131_));
 sg13g2_mux2_1 _05765_ (.A0(net265),
    .A1(\cordic_inst.cordic_state[54] ),
    .S(net1028),
    .X(_00132_));
 sg13g2_mux2_1 _05766_ (.A0(net252),
    .A1(net1240),
    .S(net1028),
    .X(_00133_));
 sg13g2_nand2b_1 _05767_ (.Y(_00391_),
    .B(net439),
    .A_N(net1318));
 sg13g2_nand3_1 _05768_ (.B(_04890_),
    .C(net440),
    .A(net1513),
    .Y(_00134_));
 sg13g2_nor2_1 _05769_ (.A(net1268),
    .B(net1273),
    .Y(_00392_));
 sg13g2_or2_1 _05770_ (.X(_00393_),
    .B(net1272),
    .A(net1266));
 sg13g2_nand4_1 _05771_ (.B(_04796_),
    .C(_04915_),
    .A(net1259),
    .Y(_00394_),
    .D(_00392_));
 sg13g2_a21oi_1 _05772_ (.A1(net432),
    .A2(_00394_),
    .Y(_00395_),
    .B1(_04906_));
 sg13g2_nor2_1 _05773_ (.A(net1480),
    .B(net433),
    .Y(_00135_));
 sg13g2_o21ai_1 _05774_ (.B1(_04796_),
    .Y(_00396_),
    .A1(_04797_),
    .A2(_00394_));
 sg13g2_nor2b_1 _05775_ (.A(_04907_),
    .B_N(net493),
    .Y(_00136_));
 sg13g2_and2_1 _05776_ (.A(_04890_),
    .B(net1075),
    .X(_00397_));
 sg13g2_nand2_1 _05777_ (.Y(_00398_),
    .A(_04890_),
    .B(net1075));
 sg13g2_nand2_1 _05778_ (.Y(_00399_),
    .A(net1320),
    .B(net1407));
 sg13g2_nand2_1 _05779_ (.Y(_00400_),
    .A(\cordic_atan2_result[0] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ));
 sg13g2_xnor2_1 _05780_ (.Y(_00401_),
    .A(net413),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ));
 sg13g2_o21ai_1 _05781_ (.B1(_00399_),
    .Y(_00402_),
    .A1(_04911_),
    .A2(_00401_));
 sg13g2_a22oi_1 _05782_ (.Y(_00403_),
    .B1(net1048),
    .B2(_00402_),
    .A2(net1089),
    .A1(net413));
 sg13g2_nor2_1 _05783_ (.A(net1487),
    .B(net414),
    .Y(_00142_));
 sg13g2_nand2b_2 _05784_ (.Y(_00404_),
    .B(\cordic_atan2_result[23] ),
    .A_N(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ));
 sg13g2_nor4_1 _05785_ (.A(net1243),
    .B(net1244),
    .C(net1245),
    .D(net1246),
    .Y(_00405_));
 sg13g2_nor3_1 _05786_ (.A(\cordic_inst.cordic_state[54] ),
    .B(\cordic_inst.cordic_state[53] ),
    .C(\cordic_inst.cordic_state[52] ),
    .Y(_00406_));
 sg13g2_nor3_1 _05787_ (.A(\cordic_inst.cordic_state[34] ),
    .B(\cordic_inst.cordic_state[33] ),
    .C(\cordic_inst.cordic_state[32] ),
    .Y(_00407_));
 sg13g2_nor4_1 _05788_ (.A(\cordic_inst.cordic_state[38] ),
    .B(\cordic_inst.cordic_state[37] ),
    .C(\cordic_inst.cordic_state[36] ),
    .D(\cordic_inst.cordic_state[35] ),
    .Y(_00408_));
 sg13g2_nor4_1 _05789_ (.A(net1251),
    .B(\cordic_inst.cordic_state[41] ),
    .C(\cordic_inst.cordic_state[40] ),
    .D(\cordic_inst.cordic_state[39] ),
    .Y(_00409_));
 sg13g2_nor4_1 _05790_ (.A(net1247),
    .B(\cordic_inst.cordic_state[45] ),
    .C(\cordic_inst.cordic_state[44] ),
    .D(\cordic_inst.cordic_state[43] ),
    .Y(_00410_));
 sg13g2_nand4_1 _05791_ (.B(_00406_),
    .C(_00407_),
    .A(_00405_),
    .Y(_00411_),
    .D(_00408_));
 sg13g2_nand3b_1 _05792_ (.B(_00409_),
    .C(_00410_),
    .Y(_00412_),
    .A_N(net1242));
 sg13g2_nor2b_1 _05793_ (.A(net1240),
    .B_N(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .Y(_00413_));
 sg13g2_o21ai_1 _05794_ (.B1(_00413_),
    .Y(_00414_),
    .A1(_00411_),
    .A2(_00412_));
 sg13g2_and2_1 _05795_ (.A(_00404_),
    .B(_00414_),
    .X(_00415_));
 sg13g2_nand2_2 _05796_ (.Y(_00416_),
    .A(_00404_),
    .B(_00414_));
 sg13g2_nand3_1 _05797_ (.B(_00404_),
    .C(_00414_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .Y(_00417_));
 sg13g2_xor2_1 _05798_ (.B(_00417_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .X(_00418_));
 sg13g2_nand2b_1 _05799_ (.Y(_00419_),
    .B(\cordic_atan2_result[1] ),
    .A_N(_00418_));
 sg13g2_nor2b_1 _05800_ (.A(\cordic_atan2_result[1] ),
    .B_N(_00418_),
    .Y(_00420_));
 sg13g2_xor2_1 _05801_ (.B(_00418_),
    .A(\cordic_atan2_result[1] ),
    .X(_00421_));
 sg13g2_xnor2_1 _05802_ (.Y(_00422_),
    .A(_00400_),
    .B(_00421_));
 sg13g2_a221oi_1 _05803_ (.B2(_00422_),
    .C1(net1047),
    .B1(net1096),
    .A1(net1320),
    .Y(_00423_),
    .A2(_04805_));
 sg13g2_a21oi_1 _05804_ (.A1(net434),
    .A2(net1089),
    .Y(_00424_),
    .B1(_00423_));
 sg13g2_nand2_1 _05805_ (.Y(_00143_),
    .A(net1516),
    .B(net435));
 sg13g2_nand2_1 _05806_ (.Y(_00425_),
    .A(net1320),
    .B(net1392));
 sg13g2_o21ai_1 _05807_ (.B1(_00419_),
    .Y(_00426_),
    .A1(_00400_),
    .A2(_00420_));
 sg13g2_o21ai_1 _05808_ (.B1(net1045),
    .Y(_00427_),
    .A1(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .A2(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ));
 sg13g2_xor2_1 _05809_ (.B(_00427_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .X(_00428_));
 sg13g2_nor2b_1 _05810_ (.A(_00428_),
    .B_N(\cordic_atan2_result[2] ),
    .Y(_00429_));
 sg13g2_xnor2_1 _05811_ (.Y(_00430_),
    .A(\cordic_atan2_result[2] ),
    .B(_00428_));
 sg13g2_and2_1 _05812_ (.A(_00426_),
    .B(_00430_),
    .X(_00431_));
 sg13g2_o21ai_1 _05813_ (.B1(net1096),
    .Y(_00432_),
    .A1(_00426_),
    .A2(_00430_));
 sg13g2_o21ai_1 _05814_ (.B1(_00425_),
    .Y(_00433_),
    .A1(_00431_),
    .A2(_00432_));
 sg13g2_a22oi_1 _05815_ (.Y(_00434_),
    .B1(net1048),
    .B2(_00433_),
    .A2(net1089),
    .A1(net362));
 sg13g2_nor2_1 _05816_ (.A(net1487),
    .B(_00434_),
    .Y(_00144_));
 sg13g2_nor3_1 _05817_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .C(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .Y(_00435_));
 sg13g2_nor2_1 _05818_ (.A(net1040),
    .B(_00435_),
    .Y(_00436_));
 sg13g2_xnor2_1 _05819_ (.Y(_00437_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .B(_00436_));
 sg13g2_nand2b_1 _05820_ (.Y(_00438_),
    .B(\cordic_atan2_result[3] ),
    .A_N(_00437_));
 sg13g2_xor2_1 _05821_ (.B(_00437_),
    .A(\cordic_atan2_result[3] ),
    .X(_00439_));
 sg13g2_a21oi_1 _05822_ (.A1(_00426_),
    .A2(_00430_),
    .Y(_00440_),
    .B1(_00429_));
 sg13g2_xnor2_1 _05823_ (.Y(_00441_),
    .A(_00439_),
    .B(_00440_));
 sg13g2_nand2_1 _05824_ (.Y(_00442_),
    .A(net1097),
    .B(_00441_));
 sg13g2_a21oi_1 _05825_ (.A1(net1320),
    .A2(_04807_),
    .Y(_00443_),
    .B1(net1047));
 sg13g2_a21o_1 _05826_ (.A2(net1090),
    .A1(net500),
    .B1(net1487),
    .X(_00444_));
 sg13g2_a21o_1 _05827_ (.A2(_00443_),
    .A1(_00442_),
    .B1(_00444_),
    .X(_00145_));
 sg13g2_o21ai_1 _05828_ (.B1(_00438_),
    .Y(_00445_),
    .A1(_00439_),
    .A2(_00440_));
 sg13g2_nor2b_1 _05829_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .B_N(_00435_),
    .Y(_00446_));
 sg13g2_nor2_1 _05830_ (.A(net1040),
    .B(_00446_),
    .Y(_00447_));
 sg13g2_xnor2_1 _05831_ (.Y(_00448_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .B(_00447_));
 sg13g2_nor2b_1 _05832_ (.A(_00448_),
    .B_N(\cordic_atan2_result[4] ),
    .Y(_00449_));
 sg13g2_xnor2_1 _05833_ (.Y(_00450_),
    .A(\cordic_atan2_result[4] ),
    .B(_00448_));
 sg13g2_o21ai_1 _05834_ (.B1(net1097),
    .Y(_00451_),
    .A1(_00445_),
    .A2(_00450_));
 sg13g2_a21oi_1 _05835_ (.A1(_00445_),
    .A2(_00450_),
    .Y(_00452_),
    .B1(_00451_));
 sg13g2_a21o_1 _05836_ (.A2(net1377),
    .A1(net1319),
    .B1(_00452_),
    .X(_00453_));
 sg13g2_a22oi_1 _05837_ (.Y(_00454_),
    .B1(net1048),
    .B2(_00453_),
    .A2(net1089),
    .A1(net361));
 sg13g2_nor2_1 _05838_ (.A(net1487),
    .B(_00454_),
    .Y(_00146_));
 sg13g2_a21oi_1 _05839_ (.A1(_00445_),
    .A2(_00450_),
    .Y(_00455_),
    .B1(_00449_));
 sg13g2_nor2b_1 _05840_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .B_N(_00446_),
    .Y(_00456_));
 sg13g2_nor2_1 _05841_ (.A(net1040),
    .B(_00456_),
    .Y(_00457_));
 sg13g2_xor2_1 _05842_ (.B(_00457_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .X(_00458_));
 sg13g2_nand2_1 _05843_ (.Y(_00459_),
    .A(\cordic_atan2_result[5] ),
    .B(_00458_));
 sg13g2_xnor2_1 _05844_ (.Y(_00460_),
    .A(\cordic_atan2_result[5] ),
    .B(_00458_));
 sg13g2_xnor2_1 _05845_ (.Y(_00461_),
    .A(_00455_),
    .B(_00460_));
 sg13g2_a221oi_1 _05846_ (.B2(_00461_),
    .C1(net1047),
    .B1(net1096),
    .A1(net1319),
    .Y(_00462_),
    .A2(_04809_));
 sg13g2_a21oi_1 _05847_ (.A1(net398),
    .A2(net1090),
    .Y(_00463_),
    .B1(_00462_));
 sg13g2_nand2_1 _05848_ (.Y(_00147_),
    .A(net1516),
    .B(_00463_));
 sg13g2_o21ai_1 _05849_ (.B1(_00459_),
    .Y(_00464_),
    .A1(_00455_),
    .A2(_00460_));
 sg13g2_nor2b_1 _05850_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .B_N(_00456_),
    .Y(_00465_));
 sg13g2_nor2_1 _05851_ (.A(net1040),
    .B(_00465_),
    .Y(_00466_));
 sg13g2_xnor2_1 _05852_ (.Y(_00467_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .B(_00466_));
 sg13g2_nor2b_1 _05853_ (.A(_00467_),
    .B_N(\cordic_atan2_result[6] ),
    .Y(_00468_));
 sg13g2_xnor2_1 _05854_ (.Y(_00469_),
    .A(\cordic_atan2_result[6] ),
    .B(_00467_));
 sg13g2_o21ai_1 _05855_ (.B1(net1097),
    .Y(_00470_),
    .A1(_00464_),
    .A2(_00469_));
 sg13g2_a21oi_1 _05856_ (.A1(_00464_),
    .A2(_00469_),
    .Y(_00471_),
    .B1(_00470_));
 sg13g2_a21o_1 _05857_ (.A2(net1363),
    .A1(net1319),
    .B1(_00471_),
    .X(_00472_));
 sg13g2_a22oi_1 _05858_ (.Y(_00473_),
    .B1(net1048),
    .B2(_00472_),
    .A2(net1090),
    .A1(net376));
 sg13g2_nor2_1 _05859_ (.A(net1487),
    .B(_00473_),
    .Y(_00148_));
 sg13g2_a21oi_1 _05860_ (.A1(_00464_),
    .A2(_00469_),
    .Y(_00474_),
    .B1(_00468_));
 sg13g2_nor2b_1 _05861_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .B_N(_00465_),
    .Y(_00475_));
 sg13g2_nor2_1 _05862_ (.A(net1040),
    .B(_00475_),
    .Y(_00476_));
 sg13g2_xor2_1 _05863_ (.B(_00476_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ),
    .X(_00477_));
 sg13g2_nand2_1 _05864_ (.Y(_00478_),
    .A(\cordic_atan2_result[7] ),
    .B(_00477_));
 sg13g2_xnor2_1 _05865_ (.Y(_00479_),
    .A(\cordic_atan2_result[7] ),
    .B(_00477_));
 sg13g2_xnor2_1 _05866_ (.Y(_00480_),
    .A(_00474_),
    .B(_00479_));
 sg13g2_a221oi_1 _05867_ (.B2(_00480_),
    .C1(net1047),
    .B1(net1096),
    .A1(net1319),
    .Y(_00481_),
    .A2(_04810_));
 sg13g2_a21oi_1 _05868_ (.A1(net400),
    .A2(net1090),
    .Y(_00482_),
    .B1(_00481_));
 sg13g2_nand2_1 _05869_ (.Y(_00149_),
    .A(net1516),
    .B(_00482_));
 sg13g2_nand2_1 _05870_ (.Y(_00483_),
    .A(net1319),
    .B(net1473));
 sg13g2_o21ai_1 _05871_ (.B1(_00478_),
    .Y(_00484_),
    .A1(_00474_),
    .A2(_00479_));
 sg13g2_nand2b_1 _05872_ (.Y(_00485_),
    .B(_00475_),
    .A_N(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ));
 sg13g2_nand2_1 _05873_ (.Y(_00486_),
    .A(net1045),
    .B(_00485_));
 sg13g2_xor2_1 _05874_ (.B(_00486_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .X(_00487_));
 sg13g2_nor2b_1 _05875_ (.A(_00487_),
    .B_N(\cordic_atan2_result[8] ),
    .Y(_00488_));
 sg13g2_xnor2_1 _05876_ (.Y(_00489_),
    .A(\cordic_atan2_result[8] ),
    .B(_00487_));
 sg13g2_and2_1 _05877_ (.A(_00484_),
    .B(_00489_),
    .X(_00490_));
 sg13g2_o21ai_1 _05878_ (.B1(net1096),
    .Y(_00491_),
    .A1(_00484_),
    .A2(_00489_));
 sg13g2_o21ai_1 _05879_ (.B1(_00483_),
    .Y(_00492_),
    .A1(_00490_),
    .A2(_00491_));
 sg13g2_a22oi_1 _05880_ (.Y(_00493_),
    .B1(net1048),
    .B2(_00492_),
    .A2(net1089),
    .A1(net351));
 sg13g2_nor2_1 _05881_ (.A(net1487),
    .B(_00493_),
    .Y(_00150_));
 sg13g2_a21oi_1 _05882_ (.A1(_00484_),
    .A2(_00489_),
    .Y(_00494_),
    .B1(_00488_));
 sg13g2_o21ai_1 _05883_ (.B1(net1045),
    .Y(_00495_),
    .A1(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .A2(_00485_));
 sg13g2_xor2_1 _05884_ (.B(_00495_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .X(_00496_));
 sg13g2_inv_1 _05885_ (.Y(_00497_),
    .A(_00496_));
 sg13g2_nand2b_1 _05886_ (.Y(_00498_),
    .B(_00496_),
    .A_N(\cordic_atan2_result[9] ));
 sg13g2_inv_1 _05887_ (.Y(_00499_),
    .A(_00498_));
 sg13g2_xor2_1 _05888_ (.B(_00496_),
    .A(\cordic_atan2_result[9] ),
    .X(_00500_));
 sg13g2_xnor2_1 _05889_ (.Y(_00501_),
    .A(_00494_),
    .B(_00500_));
 sg13g2_a221oi_1 _05890_ (.B2(_00501_),
    .C1(net1047),
    .B1(net1096),
    .A1(net1319),
    .Y(_00502_),
    .A2(_04812_));
 sg13g2_a21oi_1 _05891_ (.A1(net437),
    .A2(net1089),
    .Y(_00503_),
    .B1(_00502_));
 sg13g2_nand2_1 _05892_ (.Y(_00151_),
    .A(net1518),
    .B(net438));
 sg13g2_nand2_1 _05893_ (.Y(_00504_),
    .A(net1319),
    .B(net1464));
 sg13g2_nor3_1 _05894_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .C(_00485_),
    .Y(_00505_));
 sg13g2_nor2_1 _05895_ (.A(_00416_),
    .B(_00505_),
    .Y(_00506_));
 sg13g2_xnor2_1 _05896_ (.Y(_00507_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ),
    .B(_00506_));
 sg13g2_nor2b_1 _05897_ (.A(_00507_),
    .B_N(\cordic_atan2_result[10] ),
    .Y(_00508_));
 sg13g2_xnor2_1 _05898_ (.Y(_00509_),
    .A(\cordic_atan2_result[10] ),
    .B(_00507_));
 sg13g2_inv_1 _05899_ (.Y(_00510_),
    .A(_00509_));
 sg13g2_a221oi_1 _05900_ (.B2(\cordic_atan2_result[9] ),
    .C1(_00488_),
    .B1(_00497_),
    .A1(_00484_),
    .Y(_00511_),
    .A2(_00489_));
 sg13g2_nor3_1 _05901_ (.A(_00499_),
    .B(_00510_),
    .C(_00511_),
    .Y(_00512_));
 sg13g2_o21ai_1 _05902_ (.B1(_00510_),
    .Y(_00513_),
    .A1(_00499_),
    .A2(_00511_));
 sg13g2_nand2_1 _05903_ (.Y(_00514_),
    .A(net1096),
    .B(_00513_));
 sg13g2_o21ai_1 _05904_ (.B1(_00504_),
    .Y(_00515_),
    .A1(_00512_),
    .A2(_00514_));
 sg13g2_a22oi_1 _05905_ (.Y(_00516_),
    .B1(_00397_),
    .B2(_00515_),
    .A2(net1089),
    .A1(net380));
 sg13g2_nor2_1 _05906_ (.A(net1487),
    .B(_00516_),
    .Y(_00152_));
 sg13g2_nor2_1 _05907_ (.A(_00508_),
    .B(_00512_),
    .Y(_00517_));
 sg13g2_nand2b_1 _05908_ (.Y(_00518_),
    .B(_00505_),
    .A_N(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ));
 sg13g2_nand2_1 _05909_ (.Y(_00519_),
    .A(net1045),
    .B(_00518_));
 sg13g2_xor2_1 _05910_ (.B(_00519_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .X(_00520_));
 sg13g2_nor2b_1 _05911_ (.A(_00520_),
    .B_N(\cordic_atan2_result[11] ),
    .Y(_00521_));
 sg13g2_nor2b_1 _05912_ (.A(\cordic_atan2_result[11] ),
    .B_N(_00520_),
    .Y(_00522_));
 sg13g2_inv_1 _05913_ (.Y(_00523_),
    .A(_00522_));
 sg13g2_nor2_1 _05914_ (.A(_00521_),
    .B(_00522_),
    .Y(_00524_));
 sg13g2_xor2_1 _05915_ (.B(_00524_),
    .A(_00517_),
    .X(_00525_));
 sg13g2_a221oi_1 _05916_ (.B2(_00525_),
    .C1(net1047),
    .B1(net1096),
    .A1(net1319),
    .Y(_00526_),
    .A2(_04814_));
 sg13g2_a21oi_1 _05917_ (.A1(net405),
    .A2(net1089),
    .Y(_00527_),
    .B1(_00526_));
 sg13g2_nand2_1 _05918_ (.Y(_00153_),
    .A(net1516),
    .B(_00527_));
 sg13g2_nor2_2 _05919_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .B(_00518_),
    .Y(_00528_));
 sg13g2_nor2_2 _05920_ (.A(_00416_),
    .B(_00528_),
    .Y(_00529_));
 sg13g2_and2_1 _05921_ (.A(\cordic_atan2_result[12] ),
    .B(_00529_),
    .X(_00530_));
 sg13g2_xnor2_1 _05922_ (.Y(_00531_),
    .A(\cordic_atan2_result[12] ),
    .B(_00529_));
 sg13g2_inv_1 _05923_ (.Y(_00532_),
    .A(_00531_));
 sg13g2_or3_1 _05924_ (.A(_00508_),
    .B(_00512_),
    .C(_00521_),
    .X(_00533_));
 sg13g2_a21oi_1 _05925_ (.A1(_00523_),
    .A2(_00533_),
    .Y(_00534_),
    .B1(_00532_));
 sg13g2_and3_2 _05926_ (.X(_00535_),
    .A(_00523_),
    .B(_00532_),
    .C(_00533_));
 sg13g2_nor3_1 _05927_ (.A(_04911_),
    .B(_00534_),
    .C(_00535_),
    .Y(_00536_));
 sg13g2_a21oi_1 _05928_ (.A1(net1321),
    .A2(net1453),
    .Y(_00537_),
    .B1(_00536_));
 sg13g2_nor2_1 _05929_ (.A(net1047),
    .B(_00537_),
    .Y(_00538_));
 sg13g2_a21oi_1 _05930_ (.A1(net372),
    .A2(net1091),
    .Y(_00539_),
    .B1(_00538_));
 sg13g2_nor2_1 _05931_ (.A(net1483),
    .B(net373),
    .Y(_00154_));
 sg13g2_nor2_1 _05932_ (.A(_00530_),
    .B(_00535_),
    .Y(_00540_));
 sg13g2_nor2_1 _05933_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .B(_00529_),
    .Y(_00541_));
 sg13g2_nand2_1 _05934_ (.Y(_00542_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .B(net1045));
 sg13g2_nor2_1 _05935_ (.A(_00528_),
    .B(_00542_),
    .Y(_00543_));
 sg13g2_nor2_1 _05936_ (.A(_00541_),
    .B(_00543_),
    .Y(_00544_));
 sg13g2_or2_1 _05937_ (.X(_00545_),
    .B(_00544_),
    .A(\cordic_atan2_result[13] ));
 sg13g2_nand2_1 _05938_ (.Y(_00546_),
    .A(\cordic_atan2_result[13] ),
    .B(_00544_));
 sg13g2_nand2_1 _05939_ (.Y(_00547_),
    .A(_00545_),
    .B(_00546_));
 sg13g2_xor2_1 _05940_ (.B(_00547_),
    .A(_00540_),
    .X(_00548_));
 sg13g2_a21oi_1 _05941_ (.A1(net1321),
    .A2(_04816_),
    .Y(_00549_),
    .B1(net1046));
 sg13g2_o21ai_1 _05942_ (.B1(_00549_),
    .Y(_00550_),
    .A1(_04911_),
    .A2(_00548_));
 sg13g2_a21oi_1 _05943_ (.A1(net401),
    .A2(net1092),
    .Y(_00551_),
    .B1(net1483));
 sg13g2_nand2_1 _05944_ (.Y(_00155_),
    .A(_00550_),
    .B(_00551_));
 sg13g2_o21ai_1 _05945_ (.B1(_00542_),
    .Y(_00552_),
    .A1(_00416_),
    .A2(_00528_));
 sg13g2_nand2_1 _05946_ (.Y(_00553_),
    .A(\cordic_atan2_result[14] ),
    .B(_00552_));
 sg13g2_xor2_1 _05947_ (.B(net1020),
    .A(\cordic_atan2_result[14] ),
    .X(_00554_));
 sg13g2_inv_1 _05948_ (.Y(_00555_),
    .A(_00554_));
 sg13g2_o21ai_1 _05949_ (.B1(_00545_),
    .Y(_00556_),
    .A1(_00530_),
    .A2(_00535_));
 sg13g2_and3_1 _05950_ (.X(_00557_),
    .A(_00546_),
    .B(_00555_),
    .C(_00556_));
 sg13g2_a21o_1 _05951_ (.A2(_00556_),
    .A1(_00546_),
    .B1(_00555_),
    .X(_00558_));
 sg13g2_nor2_1 _05952_ (.A(_04911_),
    .B(_00557_),
    .Y(_00559_));
 sg13g2_a22oi_1 _05953_ (.Y(_00560_),
    .B1(_00558_),
    .B2(_00559_),
    .A2(net1443),
    .A1(net1321));
 sg13g2_nor2_1 _05954_ (.A(net1046),
    .B(_00560_),
    .Y(_00561_));
 sg13g2_a21oi_1 _05955_ (.A1(net321),
    .A2(net1092),
    .Y(_00562_),
    .B1(_00561_));
 sg13g2_nor2_1 _05956_ (.A(net1482),
    .B(net322),
    .Y(_00156_));
 sg13g2_and2_1 _05957_ (.A(_00553_),
    .B(_00558_),
    .X(_00563_));
 sg13g2_nor2b_2 _05958_ (.A(_00541_),
    .B_N(_00542_),
    .Y(_00564_));
 sg13g2_nor2_1 _05959_ (.A(\cordic_atan2_result[15] ),
    .B(net1019),
    .Y(_00565_));
 sg13g2_nand2_1 _05960_ (.Y(_00566_),
    .A(\cordic_atan2_result[15] ),
    .B(_00564_));
 sg13g2_nand2b_1 _05961_ (.Y(_00567_),
    .B(_00566_),
    .A_N(_00565_));
 sg13g2_xnor2_1 _05962_ (.Y(_00568_),
    .A(_00563_),
    .B(_00567_));
 sg13g2_a221oi_1 _05963_ (.B2(_00568_),
    .C1(net1046),
    .B1(net1098),
    .A1(net1321),
    .Y(_00569_),
    .A2(_04817_));
 sg13g2_a21oi_1 _05964_ (.A1(net409),
    .A2(net1092),
    .Y(_00570_),
    .B1(_00569_));
 sg13g2_nand2_1 _05965_ (.Y(_00157_),
    .A(net1509),
    .B(net410));
 sg13g2_nand2_1 _05966_ (.Y(_00571_),
    .A(net1321),
    .B(net1434));
 sg13g2_and2_1 _05967_ (.A(\cordic_atan2_result[16] ),
    .B(_00552_),
    .X(_00572_));
 sg13g2_xor2_1 _05968_ (.B(_00552_),
    .A(\cordic_atan2_result[16] ),
    .X(_00573_));
 sg13g2_a21oi_1 _05969_ (.A1(_00563_),
    .A2(_00566_),
    .Y(_00574_),
    .B1(_00565_));
 sg13g2_and2_1 _05970_ (.A(_00573_),
    .B(_00574_),
    .X(_00575_));
 sg13g2_o21ai_1 _05971_ (.B1(net1098),
    .Y(_00576_),
    .A1(_00573_),
    .A2(_00574_));
 sg13g2_o21ai_1 _05972_ (.B1(_00571_),
    .Y(_00577_),
    .A1(_00575_),
    .A2(_00576_));
 sg13g2_a22oi_1 _05973_ (.Y(_00578_),
    .B1(net1048),
    .B2(_00577_),
    .A2(net1092),
    .A1(net403));
 sg13g2_nor2_1 _05974_ (.A(net1484),
    .B(net404),
    .Y(_00158_));
 sg13g2_nor2_1 _05975_ (.A(_00572_),
    .B(_00575_),
    .Y(_00579_));
 sg13g2_nor2_1 _05976_ (.A(\cordic_atan2_result[17] ),
    .B(net1019),
    .Y(_00580_));
 sg13g2_xnor2_1 _05977_ (.Y(_00581_),
    .A(\cordic_atan2_result[17] ),
    .B(net1019));
 sg13g2_xnor2_1 _05978_ (.Y(_00582_),
    .A(_00579_),
    .B(_00581_));
 sg13g2_a221oi_1 _05979_ (.B2(_00582_),
    .C1(net1046),
    .B1(net1098),
    .A1(net1317),
    .Y(_00583_),
    .A2(_04818_));
 sg13g2_a21oi_1 _05980_ (.A1(net448),
    .A2(net1092),
    .Y(_00584_),
    .B1(_00583_));
 sg13g2_nand2_1 _05981_ (.Y(_00159_),
    .A(net1508),
    .B(net449));
 sg13g2_nand2_1 _05982_ (.Y(_00585_),
    .A(\cordic_atan2_result[18] ),
    .B(net1020));
 sg13g2_nor2_1 _05983_ (.A(\cordic_atan2_result[18] ),
    .B(net1020),
    .Y(_00586_));
 sg13g2_xor2_1 _05984_ (.B(net1020),
    .A(\cordic_atan2_result[18] ),
    .X(_00587_));
 sg13g2_a221oi_1 _05985_ (.B2(_00574_),
    .C1(_00572_),
    .B1(_00573_),
    .A1(\cordic_atan2_result[17] ),
    .Y(_00588_),
    .A2(net1019));
 sg13g2_or2_1 _05986_ (.X(_00589_),
    .B(_00588_),
    .A(_00580_));
 sg13g2_inv_1 _05987_ (.Y(_00590_),
    .A(_00589_));
 sg13g2_o21ai_1 _05988_ (.B1(net1098),
    .Y(_00591_),
    .A1(_00587_),
    .A2(_00590_));
 sg13g2_a21oi_1 _05989_ (.A1(_00587_),
    .A2(_00590_),
    .Y(_00592_),
    .B1(_00591_));
 sg13g2_a21o_1 _05990_ (.A2(net1426),
    .A1(net1317),
    .B1(_00592_),
    .X(_00593_));
 sg13g2_a22oi_1 _05991_ (.Y(_00594_),
    .B1(net1048),
    .B2(_00593_),
    .A2(net1088),
    .A1(net425));
 sg13g2_nor2_1 _05992_ (.A(net1482),
    .B(net426),
    .Y(_00160_));
 sg13g2_o21ai_1 _05993_ (.B1(_00585_),
    .Y(_00595_),
    .A1(_00586_),
    .A2(_00589_));
 sg13g2_and2_1 _05994_ (.A(\cordic_atan2_result[19] ),
    .B(net1019),
    .X(_00596_));
 sg13g2_or2_1 _05995_ (.X(_00597_),
    .B(net1019),
    .A(\cordic_atan2_result[19] ));
 sg13g2_nor2b_1 _05996_ (.A(_00596_),
    .B_N(_00597_),
    .Y(_00598_));
 sg13g2_xnor2_1 _05997_ (.Y(_00599_),
    .A(_00595_),
    .B(_00598_));
 sg13g2_a221oi_1 _05998_ (.B2(_00599_),
    .C1(net1046),
    .B1(net1098),
    .A1(net1317),
    .Y(_00600_),
    .A2(_04819_));
 sg13g2_a21oi_1 _05999_ (.A1(net395),
    .A2(net1088),
    .Y(_00601_),
    .B1(_00600_));
 sg13g2_nand2_1 _06000_ (.Y(_00161_),
    .A(net1506),
    .B(net396));
 sg13g2_nand2_1 _06001_ (.Y(_00602_),
    .A(net1317),
    .B(net1420));
 sg13g2_nand2_1 _06002_ (.Y(_00603_),
    .A(\cordic_atan2_result[20] ),
    .B(net1020));
 sg13g2_xor2_1 _06003_ (.B(net1020),
    .A(\cordic_atan2_result[20] ),
    .X(_00604_));
 sg13g2_inv_1 _06004_ (.Y(_00605_),
    .A(_00604_));
 sg13g2_a21oi_1 _06005_ (.A1(_00595_),
    .A2(_00597_),
    .Y(_00606_),
    .B1(_00596_));
 sg13g2_a21oi_1 _06006_ (.A1(_00605_),
    .A2(_00606_),
    .Y(_00607_),
    .B1(_04911_));
 sg13g2_o21ai_1 _06007_ (.B1(_00607_),
    .Y(_00608_),
    .A1(_00605_),
    .A2(_00606_));
 sg13g2_a21oi_1 _06008_ (.A1(_00602_),
    .A2(_00608_),
    .Y(_00609_),
    .B1(net1046));
 sg13g2_a21oi_1 _06009_ (.A1(net349),
    .A2(net1088),
    .Y(_00610_),
    .B1(_00609_));
 sg13g2_nor2_1 _06010_ (.A(net1482),
    .B(net350),
    .Y(_00162_));
 sg13g2_o21ai_1 _06011_ (.B1(_00603_),
    .Y(_00611_),
    .A1(_00605_),
    .A2(_00606_));
 sg13g2_and2_1 _06012_ (.A(\cordic_atan2_result[21] ),
    .B(net1019),
    .X(_00612_));
 sg13g2_or2_1 _06013_ (.X(_00613_),
    .B(net1019),
    .A(\cordic_atan2_result[21] ));
 sg13g2_nor2b_1 _06014_ (.A(_00612_),
    .B_N(_00613_),
    .Y(_00614_));
 sg13g2_xnor2_1 _06015_ (.Y(_00615_),
    .A(_00611_),
    .B(_00614_));
 sg13g2_a221oi_1 _06016_ (.B2(_00615_),
    .C1(net1046),
    .B1(net1098),
    .A1(net1317),
    .Y(_00616_),
    .A2(_04820_));
 sg13g2_a21oi_1 _06017_ (.A1(net389),
    .A2(net1088),
    .Y(_00617_),
    .B1(_00616_));
 sg13g2_nand2_1 _06018_ (.Y(_00163_),
    .A(net1507),
    .B(net390));
 sg13g2_nand2_1 _06019_ (.Y(_00618_),
    .A(net1317),
    .B(net1414));
 sg13g2_xnor2_1 _06020_ (.Y(_00619_),
    .A(\cordic_atan2_result[22] ),
    .B(net1020));
 sg13g2_a21oi_1 _06021_ (.A1(_00611_),
    .A2(_00613_),
    .Y(_00620_),
    .B1(_00612_));
 sg13g2_nor2_1 _06022_ (.A(_00619_),
    .B(_00620_),
    .Y(_00621_));
 sg13g2_a21o_1 _06023_ (.A2(_00620_),
    .A1(_00619_),
    .B1(_04911_),
    .X(_00622_));
 sg13g2_o21ai_1 _06024_ (.B1(_00618_),
    .Y(_00623_),
    .A1(_00621_),
    .A2(_00622_));
 sg13g2_a22oi_1 _06025_ (.Y(_00624_),
    .B1(net1048),
    .B2(_00623_),
    .A2(net1088),
    .A1(net421));
 sg13g2_nor2_1 _06026_ (.A(net1483),
    .B(net422),
    .Y(_00164_));
 sg13g2_a21oi_1 _06027_ (.A1(net421),
    .A2(net1020),
    .Y(_00625_),
    .B1(_00621_));
 sg13g2_xor2_1 _06028_ (.B(_00564_),
    .A(net458),
    .X(_00626_));
 sg13g2_xnor2_1 _06029_ (.Y(_00627_),
    .A(_00625_),
    .B(_00626_));
 sg13g2_a21oi_1 _06030_ (.A1(net1317),
    .A2(_04822_),
    .Y(_00628_),
    .B1(net1046));
 sg13g2_o21ai_1 _06031_ (.B1(_00628_),
    .Y(_00629_),
    .A1(_04911_),
    .A2(_00627_));
 sg13g2_a21oi_1 _06032_ (.A1(net458),
    .A2(net1088),
    .Y(_00630_),
    .B1(net1482));
 sg13g2_nand2_1 _06033_ (.Y(_00165_),
    .A(_00629_),
    .B(_00630_));
 sg13g2_mux4_1 _06034_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[68] ),
    .A1(\cordic_inst.cordic_state[69] ),
    .A2(\cordic_inst.cordic_state[70] ),
    .A3(\cordic_inst.cordic_state[71] ),
    .S1(net1277),
    .X(_00631_));
 sg13g2_mux4_1 _06035_ (.S0(net1288),
    .A0(\cordic_inst.cordic_state[64] ),
    .A1(\cordic_inst.cordic_state[65] ),
    .A2(\cordic_inst.cordic_state[66] ),
    .A3(net1236),
    .S1(net1279),
    .X(_00632_));
 sg13g2_mux2_1 _06036_ (.A0(_00631_),
    .A1(_00632_),
    .S(net1133),
    .X(_00633_));
 sg13g2_nand2b_1 _06037_ (.Y(_00634_),
    .B(\cordic_inst.cordic_state[56] ),
    .A_N(net1289));
 sg13g2_a21oi_1 _06038_ (.A1(\cordic_inst.cordic_state[57] ),
    .A2(net1289),
    .Y(_00635_),
    .B1(net1279));
 sg13g2_mux2_1 _06039_ (.A0(\cordic_inst.cordic_state[58] ),
    .A1(\cordic_inst.cordic_state[59] ),
    .S(net1289),
    .X(_00636_));
 sg13g2_a21oi_1 _06040_ (.A1(_00634_),
    .A2(_00635_),
    .Y(_00637_),
    .B1(net1120));
 sg13g2_o21ai_1 _06041_ (.B1(_00637_),
    .Y(_00638_),
    .A1(net1131),
    .A2(_00636_));
 sg13g2_nor2_2 _06042_ (.A(net1267),
    .B(net1133),
    .Y(_00639_));
 sg13g2_nand2b_2 _06043_ (.Y(_00640_),
    .B(net1269),
    .A_N(net1264));
 sg13g2_mux2_1 _06044_ (.A0(\cordic_inst.cordic_state[62] ),
    .A1(\cordic_inst.cordic_state[63] ),
    .S(net1289),
    .X(_00641_));
 sg13g2_mux2_1 _06045_ (.A0(\cordic_inst.cordic_state[60] ),
    .A1(\cordic_inst.cordic_state[61] ),
    .S(net1289),
    .X(_00642_));
 sg13g2_mux2_1 _06046_ (.A0(_00641_),
    .A1(_00642_),
    .S(net1131),
    .X(_00643_));
 sg13g2_a22oi_1 _06047_ (.Y(_00644_),
    .B1(_00639_),
    .B2(_00643_),
    .A2(_00633_),
    .A1(net1266));
 sg13g2_a21o_1 _06048_ (.A2(_00644_),
    .A1(_00638_),
    .B1(net1257),
    .X(_00645_));
 sg13g2_mux2_1 _06049_ (.A0(\cordic_inst.cordic_state[78] ),
    .A1(net1230),
    .S(net1282),
    .X(_00646_));
 sg13g2_mux4_1 _06050_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[76] ),
    .A1(net1234),
    .A2(\cordic_inst.cordic_state[78] ),
    .A3(net1232),
    .S1(net1277),
    .X(_00647_));
 sg13g2_mux4_1 _06051_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[72] ),
    .A1(net1235),
    .A2(\cordic_inst.cordic_state[74] ),
    .A3(\cordic_inst.cordic_state[75] ),
    .S1(net1278),
    .X(_00648_));
 sg13g2_mux2_1 _06052_ (.A0(_00647_),
    .A1(_00648_),
    .S(net1133),
    .X(_00649_));
 sg13g2_and2_1 _06053_ (.A(net1135),
    .B(_00649_),
    .X(_00650_));
 sg13g2_nor2_2 _06054_ (.A(_04783_),
    .B(net1139),
    .Y(_00651_));
 sg13g2_nand2_1 _06055_ (.Y(_00652_),
    .A(_04929_),
    .B(_00651_));
 sg13g2_a22oi_1 _06056_ (.Y(_00653_),
    .B1(_00651_),
    .B2(_04929_),
    .A2(_00650_),
    .A1(net1256));
 sg13g2_and2_1 _06057_ (.A(_00645_),
    .B(_00653_),
    .X(_00654_));
 sg13g2_nor2_1 _06058_ (.A(\cordic_inst.cordic_state[32] ),
    .B(_00654_),
    .Y(_00655_));
 sg13g2_xor2_1 _06059_ (.B(_00654_),
    .A(net463),
    .X(_00656_));
 sg13g2_a221oi_1 _06060_ (.B2(net1408),
    .C1(net1085),
    .B1(net1125),
    .A1(net1310),
    .Y(_00657_),
    .A2(net1227));
 sg13g2_o21ai_1 _06061_ (.B1(_00657_),
    .Y(_00658_),
    .A1(net1049),
    .A2(_00656_));
 sg13g2_o21ai_1 _06062_ (.B1(_00658_),
    .Y(_00659_),
    .A1(net463),
    .A2(net1076));
 sg13g2_nor2_1 _06063_ (.A(net1480),
    .B(_00659_),
    .Y(_00166_));
 sg13g2_mux2_1 _06064_ (.A0(net1234),
    .A1(\cordic_inst.cordic_state[78] ),
    .S(net1286),
    .X(_00660_));
 sg13g2_nor2b_2 _06065_ (.A(net1286),
    .B_N(net1276),
    .Y(_00661_));
 sg13g2_a22oi_1 _06066_ (.Y(_00662_),
    .B1(_00661_),
    .B2(net1231),
    .A2(_00660_),
    .A1(net1129));
 sg13g2_a221oi_1 _06067_ (.B2(net1231),
    .C1(net1132),
    .B1(_00661_),
    .A1(net1129),
    .Y(_00663_),
    .A2(_00660_));
 sg13g2_mux4_1 _06068_ (.S0(net1287),
    .A0(net1235),
    .A1(\cordic_inst.cordic_state[74] ),
    .A2(\cordic_inst.cordic_state[75] ),
    .A3(\cordic_inst.cordic_state[76] ),
    .S1(net1277),
    .X(_00664_));
 sg13g2_nor2_1 _06069_ (.A(net1271),
    .B(_00664_),
    .Y(_00665_));
 sg13g2_or3_1 _06070_ (.A(net1262),
    .B(_00663_),
    .C(_00665_),
    .X(_00666_));
 sg13g2_mux4_1 _06071_ (.S0(net1288),
    .A0(\cordic_inst.cordic_state[65] ),
    .A1(\cordic_inst.cordic_state[66] ),
    .A2(net1236),
    .A3(\cordic_inst.cordic_state[68] ),
    .S1(net1277),
    .X(_00667_));
 sg13g2_mux4_1 _06072_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[69] ),
    .A1(\cordic_inst.cordic_state[70] ),
    .A2(\cordic_inst.cordic_state[71] ),
    .A3(\cordic_inst.cordic_state[72] ),
    .S1(net1277),
    .X(_00668_));
 sg13g2_mux2_1 _06073_ (.A0(_00667_),
    .A1(_00668_),
    .S(net1272),
    .X(_00669_));
 sg13g2_mux4_1 _06074_ (.S0(net1289),
    .A0(\cordic_inst.cordic_state[61] ),
    .A1(\cordic_inst.cordic_state[62] ),
    .A2(\cordic_inst.cordic_state[63] ),
    .A3(\cordic_inst.cordic_state[64] ),
    .S1(net1279),
    .X(_00670_));
 sg13g2_mux4_1 _06075_ (.S0(net1290),
    .A0(\cordic_inst.cordic_state[57] ),
    .A1(\cordic_inst.cordic_state[58] ),
    .A2(\cordic_inst.cordic_state[59] ),
    .A3(\cordic_inst.cordic_state[60] ),
    .S1(net1279),
    .X(_00671_));
 sg13g2_mux4_1 _06076_ (.S0(net1272),
    .A0(_00667_),
    .A1(_00668_),
    .A2(_00671_),
    .A3(_00670_),
    .S1(net1136),
    .X(_00672_));
 sg13g2_nor2_1 _06077_ (.A(net1259),
    .B(_00672_),
    .Y(_00673_));
 sg13g2_a21o_1 _06078_ (.A2(_00666_),
    .A1(net1256),
    .B1(_00673_),
    .X(_00674_));
 sg13g2_and2_1 _06079_ (.A(_00652_),
    .B(_00674_),
    .X(_00675_));
 sg13g2_a21oi_1 _06080_ (.A1(_00645_),
    .A2(_00653_),
    .Y(_00676_),
    .B1(net1039));
 sg13g2_xor2_1 _06081_ (.B(_00676_),
    .A(_00675_),
    .X(_00677_));
 sg13g2_nand2_1 _06082_ (.Y(_00678_),
    .A(\cordic_inst.cordic_state[33] ),
    .B(_00677_));
 sg13g2_nor2_1 _06083_ (.A(\cordic_inst.cordic_state[33] ),
    .B(_00677_),
    .Y(_00679_));
 sg13g2_xnor2_1 _06084_ (.Y(_00680_),
    .A(\cordic_inst.cordic_state[33] ),
    .B(_00677_));
 sg13g2_xnor2_1 _06085_ (.Y(_00681_),
    .A(_00655_),
    .B(_00680_));
 sg13g2_a221oi_1 _06086_ (.B2(net1402),
    .C1(net1084),
    .B1(net1125),
    .A1(net1307),
    .Y(_00682_),
    .A2(net1223));
 sg13g2_o21ai_1 _06087_ (.B1(_00682_),
    .Y(_00683_),
    .A1(_04906_),
    .A2(_00681_));
 sg13g2_o21ai_1 _06088_ (.B1(_00683_),
    .Y(_00684_),
    .A1(net502),
    .A2(net1073));
 sg13g2_nand2_1 _06089_ (.Y(_00167_),
    .A(net1504),
    .B(_00684_));
 sg13g2_mux4_1 _06090_ (.S0(net1288),
    .A0(\cordic_inst.cordic_state[70] ),
    .A1(\cordic_inst.cordic_state[71] ),
    .A2(\cordic_inst.cordic_state[72] ),
    .A3(net1235),
    .S1(net1278),
    .X(_00685_));
 sg13g2_mux4_1 _06091_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[66] ),
    .A1(net1236),
    .A2(\cordic_inst.cordic_state[68] ),
    .A3(\cordic_inst.cordic_state[69] ),
    .S1(net1278),
    .X(_00686_));
 sg13g2_mux2_1 _06092_ (.A0(_00685_),
    .A1(_00686_),
    .S(net1133),
    .X(_00687_));
 sg13g2_nand2b_1 _06093_ (.Y(_00688_),
    .B(net1262),
    .A_N(_00687_));
 sg13g2_nand2_1 _06094_ (.Y(_00689_),
    .A(net1131),
    .B(_00636_));
 sg13g2_a21oi_1 _06095_ (.A1(net1279),
    .A2(_00642_),
    .Y(_00690_),
    .B1(net1120));
 sg13g2_mux4_1 _06096_ (.S0(net1289),
    .A0(\cordic_inst.cordic_state[62] ),
    .A1(\cordic_inst.cordic_state[63] ),
    .A2(\cordic_inst.cordic_state[64] ),
    .A3(\cordic_inst.cordic_state[65] ),
    .S1(net1279),
    .X(_00691_));
 sg13g2_o21ai_1 _06097_ (.B1(net1140),
    .Y(_00692_),
    .A1(_00640_),
    .A2(_00691_));
 sg13g2_a21oi_1 _06098_ (.A1(_00689_),
    .A2(_00690_),
    .Y(_00693_),
    .B1(_00692_));
 sg13g2_a21o_2 _06099_ (.A2(_04936_),
    .A1(net1135),
    .B1(net1121),
    .X(_00694_));
 sg13g2_nor3_1 _06100_ (.A(_04783_),
    .B(net1139),
    .C(_00694_),
    .Y(_00695_));
 sg13g2_mux4_1 _06101_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[74] ),
    .A1(\cordic_inst.cordic_state[75] ),
    .A2(\cordic_inst.cordic_state[76] ),
    .A3(net1234),
    .S1(net1277),
    .X(_00696_));
 sg13g2_a21oi_1 _06102_ (.A1(net1129),
    .A2(_00646_),
    .Y(_00697_),
    .B1(net1132));
 sg13g2_nor2_1 _06103_ (.A(net1271),
    .B(_00696_),
    .Y(_00698_));
 sg13g2_nor3_1 _06104_ (.A(net1262),
    .B(_00697_),
    .C(_00698_),
    .Y(_00699_));
 sg13g2_a221oi_1 _06105_ (.B2(net1256),
    .C1(_00695_),
    .B1(_00699_),
    .A1(_00688_),
    .Y(_00700_),
    .A2(_00693_));
 sg13g2_a21o_1 _06106_ (.A2(_00674_),
    .A1(_00654_),
    .B1(net1038),
    .X(_00701_));
 sg13g2_xor2_1 _06107_ (.B(_00701_),
    .A(_00700_),
    .X(_00702_));
 sg13g2_nor2_1 _06108_ (.A(_04791_),
    .B(_00702_),
    .Y(_00703_));
 sg13g2_xnor2_1 _06109_ (.Y(_00704_),
    .A(\cordic_inst.cordic_state[34] ),
    .B(_00702_));
 sg13g2_o21ai_1 _06110_ (.B1(_00678_),
    .Y(_00705_),
    .A1(_00655_),
    .A2(_00679_));
 sg13g2_a21oi_1 _06111_ (.A1(_00704_),
    .A2(_00705_),
    .Y(_00706_),
    .B1(_04913_));
 sg13g2_o21ai_1 _06112_ (.B1(_00706_),
    .Y(_00707_),
    .A1(_00704_),
    .A2(_00705_));
 sg13g2_a21oi_1 _06113_ (.A1(net1314),
    .A2(net1394),
    .Y(_00708_),
    .B1(net1306));
 sg13g2_a221oi_1 _06114_ (.B2(_00708_),
    .C1(net1085),
    .B1(_00707_),
    .A1(net1306),
    .Y(_00709_),
    .A2(_04824_));
 sg13g2_a21oi_1 _06115_ (.A1(net179),
    .A2(net1085),
    .Y(_00710_),
    .B1(_00709_));
 sg13g2_nor2_1 _06116_ (.A(net1477),
    .B(_00710_),
    .Y(_00168_));
 sg13g2_a21oi_1 _06117_ (.A1(_00704_),
    .A2(_00705_),
    .Y(_00711_),
    .B1(_00703_));
 sg13g2_mux4_1 _06118_ (.S0(net1288),
    .A0(\cordic_inst.cordic_state[71] ),
    .A1(\cordic_inst.cordic_state[72] ),
    .A2(net1235),
    .A3(\cordic_inst.cordic_state[74] ),
    .S1(net1278),
    .X(_00712_));
 sg13g2_mux4_1 _06119_ (.S0(net1288),
    .A0(net1236),
    .A1(\cordic_inst.cordic_state[68] ),
    .A2(\cordic_inst.cordic_state[69] ),
    .A3(\cordic_inst.cordic_state[70] ),
    .S1(net1277),
    .X(_00713_));
 sg13g2_mux2_1 _06120_ (.A0(_00712_),
    .A1(_00713_),
    .S(net1133),
    .X(_00714_));
 sg13g2_mux4_1 _06121_ (.S0(net1290),
    .A0(\cordic_inst.cordic_state[59] ),
    .A1(\cordic_inst.cordic_state[60] ),
    .A2(\cordic_inst.cordic_state[61] ),
    .A3(\cordic_inst.cordic_state[62] ),
    .S1(net1279),
    .X(_00715_));
 sg13g2_and2_1 _06122_ (.A(net1122),
    .B(_00715_),
    .X(_00716_));
 sg13g2_mux4_1 _06123_ (.S0(net1289),
    .A0(\cordic_inst.cordic_state[63] ),
    .A1(\cordic_inst.cordic_state[64] ),
    .A2(\cordic_inst.cordic_state[65] ),
    .A3(\cordic_inst.cordic_state[66] ),
    .S1(net1280),
    .X(_00717_));
 sg13g2_a221oi_1 _06124_ (.B2(_00639_),
    .C1(_00716_),
    .B1(_00717_),
    .A1(net1266),
    .Y(_00718_),
    .A2(_00714_));
 sg13g2_mux4_1 _06125_ (.S0(net1287),
    .A0(\cordic_inst.cordic_state[75] ),
    .A1(\cordic_inst.cordic_state[76] ),
    .A2(net1234),
    .A3(\cordic_inst.cordic_state[78] ),
    .S1(net1277),
    .X(_00719_));
 sg13g2_nand2_1 _06126_ (.Y(_00720_),
    .A(_04794_),
    .B(_00719_));
 sg13g2_nand3_1 _06127_ (.B(net1271),
    .C(_04936_),
    .A(net1232),
    .Y(_00721_));
 sg13g2_a21oi_1 _06128_ (.A1(_00720_),
    .A2(_00721_),
    .Y(_00722_),
    .B1(net1262));
 sg13g2_a21oi_1 _06129_ (.A1(net1253),
    .A2(_00722_),
    .Y(_00723_),
    .B1(_00695_));
 sg13g2_o21ai_1 _06130_ (.B1(_00723_),
    .Y(_00724_),
    .A1(net1256),
    .A2(_00718_));
 sg13g2_nand4_1 _06131_ (.B(_00653_),
    .C(_00674_),
    .A(_00645_),
    .Y(_00725_),
    .D(_00700_));
 sg13g2_nand2_1 _06132_ (.Y(_00726_),
    .A(net1043),
    .B(_00725_));
 sg13g2_xor2_1 _06133_ (.B(_00726_),
    .A(_00724_),
    .X(_00727_));
 sg13g2_nand2_1 _06134_ (.Y(_00728_),
    .A(\cordic_inst.cordic_state[35] ),
    .B(_00727_));
 sg13g2_xnor2_1 _06135_ (.Y(_00729_),
    .A(\cordic_inst.cordic_state[35] ),
    .B(_00727_));
 sg13g2_xor2_1 _06136_ (.B(_00729_),
    .A(_00711_),
    .X(_00730_));
 sg13g2_o21ai_1 _06137_ (.B1(_04887_),
    .Y(_00731_),
    .A1(_04909_),
    .A2(_00730_));
 sg13g2_a21oi_1 _06138_ (.A1(net1314),
    .A2(net1386),
    .Y(_00732_),
    .B1(net1306));
 sg13g2_a221oi_1 _06139_ (.B2(_00732_),
    .C1(net1086),
    .B1(_00731_),
    .A1(net1306),
    .Y(_00733_),
    .A2(_04825_));
 sg13g2_a21oi_1 _06140_ (.A1(net473),
    .A2(net1082),
    .Y(_00734_),
    .B1(_00733_));
 sg13g2_nand2_1 _06141_ (.Y(_00169_),
    .A(net1495),
    .B(_00734_));
 sg13g2_mux2_1 _06142_ (.A0(_00631_),
    .A1(_00648_),
    .S(net1272),
    .X(_00735_));
 sg13g2_and2_1 _06143_ (.A(net1122),
    .B(_00643_),
    .X(_00736_));
 sg13g2_a221oi_1 _06144_ (.B2(net1266),
    .C1(_00736_),
    .B1(_00735_),
    .A1(_00632_),
    .Y(_00737_),
    .A2(_00639_));
 sg13g2_and2_1 _06145_ (.A(net1121),
    .B(_00647_),
    .X(_00738_));
 sg13g2_nand2_2 _06146_ (.Y(_00739_),
    .A(_04916_),
    .B(net1121));
 sg13g2_a22oi_1 _06147_ (.Y(_00740_),
    .B1(_00739_),
    .B2(_00651_),
    .A2(_00738_),
    .A1(net1255));
 sg13g2_o21ai_1 _06148_ (.B1(_00740_),
    .Y(_00741_),
    .A1(net1255),
    .A2(_00737_));
 sg13g2_o21ai_1 _06149_ (.B1(net1043),
    .Y(_00742_),
    .A1(_00724_),
    .A2(_00725_));
 sg13g2_xor2_1 _06150_ (.B(_00742_),
    .A(_00741_),
    .X(_00743_));
 sg13g2_and2_1 _06151_ (.A(\cordic_inst.cordic_state[36] ),
    .B(_00743_),
    .X(_00744_));
 sg13g2_xnor2_1 _06152_ (.Y(_00745_),
    .A(\cordic_inst.cordic_state[36] ),
    .B(_00743_));
 sg13g2_inv_1 _06153_ (.Y(_00746_),
    .A(_00745_));
 sg13g2_o21ai_1 _06154_ (.B1(_00728_),
    .Y(_00747_),
    .A1(_00711_),
    .A2(_00729_));
 sg13g2_a21oi_1 _06155_ (.A1(_00746_),
    .A2(_00747_),
    .Y(_00748_),
    .B1(_04913_));
 sg13g2_o21ai_1 _06156_ (.B1(_00748_),
    .Y(_00749_),
    .A1(_00746_),
    .A2(_00747_));
 sg13g2_a21oi_1 _06157_ (.A1(net1314),
    .A2(net1378),
    .Y(_00750_),
    .B1(net1306));
 sg13g2_a221oi_1 _06158_ (.B2(_00750_),
    .C1(net1086),
    .B1(_00749_),
    .A1(net1306),
    .Y(_00751_),
    .A2(_04826_));
 sg13g2_a21oi_1 _06159_ (.A1(net423),
    .A2(net1082),
    .Y(_00752_),
    .B1(_00751_));
 sg13g2_nor2_1 _06160_ (.A(net1477),
    .B(_00752_),
    .Y(_00170_));
 sg13g2_a21oi_1 _06161_ (.A1(_00746_),
    .A2(_00747_),
    .Y(_00753_),
    .B1(_00744_));
 sg13g2_mux2_1 _06162_ (.A0(_00664_),
    .A1(_00668_),
    .S(_04794_),
    .X(_00754_));
 sg13g2_nor2_1 _06163_ (.A(net1120),
    .B(_00670_),
    .Y(_00755_));
 sg13g2_nor2_1 _06164_ (.A(_00640_),
    .B(_00667_),
    .Y(_00756_));
 sg13g2_o21ai_1 _06165_ (.B1(net1138),
    .Y(_00757_),
    .A1(net1136),
    .A2(_00754_));
 sg13g2_nor3_1 _06166_ (.A(_00755_),
    .B(_00756_),
    .C(_00757_),
    .Y(_00758_));
 sg13g2_nor2_1 _06167_ (.A(net1119),
    .B(_00662_),
    .Y(_00759_));
 sg13g2_a221oi_1 _06168_ (.B2(net1255),
    .C1(_00758_),
    .B1(_00759_),
    .A1(_00651_),
    .Y(_00760_),
    .A2(_00739_));
 sg13g2_nor3_1 _06169_ (.A(_00724_),
    .B(_00725_),
    .C(_00741_),
    .Y(_00761_));
 sg13g2_nor2_1 _06170_ (.A(net1038),
    .B(_00761_),
    .Y(_00762_));
 sg13g2_xor2_1 _06171_ (.B(_00762_),
    .A(_00760_),
    .X(_00763_));
 sg13g2_nand2_1 _06172_ (.Y(_00764_),
    .A(\cordic_inst.cordic_state[37] ),
    .B(_00763_));
 sg13g2_xnor2_1 _06173_ (.Y(_00765_),
    .A(\cordic_inst.cordic_state[37] ),
    .B(_00763_));
 sg13g2_xnor2_1 _06174_ (.Y(_00766_),
    .A(_00753_),
    .B(_00765_));
 sg13g2_nand2_1 _06175_ (.Y(_00767_),
    .A(net1107),
    .B(_00766_));
 sg13g2_a221oi_1 _06176_ (.B2(_00767_),
    .C1(net1305),
    .B1(_04887_),
    .A1(net1314),
    .Y(_00768_),
    .A2(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ));
 sg13g2_o21ai_1 _06177_ (.B1(net1076),
    .Y(_00769_),
    .A1(net1128),
    .A2(net1204));
 sg13g2_a21oi_1 _06178_ (.A1(net474),
    .A2(net1082),
    .Y(_00770_),
    .B1(net1477));
 sg13g2_o21ai_1 _06179_ (.B1(_00770_),
    .Y(_00171_),
    .A1(_00768_),
    .A2(_00769_));
 sg13g2_o21ai_1 _06180_ (.B1(_00764_),
    .Y(_00771_),
    .A1(_00753_),
    .A2(_00765_));
 sg13g2_nand2_1 _06181_ (.Y(_00772_),
    .A(_00760_),
    .B(_00761_));
 sg13g2_nand2_1 _06182_ (.Y(_00773_),
    .A(net1043),
    .B(_00772_));
 sg13g2_mux2_1 _06183_ (.A0(_00685_),
    .A1(_00696_),
    .S(net1271),
    .X(_00774_));
 sg13g2_or2_1 _06184_ (.X(_00775_),
    .B(_00774_),
    .A(net1135));
 sg13g2_nand3_1 _06185_ (.B(net1121),
    .C(_00646_),
    .A(net1129),
    .Y(_00776_));
 sg13g2_nand2_1 _06186_ (.Y(_00777_),
    .A(net1132),
    .B(_04936_));
 sg13g2_nand2_2 _06187_ (.Y(_00778_),
    .A(_04936_),
    .B(net1121));
 sg13g2_nor2_1 _06188_ (.A(net1138),
    .B(_00776_),
    .Y(_00779_));
 sg13g2_a21oi_1 _06189_ (.A1(_00651_),
    .A2(_00778_),
    .Y(_00780_),
    .B1(_00779_));
 sg13g2_o21ai_1 _06190_ (.B1(net1140),
    .Y(_00781_),
    .A1(net1119),
    .A2(_00691_));
 sg13g2_o21ai_1 _06191_ (.B1(_00775_),
    .Y(_00782_),
    .A1(_00640_),
    .A2(_00686_));
 sg13g2_o21ai_1 _06192_ (.B1(_00780_),
    .Y(_00783_),
    .A1(_00781_),
    .A2(_00782_));
 sg13g2_inv_1 _06193_ (.Y(_00784_),
    .A(_00783_));
 sg13g2_xnor2_1 _06194_ (.Y(_00785_),
    .A(_00773_),
    .B(_00784_));
 sg13g2_nand2_1 _06195_ (.Y(_00786_),
    .A(\cordic_inst.cordic_state[38] ),
    .B(_00785_));
 sg13g2_inv_1 _06196_ (.Y(_00787_),
    .A(_00786_));
 sg13g2_xor2_1 _06197_ (.B(_00785_),
    .A(\cordic_inst.cordic_state[38] ),
    .X(_00788_));
 sg13g2_and2_1 _06198_ (.A(_00771_),
    .B(_00788_),
    .X(_00789_));
 sg13g2_o21ai_1 _06199_ (.B1(net1094),
    .Y(_00790_),
    .A1(_00771_),
    .A2(_00788_));
 sg13g2_a21oi_1 _06200_ (.A1(net1314),
    .A2(net1359),
    .Y(_00791_),
    .B1(net1305));
 sg13g2_o21ai_1 _06201_ (.B1(_00791_),
    .Y(_00792_),
    .A1(_00789_),
    .A2(_00790_));
 sg13g2_o21ai_1 _06202_ (.B1(_00792_),
    .Y(_00793_),
    .A1(net1127),
    .A2(net1195));
 sg13g2_o21ai_1 _06203_ (.B1(net1493),
    .Y(_00794_),
    .A1(net467),
    .A2(net1073));
 sg13g2_a21oi_1 _06204_ (.A1(net1074),
    .A2(_00793_),
    .Y(_00172_),
    .B1(_00794_));
 sg13g2_a21oi_1 _06205_ (.A1(_00771_),
    .A2(_00788_),
    .Y(_00795_),
    .B1(_00787_));
 sg13g2_mux2_1 _06206_ (.A0(_00712_),
    .A1(_00719_),
    .S(net1271),
    .X(_00796_));
 sg13g2_nor2_1 _06207_ (.A(net1136),
    .B(_00796_),
    .Y(_00797_));
 sg13g2_o21ai_1 _06208_ (.B1(net1140),
    .Y(_00798_),
    .A1(net1120),
    .A2(_00717_));
 sg13g2_nor2_1 _06209_ (.A(_00640_),
    .B(_00713_),
    .Y(_00799_));
 sg13g2_nor3_1 _06210_ (.A(_00797_),
    .B(_00798_),
    .C(_00799_),
    .Y(_00800_));
 sg13g2_nor2_1 _06211_ (.A(_00651_),
    .B(_00800_),
    .Y(_00801_));
 sg13g2_o21ai_1 _06212_ (.B1(net1043),
    .Y(_00802_),
    .A1(_00772_),
    .A2(_00783_));
 sg13g2_xor2_1 _06213_ (.B(_00802_),
    .A(_00801_),
    .X(_00803_));
 sg13g2_nand2b_1 _06214_ (.Y(_00804_),
    .B(\cordic_inst.cordic_state[39] ),
    .A_N(_00803_));
 sg13g2_xnor2_1 _06215_ (.Y(_00805_),
    .A(_04790_),
    .B(_00803_));
 sg13g2_xnor2_1 _06216_ (.Y(_00806_),
    .A(_00795_),
    .B(_00805_));
 sg13g2_a22oi_1 _06217_ (.Y(_00807_),
    .B1(_04902_),
    .B2(net1357),
    .A2(net1193),
    .A1(net1305));
 sg13g2_o21ai_1 _06218_ (.B1(_00807_),
    .Y(_00808_),
    .A1(_04906_),
    .A2(_00806_));
 sg13g2_a21oi_1 _06219_ (.A1(net1074),
    .A2(_00808_),
    .Y(_00809_),
    .B1(net1477));
 sg13g2_o21ai_1 _06220_ (.B1(_00809_),
    .Y(_00173_),
    .A1(_04790_),
    .A2(net1074));
 sg13g2_o21ai_1 _06221_ (.B1(_00804_),
    .Y(_00810_),
    .A1(_00795_),
    .A2(_00805_));
 sg13g2_nand4_1 _06222_ (.B(_00761_),
    .C(_00784_),
    .A(_00760_),
    .Y(_00811_),
    .D(_00801_));
 sg13g2_nand2_1 _06223_ (.Y(_00812_),
    .A(net1043),
    .B(_00811_));
 sg13g2_nor2_1 _06224_ (.A(net1265),
    .B(_00633_),
    .Y(_00813_));
 sg13g2_or2_1 _06225_ (.X(_00814_),
    .B(_00649_),
    .A(net1134));
 sg13g2_nor2_1 _06226_ (.A(net1258),
    .B(_00813_),
    .Y(_00815_));
 sg13g2_a21oi_1 _06227_ (.A1(_00814_),
    .A2(_00815_),
    .Y(_00816_),
    .B1(_00651_));
 sg13g2_xnor2_1 _06228_ (.Y(_00817_),
    .A(_00812_),
    .B(_00816_));
 sg13g2_nand2_1 _06229_ (.Y(_00818_),
    .A(\cordic_inst.cordic_state[40] ),
    .B(_00817_));
 sg13g2_inv_1 _06230_ (.Y(_00819_),
    .A(_00818_));
 sg13g2_xor2_1 _06231_ (.B(_00817_),
    .A(\cordic_inst.cordic_state[40] ),
    .X(_00820_));
 sg13g2_o21ai_1 _06232_ (.B1(net1094),
    .Y(_00821_),
    .A1(_00810_),
    .A2(_00820_));
 sg13g2_a21o_1 _06233_ (.A2(_00820_),
    .A1(_00810_),
    .B1(_00821_),
    .X(_00822_));
 sg13g2_a21oi_1 _06234_ (.A1(net1314),
    .A2(net1474),
    .Y(_00823_),
    .B1(net1305));
 sg13g2_a22oi_1 _06235_ (.Y(_00824_),
    .B1(_00822_),
    .B2(_00823_),
    .A2(_04830_),
    .A1(net1306));
 sg13g2_nor2_1 _06236_ (.A(net1082),
    .B(_00824_),
    .Y(_00825_));
 sg13g2_o21ai_1 _06237_ (.B1(net1493),
    .Y(_00826_),
    .A1(net479),
    .A2(net1074));
 sg13g2_nor2_1 _06238_ (.A(_00825_),
    .B(_00826_),
    .Y(_00174_));
 sg13g2_a21oi_1 _06239_ (.A1(_00810_),
    .A2(_00820_),
    .Y(_00827_),
    .B1(_00819_));
 sg13g2_a21oi_2 _06240_ (.B1(net1253),
    .Y(_00828_),
    .A2(net1269),
    .A1(net1260));
 sg13g2_a21oi_2 _06241_ (.B1(_00828_),
    .Y(_00829_),
    .A2(net1129),
    .A1(net1139));
 sg13g2_nand2_1 _06242_ (.Y(_00830_),
    .A(net1232),
    .B(_00829_));
 sg13g2_nor2_1 _06243_ (.A(net1266),
    .B(_00669_),
    .Y(_00831_));
 sg13g2_o21ai_1 _06244_ (.B1(net1262),
    .Y(_00832_),
    .A1(_00663_),
    .A2(_00665_));
 sg13g2_nand2_1 _06245_ (.Y(_00833_),
    .A(net1138),
    .B(_00832_));
 sg13g2_o21ai_1 _06246_ (.B1(_00830_),
    .Y(_00834_),
    .A1(_00831_),
    .A2(_00833_));
 sg13g2_a21o_1 _06247_ (.A2(_00815_),
    .A1(_00814_),
    .B1(_00811_),
    .X(_00835_));
 sg13g2_nand2_1 _06248_ (.Y(_00836_),
    .A(net1043),
    .B(_00835_));
 sg13g2_xor2_1 _06249_ (.B(_00836_),
    .A(_00834_),
    .X(_00837_));
 sg13g2_nand2_1 _06250_ (.Y(_00838_),
    .A(\cordic_inst.cordic_state[41] ),
    .B(_00837_));
 sg13g2_xnor2_1 _06251_ (.Y(_00839_),
    .A(\cordic_inst.cordic_state[41] ),
    .B(_00837_));
 sg13g2_xnor2_1 _06252_ (.Y(_00840_),
    .A(_00827_),
    .B(_00839_));
 sg13g2_a22oi_1 _06253_ (.Y(_00841_),
    .B1(net1124),
    .B2(net1466),
    .A2(net1177),
    .A1(net1305));
 sg13g2_o21ai_1 _06254_ (.B1(_00841_),
    .Y(_00842_),
    .A1(_04906_),
    .A2(_00840_));
 sg13g2_a21oi_1 _06255_ (.A1(net1074),
    .A2(_00842_),
    .Y(_00843_),
    .B1(net1477));
 sg13g2_o21ai_1 _06256_ (.B1(_00843_),
    .Y(_00175_),
    .A1(_04789_),
    .A2(net1074));
 sg13g2_o21ai_1 _06257_ (.B1(_00838_),
    .Y(_00844_),
    .A1(_00827_),
    .A2(_00839_));
 sg13g2_nor2_1 _06258_ (.A(net1262),
    .B(_00687_),
    .Y(_00845_));
 sg13g2_o21ai_1 _06259_ (.B1(net1262),
    .Y(_00846_),
    .A1(_00697_),
    .A2(_00698_));
 sg13g2_nor2_1 _06260_ (.A(net1253),
    .B(_00845_),
    .Y(_00847_));
 sg13g2_a22oi_1 _06261_ (.Y(_00848_),
    .B1(_00846_),
    .B2(_00847_),
    .A2(_00829_),
    .A1(net1231));
 sg13g2_nor2_1 _06262_ (.A(_00834_),
    .B(_00835_),
    .Y(_00849_));
 sg13g2_nor2_1 _06263_ (.A(net1039),
    .B(_00849_),
    .Y(_00850_));
 sg13g2_xnor2_1 _06264_ (.Y(_00851_),
    .A(_00848_),
    .B(_00850_));
 sg13g2_nor2b_1 _06265_ (.A(_00851_),
    .B_N(net1251),
    .Y(_00852_));
 sg13g2_xnor2_1 _06266_ (.Y(_00853_),
    .A(net1251),
    .B(_00851_));
 sg13g2_o21ai_1 _06267_ (.B1(net1094),
    .Y(_00854_),
    .A1(_00844_),
    .A2(_00853_));
 sg13g2_a21o_1 _06268_ (.A2(_00853_),
    .A1(_00844_),
    .B1(_00854_),
    .X(_00855_));
 sg13g2_a21oi_1 _06269_ (.A1(net1314),
    .A2(net1461),
    .Y(_00856_),
    .B1(net1305));
 sg13g2_a221oi_1 _06270_ (.B2(_00856_),
    .C1(net1082),
    .B1(_00855_),
    .A1(net1305),
    .Y(_00857_),
    .A2(_04832_));
 sg13g2_a21oi_1 _06271_ (.A1(net1251),
    .A2(net1082),
    .Y(_00858_),
    .B1(_00857_));
 sg13g2_nor2_1 _06272_ (.A(net1481),
    .B(_00858_),
    .Y(_00176_));
 sg13g2_nor2_2 _06273_ (.A(_04814_),
    .B(_04903_),
    .Y(_00859_));
 sg13g2_a21oi_1 _06274_ (.A1(_00844_),
    .A2(_00853_),
    .Y(_00860_),
    .B1(_00852_));
 sg13g2_a21oi_1 _06275_ (.A1(net1138),
    .A2(_04936_),
    .Y(_00861_),
    .B1(_00828_));
 sg13g2_nand2_1 _06276_ (.Y(_00862_),
    .A(net1231),
    .B(_00861_));
 sg13g2_nand3_1 _06277_ (.B(_00720_),
    .C(_00721_),
    .A(net1262),
    .Y(_00863_));
 sg13g2_o21ai_1 _06278_ (.B1(_00863_),
    .Y(_00864_),
    .A1(net1263),
    .A2(_00714_));
 sg13g2_o21ai_1 _06279_ (.B1(_00862_),
    .Y(_00865_),
    .A1(net1254),
    .A2(_00864_));
 sg13g2_nand2_1 _06280_ (.Y(_00866_),
    .A(_00848_),
    .B(_00849_));
 sg13g2_nand2_1 _06281_ (.Y(_00867_),
    .A(net1041),
    .B(_00866_));
 sg13g2_xor2_1 _06282_ (.B(_00867_),
    .A(_00865_),
    .X(_00868_));
 sg13g2_nor2_1 _06283_ (.A(net1250),
    .B(_00868_),
    .Y(_00869_));
 sg13g2_xnor2_1 _06284_ (.Y(_00870_),
    .A(net1250),
    .B(_00868_));
 sg13g2_xor2_1 _06285_ (.B(_00870_),
    .A(_00860_),
    .X(_00871_));
 sg13g2_a221oi_1 _06286_ (.B2(_00871_),
    .C1(_00859_),
    .B1(net1109),
    .A1(net1305),
    .Y(_00872_),
    .A2(net1168));
 sg13g2_a21oi_1 _06287_ (.A1(net1250),
    .A2(net1082),
    .Y(_00873_),
    .B1(net1476));
 sg13g2_o21ai_1 _06288_ (.B1(_00873_),
    .Y(_00177_),
    .A1(net1082),
    .A2(_00872_));
 sg13g2_a21oi_1 _06289_ (.A1(net1260),
    .A2(_04925_),
    .Y(_00874_),
    .B1(net1253));
 sg13g2_nor2_1 _06290_ (.A(_04783_),
    .B(_00874_),
    .Y(_00875_));
 sg13g2_mux2_1 _06291_ (.A0(_00647_),
    .A1(_00735_),
    .S(net1135),
    .X(_00876_));
 sg13g2_a21o_1 _06292_ (.A2(_00876_),
    .A1(_00828_),
    .B1(_00875_),
    .X(_00877_));
 sg13g2_o21ai_1 _06293_ (.B1(net1042),
    .Y(_00878_),
    .A1(_00865_),
    .A2(_00866_));
 sg13g2_inv_1 _06294_ (.Y(_00879_),
    .A(_00878_));
 sg13g2_xor2_1 _06295_ (.B(_00878_),
    .A(_00877_),
    .X(_00880_));
 sg13g2_and2_1 _06296_ (.A(net1249),
    .B(_00880_),
    .X(_00881_));
 sg13g2_xnor2_1 _06297_ (.Y(_00882_),
    .A(net1249),
    .B(_00880_));
 sg13g2_a221oi_1 _06298_ (.B2(net1250),
    .C1(_00852_),
    .B1(_00868_),
    .A1(_00844_),
    .Y(_00883_),
    .A2(_00853_));
 sg13g2_nor3_1 _06299_ (.A(_00869_),
    .B(_00882_),
    .C(_00883_),
    .Y(_00884_));
 sg13g2_o21ai_1 _06300_ (.B1(_00882_),
    .Y(_00885_),
    .A1(_00869_),
    .A2(_00883_));
 sg13g2_nand3b_1 _06301_ (.B(_00885_),
    .C(net1094),
    .Y(_00886_),
    .A_N(_00884_));
 sg13g2_a21oi_1 _06302_ (.A1(net1312),
    .A2(net1452),
    .Y(_00887_),
    .B1(net1303));
 sg13g2_a221oi_1 _06303_ (.B2(_00887_),
    .C1(net1080),
    .B1(_00886_),
    .A1(net1303),
    .Y(_00888_),
    .A2(_04833_));
 sg13g2_a21oi_1 _06304_ (.A1(net1249),
    .A2(net1080),
    .Y(_00889_),
    .B1(_00888_));
 sg13g2_nor2_1 _06305_ (.A(net1476),
    .B(_00889_),
    .Y(_00178_));
 sg13g2_o21ai_1 _06306_ (.B1(_00828_),
    .Y(_00890_),
    .A1(net1260),
    .A2(_00754_));
 sg13g2_a21o_1 _06307_ (.A2(_00662_),
    .A1(net1260),
    .B1(_00890_),
    .X(_00891_));
 sg13g2_nor2b_1 _06308_ (.A(_00875_),
    .B_N(_00891_),
    .Y(_00892_));
 sg13g2_a21oi_1 _06309_ (.A1(net1042),
    .A2(_00877_),
    .Y(_00893_),
    .B1(_00879_));
 sg13g2_xnor2_1 _06310_ (.Y(_00894_),
    .A(_00892_),
    .B(_00893_));
 sg13g2_nand2_1 _06311_ (.Y(_00895_),
    .A(net1248),
    .B(_00894_));
 sg13g2_xnor2_1 _06312_ (.Y(_00896_),
    .A(net1248),
    .B(_00894_));
 sg13g2_inv_1 _06313_ (.Y(_00897_),
    .A(_00896_));
 sg13g2_or3_1 _06314_ (.A(_00881_),
    .B(_00884_),
    .C(_00897_),
    .X(_00898_));
 sg13g2_or4_1 _06315_ (.A(_00869_),
    .B(_00882_),
    .C(_00883_),
    .D(_00896_),
    .X(_00899_));
 sg13g2_nand2_1 _06316_ (.Y(_00900_),
    .A(_00881_),
    .B(_00897_));
 sg13g2_nand4_1 _06317_ (.B(_00898_),
    .C(_00899_),
    .A(net1109),
    .Y(_00901_),
    .D(_00900_));
 sg13g2_a22oi_1 _06318_ (.Y(_00902_),
    .B1(net1124),
    .B2(net1446),
    .A2(net1157),
    .A1(net1303));
 sg13g2_a21oi_1 _06319_ (.A1(_00901_),
    .A2(_00902_),
    .Y(_00903_),
    .B1(net1080));
 sg13g2_a21oi_1 _06320_ (.A1(net1248),
    .A2(net1080),
    .Y(_00904_),
    .B1(_00903_));
 sg13g2_nand2_1 _06321_ (.Y(_00179_),
    .A(net1489),
    .B(_00904_));
 sg13g2_and2_1 _06322_ (.A(_00895_),
    .B(_00900_),
    .X(_00905_));
 sg13g2_a21oi_1 _06323_ (.A1(net1260),
    .A2(_00777_),
    .Y(_00906_),
    .B1(net1252));
 sg13g2_nand2b_1 _06324_ (.Y(_00907_),
    .B(net1230),
    .A_N(_00906_));
 sg13g2_a21oi_1 _06325_ (.A1(net1130),
    .A2(_00646_),
    .Y(_00908_),
    .B1(net1134));
 sg13g2_o21ai_1 _06326_ (.B1(_00828_),
    .Y(_00909_),
    .A1(net1260),
    .A2(_00774_));
 sg13g2_o21ai_1 _06327_ (.B1(_00907_),
    .Y(_00910_),
    .A1(_00908_),
    .A2(_00909_));
 sg13g2_nor2_1 _06328_ (.A(net1038),
    .B(_00891_),
    .Y(_00911_));
 sg13g2_nor2b_1 _06329_ (.A(_00911_),
    .B_N(_00893_),
    .Y(_00912_));
 sg13g2_xor2_1 _06330_ (.B(_00912_),
    .A(_00910_),
    .X(_00913_));
 sg13g2_and2_1 _06331_ (.A(net1247),
    .B(_00913_),
    .X(_00914_));
 sg13g2_xnor2_1 _06332_ (.Y(_00915_),
    .A(net1247),
    .B(_00913_));
 sg13g2_a21oi_1 _06333_ (.A1(_00899_),
    .A2(_00905_),
    .Y(_00916_),
    .B1(_00915_));
 sg13g2_nand3_1 _06334_ (.B(_00905_),
    .C(_00915_),
    .A(_00899_),
    .Y(_00917_));
 sg13g2_nand2_1 _06335_ (.Y(_00918_),
    .A(net1094),
    .B(_00917_));
 sg13g2_a21oi_1 _06336_ (.A1(net1313),
    .A2(net1441),
    .Y(_00919_),
    .B1(net1303));
 sg13g2_o21ai_1 _06337_ (.B1(_00919_),
    .Y(_00920_),
    .A1(_00916_),
    .A2(_00918_));
 sg13g2_a21oi_1 _06338_ (.A1(net1301),
    .A2(_04834_),
    .Y(_00921_),
    .B1(net1078));
 sg13g2_a22oi_1 _06339_ (.Y(_00922_),
    .B1(_00920_),
    .B2(_00921_),
    .A2(net1080),
    .A1(net1247));
 sg13g2_nor2_1 _06340_ (.A(net1476),
    .B(_00922_),
    .Y(_00180_));
 sg13g2_nor2_1 _06341_ (.A(net1134),
    .B(_00777_),
    .Y(_00923_));
 sg13g2_a22oi_1 _06342_ (.Y(_00924_),
    .B1(_00923_),
    .B2(net1231),
    .A2(_00796_),
    .A1(net1134));
 sg13g2_o21ai_1 _06343_ (.B1(_00907_),
    .Y(_00925_),
    .A1(net1252),
    .A2(_00924_));
 sg13g2_nand2_1 _06344_ (.Y(_00926_),
    .A(net1041),
    .B(_00910_));
 sg13g2_nand2_1 _06345_ (.Y(_00927_),
    .A(_00912_),
    .B(_00926_));
 sg13g2_xor2_1 _06346_ (.B(_00927_),
    .A(_00925_),
    .X(_00928_));
 sg13g2_nor2b_1 _06347_ (.A(_00928_),
    .B_N(net1246),
    .Y(_00929_));
 sg13g2_inv_1 _06348_ (.Y(_00930_),
    .A(_00929_));
 sg13g2_xnor2_1 _06349_ (.Y(_00931_),
    .A(net1246),
    .B(_00928_));
 sg13g2_or3_1 _06350_ (.A(_00914_),
    .B(_00916_),
    .C(_00931_),
    .X(_00932_));
 sg13g2_o21ai_1 _06351_ (.B1(_00931_),
    .Y(_00933_),
    .A1(_00914_),
    .A2(_00916_));
 sg13g2_nand3_1 _06352_ (.B(_00932_),
    .C(_00933_),
    .A(net1109),
    .Y(_00934_));
 sg13g2_a22oi_1 _06353_ (.Y(_00935_),
    .B1(net1124),
    .B2(net1436),
    .A2(net1145),
    .A1(net1301));
 sg13g2_a21oi_1 _06354_ (.A1(_00934_),
    .A2(_00935_),
    .Y(_00936_),
    .B1(net1079));
 sg13g2_a21oi_1 _06355_ (.A1(net1246),
    .A2(net1079),
    .Y(_00937_),
    .B1(_00936_));
 sg13g2_nand2_1 _06356_ (.Y(_00181_),
    .A(net1490),
    .B(_00937_));
 sg13g2_nor2_2 _06357_ (.A(net1254),
    .B(_04929_),
    .Y(_00938_));
 sg13g2_inv_1 _06358_ (.Y(_00939_),
    .A(_00938_));
 sg13g2_nand2_1 _06359_ (.Y(_00940_),
    .A(net1139),
    .B(_00650_));
 sg13g2_o21ai_1 _06360_ (.B1(_00940_),
    .Y(_00941_),
    .A1(_04783_),
    .A2(_00938_));
 sg13g2_a21o_1 _06361_ (.A2(_00925_),
    .A1(net1041),
    .B1(_00927_),
    .X(_00942_));
 sg13g2_xnor2_1 _06362_ (.Y(_00943_),
    .A(_00941_),
    .B(_00942_));
 sg13g2_and2_1 _06363_ (.A(net1245),
    .B(_00943_),
    .X(_00944_));
 sg13g2_xor2_1 _06364_ (.B(_00943_),
    .A(net1245),
    .X(_00945_));
 sg13g2_inv_1 _06365_ (.Y(_00946_),
    .A(_00945_));
 sg13g2_a21oi_1 _06366_ (.A1(_00930_),
    .A2(_00933_),
    .Y(_00947_),
    .B1(_00946_));
 sg13g2_nand3_1 _06367_ (.B(_00933_),
    .C(_00946_),
    .A(_00930_),
    .Y(_00948_));
 sg13g2_nand2_1 _06368_ (.Y(_00949_),
    .A(net1094),
    .B(_00948_));
 sg13g2_a21oi_1 _06369_ (.A1(net1312),
    .A2(net1432),
    .Y(_00950_),
    .B1(net1302));
 sg13g2_o21ai_1 _06370_ (.B1(_00950_),
    .Y(_00951_),
    .A1(_00947_),
    .A2(_00949_));
 sg13g2_a21oi_1 _06371_ (.A1(net1301),
    .A2(_04835_),
    .Y(_00952_),
    .B1(net1078));
 sg13g2_a22oi_1 _06372_ (.Y(_00953_),
    .B1(_00951_),
    .B2(_00952_),
    .A2(net1078),
    .A1(net1245));
 sg13g2_nor2_1 _06373_ (.A(net1476),
    .B(_00953_),
    .Y(_00182_));
 sg13g2_nor2_1 _06374_ (.A(_00944_),
    .B(_00947_),
    .Y(_00954_));
 sg13g2_nor2_1 _06375_ (.A(net1252),
    .B(_00666_),
    .Y(_00955_));
 sg13g2_a21oi_1 _06376_ (.A1(net1230),
    .A2(_00939_),
    .Y(_00956_),
    .B1(_00955_));
 sg13g2_a21o_1 _06377_ (.A2(_00941_),
    .A1(net1041),
    .B1(_00942_),
    .X(_00957_));
 sg13g2_xor2_1 _06378_ (.B(_00957_),
    .A(_00956_),
    .X(_00958_));
 sg13g2_nor2_1 _06379_ (.A(net1244),
    .B(_00958_),
    .Y(_00959_));
 sg13g2_nand2_1 _06380_ (.Y(_00960_),
    .A(net1244),
    .B(_00958_));
 sg13g2_inv_1 _06381_ (.Y(_00961_),
    .A(_00960_));
 sg13g2_nor2_1 _06382_ (.A(_00959_),
    .B(_00961_),
    .Y(_00962_));
 sg13g2_xnor2_1 _06383_ (.Y(_00963_),
    .A(_00954_),
    .B(_00962_));
 sg13g2_o21ai_1 _06384_ (.B1(_04887_),
    .Y(_00964_),
    .A1(_04909_),
    .A2(_00963_));
 sg13g2_a21oi_1 _06385_ (.A1(net1312),
    .A2(net1428),
    .Y(_00965_),
    .B1(net1302));
 sg13g2_a221oi_1 _06386_ (.B2(_00965_),
    .C1(net1081),
    .B1(_00964_),
    .A1(net1302),
    .Y(_00966_),
    .A2(_04836_));
 sg13g2_a21oi_1 _06387_ (.A1(net1244),
    .A2(net1078),
    .Y(_00967_),
    .B1(_00966_));
 sg13g2_nand2_1 _06388_ (.Y(_00183_),
    .A(net1489),
    .B(_00967_));
 sg13g2_nand2_2 _06389_ (.Y(_00968_),
    .A(net1137),
    .B(_00694_));
 sg13g2_a22oi_1 _06390_ (.Y(_00969_),
    .B1(_00968_),
    .B2(net1230),
    .A2(_00699_),
    .A1(net1137));
 sg13g2_a21oi_1 _06391_ (.A1(net1041),
    .A2(_00955_),
    .Y(_00970_),
    .B1(_00957_));
 sg13g2_xnor2_1 _06392_ (.Y(_00971_),
    .A(_00969_),
    .B(_00970_));
 sg13g2_and2_1 _06393_ (.A(net1243),
    .B(_00971_),
    .X(_00972_));
 sg13g2_xor2_1 _06394_ (.B(_00971_),
    .A(net1243),
    .X(_00973_));
 sg13g2_inv_1 _06395_ (.Y(_00974_),
    .A(_00973_));
 sg13g2_nor3_1 _06396_ (.A(_00944_),
    .B(_00947_),
    .C(_00961_),
    .Y(_00975_));
 sg13g2_nor3_1 _06397_ (.A(_00959_),
    .B(_00974_),
    .C(_00975_),
    .Y(_00976_));
 sg13g2_o21ai_1 _06398_ (.B1(_00974_),
    .Y(_00977_),
    .A1(_00959_),
    .A2(_00975_));
 sg13g2_nand2_1 _06399_ (.Y(_00978_),
    .A(net1094),
    .B(_00977_));
 sg13g2_a21oi_1 _06400_ (.A1(net1312),
    .A2(net1424),
    .Y(_00979_),
    .B1(net1301));
 sg13g2_o21ai_1 _06401_ (.B1(_00979_),
    .Y(_00980_),
    .A1(_00976_),
    .A2(_00978_));
 sg13g2_o21ai_1 _06402_ (.B1(_00980_),
    .Y(_00981_),
    .A1(net1127),
    .A2(net1337));
 sg13g2_nand2_1 _06403_ (.Y(_00982_),
    .A(net1243),
    .B(net1078));
 sg13g2_a21oi_1 _06404_ (.A1(_00981_),
    .A2(_00982_),
    .Y(_00184_),
    .B1(net1476));
 sg13g2_or2_1 _06405_ (.X(_00983_),
    .B(_00976_),
    .A(_00972_));
 sg13g2_and2_1 _06406_ (.A(net1137),
    .B(_00722_),
    .X(_00984_));
 sg13g2_a21oi_1 _06407_ (.A1(net1233),
    .A2(_00968_),
    .Y(_00985_),
    .B1(_00984_));
 sg13g2_a21oi_1 _06408_ (.A1(_00969_),
    .A2(_00970_),
    .Y(_00986_),
    .B1(net1038));
 sg13g2_xor2_1 _06409_ (.B(_00986_),
    .A(_00985_),
    .X(_00987_));
 sg13g2_or2_1 _06410_ (.X(_00988_),
    .B(_00987_),
    .A(net1242));
 sg13g2_xor2_1 _06411_ (.B(_00987_),
    .A(net1242),
    .X(_00989_));
 sg13g2_o21ai_1 _06412_ (.B1(net1109),
    .Y(_00990_),
    .A1(_00983_),
    .A2(_00989_));
 sg13g2_a21oi_1 _06413_ (.A1(net1242),
    .A2(_00987_),
    .Y(_00991_),
    .B1(_00972_));
 sg13g2_nand2b_1 _06414_ (.Y(_00992_),
    .B(_00991_),
    .A_N(_00976_));
 sg13g2_a21oi_1 _06415_ (.A1(_00983_),
    .A2(_00989_),
    .Y(_00993_),
    .B1(_00990_));
 sg13g2_a221oi_1 _06416_ (.B2(net1421),
    .C1(_00993_),
    .B1(net1124),
    .A1(net1301),
    .Y(_00994_),
    .A2(net1335));
 sg13g2_a21oi_1 _06417_ (.A1(net1242),
    .A2(net1078),
    .Y(_00995_),
    .B1(net1476));
 sg13g2_o21ai_1 _06418_ (.B1(_00995_),
    .Y(_00185_),
    .A1(net1078),
    .A2(_00994_));
 sg13g2_nand3_1 _06419_ (.B(_04916_),
    .C(net1121),
    .A(net1137),
    .Y(_00996_));
 sg13g2_nand2_1 _06420_ (.Y(_00997_),
    .A(net1230),
    .B(_00996_));
 sg13g2_nand2_1 _06421_ (.Y(_00998_),
    .A(net1137),
    .B(_00738_));
 sg13g2_nand2_1 _06422_ (.Y(_00999_),
    .A(_00997_),
    .B(_00998_));
 sg13g2_a21oi_1 _06423_ (.A1(net1041),
    .A2(_00984_),
    .Y(_01000_),
    .B1(_00986_));
 sg13g2_nand2b_1 _06424_ (.Y(_01001_),
    .B(_01000_),
    .A_N(_00999_));
 sg13g2_xor2_1 _06425_ (.B(_01000_),
    .A(_00999_),
    .X(_01002_));
 sg13g2_nand2_1 _06426_ (.Y(_01003_),
    .A(net1241),
    .B(_01002_));
 sg13g2_xor2_1 _06427_ (.B(_01002_),
    .A(net1241),
    .X(_01004_));
 sg13g2_a21oi_1 _06428_ (.A1(_00988_),
    .A2(_00992_),
    .Y(_01005_),
    .B1(_01004_));
 sg13g2_and3_1 _06429_ (.X(_01006_),
    .A(_00988_),
    .B(_00992_),
    .C(_01004_));
 sg13g2_or3_1 _06430_ (.A(_04913_),
    .B(_01005_),
    .C(_01006_),
    .X(_01007_));
 sg13g2_a21oi_1 _06431_ (.A1(net1312),
    .A2(net1418),
    .Y(_01008_),
    .B1(net1301));
 sg13g2_o21ai_1 _06432_ (.B1(net1073),
    .Y(_01009_),
    .A1(net1127),
    .A2(net1332));
 sg13g2_a21oi_1 _06433_ (.A1(_01007_),
    .A2(_01008_),
    .Y(_01010_),
    .B1(_01009_));
 sg13g2_a21oi_1 _06434_ (.A1(net1241),
    .A2(net1078),
    .Y(_01011_),
    .B1(_01010_));
 sg13g2_nor2_1 _06435_ (.A(net1476),
    .B(_01011_),
    .Y(_00186_));
 sg13g2_a22oi_1 _06436_ (.Y(_01012_),
    .B1(_00996_),
    .B2(net1230),
    .A2(_00759_),
    .A1(net1137));
 sg13g2_nand2_1 _06437_ (.Y(_01013_),
    .A(net1041),
    .B(_01001_));
 sg13g2_xnor2_1 _06438_ (.Y(_01014_),
    .A(_01012_),
    .B(_01013_));
 sg13g2_or2_1 _06439_ (.X(_01015_),
    .B(_01014_),
    .A(\cordic_inst.cordic_state[53] ));
 sg13g2_nand2_1 _06440_ (.Y(_01016_),
    .A(\cordic_inst.cordic_state[53] ),
    .B(_01014_));
 sg13g2_nand2_1 _06441_ (.Y(_01017_),
    .A(_01015_),
    .B(_01016_));
 sg13g2_a21oi_1 _06442_ (.A1(net1241),
    .A2(_01002_),
    .Y(_01018_),
    .B1(_01006_));
 sg13g2_nand2_1 _06443_ (.Y(_01019_),
    .A(_01003_),
    .B(_01016_));
 sg13g2_xnor2_1 _06444_ (.Y(_01020_),
    .A(_01017_),
    .B(_01018_));
 sg13g2_a21oi_1 _06445_ (.A1(net1107),
    .A2(_01020_),
    .Y(_01021_),
    .B1(_04906_));
 sg13g2_a221oi_1 _06446_ (.B2(net1415),
    .C1(_01021_),
    .B1(net1124),
    .A1(net1301),
    .Y(_01022_),
    .A2(net1330));
 sg13g2_nor2_1 _06447_ (.A(net488),
    .B(net1073),
    .Y(_01023_));
 sg13g2_o21ai_1 _06448_ (.B1(net1489),
    .Y(_00187_),
    .A1(_01022_),
    .A2(_01023_));
 sg13g2_o21ai_1 _06449_ (.B1(net1230),
    .Y(_01024_),
    .A1(net1252),
    .A2(_00778_));
 sg13g2_o21ai_1 _06450_ (.B1(_01024_),
    .Y(_01025_),
    .A1(net1252),
    .A2(_00776_));
 sg13g2_o21ai_1 _06451_ (.B1(_01013_),
    .Y(_01026_),
    .A1(net1038),
    .A2(_01012_));
 sg13g2_xnor2_1 _06452_ (.Y(_01027_),
    .A(_01025_),
    .B(_01026_));
 sg13g2_nand2_1 _06453_ (.Y(_01028_),
    .A(\cordic_inst.cordic_state[54] ),
    .B(_01027_));
 sg13g2_xnor2_1 _06454_ (.Y(_01029_),
    .A(\cordic_inst.cordic_state[54] ),
    .B(_01027_));
 sg13g2_o21ai_1 _06455_ (.B1(_01015_),
    .Y(_01030_),
    .A1(_01006_),
    .A2(_01019_));
 sg13g2_nor2_1 _06456_ (.A(_01029_),
    .B(_01030_),
    .Y(_01031_));
 sg13g2_a21o_1 _06457_ (.A2(_01030_),
    .A1(_01029_),
    .B1(_04913_),
    .X(_01032_));
 sg13g2_a21oi_1 _06458_ (.A1(net1312),
    .A2(net1413),
    .Y(_01033_),
    .B1(net1302));
 sg13g2_o21ai_1 _06459_ (.B1(_01033_),
    .Y(_01034_),
    .A1(_01031_),
    .A2(_01032_));
 sg13g2_a21oi_1 _06460_ (.A1(net1302),
    .A2(_04837_),
    .Y(_01035_),
    .B1(net1079));
 sg13g2_a22oi_1 _06461_ (.Y(_01036_),
    .B1(_01034_),
    .B2(_01035_),
    .A2(net1079),
    .A1(net496));
 sg13g2_nor2_1 _06462_ (.A(net1476),
    .B(_01036_),
    .Y(_00188_));
 sg13g2_o21ai_1 _06463_ (.B1(_01028_),
    .Y(_01037_),
    .A1(_01029_),
    .A2(_01030_));
 sg13g2_o21ai_1 _06464_ (.B1(net1041),
    .Y(_01038_),
    .A1(_01025_),
    .A2(_01026_));
 sg13g2_xor2_1 _06465_ (.B(net1239),
    .A(net1233),
    .X(_01039_));
 sg13g2_xnor2_1 _06466_ (.Y(_01040_),
    .A(_01038_),
    .B(_01039_));
 sg13g2_and2_1 _06467_ (.A(_01037_),
    .B(_01040_),
    .X(_01041_));
 sg13g2_o21ai_1 _06468_ (.B1(net1107),
    .Y(_01042_),
    .A1(_01037_),
    .A2(_01040_));
 sg13g2_o21ai_1 _06469_ (.B1(net1109),
    .Y(_01043_),
    .A1(_01041_),
    .A2(_01042_));
 sg13g2_a22oi_1 _06470_ (.Y(_01044_),
    .B1(net1124),
    .B2(net1410),
    .A2(net1325),
    .A1(net1302));
 sg13g2_a21oi_1 _06471_ (.A1(_01043_),
    .A2(_01044_),
    .Y(_01045_),
    .B1(net1081));
 sg13g2_a21oi_1 _06472_ (.A1(net1239),
    .A2(net1079),
    .Y(_01046_),
    .B1(_01045_));
 sg13g2_nand2_1 _06473_ (.Y(_00189_),
    .A(net1489),
    .B(_01046_));
 sg13g2_nand2_1 _06474_ (.Y(_01047_),
    .A(net415),
    .B(net1085));
 sg13g2_mux4_1 _06475_ (.S0(net1283),
    .A0(net1249),
    .A1(net1248),
    .A2(net1247),
    .A3(net1246),
    .S1(net1274),
    .X(_01048_));
 sg13g2_mux2_1 _06476_ (.A0(\cordic_inst.cordic_state[40] ),
    .A1(\cordic_inst.cordic_state[41] ),
    .S(net1284),
    .X(_01049_));
 sg13g2_mux4_1 _06477_ (.S0(net1284),
    .A0(\cordic_inst.cordic_state[40] ),
    .A1(\cordic_inst.cordic_state[41] ),
    .A2(net1251),
    .A3(net1250),
    .S1(net1274),
    .X(_01050_));
 sg13g2_mux2_1 _06478_ (.A0(_01048_),
    .A1(_01050_),
    .S(net1133),
    .X(_01051_));
 sg13g2_nor2b_1 _06479_ (.A(net1290),
    .B_N(\cordic_inst.cordic_state[32] ),
    .Y(_01052_));
 sg13g2_a21oi_1 _06480_ (.A1(\cordic_inst.cordic_state[33] ),
    .A2(net1290),
    .Y(_01053_),
    .B1(_01052_));
 sg13g2_mux2_1 _06481_ (.A0(\cordic_inst.cordic_state[34] ),
    .A1(\cordic_inst.cordic_state[35] ),
    .S(net1290),
    .X(_01054_));
 sg13g2_o21ai_1 _06482_ (.B1(net1122),
    .Y(_01055_),
    .A1(net1131),
    .A2(_01054_));
 sg13g2_a21o_1 _06483_ (.A2(_01053_),
    .A1(net1131),
    .B1(_01055_),
    .X(_01056_));
 sg13g2_mux2_1 _06484_ (.A0(\cordic_inst.cordic_state[38] ),
    .A1(\cordic_inst.cordic_state[39] ),
    .S(net1283),
    .X(_01057_));
 sg13g2_mux2_1 _06485_ (.A0(\cordic_inst.cordic_state[36] ),
    .A1(\cordic_inst.cordic_state[37] ),
    .S(net1285),
    .X(_01058_));
 sg13g2_mux2_1 _06486_ (.A0(_01057_),
    .A1(_01058_),
    .S(net1130),
    .X(_01059_));
 sg13g2_a22oi_1 _06487_ (.Y(_01060_),
    .B1(_01059_),
    .B2(_00639_),
    .A2(_01051_),
    .A1(net1264));
 sg13g2_nand2_1 _06488_ (.Y(_01061_),
    .A(_01056_),
    .B(_01060_));
 sg13g2_a21oi_1 _06489_ (.A1(_01056_),
    .A2(_01060_),
    .Y(_01062_),
    .B1(net1257));
 sg13g2_mux4_1 _06490_ (.S0(net1282),
    .A0(net1245),
    .A1(net1244),
    .A2(net1243),
    .A3(net1242),
    .S1(net1276),
    .X(_01063_));
 sg13g2_mux2_1 _06491_ (.A0(\cordic_inst.cordic_state[54] ),
    .A1(net1237),
    .S(net1286),
    .X(_01064_));
 sg13g2_mux4_1 _06492_ (.S0(net1282),
    .A0(net1241),
    .A1(\cordic_inst.cordic_state[53] ),
    .A2(\cordic_inst.cordic_state[54] ),
    .A3(net1237),
    .S1(net1276),
    .X(_01065_));
 sg13g2_mux2_1 _06493_ (.A0(_01063_),
    .A1(_01065_),
    .S(net1269),
    .X(_01066_));
 sg13g2_and2_1 _06494_ (.A(net1136),
    .B(_01066_),
    .X(_01067_));
 sg13g2_and2_1 _06495_ (.A(net1237),
    .B(net1256),
    .X(_01068_));
 sg13g2_nand2_1 _06496_ (.Y(_01069_),
    .A(net1238),
    .B(net1256));
 sg13g2_a21oi_1 _06497_ (.A1(net1136),
    .A2(_04917_),
    .Y(_01070_),
    .B1(_01069_));
 sg13g2_a21o_2 _06498_ (.A2(_01067_),
    .A1(net1257),
    .B1(_01070_),
    .X(_01071_));
 sg13g2_o21ai_1 _06499_ (.B1(\cordic_inst.cordic_state[56] ),
    .Y(_01072_),
    .A1(_01062_),
    .A2(_01071_));
 sg13g2_nor3_1 _06500_ (.A(\cordic_inst.cordic_state[56] ),
    .B(_01062_),
    .C(_01071_),
    .Y(_01073_));
 sg13g2_nand3b_1 _06501_ (.B(net1107),
    .C(_01072_),
    .Y(_01074_),
    .A_N(_01073_));
 sg13g2_a22oi_1 _06502_ (.Y(_01075_),
    .B1(net1108),
    .B2(_01074_),
    .A2(_04804_),
    .A1(net1310));
 sg13g2_o21ai_1 _06503_ (.B1(_01075_),
    .Y(_01076_),
    .A1(net1227),
    .A2(_04903_));
 sg13g2_a21oi_1 _06504_ (.A1(_01047_),
    .A2(_01076_),
    .Y(_00190_),
    .B1(net1479));
 sg13g2_nor2b_1 _06505_ (.A(net1283),
    .B_N(\cordic_inst.cordic_state[41] ),
    .Y(_01077_));
 sg13g2_a21oi_1 _06506_ (.A1(net1251),
    .A2(net1284),
    .Y(_01078_),
    .B1(_01077_));
 sg13g2_mux4_1 _06507_ (.S0(net1284),
    .A0(\cordic_inst.cordic_state[41] ),
    .A1(net1251),
    .A2(net1250),
    .A3(net1249),
    .S1(net1275),
    .X(_01079_));
 sg13g2_mux4_1 _06508_ (.S0(net1283),
    .A0(net1248),
    .A1(net1247),
    .A2(\cordic_inst.cordic_state[47] ),
    .A3(net1245),
    .S1(net1275),
    .X(_01080_));
 sg13g2_mux2_1 _06509_ (.A0(_01079_),
    .A1(_01080_),
    .S(net1270),
    .X(_01081_));
 sg13g2_and2_1 _06510_ (.A(net1265),
    .B(_01081_),
    .X(_01082_));
 sg13g2_nand2b_1 _06511_ (.Y(_01083_),
    .B(\cordic_inst.cordic_state[33] ),
    .A_N(net1290));
 sg13g2_a21oi_1 _06512_ (.A1(\cordic_inst.cordic_state[34] ),
    .A2(net1290),
    .Y(_01084_),
    .B1(net1279));
 sg13g2_nand2b_1 _06513_ (.Y(_01085_),
    .B(net1285),
    .A_N(\cordic_inst.cordic_state[36] ));
 sg13g2_o21ai_1 _06514_ (.B1(_01085_),
    .Y(_01086_),
    .A1(\cordic_inst.cordic_state[35] ),
    .A2(net1285));
 sg13g2_a221oi_1 _06515_ (.B2(net1275),
    .C1(net1119),
    .B1(_01086_),
    .A1(_01083_),
    .Y(_01087_),
    .A2(_01084_));
 sg13g2_mux2_1 _06516_ (.A0(\cordic_inst.cordic_state[39] ),
    .A1(\cordic_inst.cordic_state[40] ),
    .S(net1284),
    .X(_01088_));
 sg13g2_mux2_1 _06517_ (.A0(\cordic_inst.cordic_state[37] ),
    .A1(\cordic_inst.cordic_state[38] ),
    .S(net1285),
    .X(_01089_));
 sg13g2_mux2_1 _06518_ (.A0(_01088_),
    .A1(_01089_),
    .S(net1130),
    .X(_01090_));
 sg13g2_and2_1 _06519_ (.A(_00639_),
    .B(_01090_),
    .X(_01091_));
 sg13g2_or4_1 _06520_ (.A(net1258),
    .B(_01082_),
    .C(_01087_),
    .D(_01091_),
    .X(_01092_));
 sg13g2_mux2_1 _06521_ (.A0(net1242),
    .A1(net1241),
    .S(net1282),
    .X(_01093_));
 sg13g2_mux4_1 _06522_ (.S0(net1283),
    .A0(net1244),
    .A1(net1243),
    .A2(\cordic_inst.cordic_state[51] ),
    .A3(\cordic_inst.cordic_state[52] ),
    .S1(net1274),
    .X(_01094_));
 sg13g2_mux2_1 _06523_ (.A0(\cordic_inst.cordic_state[53] ),
    .A1(\cordic_inst.cordic_state[54] ),
    .S(net1282),
    .X(_01095_));
 sg13g2_a22oi_1 _06524_ (.Y(_01096_),
    .B1(_01095_),
    .B2(net1129),
    .A2(_00661_),
    .A1(net1237));
 sg13g2_nor2_1 _06525_ (.A(net1269),
    .B(_01094_),
    .Y(_01097_));
 sg13g2_a21o_2 _06526_ (.A2(_01096_),
    .A1(net1269),
    .B1(_01097_),
    .X(_01098_));
 sg13g2_o21ai_1 _06527_ (.B1(net1257),
    .Y(_01099_),
    .A1(net1266),
    .A2(_01098_));
 sg13g2_a21oi_1 _06528_ (.A1(_01092_),
    .A2(_01099_),
    .Y(_01100_),
    .B1(_01070_));
 sg13g2_o21ai_1 _06529_ (.B1(net1044),
    .Y(_01101_),
    .A1(_01062_),
    .A2(_01071_));
 sg13g2_xor2_1 _06530_ (.B(_01101_),
    .A(_01100_),
    .X(_01102_));
 sg13g2_nand2_1 _06531_ (.Y(_01103_),
    .A(\cordic_inst.cordic_state[57] ),
    .B(_01102_));
 sg13g2_xnor2_1 _06532_ (.Y(_01104_),
    .A(\cordic_inst.cordic_state[57] ),
    .B(_01102_));
 sg13g2_xor2_1 _06533_ (.B(_01104_),
    .A(_01072_),
    .X(_01105_));
 sg13g2_a221oi_1 _06534_ (.B2(net1125),
    .C1(net1083),
    .B1(_04823_),
    .A1(net1310),
    .Y(_01106_),
    .A2(_04805_));
 sg13g2_o21ai_1 _06535_ (.B1(_01106_),
    .Y(_01107_),
    .A1(net1049),
    .A2(_01105_));
 sg13g2_a21oi_1 _06536_ (.A1(net483),
    .A2(net1085),
    .Y(_01108_),
    .B1(net1480));
 sg13g2_nand2_1 _06537_ (.Y(_00191_),
    .A(_01107_),
    .B(_01108_));
 sg13g2_o21ai_1 _06538_ (.B1(_01103_),
    .Y(_01109_),
    .A1(_01072_),
    .A2(_01104_));
 sg13g2_mux4_1 _06539_ (.S0(net1283),
    .A0(net1247),
    .A1(net1246),
    .A2(\cordic_inst.cordic_state[48] ),
    .A3(\cordic_inst.cordic_state[49] ),
    .S1(net1274),
    .X(_01110_));
 sg13g2_mux4_1 _06540_ (.S0(net1283),
    .A0(net1251),
    .A1(net1250),
    .A2(net1249),
    .A3(net1248),
    .S1(net1274),
    .X(_01111_));
 sg13g2_mux2_1 _06541_ (.A0(_01110_),
    .A1(_01111_),
    .S(net1133),
    .X(_01112_));
 sg13g2_nand2b_1 _06542_ (.Y(_01113_),
    .B(net1264),
    .A_N(_01112_));
 sg13g2_nand2_1 _06543_ (.Y(_01114_),
    .A(net1131),
    .B(_01054_));
 sg13g2_a21oi_1 _06544_ (.A1(net1275),
    .A2(_01058_),
    .Y(_01115_),
    .B1(net1119));
 sg13g2_mux2_1 _06545_ (.A0(_01049_),
    .A1(_01057_),
    .S(net1130),
    .X(_01116_));
 sg13g2_inv_1 _06546_ (.Y(_01117_),
    .A(_01116_));
 sg13g2_a221oi_1 _06547_ (.B2(_00639_),
    .C1(net1258),
    .B1(_01117_),
    .A1(_01114_),
    .Y(_01118_),
    .A2(_01115_));
 sg13g2_nor2_1 _06548_ (.A(_00694_),
    .B(_01069_),
    .Y(_01119_));
 sg13g2_mux4_1 _06549_ (.S0(net1283),
    .A0(\cordic_inst.cordic_state[50] ),
    .A1(\cordic_inst.cordic_state[51] ),
    .A2(net1241),
    .A3(\cordic_inst.cordic_state[53] ),
    .S1(net1274),
    .X(_01120_));
 sg13g2_nand2_1 _06550_ (.Y(_01121_),
    .A(net1132),
    .B(_01120_));
 sg13g2_nand2_1 _06551_ (.Y(_01122_),
    .A(net1129),
    .B(_01064_));
 sg13g2_o21ai_1 _06552_ (.B1(_01121_),
    .Y(_01123_),
    .A1(net1132),
    .A2(_01122_));
 sg13g2_and2_1 _06553_ (.A(net1135),
    .B(_01123_),
    .X(_01124_));
 sg13g2_a221oi_1 _06554_ (.B2(net1255),
    .C1(_01119_),
    .B1(_01124_),
    .A1(_01113_),
    .Y(_01125_),
    .A2(_01118_));
 sg13g2_a221oi_1 _06555_ (.B2(_01099_),
    .C1(_01071_),
    .B1(_01092_),
    .A1(net1140),
    .Y(_01126_),
    .A2(_01061_));
 sg13g2_nor2_1 _06556_ (.A(net1039),
    .B(_01126_),
    .Y(_01127_));
 sg13g2_xnor2_1 _06557_ (.Y(_01128_),
    .A(_01125_),
    .B(_01127_));
 sg13g2_and2_1 _06558_ (.A(\cordic_inst.cordic_state[58] ),
    .B(_01128_),
    .X(_01129_));
 sg13g2_xor2_1 _06559_ (.B(_01128_),
    .A(\cordic_inst.cordic_state[58] ),
    .X(_01130_));
 sg13g2_a21oi_1 _06560_ (.A1(_01109_),
    .A2(_01130_),
    .Y(_01131_),
    .B1(_04909_));
 sg13g2_o21ai_1 _06561_ (.B1(_01131_),
    .Y(_01132_),
    .A1(_01109_),
    .A2(_01130_));
 sg13g2_nand2_1 _06562_ (.Y(_01133_),
    .A(_04824_),
    .B(net1126));
 sg13g2_a22oi_1 _06563_ (.Y(_01134_),
    .B1(net1108),
    .B2(_01132_),
    .A2(_04806_),
    .A1(net1309));
 sg13g2_a22oi_1 _06564_ (.Y(_01135_),
    .B1(_01133_),
    .B2(_01134_),
    .A2(net1087),
    .A1(net472));
 sg13g2_nor2_1 _06565_ (.A(net1484),
    .B(_01135_),
    .Y(_00192_));
 sg13g2_a21oi_1 _06566_ (.A1(_01109_),
    .A2(_01130_),
    .Y(_01136_),
    .B1(_01129_));
 sg13g2_mux4_1 _06567_ (.S0(net1282),
    .A0(net1246),
    .A1(net1245),
    .A2(net1244),
    .A3(net1243),
    .S1(net1276),
    .X(_01137_));
 sg13g2_mux4_1 _06568_ (.S0(net1282),
    .A0(net1250),
    .A1(net1249),
    .A2(net1248),
    .A3(net1247),
    .S1(net1276),
    .X(_01138_));
 sg13g2_mux2_1 _06569_ (.A0(_01137_),
    .A1(_01138_),
    .S(net1132),
    .X(_01139_));
 sg13g2_nand2b_1 _06570_ (.Y(_01140_),
    .B(net1264),
    .A_N(_01139_));
 sg13g2_a21oi_1 _06571_ (.A1(net1275),
    .A2(_01089_),
    .Y(_01141_),
    .B1(net1119));
 sg13g2_o21ai_1 _06572_ (.B1(_01141_),
    .Y(_01142_),
    .A1(net1275),
    .A2(_01086_));
 sg13g2_nor2_1 _06573_ (.A(net1274),
    .B(_01088_),
    .Y(_01143_));
 sg13g2_a21oi_1 _06574_ (.A1(net1275),
    .A2(_01078_),
    .Y(_01144_),
    .B1(_01143_));
 sg13g2_or2_1 _06575_ (.X(_01145_),
    .B(_01144_),
    .A(_00640_));
 sg13g2_nand4_1 _06576_ (.B(_01140_),
    .C(_01142_),
    .A(net1139),
    .Y(_01146_),
    .D(_01145_));
 sg13g2_nand3_1 _06577_ (.B(net1269),
    .C(_04936_),
    .A(net1237),
    .Y(_01147_));
 sg13g2_mux2_1 _06578_ (.A0(_01093_),
    .A1(_01095_),
    .S(net1276),
    .X(_01148_));
 sg13g2_nand2_1 _06579_ (.Y(_01149_),
    .A(net1132),
    .B(_01148_));
 sg13g2_a21oi_1 _06580_ (.A1(_01147_),
    .A2(_01149_),
    .Y(_01150_),
    .B1(net1260));
 sg13g2_a21oi_1 _06581_ (.A1(net1255),
    .A2(_01150_),
    .Y(_01151_),
    .B1(_01119_));
 sg13g2_and2_1 _06582_ (.A(_01146_),
    .B(_01151_),
    .X(_01152_));
 sg13g2_and2_1 _06583_ (.A(_01125_),
    .B(_01126_),
    .X(_01153_));
 sg13g2_nor2_1 _06584_ (.A(net1039),
    .B(_01153_),
    .Y(_01154_));
 sg13g2_xnor2_1 _06585_ (.Y(_01155_),
    .A(_01152_),
    .B(_01154_));
 sg13g2_nand2_1 _06586_ (.Y(_01156_),
    .A(\cordic_inst.cordic_state[59] ),
    .B(_01155_));
 sg13g2_xnor2_1 _06587_ (.Y(_01157_),
    .A(\cordic_inst.cordic_state[59] ),
    .B(_01155_));
 sg13g2_xnor2_1 _06588_ (.Y(_01158_),
    .A(_01136_),
    .B(_01157_));
 sg13g2_nand2_1 _06589_ (.Y(_01159_),
    .A(net1107),
    .B(_01158_));
 sg13g2_a221oi_1 _06590_ (.B2(_01159_),
    .C1(net1309),
    .B1(_04887_),
    .A1(net1315),
    .Y(_01160_),
    .A2(net1213));
 sg13g2_o21ai_1 _06591_ (.B1(net1075),
    .Y(_01161_),
    .A1(net1128),
    .A2(net1386));
 sg13g2_a21oi_1 _06592_ (.A1(net485),
    .A2(net1088),
    .Y(_01162_),
    .B1(net1479));
 sg13g2_o21ai_1 _06593_ (.B1(_01162_),
    .Y(_00193_),
    .A1(_01160_),
    .A2(_01161_));
 sg13g2_o21ai_1 _06594_ (.B1(_01156_),
    .Y(_01163_),
    .A1(_01136_),
    .A2(_01157_));
 sg13g2_mux2_1 _06595_ (.A0(_01048_),
    .A1(_01063_),
    .S(net1270),
    .X(_01164_));
 sg13g2_nor2_1 _06596_ (.A(net1119),
    .B(_01059_),
    .Y(_01165_));
 sg13g2_nor2_1 _06597_ (.A(_00640_),
    .B(_01050_),
    .Y(_01166_));
 sg13g2_o21ai_1 _06598_ (.B1(net1139),
    .Y(_01167_),
    .A1(net1134),
    .A2(_01164_));
 sg13g2_nor3_1 _06599_ (.A(_01165_),
    .B(_01166_),
    .C(_01167_),
    .Y(_01168_));
 sg13g2_nand2_1 _06600_ (.Y(_01169_),
    .A(net1121),
    .B(_01065_));
 sg13g2_inv_1 _06601_ (.Y(_01170_),
    .A(_01169_));
 sg13g2_a221oi_1 _06602_ (.B2(net1255),
    .C1(_01168_),
    .B1(_01170_),
    .A1(_00739_),
    .Y(_01171_),
    .A2(_01068_));
 sg13g2_a21oi_1 _06603_ (.A1(_01152_),
    .A2(_01153_),
    .Y(_01172_),
    .B1(net1039));
 sg13g2_xnor2_1 _06604_ (.Y(_01173_),
    .A(_01171_),
    .B(_01172_));
 sg13g2_and2_1 _06605_ (.A(\cordic_inst.cordic_state[60] ),
    .B(_01173_),
    .X(_01174_));
 sg13g2_xor2_1 _06606_ (.B(_01173_),
    .A(\cordic_inst.cordic_state[60] ),
    .X(_01175_));
 sg13g2_and2_1 _06607_ (.A(_01163_),
    .B(_01175_),
    .X(_01176_));
 sg13g2_o21ai_1 _06608_ (.B1(_04908_),
    .Y(_01177_),
    .A1(_01163_),
    .A2(_01175_));
 sg13g2_o21ai_1 _06609_ (.B1(net1108),
    .Y(_01178_),
    .A1(_01176_),
    .A2(_01177_));
 sg13g2_a22oi_1 _06610_ (.Y(_01179_),
    .B1(_04826_),
    .B2(net1125),
    .A2(_04808_),
    .A1(net1309));
 sg13g2_a22oi_1 _06611_ (.Y(_01180_),
    .B1(_01178_),
    .B2(_01179_),
    .A2(net1087),
    .A1(net481));
 sg13g2_nor2_1 _06612_ (.A(net1479),
    .B(net482),
    .Y(_00194_));
 sg13g2_a21oi_1 _06613_ (.A1(_01163_),
    .A2(_01175_),
    .Y(_01181_),
    .B1(_01174_));
 sg13g2_mux2_1 _06614_ (.A0(_01080_),
    .A1(_01094_),
    .S(net1270),
    .X(_01182_));
 sg13g2_nand2_1 _06615_ (.Y(_01183_),
    .A(net1264),
    .B(_01182_));
 sg13g2_a22oi_1 _06616_ (.Y(_01184_),
    .B1(_01090_),
    .B2(net1122),
    .A2(_01079_),
    .A1(_00639_));
 sg13g2_nand2_1 _06617_ (.Y(_01185_),
    .A(_01183_),
    .B(_01184_));
 sg13g2_nand2b_1 _06618_ (.Y(_01186_),
    .B(net1121),
    .A_N(_01096_));
 sg13g2_a22oi_1 _06619_ (.Y(_01187_),
    .B1(_01185_),
    .B2(net1139),
    .A2(_01068_),
    .A1(_00739_));
 sg13g2_o21ai_1 _06620_ (.B1(_01187_),
    .Y(_01188_),
    .A1(net1139),
    .A2(_01186_));
 sg13g2_nand3_1 _06621_ (.B(_01153_),
    .C(_01171_),
    .A(_01152_),
    .Y(_01189_));
 sg13g2_nand2_1 _06622_ (.Y(_01190_),
    .A(net1044),
    .B(_01189_));
 sg13g2_xnor2_1 _06623_ (.Y(_01191_),
    .A(_01188_),
    .B(_01190_));
 sg13g2_nand2_1 _06624_ (.Y(_01192_),
    .A(\cordic_inst.cordic_state[61] ),
    .B(_01191_));
 sg13g2_xnor2_1 _06625_ (.Y(_01193_),
    .A(\cordic_inst.cordic_state[61] ),
    .B(_01191_));
 sg13g2_xor2_1 _06626_ (.B(_01193_),
    .A(_01181_),
    .X(_01194_));
 sg13g2_a221oi_1 _06627_ (.B2(net1125),
    .C1(net1087),
    .B1(_04827_),
    .A1(net1310),
    .Y(_01195_),
    .A2(_04809_));
 sg13g2_o21ai_1 _06628_ (.B1(_01195_),
    .Y(_01196_),
    .A1(net1049),
    .A2(_01194_));
 sg13g2_a21oi_1 _06629_ (.A1(net490),
    .A2(net1087),
    .Y(_01197_),
    .B1(net1479));
 sg13g2_nand2_1 _06630_ (.Y(_00195_),
    .A(_01196_),
    .B(_01197_));
 sg13g2_o21ai_1 _06631_ (.B1(_01192_),
    .Y(_01198_),
    .A1(_01181_),
    .A2(_01193_));
 sg13g2_mux2_1 _06632_ (.A0(_01110_),
    .A1(_01120_),
    .S(net1270),
    .X(_01199_));
 sg13g2_inv_1 _06633_ (.Y(_01200_),
    .A(_01199_));
 sg13g2_o21ai_1 _06634_ (.B1(net1140),
    .Y(_01201_),
    .A1(_00640_),
    .A2(_01111_));
 sg13g2_a221oi_1 _06635_ (.B2(net1264),
    .C1(_01201_),
    .B1(_01200_),
    .A1(net1122),
    .Y(_01202_),
    .A2(_01117_));
 sg13g2_nor2_1 _06636_ (.A(net1119),
    .B(_01122_),
    .Y(_01203_));
 sg13g2_inv_1 _06637_ (.Y(_01204_),
    .A(_01203_));
 sg13g2_a221oi_1 _06638_ (.B2(net1255),
    .C1(_01202_),
    .B1(_01203_),
    .A1(_00778_),
    .Y(_01205_),
    .A2(_01068_));
 sg13g2_nor2_1 _06639_ (.A(_01188_),
    .B(_01189_),
    .Y(_01206_));
 sg13g2_nor2_1 _06640_ (.A(net1039),
    .B(_01206_),
    .Y(_01207_));
 sg13g2_xnor2_1 _06641_ (.Y(_01208_),
    .A(_01205_),
    .B(_01207_));
 sg13g2_and2_1 _06642_ (.A(\cordic_inst.cordic_state[62] ),
    .B(_01208_),
    .X(_01209_));
 sg13g2_xor2_1 _06643_ (.B(_01208_),
    .A(\cordic_inst.cordic_state[62] ),
    .X(_01210_));
 sg13g2_and2_1 _06644_ (.A(_01198_),
    .B(_01210_),
    .X(_01211_));
 sg13g2_o21ai_1 _06645_ (.B1(net1095),
    .Y(_01212_),
    .A1(_01198_),
    .A2(_01210_));
 sg13g2_a21oi_1 _06646_ (.A1(net1316),
    .A2(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .Y(_01213_),
    .B1(net1310));
 sg13g2_o21ai_1 _06647_ (.B1(_01213_),
    .Y(_01214_),
    .A1(_01211_),
    .A2(_01212_));
 sg13g2_o21ai_1 _06648_ (.B1(_01214_),
    .Y(_01215_),
    .A1(net1128),
    .A2(net1359));
 sg13g2_nand2_1 _06649_ (.Y(_01216_),
    .A(net460),
    .B(net1085));
 sg13g2_a21oi_1 _06650_ (.A1(_01215_),
    .A2(_01216_),
    .Y(_00196_),
    .B1(net1479));
 sg13g2_a21oi_1 _06651_ (.A1(_01198_),
    .A2(_01210_),
    .Y(_01217_),
    .B1(_01209_));
 sg13g2_mux2_1 _06652_ (.A0(_01137_),
    .A1(_01148_),
    .S(net1269),
    .X(_01218_));
 sg13g2_nand2b_1 _06653_ (.Y(_01219_),
    .B(net1261),
    .A_N(_01218_));
 sg13g2_nor2_1 _06654_ (.A(_00640_),
    .B(_01138_),
    .Y(_01220_));
 sg13g2_o21ai_1 _06655_ (.B1(net1140),
    .Y(_01221_),
    .A1(net1119),
    .A2(_01144_));
 sg13g2_nor2_1 _06656_ (.A(_01220_),
    .B(_01221_),
    .Y(_01222_));
 sg13g2_a21oi_2 _06657_ (.B1(_01068_),
    .Y(_01223_),
    .A2(_01222_),
    .A1(_01219_));
 sg13g2_a21oi_1 _06658_ (.A1(_01205_),
    .A2(_01206_),
    .Y(_01224_),
    .B1(net1040));
 sg13g2_xnor2_1 _06659_ (.Y(_01225_),
    .A(_01223_),
    .B(_01224_));
 sg13g2_nand2_1 _06660_ (.Y(_01226_),
    .A(\cordic_inst.cordic_state[63] ),
    .B(_01225_));
 sg13g2_xnor2_1 _06661_ (.Y(_01227_),
    .A(\cordic_inst.cordic_state[63] ),
    .B(_01225_));
 sg13g2_xor2_1 _06662_ (.B(_01227_),
    .A(_01217_),
    .X(_01228_));
 sg13g2_a221oi_1 _06663_ (.B2(net1126),
    .C1(net1087),
    .B1(_04829_),
    .A1(net1309),
    .Y(_01229_),
    .A2(_04810_));
 sg13g2_o21ai_1 _06664_ (.B1(_01229_),
    .Y(_01230_),
    .A1(net1049),
    .A2(_01228_));
 sg13g2_a21oi_1 _06665_ (.A1(net495),
    .A2(net1087),
    .Y(_01231_),
    .B1(net1479));
 sg13g2_nand2_1 _06666_ (.Y(_00197_),
    .A(_01230_),
    .B(_01231_));
 sg13g2_o21ai_1 _06667_ (.B1(_01226_),
    .Y(_01232_),
    .A1(_01217_),
    .A2(_01227_));
 sg13g2_or2_1 _06668_ (.X(_01233_),
    .B(_01066_),
    .A(net1136));
 sg13g2_nor2_1 _06669_ (.A(net1265),
    .B(_01051_),
    .Y(_01234_));
 sg13g2_nor2_1 _06670_ (.A(net1256),
    .B(_01234_),
    .Y(_01235_));
 sg13g2_a21oi_1 _06671_ (.A1(_01233_),
    .A2(_01235_),
    .Y(_01236_),
    .B1(_01068_));
 sg13g2_nand3_1 _06672_ (.B(_01206_),
    .C(_01223_),
    .A(_01205_),
    .Y(_01237_));
 sg13g2_nand2_1 _06673_ (.Y(_01238_),
    .A(net1044),
    .B(_01237_));
 sg13g2_xor2_1 _06674_ (.B(_01238_),
    .A(_01236_),
    .X(_01239_));
 sg13g2_and2_1 _06675_ (.A(\cordic_inst.cordic_state[64] ),
    .B(_01239_),
    .X(_01240_));
 sg13g2_xor2_1 _06676_ (.B(_01239_),
    .A(\cordic_inst.cordic_state[64] ),
    .X(_01241_));
 sg13g2_and2_1 _06677_ (.A(_01232_),
    .B(_01241_),
    .X(_01242_));
 sg13g2_o21ai_1 _06678_ (.B1(net1107),
    .Y(_01243_),
    .A1(_01232_),
    .A2(_01241_));
 sg13g2_o21ai_1 _06679_ (.B1(_04905_),
    .Y(_01244_),
    .A1(_01242_),
    .A2(_01243_));
 sg13g2_a22oi_1 _06680_ (.Y(_01245_),
    .B1(_04830_),
    .B2(net1125),
    .A2(_04811_),
    .A1(net1309));
 sg13g2_a22oi_1 _06681_ (.Y(_01246_),
    .B1(_01244_),
    .B2(_01245_),
    .A2(net1087),
    .A1(net487));
 sg13g2_nor2_1 _06682_ (.A(net1479),
    .B(_01246_),
    .Y(_00198_));
 sg13g2_a21oi_1 _06683_ (.A1(_01232_),
    .A2(_01241_),
    .Y(_01247_),
    .B1(_01240_));
 sg13g2_o21ai_1 _06684_ (.B1(net1140),
    .Y(_01248_),
    .A1(net1265),
    .A2(_01081_));
 sg13g2_a21oi_2 _06685_ (.B1(_01248_),
    .Y(_01249_),
    .A2(_01098_),
    .A1(net1265));
 sg13g2_a21oi_1 _06686_ (.A1(net1238),
    .A2(_00829_),
    .Y(_01250_),
    .B1(_01249_));
 sg13g2_a21o_1 _06687_ (.A2(_01235_),
    .A1(_01233_),
    .B1(_01237_),
    .X(_01251_));
 sg13g2_nand2_1 _06688_ (.Y(_01252_),
    .A(net1044),
    .B(_01251_));
 sg13g2_xor2_1 _06689_ (.B(_01252_),
    .A(_01250_),
    .X(_01253_));
 sg13g2_nand2_1 _06690_ (.Y(_01254_),
    .A(\cordic_inst.cordic_state[65] ),
    .B(_01253_));
 sg13g2_xnor2_1 _06691_ (.Y(_01255_),
    .A(\cordic_inst.cordic_state[65] ),
    .B(_01253_));
 sg13g2_xnor2_1 _06692_ (.Y(_01256_),
    .A(_01247_),
    .B(_01255_));
 sg13g2_a22oi_1 _06693_ (.Y(_01257_),
    .B1(net1177),
    .B2(net1125),
    .A2(net1466),
    .A1(net1310));
 sg13g2_o21ai_1 _06694_ (.B1(_01257_),
    .Y(_01258_),
    .A1(_04906_),
    .A2(_01256_));
 sg13g2_a21oi_1 _06695_ (.A1(net1076),
    .A2(_01258_),
    .Y(_01259_),
    .B1(net1481));
 sg13g2_o21ai_1 _06696_ (.B1(_01259_),
    .Y(_00199_),
    .A1(_04788_),
    .A2(net1076));
 sg13g2_o21ai_1 _06697_ (.B1(_01254_),
    .Y(_01260_),
    .A1(_01247_),
    .A2(_01255_));
 sg13g2_or2_1 _06698_ (.X(_01261_),
    .B(_01123_),
    .A(net1135));
 sg13g2_nor2_1 _06699_ (.A(net1264),
    .B(_01112_),
    .Y(_01262_));
 sg13g2_nor2_1 _06700_ (.A(net1255),
    .B(_01262_),
    .Y(_01263_));
 sg13g2_a22oi_1 _06701_ (.Y(_01264_),
    .B1(_01261_),
    .B2(_01263_),
    .A2(_00829_),
    .A1(net1238));
 sg13g2_inv_1 _06702_ (.Y(_01265_),
    .A(_01264_));
 sg13g2_o21ai_1 _06703_ (.B1(net1044),
    .Y(_01266_),
    .A1(_01249_),
    .A2(_01251_));
 sg13g2_xnor2_1 _06704_ (.Y(_01267_),
    .A(_01265_),
    .B(_01266_));
 sg13g2_and2_1 _06705_ (.A(\cordic_inst.cordic_state[66] ),
    .B(_01267_),
    .X(_01268_));
 sg13g2_xnor2_1 _06706_ (.Y(_01269_),
    .A(\cordic_inst.cordic_state[66] ),
    .B(_01267_));
 sg13g2_inv_2 _06707_ (.Y(_01270_),
    .A(_01269_));
 sg13g2_o21ai_1 _06708_ (.B1(net1095),
    .Y(_01271_),
    .A1(_01260_),
    .A2(_01270_));
 sg13g2_a21o_1 _06709_ (.A2(_01270_),
    .A1(_01260_),
    .B1(_01271_),
    .X(_01272_));
 sg13g2_a21oi_1 _06710_ (.A1(net1315),
    .A2(net1173),
    .Y(_01273_),
    .B1(net1308));
 sg13g2_a22oi_1 _06711_ (.Y(_01274_),
    .B1(_01272_),
    .B2(_01273_),
    .A2(_04813_),
    .A1(net1307));
 sg13g2_o21ai_1 _06712_ (.B1(net1499),
    .Y(_01275_),
    .A1(net1083),
    .A2(_01274_));
 sg13g2_a21oi_1 _06713_ (.A1(_04787_),
    .A2(net1083),
    .Y(_00200_),
    .B1(_01275_));
 sg13g2_a21oi_1 _06714_ (.A1(_01260_),
    .A2(_01270_),
    .Y(_01276_),
    .B1(_01268_));
 sg13g2_nand3_1 _06715_ (.B(_01147_),
    .C(_01149_),
    .A(net1261),
    .Y(_01277_));
 sg13g2_nor2_1 _06716_ (.A(net1264),
    .B(_01139_),
    .Y(_01278_));
 sg13g2_nor2_1 _06717_ (.A(net1253),
    .B(_01278_),
    .Y(_01279_));
 sg13g2_a22oi_1 _06718_ (.Y(_01280_),
    .B1(_01277_),
    .B2(_01279_),
    .A2(_00861_),
    .A1(net1237));
 sg13g2_nor3_1 _06719_ (.A(_01249_),
    .B(_01251_),
    .C(_01265_),
    .Y(_01281_));
 sg13g2_nor2_1 _06720_ (.A(net1039),
    .B(_01281_),
    .Y(_01282_));
 sg13g2_xor2_1 _06721_ (.B(_01282_),
    .A(_01280_),
    .X(_01283_));
 sg13g2_inv_1 _06722_ (.Y(_01284_),
    .A(_01283_));
 sg13g2_nor2_1 _06723_ (.A(net1236),
    .B(_01284_),
    .Y(_01285_));
 sg13g2_xnor2_1 _06724_ (.Y(_01286_),
    .A(net1236),
    .B(_01283_));
 sg13g2_a221oi_1 _06725_ (.B2(net1236),
    .C1(_01268_),
    .B1(_01284_),
    .A1(_01260_),
    .Y(_01287_),
    .A2(_01270_));
 sg13g2_nand2_1 _06726_ (.Y(_01288_),
    .A(_01276_),
    .B(_01286_));
 sg13g2_nor2_1 _06727_ (.A(_01276_),
    .B(_01286_),
    .Y(_01289_));
 sg13g2_nor2_1 _06728_ (.A(net1049),
    .B(_01289_),
    .Y(_01290_));
 sg13g2_o21ai_1 _06729_ (.B1(net1075),
    .Y(_01291_),
    .A1(net1168),
    .A2(_04903_));
 sg13g2_a221oi_1 _06730_ (.B2(_01290_),
    .C1(_01291_),
    .B1(_01288_),
    .A1(net1310),
    .Y(_01292_),
    .A2(_04814_));
 sg13g2_a21oi_1 _06731_ (.A1(net1236),
    .A2(net1086),
    .Y(_01293_),
    .B1(_01292_));
 sg13g2_nand2_1 _06732_ (.Y(_00201_),
    .A(net1499),
    .B(_01293_));
 sg13g2_nand2b_1 _06733_ (.Y(_01294_),
    .B(net1238),
    .A_N(_00874_));
 sg13g2_nor2_1 _06734_ (.A(net1134),
    .B(_01065_),
    .Y(_01295_));
 sg13g2_o21ai_1 _06735_ (.B1(_00828_),
    .Y(_01296_),
    .A1(net1261),
    .A2(_01164_));
 sg13g2_o21ai_1 _06736_ (.B1(_01294_),
    .Y(_01297_),
    .A1(_01295_),
    .A2(_01296_));
 sg13g2_a21oi_1 _06737_ (.A1(_01280_),
    .A2(_01281_),
    .Y(_01298_),
    .B1(net1040));
 sg13g2_xnor2_1 _06738_ (.Y(_01299_),
    .A(_01297_),
    .B(_01298_));
 sg13g2_nor2b_1 _06739_ (.A(_01299_),
    .B_N(\cordic_inst.cordic_state[68] ),
    .Y(_01300_));
 sg13g2_xor2_1 _06740_ (.B(_01299_),
    .A(\cordic_inst.cordic_state[68] ),
    .X(_01301_));
 sg13g2_nor3_1 _06741_ (.A(_01285_),
    .B(_01287_),
    .C(_01301_),
    .Y(_01302_));
 sg13g2_o21ai_1 _06742_ (.B1(_01301_),
    .Y(_01303_),
    .A1(_01285_),
    .A2(_01287_));
 sg13g2_nand2_1 _06743_ (.Y(_01304_),
    .A(net1094),
    .B(_01303_));
 sg13g2_a21oi_1 _06744_ (.A1(net1315),
    .A2(net1162),
    .Y(_01305_),
    .B1(net1308));
 sg13g2_o21ai_1 _06745_ (.B1(_01305_),
    .Y(_01306_),
    .A1(_01302_),
    .A2(_01304_));
 sg13g2_a21oi_1 _06746_ (.A1(net1308),
    .A2(_04815_),
    .Y(_01307_),
    .B1(net1085));
 sg13g2_a22oi_1 _06747_ (.Y(_01308_),
    .B1(_01306_),
    .B2(_01307_),
    .A2(net1083),
    .A1(net476));
 sg13g2_nor2_1 _06748_ (.A(net1478),
    .B(_01308_),
    .Y(_00202_));
 sg13g2_nor2_1 _06749_ (.A(_01300_),
    .B(_01302_),
    .Y(_01309_));
 sg13g2_o21ai_1 _06750_ (.B1(_00828_),
    .Y(_01310_),
    .A1(net1261),
    .A2(_01182_));
 sg13g2_a21o_1 _06751_ (.A2(_01096_),
    .A1(net1260),
    .B1(_01310_),
    .X(_01311_));
 sg13g2_nand2_1 _06752_ (.Y(_01312_),
    .A(_01294_),
    .B(_01311_));
 sg13g2_a21oi_1 _06753_ (.A1(net1044),
    .A2(_01297_),
    .Y(_01313_),
    .B1(_01298_));
 sg13g2_xor2_1 _06754_ (.B(_01313_),
    .A(_01312_),
    .X(_01314_));
 sg13g2_nor2b_1 _06755_ (.A(\cordic_inst.cordic_state[69] ),
    .B_N(_01314_),
    .Y(_01315_));
 sg13g2_nor2b_1 _06756_ (.A(_01314_),
    .B_N(\cordic_inst.cordic_state[69] ),
    .Y(_01316_));
 sg13g2_nor2_1 _06757_ (.A(_01315_),
    .B(_01316_),
    .Y(_01317_));
 sg13g2_xnor2_1 _06758_ (.Y(_01318_),
    .A(_01309_),
    .B(_01317_));
 sg13g2_nand2_1 _06759_ (.Y(_01319_),
    .A(net1108),
    .B(_01318_));
 sg13g2_a22oi_1 _06760_ (.Y(_01320_),
    .B1(net1158),
    .B2(net1126),
    .A2(net1447),
    .A1(net1307));
 sg13g2_a21oi_1 _06761_ (.A1(_01319_),
    .A2(_01320_),
    .Y(_01321_),
    .B1(net1083));
 sg13g2_a21oi_1 _06762_ (.A1(net466),
    .A2(net1083),
    .Y(_01322_),
    .B1(_01321_));
 sg13g2_nand2_1 _06763_ (.Y(_00203_),
    .A(net1500),
    .B(_01322_));
 sg13g2_nand2b_1 _06764_ (.Y(_01323_),
    .B(net1239),
    .A_N(_00906_));
 sg13g2_a21oi_1 _06765_ (.A1(net1129),
    .A2(_01064_),
    .Y(_01324_),
    .B1(net1134));
 sg13g2_o21ai_1 _06766_ (.B1(_00828_),
    .Y(_01325_),
    .A1(net1261),
    .A2(_01199_));
 sg13g2_o21ai_1 _06767_ (.B1(_01323_),
    .Y(_01326_),
    .A1(_01324_),
    .A2(_01325_));
 sg13g2_nor2_1 _06768_ (.A(net1038),
    .B(_01311_),
    .Y(_01327_));
 sg13g2_nor2b_1 _06769_ (.A(_01327_),
    .B_N(_01313_),
    .Y(_01328_));
 sg13g2_xnor2_1 _06770_ (.Y(_01329_),
    .A(_01326_),
    .B(_01328_));
 sg13g2_and2_1 _06771_ (.A(\cordic_inst.cordic_state[70] ),
    .B(_01329_),
    .X(_01330_));
 sg13g2_inv_1 _06772_ (.Y(_01331_),
    .A(_01330_));
 sg13g2_xnor2_1 _06773_ (.Y(_01332_),
    .A(\cordic_inst.cordic_state[70] ),
    .B(_01329_));
 sg13g2_nor3_1 _06774_ (.A(_01300_),
    .B(_01302_),
    .C(_01316_),
    .Y(_01333_));
 sg13g2_o21ai_1 _06775_ (.B1(_01332_),
    .Y(_01334_),
    .A1(_01315_),
    .A2(_01333_));
 sg13g2_or3_1 _06776_ (.A(_01315_),
    .B(_01332_),
    .C(_01333_),
    .X(_01335_));
 sg13g2_and2_1 _06777_ (.A(net1095),
    .B(_01335_),
    .X(_01336_));
 sg13g2_a221oi_1 _06778_ (.B2(_01336_),
    .C1(net1307),
    .B1(_01334_),
    .A1(net1315),
    .Y(_01337_),
    .A2(net1152));
 sg13g2_o21ai_1 _06779_ (.B1(net1075),
    .Y(_01338_),
    .A1(net1128),
    .A2(net1442));
 sg13g2_nor2_1 _06780_ (.A(_01337_),
    .B(_01338_),
    .Y(_01339_));
 sg13g2_a21oi_1 _06781_ (.A1(net455),
    .A2(net1083),
    .Y(_01340_),
    .B1(_01339_));
 sg13g2_nor2_1 _06782_ (.A(net1478),
    .B(_01340_),
    .Y(_00204_));
 sg13g2_a22oi_1 _06783_ (.Y(_01341_),
    .B1(_01218_),
    .B2(net1134),
    .A2(_00923_),
    .A1(net1237));
 sg13g2_o21ai_1 _06784_ (.B1(_01323_),
    .Y(_01342_),
    .A1(net1252),
    .A2(_01341_));
 sg13g2_nand2_1 _06785_ (.Y(_01343_),
    .A(net1042),
    .B(_01326_));
 sg13g2_nand2_1 _06786_ (.Y(_01344_),
    .A(_01328_),
    .B(_01343_));
 sg13g2_xnor2_1 _06787_ (.Y(_01345_),
    .A(_01342_),
    .B(_01344_));
 sg13g2_nor2_1 _06788_ (.A(_04786_),
    .B(_01345_),
    .Y(_01346_));
 sg13g2_xnor2_1 _06789_ (.Y(_01347_),
    .A(\cordic_inst.cordic_state[71] ),
    .B(_01345_));
 sg13g2_inv_1 _06790_ (.Y(_01348_),
    .A(_01347_));
 sg13g2_nand3_1 _06791_ (.B(_01335_),
    .C(_01348_),
    .A(_01331_),
    .Y(_01349_));
 sg13g2_a21oi_1 _06792_ (.A1(_01331_),
    .A2(_01335_),
    .Y(_01350_),
    .B1(_01348_));
 sg13g2_nand2_1 _06793_ (.Y(_01351_),
    .A(net1108),
    .B(_01349_));
 sg13g2_a22oi_1 _06794_ (.Y(_01352_),
    .B1(net1146),
    .B2(net1126),
    .A2(net1437),
    .A1(net1307));
 sg13g2_o21ai_1 _06795_ (.B1(_01352_),
    .Y(_01353_),
    .A1(_01350_),
    .A2(_01351_));
 sg13g2_a21oi_1 _06796_ (.A1(net1075),
    .A2(_01353_),
    .Y(_01354_),
    .B1(net1478));
 sg13g2_o21ai_1 _06797_ (.B1(_01354_),
    .Y(_00205_),
    .A1(_04786_),
    .A2(net1075));
 sg13g2_nor2b_1 _06798_ (.A(_00938_),
    .B_N(net1239),
    .Y(_01355_));
 sg13g2_a21oi_1 _06799_ (.A1(net1138),
    .A2(_01067_),
    .Y(_01356_),
    .B1(_01355_));
 sg13g2_a21oi_1 _06800_ (.A1(net1044),
    .A2(_01342_),
    .Y(_01357_),
    .B1(_01344_));
 sg13g2_xnor2_1 _06801_ (.Y(_01358_),
    .A(_01356_),
    .B(_01357_));
 sg13g2_nor2b_1 _06802_ (.A(_01358_),
    .B_N(\cordic_inst.cordic_state[72] ),
    .Y(_01359_));
 sg13g2_xnor2_1 _06803_ (.Y(_01360_),
    .A(\cordic_inst.cordic_state[72] ),
    .B(_01358_));
 sg13g2_nor2_1 _06804_ (.A(_01346_),
    .B(_01350_),
    .Y(_01361_));
 sg13g2_nor2b_1 _06805_ (.A(_01361_),
    .B_N(_01360_),
    .Y(_01362_));
 sg13g2_o21ai_1 _06806_ (.B1(_01360_),
    .Y(_01363_),
    .A1(_01346_),
    .A2(_01350_));
 sg13g2_nand2b_1 _06807_ (.Y(_01364_),
    .B(_01361_),
    .A_N(_01360_));
 sg13g2_nand3_1 _06808_ (.B(_01363_),
    .C(_01364_),
    .A(net1095),
    .Y(_01365_));
 sg13g2_a21oi_1 _06809_ (.A1(net1315),
    .A2(net1351),
    .Y(_01366_),
    .B1(net1307));
 sg13g2_o21ai_1 _06810_ (.B1(net1075),
    .Y(_01367_),
    .A1(net1128),
    .A2(net1433));
 sg13g2_a21oi_1 _06811_ (.A1(_01365_),
    .A2(_01366_),
    .Y(_01368_),
    .B1(_01367_));
 sg13g2_a21oi_1 _06812_ (.A1(net430),
    .A2(net1083),
    .Y(_01369_),
    .B1(_01368_));
 sg13g2_nor2_1 _06813_ (.A(net1478),
    .B(net431),
    .Y(_00206_));
 sg13g2_nor3_1 _06814_ (.A(net1254),
    .B(net1266),
    .C(_01098_),
    .Y(_01370_));
 sg13g2_nor2_1 _06815_ (.A(_01355_),
    .B(_01370_),
    .Y(_01371_));
 sg13g2_o21ai_1 _06816_ (.B1(_01357_),
    .Y(_01372_),
    .A1(net1038),
    .A2(_01356_));
 sg13g2_xnor2_1 _06817_ (.Y(_01373_),
    .A(_01371_),
    .B(_01372_));
 sg13g2_inv_1 _06818_ (.Y(_01374_),
    .A(_01373_));
 sg13g2_nor2_1 _06819_ (.A(net1235),
    .B(_01373_),
    .Y(_01375_));
 sg13g2_xnor2_1 _06820_ (.Y(_01376_),
    .A(net1235),
    .B(_01373_));
 sg13g2_nor2_1 _06821_ (.A(_01359_),
    .B(_01362_),
    .Y(_01377_));
 sg13g2_o21ai_1 _06822_ (.B1(net1109),
    .Y(_01378_),
    .A1(_01376_),
    .A2(_01377_));
 sg13g2_a21o_1 _06823_ (.A2(_01377_),
    .A1(_01376_),
    .B1(_01378_),
    .X(_01379_));
 sg13g2_a221oi_1 _06824_ (.B2(net1124),
    .C1(net1084),
    .B1(net1343),
    .A1(net1304),
    .Y(_01380_),
    .A2(net1429));
 sg13g2_a22oi_1 _06825_ (.Y(_01381_),
    .B1(_01379_),
    .B2(_01380_),
    .A2(net1084),
    .A1(_04785_));
 sg13g2_nand2b_1 _06826_ (.Y(_00207_),
    .B(net1500),
    .A_N(_01381_));
 sg13g2_a22oi_1 _06827_ (.Y(_01382_),
    .B1(_01124_),
    .B2(net1137),
    .A2(_00968_),
    .A1(net1239));
 sg13g2_a21oi_1 _06828_ (.A1(net1042),
    .A2(_01370_),
    .Y(_01383_),
    .B1(_01372_));
 sg13g2_or2_1 _06829_ (.X(_01384_),
    .B(_01383_),
    .A(_01382_));
 sg13g2_nand2_2 _06830_ (.Y(_01385_),
    .A(_01382_),
    .B(_01383_));
 sg13g2_and3_1 _06831_ (.X(_01386_),
    .A(\cordic_inst.cordic_state[74] ),
    .B(_01384_),
    .C(_01385_));
 sg13g2_a21oi_1 _06832_ (.A1(_01384_),
    .A2(_01385_),
    .Y(_01387_),
    .B1(\cordic_inst.cordic_state[74] ));
 sg13g2_or2_1 _06833_ (.X(_01388_),
    .B(_01387_),
    .A(_01386_));
 sg13g2_a21oi_1 _06834_ (.A1(net1235),
    .A2(_01373_),
    .Y(_01389_),
    .B1(_01359_));
 sg13g2_a21o_1 _06835_ (.A2(_01389_),
    .A1(_01363_),
    .B1(_01375_),
    .X(_01390_));
 sg13g2_a221oi_1 _06836_ (.B2(_01363_),
    .C1(_01388_),
    .B1(_01389_),
    .A1(_04785_),
    .Y(_01391_),
    .A2(_01374_));
 sg13g2_a21oi_1 _06837_ (.A1(_01388_),
    .A2(_01390_),
    .Y(_01392_),
    .B1(_04913_));
 sg13g2_nand2b_1 _06838_ (.Y(_01393_),
    .B(_01392_),
    .A_N(_01391_));
 sg13g2_a21oi_1 _06839_ (.A1(net1313),
    .A2(net1338),
    .Y(_01394_),
    .B1(net1304));
 sg13g2_o21ai_1 _06840_ (.B1(net1073),
    .Y(_01395_),
    .A1(net1127),
    .A2(net1424));
 sg13g2_a21oi_1 _06841_ (.A1(_01393_),
    .A2(_01394_),
    .Y(_01396_),
    .B1(_01395_));
 sg13g2_a21oi_1 _06842_ (.A1(net454),
    .A2(net1084),
    .Y(_01397_),
    .B1(_01396_));
 sg13g2_nor2_1 _06843_ (.A(net1477),
    .B(_01397_),
    .Y(_00208_));
 sg13g2_nor2_1 _06844_ (.A(_01386_),
    .B(_01391_),
    .Y(_01398_));
 sg13g2_nand2_1 _06845_ (.Y(_01399_),
    .A(net1042),
    .B(_01385_));
 sg13g2_and2_1 _06846_ (.A(net1137),
    .B(_01150_),
    .X(_01400_));
 sg13g2_a21oi_1 _06847_ (.A1(net1239),
    .A2(_00968_),
    .Y(_01401_),
    .B1(_01400_));
 sg13g2_xnor2_1 _06848_ (.Y(_01402_),
    .A(_01399_),
    .B(_01401_));
 sg13g2_nand2b_1 _06849_ (.Y(_01403_),
    .B(_01402_),
    .A_N(\cordic_inst.cordic_state[75] ));
 sg13g2_nand2b_1 _06850_ (.Y(_01404_),
    .B(\cordic_inst.cordic_state[75] ),
    .A_N(_01402_));
 sg13g2_nand2_1 _06851_ (.Y(_01405_),
    .A(_01403_),
    .B(_01404_));
 sg13g2_nand2b_1 _06852_ (.Y(_01406_),
    .B(_01404_),
    .A_N(_01386_));
 sg13g2_xnor2_1 _06853_ (.Y(_01407_),
    .A(_01398_),
    .B(_01405_));
 sg13g2_nand2b_1 _06854_ (.Y(_01408_),
    .B(net1109),
    .A_N(_01407_));
 sg13g2_a22oi_1 _06855_ (.Y(_01409_),
    .B1(net1335),
    .B2(net1126),
    .A2(net1421),
    .A1(net1307));
 sg13g2_a21oi_1 _06856_ (.A1(_01408_),
    .A2(_01409_),
    .Y(_01410_),
    .B1(net1084));
 sg13g2_a21oi_1 _06857_ (.A1(net480),
    .A2(net1084),
    .Y(_01411_),
    .B1(_01410_));
 sg13g2_nand2_1 _06858_ (.Y(_00209_),
    .A(net1500),
    .B(_01411_));
 sg13g2_nand2_1 _06859_ (.Y(_01412_),
    .A(net1239),
    .B(_00996_));
 sg13g2_o21ai_1 _06860_ (.B1(_01412_),
    .Y(_01413_),
    .A1(net1252),
    .A2(_01169_));
 sg13g2_inv_1 _06861_ (.Y(_01414_),
    .A(_01413_));
 sg13g2_o21ai_1 _06862_ (.B1(net1043),
    .Y(_01415_),
    .A1(_01385_),
    .A2(_01400_));
 sg13g2_xnor2_1 _06863_ (.Y(_01416_),
    .A(_01413_),
    .B(_01415_));
 sg13g2_nand2_1 _06864_ (.Y(_01417_),
    .A(\cordic_inst.cordic_state[76] ),
    .B(_01416_));
 sg13g2_xnor2_1 _06865_ (.Y(_01418_),
    .A(\cordic_inst.cordic_state[76] ),
    .B(_01416_));
 sg13g2_o21ai_1 _06866_ (.B1(_01403_),
    .Y(_01419_),
    .A1(_01391_),
    .A2(_01406_));
 sg13g2_or2_1 _06867_ (.X(_01420_),
    .B(_01419_),
    .A(_01418_));
 sg13g2_a21oi_1 _06868_ (.A1(_01418_),
    .A2(_01419_),
    .Y(_01421_),
    .B1(_04913_));
 sg13g2_a221oi_1 _06869_ (.B2(_01421_),
    .C1(net1304),
    .B1(_01420_),
    .A1(net1313),
    .Y(_01422_),
    .A2(net1332));
 sg13g2_nor2_1 _06870_ (.A(net1127),
    .B(net1418),
    .Y(_01423_));
 sg13g2_nand2_1 _06871_ (.Y(_01424_),
    .A(net509),
    .B(net1084));
 sg13g2_o21ai_1 _06872_ (.B1(_01424_),
    .Y(_01425_),
    .A1(_01422_),
    .A2(_01423_));
 sg13g2_and2_1 _06873_ (.A(net1490),
    .B(_01425_),
    .X(_00210_));
 sg13g2_nand2_1 _06874_ (.Y(_01426_),
    .A(_01417_),
    .B(_01420_));
 sg13g2_a21oi_1 _06875_ (.A1(_01414_),
    .A2(_01415_),
    .Y(_01427_),
    .B1(net1038));
 sg13g2_o21ai_1 _06876_ (.B1(_01412_),
    .Y(_01428_),
    .A1(net1252),
    .A2(_01186_));
 sg13g2_xor2_1 _06877_ (.B(_01428_),
    .A(_01427_),
    .X(_01429_));
 sg13g2_or2_1 _06878_ (.X(_01430_),
    .B(_01429_),
    .A(net1234));
 sg13g2_and2_1 _06879_ (.A(net1234),
    .B(_01429_),
    .X(_01431_));
 sg13g2_xnor2_1 _06880_ (.Y(_01432_),
    .A(net1234),
    .B(_01429_));
 sg13g2_xnor2_1 _06881_ (.Y(_01433_),
    .A(_01426_),
    .B(_01432_));
 sg13g2_a22oi_1 _06882_ (.Y(_01434_),
    .B1(net1330),
    .B2(net1124),
    .A2(net1415),
    .A1(net1304));
 sg13g2_nand2_1 _06883_ (.Y(_01435_),
    .A(net1073),
    .B(_01434_));
 sg13g2_a21oi_1 _06884_ (.A1(net1109),
    .A2(_01433_),
    .Y(_01436_),
    .B1(_01435_));
 sg13g2_nor2_1 _06885_ (.A(net1234),
    .B(net1073),
    .Y(_01437_));
 sg13g2_o21ai_1 _06886_ (.B1(net1490),
    .Y(_00211_),
    .A1(_01436_),
    .A2(_01437_));
 sg13g2_o21ai_1 _06887_ (.B1(net1237),
    .Y(_01438_),
    .A1(net1253),
    .A2(_00778_));
 sg13g2_o21ai_1 _06888_ (.B1(_01438_),
    .Y(_01439_),
    .A1(net1253),
    .A2(_01204_));
 sg13g2_a21oi_1 _06889_ (.A1(net1042),
    .A2(_01428_),
    .Y(_01440_),
    .B1(_01427_));
 sg13g2_inv_1 _06890_ (.Y(_01441_),
    .A(_01440_));
 sg13g2_xnor2_1 _06891_ (.Y(_01442_),
    .A(_01439_),
    .B(_01440_));
 sg13g2_nand2_1 _06892_ (.Y(_01443_),
    .A(\cordic_inst.cordic_state[78] ),
    .B(_01442_));
 sg13g2_xnor2_1 _06893_ (.Y(_01444_),
    .A(\cordic_inst.cordic_state[78] ),
    .B(_01442_));
 sg13g2_o21ai_1 _06894_ (.B1(_01430_),
    .Y(_01445_),
    .A1(_01426_),
    .A2(_01431_));
 sg13g2_a21oi_1 _06895_ (.A1(_01444_),
    .A2(_01445_),
    .Y(_01446_),
    .B1(_04913_));
 sg13g2_o21ai_1 _06896_ (.B1(_01446_),
    .Y(_01447_),
    .A1(_01444_),
    .A2(_01445_));
 sg13g2_a21oi_1 _06897_ (.A1(net1313),
    .A2(net1327),
    .Y(_01448_),
    .B1(net1304));
 sg13g2_a22oi_1 _06898_ (.Y(_01449_),
    .B1(_01447_),
    .B2(_01448_),
    .A2(_04821_),
    .A1(net1304));
 sg13g2_o21ai_1 _06899_ (.B1(net1490),
    .Y(_01450_),
    .A1(net1081),
    .A2(_01449_));
 sg13g2_a21oi_1 _06900_ (.A1(_04784_),
    .A2(net1081),
    .Y(_00212_),
    .B1(_01450_));
 sg13g2_o21ai_1 _06901_ (.B1(_01443_),
    .Y(_01451_),
    .A1(_01444_),
    .A2(_01445_));
 sg13g2_a21oi_1 _06902_ (.A1(net1042),
    .A2(_01439_),
    .Y(_01452_),
    .B1(_01441_));
 sg13g2_xor2_1 _06903_ (.B(_01452_),
    .A(_01039_),
    .X(_01453_));
 sg13g2_a21oi_1 _06904_ (.A1(_01451_),
    .A2(_01453_),
    .Y(_01454_),
    .B1(_04909_));
 sg13g2_o21ai_1 _06905_ (.B1(_01454_),
    .Y(_01455_),
    .A1(_01451_),
    .A2(_01453_));
 sg13g2_a221oi_1 _06906_ (.B2(_01455_),
    .C1(net1302),
    .B1(_04887_),
    .A1(net1312),
    .Y(_01456_),
    .A2(net1325));
 sg13g2_o21ai_1 _06907_ (.B1(net1073),
    .Y(_01457_),
    .A1(net1127),
    .A2(net1410));
 sg13g2_a21oi_1 _06908_ (.A1(net1233),
    .A2(net1081),
    .Y(_01458_),
    .B1(net1477));
 sg13g2_o21ai_1 _06909_ (.B1(_01458_),
    .Y(_00213_),
    .A1(_01456_),
    .A2(_01457_));
 sg13g2_nor2b_1 _06910_ (.A(cordic_busy),
    .B_N(net194),
    .Y(_01459_));
 sg13g2_o21ai_1 _06911_ (.B1(net194),
    .Y(_01460_),
    .A1(\cordic_inst.result_ready ),
    .A2(cordic_busy));
 sg13g2_a21oi_1 _06912_ (.A1(net1108),
    .A2(net195),
    .Y(_00214_),
    .B1(net1484));
 sg13g2_nor4_1 _06913_ (.A(_04782_),
    .B(cordic_en_get_atan2),
    .C(cordic_en_get_sqrt),
    .D(net325),
    .Y(_01461_));
 sg13g2_a21oi_1 _06914_ (.A1(_04782_),
    .A2(_01459_),
    .Y(_01462_),
    .B1(net326));
 sg13g2_nor2_1 _06915_ (.A(_04907_),
    .B(net327),
    .Y(_00215_));
 sg13g2_nor2b_1 _06916_ (.A(_04865_),
    .B_N(net1123),
    .Y(_01463_));
 sg13g2_mux2_1 _06917_ (.A0(net1227),
    .A1(net1),
    .S(net1067),
    .X(_00216_));
 sg13g2_nand2_1 _06918_ (.Y(_01464_),
    .A(net2),
    .B(net1067));
 sg13g2_o21ai_1 _06919_ (.B1(_01464_),
    .Y(_00217_),
    .A1(_04823_),
    .A2(net1067));
 sg13g2_nand2_1 _06920_ (.Y(_01465_),
    .A(net3),
    .B(net1068));
 sg13g2_o21ai_1 _06921_ (.B1(_01465_),
    .Y(_00218_),
    .A1(_04824_),
    .A2(net1068));
 sg13g2_nand2_1 _06922_ (.Y(_01466_),
    .A(net4),
    .B(net1068));
 sg13g2_o21ai_1 _06923_ (.B1(_01466_),
    .Y(_00219_),
    .A1(_04825_),
    .A2(net1067));
 sg13g2_nand2_1 _06924_ (.Y(_01467_),
    .A(net5),
    .B(net1067));
 sg13g2_o21ai_1 _06925_ (.B1(_01467_),
    .Y(_00220_),
    .A1(_04826_),
    .A2(net1067));
 sg13g2_nand2_1 _06926_ (.Y(_01468_),
    .A(net6),
    .B(net1069));
 sg13g2_o21ai_1 _06927_ (.B1(_01468_),
    .Y(_00221_),
    .A1(_04827_),
    .A2(net1069));
 sg13g2_nand2_1 _06928_ (.Y(_01469_),
    .A(net7),
    .B(net1067));
 sg13g2_o21ai_1 _06929_ (.B1(_01469_),
    .Y(_00222_),
    .A1(_04828_),
    .A2(net1067));
 sg13g2_nand2_1 _06930_ (.Y(_01470_),
    .A(net8),
    .B(net1069));
 sg13g2_o21ai_1 _06931_ (.B1(_01470_),
    .Y(_00223_),
    .A1(_04829_),
    .A2(net1069));
 sg13g2_nand2_1 _06932_ (.Y(_01471_),
    .A(net1406),
    .B(net1192));
 sg13g2_nor3_1 _06933_ (.A(_04805_),
    .B(_04830_),
    .C(_01471_),
    .Y(_01472_));
 sg13g2_nand2_1 _06934_ (.Y(_01473_),
    .A(net1390),
    .B(net1192));
 sg13g2_and4_1 _06935_ (.A(net1406),
    .B(net1398),
    .C(net1187),
    .D(net1181),
    .X(_01474_));
 sg13g2_nand4_1 _06936_ (.B(net1398),
    .C(net1187),
    .A(net1407),
    .Y(_01475_),
    .D(net1181));
 sg13g2_a22oi_1 _06937_ (.Y(_01476_),
    .B1(net1181),
    .B2(net1407),
    .A2(net1187),
    .A1(net1398));
 sg13g2_or3_1 _06938_ (.A(_01473_),
    .B(_01474_),
    .C(_01476_),
    .X(_01477_));
 sg13g2_o21ai_1 _06939_ (.B1(_01473_),
    .Y(_01478_),
    .A1(_01474_),
    .A2(_01476_));
 sg13g2_and3_1 _06940_ (.X(_01479_),
    .A(_01472_),
    .B(_01477_),
    .C(_01478_));
 sg13g2_a21o_1 _06941_ (.A2(_01478_),
    .A1(_01477_),
    .B1(_01472_),
    .X(_01480_));
 sg13g2_nor2b_1 _06942_ (.A(_01479_),
    .B_N(_01480_),
    .Y(_01481_));
 sg13g2_nand2_1 _06943_ (.Y(_01482_),
    .A(net1370),
    .B(net1206));
 sg13g2_nand2_1 _06944_ (.Y(_01483_),
    .A(net1377),
    .B(net1199));
 sg13g2_nand2_1 _06945_ (.Y(_01484_),
    .A(net1383),
    .B(net1203));
 sg13g2_and4_1 _06946_ (.A(net1384),
    .B(net1377),
    .C(net1203),
    .D(net1199),
    .X(_01485_));
 sg13g2_a22oi_1 _06947_ (.Y(_01486_),
    .B1(net1199),
    .B2(net1384),
    .A2(net1203),
    .A1(net1376));
 sg13g2_nor3_1 _06948_ (.A(_01482_),
    .B(_01485_),
    .C(_01486_),
    .Y(_01487_));
 sg13g2_o21ai_1 _06949_ (.B1(_01482_),
    .Y(_01488_),
    .A1(_01485_),
    .A2(_01486_));
 sg13g2_nor2b_1 _06950_ (.A(_01487_),
    .B_N(_01488_),
    .Y(_01489_));
 sg13g2_a21o_1 _06951_ (.A2(_01489_),
    .A1(_01480_),
    .B1(_01479_),
    .X(_01490_));
 sg13g2_o21ai_1 _06952_ (.B1(_01475_),
    .Y(_01491_),
    .A1(_01473_),
    .A2(_01476_));
 sg13g2_nand2_1 _06953_ (.Y(_01492_),
    .A(net1384),
    .B(net1194));
 sg13g2_and4_1 _06954_ (.A(net1401),
    .B(net1391),
    .C(net1187),
    .D(net1179),
    .X(_01493_));
 sg13g2_nand4_1 _06955_ (.B(net1390),
    .C(net1186),
    .A(net1399),
    .Y(_01494_),
    .D(net1179));
 sg13g2_a22oi_1 _06956_ (.Y(_01495_),
    .B1(net1179),
    .B2(net1401),
    .A2(net1186),
    .A1(net1390));
 sg13g2_or3_1 _06957_ (.A(_01492_),
    .B(_01493_),
    .C(_01495_),
    .X(_01496_));
 sg13g2_o21ai_1 _06958_ (.B1(_01492_),
    .Y(_01497_),
    .A1(_01493_),
    .A2(_01495_));
 sg13g2_and3_1 _06959_ (.X(_01498_),
    .A(_01491_),
    .B(_01496_),
    .C(_01497_));
 sg13g2_nand3_1 _06960_ (.B(_01496_),
    .C(_01497_),
    .A(_01491_),
    .Y(_01499_));
 sg13g2_a21o_1 _06961_ (.A2(_01497_),
    .A1(_01496_),
    .B1(_01491_),
    .X(_01500_));
 sg13g2_nand2_1 _06962_ (.Y(_01501_),
    .A(net1363),
    .B(net1206));
 sg13g2_nand2_1 _06963_ (.Y(_01502_),
    .A(net1370),
    .B(net1203));
 sg13g2_or2_1 _06964_ (.X(_01503_),
    .B(_01502_),
    .A(_01483_));
 sg13g2_and2_1 _06965_ (.A(_01483_),
    .B(_01502_),
    .X(_01504_));
 sg13g2_xor2_1 _06966_ (.B(_01502_),
    .A(_01483_),
    .X(_01505_));
 sg13g2_xnor2_1 _06967_ (.Y(_01506_),
    .A(_01501_),
    .B(_01505_));
 sg13g2_nand3_1 _06968_ (.B(_01500_),
    .C(_01506_),
    .A(_01499_),
    .Y(_01507_));
 sg13g2_a21o_1 _06969_ (.A2(_01500_),
    .A1(_01499_),
    .B1(_01506_),
    .X(_01508_));
 sg13g2_and3_1 _06970_ (.X(_01509_),
    .A(_01490_),
    .B(_01507_),
    .C(_01508_));
 sg13g2_nand2_1 _06971_ (.Y(_01510_),
    .A(net1356),
    .B(net1212));
 sg13g2_nand2_1 _06972_ (.Y(_01511_),
    .A(net1362),
    .B(net1217));
 sg13g2_and4_1 _06973_ (.A(net1362),
    .B(net1356),
    .C(net1217),
    .D(net1212),
    .X(_01512_));
 sg13g2_nand2_1 _06974_ (.Y(_01513_),
    .A(net1469),
    .B(net1226));
 sg13g2_a22oi_1 _06975_ (.Y(_01514_),
    .B1(net1212),
    .B2(net1362),
    .A2(net1217),
    .A1(net1356));
 sg13g2_nor3_1 _06976_ (.A(_01512_),
    .B(_01513_),
    .C(_01514_),
    .Y(_01515_));
 sg13g2_or2_1 _06977_ (.X(_01516_),
    .B(_01515_),
    .A(_01512_));
 sg13g2_inv_1 _06978_ (.Y(_01517_),
    .A(_01516_));
 sg13g2_or2_1 _06979_ (.X(_01518_),
    .B(_01487_),
    .A(_01485_));
 sg13g2_nand2_1 _06980_ (.Y(_01519_),
    .A(net1464),
    .B(net1226));
 sg13g2_nand2_1 _06981_ (.Y(_01520_),
    .A(net1473),
    .B(net1212));
 sg13g2_nand2_1 _06982_ (.Y(_01521_),
    .A(net1473),
    .B(net1217));
 sg13g2_or2_1 _06983_ (.X(_01522_),
    .B(_01521_),
    .A(_01510_));
 sg13g2_xnor2_1 _06984_ (.Y(_01523_),
    .A(_01510_),
    .B(_01521_));
 sg13g2_xor2_1 _06985_ (.B(_01523_),
    .A(_01519_),
    .X(_01524_));
 sg13g2_nand2_1 _06986_ (.Y(_01525_),
    .A(_01518_),
    .B(_01524_));
 sg13g2_xnor2_1 _06987_ (.Y(_01526_),
    .A(_01518_),
    .B(_01524_));
 sg13g2_xnor2_1 _06988_ (.Y(_01527_),
    .A(_01517_),
    .B(_01526_));
 sg13g2_a21oi_1 _06989_ (.A1(_01507_),
    .A2(_01508_),
    .Y(_01528_),
    .B1(_01490_));
 sg13g2_or3_1 _06990_ (.A(_01509_),
    .B(_01527_),
    .C(_01528_),
    .X(_01529_));
 sg13g2_nand2b_1 _06991_ (.Y(_01530_),
    .B(_01529_),
    .A_N(_01509_));
 sg13g2_o21ai_1 _06992_ (.B1(_01525_),
    .Y(_01531_),
    .A1(_01517_),
    .A2(_01526_));
 sg13g2_nand2_1 _06993_ (.Y(_01532_),
    .A(_01530_),
    .B(_01531_));
 sg13g2_o21ai_1 _06994_ (.B1(_01522_),
    .Y(_01533_),
    .A1(_01519_),
    .A2(_01523_));
 sg13g2_inv_1 _06995_ (.Y(_01534_),
    .A(_01533_));
 sg13g2_o21ai_1 _06996_ (.B1(_01503_),
    .Y(_01535_),
    .A1(_01501_),
    .A2(_01504_));
 sg13g2_nand2_1 _06997_ (.Y(_01536_),
    .A(net1458),
    .B(net1226));
 sg13g2_nand2_1 _06998_ (.Y(_01537_),
    .A(net1469),
    .B(net1212));
 sg13g2_nand2_1 _06999_ (.Y(_01538_),
    .A(net1469),
    .B(net1217));
 sg13g2_or2_1 _07000_ (.X(_01539_),
    .B(_01537_),
    .A(_01521_));
 sg13g2_xnor2_1 _07001_ (.Y(_01540_),
    .A(_01520_),
    .B(_01538_));
 sg13g2_xor2_1 _07002_ (.B(_01540_),
    .A(_01536_),
    .X(_01541_));
 sg13g2_nand2_1 _07003_ (.Y(_01542_),
    .A(_01535_),
    .B(_01541_));
 sg13g2_xnor2_1 _07004_ (.Y(_01543_),
    .A(_01535_),
    .B(_01541_));
 sg13g2_xnor2_1 _07005_ (.Y(_01544_),
    .A(_01534_),
    .B(_01543_));
 sg13g2_a21o_1 _07006_ (.A2(_01506_),
    .A1(_01500_),
    .B1(_01498_),
    .X(_01545_));
 sg13g2_o21ai_1 _07007_ (.B1(_01494_),
    .Y(_01546_),
    .A1(_01492_),
    .A2(_01495_));
 sg13g2_nand2_1 _07008_ (.Y(_01547_),
    .A(net1376),
    .B(net1194));
 sg13g2_and4_1 _07009_ (.A(net1391),
    .B(net1384),
    .C(net1186),
    .D(net1180),
    .X(_01548_));
 sg13g2_nand4_1 _07010_ (.B(net1383),
    .C(net1186),
    .A(net1391),
    .Y(_01549_),
    .D(net1179));
 sg13g2_a22oi_1 _07011_ (.Y(_01550_),
    .B1(net1179),
    .B2(net1391),
    .A2(net1186),
    .A1(net1383));
 sg13g2_or3_1 _07012_ (.A(_01547_),
    .B(_01548_),
    .C(_01550_),
    .X(_01551_));
 sg13g2_o21ai_1 _07013_ (.B1(_01547_),
    .Y(_01552_),
    .A1(_01548_),
    .A2(_01550_));
 sg13g2_and3_1 _07014_ (.X(_01553_),
    .A(_01546_),
    .B(_01551_),
    .C(_01552_));
 sg13g2_nand3_1 _07015_ (.B(_01551_),
    .C(_01552_),
    .A(_01546_),
    .Y(_01554_));
 sg13g2_a21oi_1 _07016_ (.A1(_01551_),
    .A2(_01552_),
    .Y(_01555_),
    .B1(_01546_));
 sg13g2_nand2_1 _07017_ (.Y(_01556_),
    .A(net1356),
    .B(net1206));
 sg13g2_nand2_1 _07018_ (.Y(_01557_),
    .A(net1362),
    .B(net1199));
 sg13g2_and4_1 _07019_ (.A(net1370),
    .B(net1363),
    .C(net1203),
    .D(net1199),
    .X(_01558_));
 sg13g2_a22oi_1 _07020_ (.Y(_01559_),
    .B1(net1199),
    .B2(net1370),
    .A2(net1203),
    .A1(net1363));
 sg13g2_nor3_1 _07021_ (.A(_01556_),
    .B(_01558_),
    .C(_01559_),
    .Y(_01560_));
 sg13g2_o21ai_1 _07022_ (.B1(_01556_),
    .Y(_01561_),
    .A1(_01558_),
    .A2(_01559_));
 sg13g2_nand2b_1 _07023_ (.Y(_01562_),
    .B(_01561_),
    .A_N(_01560_));
 sg13g2_or3_1 _07024_ (.A(_01553_),
    .B(_01555_),
    .C(_01562_),
    .X(_01563_));
 sg13g2_o21ai_1 _07025_ (.B1(_01562_),
    .Y(_01564_),
    .A1(_01553_),
    .A2(_01555_));
 sg13g2_and3_1 _07026_ (.X(_01565_),
    .A(_01545_),
    .B(_01563_),
    .C(_01564_));
 sg13g2_a21oi_1 _07027_ (.A1(_01563_),
    .A2(_01564_),
    .Y(_01566_),
    .B1(_01545_));
 sg13g2_or3_1 _07028_ (.A(_01544_),
    .B(_01565_),
    .C(_01566_),
    .X(_01567_));
 sg13g2_o21ai_1 _07029_ (.B1(_01544_),
    .Y(_01568_),
    .A1(_01565_),
    .A2(_01566_));
 sg13g2_nor2_2 _07030_ (.A(_04804_),
    .B(_04832_),
    .Y(_01569_));
 sg13g2_and2_1 _07031_ (.A(net1398),
    .B(net1172),
    .X(_01570_));
 sg13g2_nand2_1 _07032_ (.Y(_01571_),
    .A(_01569_),
    .B(_01570_));
 sg13g2_a22oi_1 _07033_ (.Y(_01572_),
    .B1(net1172),
    .B2(net1406),
    .A2(net1176),
    .A1(net1398));
 sg13g2_a21oi_1 _07034_ (.A1(_01569_),
    .A2(_01570_),
    .Y(_01573_),
    .B1(_01572_));
 sg13g2_a21oi_1 _07035_ (.A1(_01567_),
    .A2(_01568_),
    .Y(_01574_),
    .B1(_01573_));
 sg13g2_and3_2 _07036_ (.X(_01575_),
    .A(_01567_),
    .B(_01568_),
    .C(_01573_));
 sg13g2_o21ai_1 _07037_ (.B1(_01527_),
    .Y(_01576_),
    .A1(_01509_),
    .A2(_01528_));
 sg13g2_nand3_1 _07038_ (.B(_01569_),
    .C(_01576_),
    .A(_01529_),
    .Y(_01577_));
 sg13g2_or3_1 _07039_ (.A(_01574_),
    .B(_01575_),
    .C(_01577_),
    .X(_01578_));
 sg13g2_o21ai_1 _07040_ (.B1(_01577_),
    .Y(_01579_),
    .A1(_01574_),
    .A2(_01575_));
 sg13g2_and4_1 _07041_ (.A(net1464),
    .B(net1220),
    .C(_01578_),
    .D(_01579_),
    .X(_01580_));
 sg13g2_nand4_1 _07042_ (.B(net1220),
    .C(_01578_),
    .A(net1464),
    .Y(_01581_),
    .D(_01579_));
 sg13g2_a22oi_1 _07043_ (.Y(_01582_),
    .B1(_01578_),
    .B2(_01579_),
    .A2(net1220),
    .A1(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ));
 sg13g2_a21o_1 _07044_ (.A2(_01576_),
    .A1(_01529_),
    .B1(_01569_),
    .X(_01583_));
 sg13g2_nor2_1 _07045_ (.A(_04812_),
    .B(_04823_),
    .Y(_01584_));
 sg13g2_nand3_1 _07046_ (.B(_01583_),
    .C(_01584_),
    .A(_01577_),
    .Y(_01585_));
 sg13g2_nor3_1 _07047_ (.A(_01580_),
    .B(_01582_),
    .C(_01585_),
    .Y(_01586_));
 sg13g2_or3_1 _07048_ (.A(_01580_),
    .B(_01582_),
    .C(_01585_),
    .X(_01587_));
 sg13g2_xor2_1 _07049_ (.B(_01531_),
    .A(_01530_),
    .X(_01588_));
 sg13g2_o21ai_1 _07050_ (.B1(_01585_),
    .Y(_01589_),
    .A1(_01580_),
    .A2(_01582_));
 sg13g2_nand3_1 _07051_ (.B(_01588_),
    .C(_01589_),
    .A(_01587_),
    .Y(_01590_));
 sg13g2_a21o_1 _07052_ (.A2(_01589_),
    .A1(_01588_),
    .B1(_01586_),
    .X(_01591_));
 sg13g2_o21ai_1 _07053_ (.B1(_01542_),
    .Y(_01592_),
    .A1(_01534_),
    .A2(_01543_));
 sg13g2_nand2b_1 _07054_ (.Y(_01593_),
    .B(_01567_),
    .A_N(_01565_));
 sg13g2_nor2b_1 _07055_ (.A(_01578_),
    .B_N(_01593_),
    .Y(_01594_));
 sg13g2_xnor2_1 _07056_ (.Y(_01595_),
    .A(_01578_),
    .B(_01593_));
 sg13g2_xor2_1 _07057_ (.B(_01595_),
    .A(_01592_),
    .X(_01596_));
 sg13g2_nor2_2 _07058_ (.A(_04806_),
    .B(_04832_),
    .Y(_01597_));
 sg13g2_nand2_1 _07059_ (.Y(_01598_),
    .A(net1406),
    .B(net1165));
 sg13g2_and3_1 _07060_ (.X(_01599_),
    .A(net1406),
    .B(net1165),
    .C(_01570_));
 sg13g2_xnor2_1 _07061_ (.Y(_01600_),
    .A(_01570_),
    .B(_01598_));
 sg13g2_xor2_1 _07062_ (.B(_01600_),
    .A(_01597_),
    .X(_01601_));
 sg13g2_nand2b_1 _07063_ (.Y(_01602_),
    .B(_01601_),
    .A_N(_01571_));
 sg13g2_xnor2_1 _07064_ (.Y(_01603_),
    .A(_01571_),
    .B(_01601_));
 sg13g2_o21ai_1 _07065_ (.B1(_01539_),
    .Y(_01604_),
    .A1(_01536_),
    .A2(_01540_));
 sg13g2_inv_1 _07066_ (.Y(_01605_),
    .A(_01604_));
 sg13g2_or2_1 _07067_ (.X(_01606_),
    .B(_01560_),
    .A(_01558_));
 sg13g2_nand2_1 _07068_ (.Y(_01607_),
    .A(net1453),
    .B(net1226));
 sg13g2_nand2_1 _07069_ (.Y(_01608_),
    .A(net1464),
    .B(net1213));
 sg13g2_nand2_1 _07070_ (.Y(_01609_),
    .A(net1464),
    .B(net1217));
 sg13g2_or2_1 _07071_ (.X(_01610_),
    .B(_01608_),
    .A(_01538_));
 sg13g2_xnor2_1 _07072_ (.Y(_01611_),
    .A(_01537_),
    .B(_01609_));
 sg13g2_xor2_1 _07073_ (.B(_01611_),
    .A(_01607_),
    .X(_01612_));
 sg13g2_nand2_1 _07074_ (.Y(_01613_),
    .A(_01606_),
    .B(_01612_));
 sg13g2_xnor2_1 _07075_ (.Y(_01614_),
    .A(_01606_),
    .B(_01612_));
 sg13g2_xnor2_1 _07076_ (.Y(_01615_),
    .A(_01605_),
    .B(_01614_));
 sg13g2_o21ai_1 _07077_ (.B1(_01554_),
    .Y(_01616_),
    .A1(_01555_),
    .A2(_01562_));
 sg13g2_nand2_1 _07078_ (.Y(_01617_),
    .A(net1473),
    .B(net1206));
 sg13g2_nand2_1 _07079_ (.Y(_01618_),
    .A(net1355),
    .B(net1204));
 sg13g2_or2_1 _07080_ (.X(_01619_),
    .B(_01618_),
    .A(_01557_));
 sg13g2_and2_1 _07081_ (.A(_01557_),
    .B(_01618_),
    .X(_01620_));
 sg13g2_xnor2_1 _07082_ (.Y(_01621_),
    .A(_01557_),
    .B(_01618_));
 sg13g2_xnor2_1 _07083_ (.Y(_01622_),
    .A(_01617_),
    .B(_01621_));
 sg13g2_o21ai_1 _07084_ (.B1(_01549_),
    .Y(_01623_),
    .A1(_01547_),
    .A2(_01550_));
 sg13g2_nand2_1 _07085_ (.Y(_01624_),
    .A(net1369),
    .B(net1192));
 sg13g2_and4_1 _07086_ (.A(net1383),
    .B(net1376),
    .C(net1185),
    .D(net1179),
    .X(_01625_));
 sg13g2_nand4_1 _07087_ (.B(net1376),
    .C(net1185),
    .A(net1383),
    .Y(_01626_),
    .D(net1179));
 sg13g2_a22oi_1 _07088_ (.Y(_01627_),
    .B1(net1179),
    .B2(net1383),
    .A2(net1185),
    .A1(net1376));
 sg13g2_or3_1 _07089_ (.A(_01624_),
    .B(_01625_),
    .C(_01627_),
    .X(_01628_));
 sg13g2_o21ai_1 _07090_ (.B1(_01624_),
    .Y(_01629_),
    .A1(_01625_),
    .A2(_01627_));
 sg13g2_and3_1 _07091_ (.X(_01630_),
    .A(_01623_),
    .B(_01628_),
    .C(_01629_));
 sg13g2_nand3_1 _07092_ (.B(_01628_),
    .C(_01629_),
    .A(_01623_),
    .Y(_01631_));
 sg13g2_a21oi_1 _07093_ (.A1(_01628_),
    .A2(_01629_),
    .Y(_01632_),
    .B1(_01623_));
 sg13g2_or3_1 _07094_ (.A(_01622_),
    .B(_01630_),
    .C(_01632_),
    .X(_01633_));
 sg13g2_o21ai_1 _07095_ (.B1(_01622_),
    .Y(_01634_),
    .A1(_01630_),
    .A2(_01632_));
 sg13g2_and3_1 _07096_ (.X(_01635_),
    .A(_01616_),
    .B(_01633_),
    .C(_01634_));
 sg13g2_a21oi_1 _07097_ (.A1(_01633_),
    .A2(_01634_),
    .Y(_01636_),
    .B1(_01616_));
 sg13g2_or3_1 _07098_ (.A(_01615_),
    .B(_01635_),
    .C(_01636_),
    .X(_01637_));
 sg13g2_o21ai_1 _07099_ (.B1(_01615_),
    .Y(_01638_),
    .A1(_01635_),
    .A2(_01636_));
 sg13g2_a21o_1 _07100_ (.A2(_01638_),
    .A1(_01637_),
    .B1(_01603_),
    .X(_01639_));
 sg13g2_and3_1 _07101_ (.X(_01640_),
    .A(_01603_),
    .B(_01637_),
    .C(_01638_));
 sg13g2_nand3_1 _07102_ (.B(_01637_),
    .C(_01638_),
    .A(_01603_),
    .Y(_01641_));
 sg13g2_nand3_1 _07103_ (.B(_01639_),
    .C(_01641_),
    .A(_01575_),
    .Y(_01642_));
 sg13g2_a21o_1 _07104_ (.A2(_01641_),
    .A1(_01639_),
    .B1(_01575_),
    .X(_01643_));
 sg13g2_and4_1 _07105_ (.A(net1458),
    .B(net1221),
    .C(_01642_),
    .D(_01643_),
    .X(_01644_));
 sg13g2_a22oi_1 _07106_ (.Y(_01645_),
    .B1(_01642_),
    .B2(_01643_),
    .A2(net1221),
    .A1(net1458));
 sg13g2_nor3_1 _07107_ (.A(_01581_),
    .B(_01644_),
    .C(_01645_),
    .Y(_01646_));
 sg13g2_or3_1 _07108_ (.A(_01581_),
    .B(_01644_),
    .C(_01645_),
    .X(_01647_));
 sg13g2_o21ai_1 _07109_ (.B1(_01581_),
    .Y(_01648_),
    .A1(_01644_),
    .A2(_01645_));
 sg13g2_nand3_1 _07110_ (.B(_01647_),
    .C(_01648_),
    .A(_01596_),
    .Y(_01649_));
 sg13g2_a21o_1 _07111_ (.A2(_01648_),
    .A1(_01647_),
    .B1(_01596_),
    .X(_01650_));
 sg13g2_and3_1 _07112_ (.X(_01651_),
    .A(_01591_),
    .B(_01649_),
    .C(_01650_));
 sg13g2_nand3_1 _07113_ (.B(_01649_),
    .C(_01650_),
    .A(_01591_),
    .Y(_01652_));
 sg13g2_a21oi_1 _07114_ (.A1(_01649_),
    .A2(_01650_),
    .Y(_01653_),
    .B1(_01591_));
 sg13g2_nor2_1 _07115_ (.A(_01651_),
    .B(_01653_),
    .Y(_01654_));
 sg13g2_xnor2_1 _07116_ (.Y(_01655_),
    .A(_01532_),
    .B(_01654_));
 sg13g2_a21o_1 _07117_ (.A2(_01583_),
    .A1(_01577_),
    .B1(_01584_),
    .X(_01656_));
 sg13g2_nand2_1 _07118_ (.Y(_01657_),
    .A(net1369),
    .B(net1217));
 sg13g2_nand2_1 _07119_ (.Y(_01658_),
    .A(net1369),
    .B(net1212));
 sg13g2_nand2_1 _07120_ (.Y(_01659_),
    .A(net1473),
    .B(net1226));
 sg13g2_xor2_1 _07121_ (.B(_01658_),
    .A(_01511_),
    .X(_01660_));
 sg13g2_nand2b_1 _07122_ (.Y(_01661_),
    .B(_01660_),
    .A_N(_01659_));
 sg13g2_o21ai_1 _07123_ (.B1(_01661_),
    .Y(_01662_),
    .A1(_01511_),
    .A2(_01658_));
 sg13g2_nand2_1 _07124_ (.Y(_01663_),
    .A(net1390),
    .B(net1199));
 sg13g2_or2_1 _07125_ (.X(_01664_),
    .B(_01663_),
    .A(_01484_));
 sg13g2_nand2_1 _07126_ (.Y(_01665_),
    .A(net1376),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ));
 sg13g2_xor2_1 _07127_ (.B(_01663_),
    .A(_01484_),
    .X(_01666_));
 sg13g2_nand2b_1 _07128_ (.Y(_01667_),
    .B(_01666_),
    .A_N(_01665_));
 sg13g2_and2_1 _07129_ (.A(_01664_),
    .B(_01667_),
    .X(_01668_));
 sg13g2_o21ai_1 _07130_ (.B1(_01513_),
    .Y(_01669_),
    .A1(_01512_),
    .A2(_01514_));
 sg13g2_nor2b_1 _07131_ (.A(_01515_),
    .B_N(_01669_),
    .Y(_01670_));
 sg13g2_nor2b_1 _07132_ (.A(_01668_),
    .B_N(_01670_),
    .Y(_01671_));
 sg13g2_xnor2_1 _07133_ (.Y(_01672_),
    .A(_01668_),
    .B(_01670_));
 sg13g2_xor2_1 _07134_ (.B(_01672_),
    .A(_01662_),
    .X(_01673_));
 sg13g2_xnor2_1 _07135_ (.Y(_01674_),
    .A(_01665_),
    .B(_01666_));
 sg13g2_a22oi_1 _07136_ (.Y(_01675_),
    .B1(net1187),
    .B2(net1406),
    .A2(net1194),
    .A1(net1398));
 sg13g2_nor2_1 _07137_ (.A(_01472_),
    .B(_01675_),
    .Y(_01676_));
 sg13g2_nand2_1 _07138_ (.Y(_01677_),
    .A(_01674_),
    .B(_01676_));
 sg13g2_xnor2_1 _07139_ (.Y(_01678_),
    .A(_01481_),
    .B(_01489_));
 sg13g2_nor2_1 _07140_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 sg13g2_xor2_1 _07141_ (.B(_01678_),
    .A(_01677_),
    .X(_01680_));
 sg13g2_xor2_1 _07142_ (.B(_01680_),
    .A(_01673_),
    .X(_01681_));
 sg13g2_nor2_1 _07143_ (.A(_04811_),
    .B(_04823_),
    .Y(_01682_));
 sg13g2_and4_1 _07144_ (.A(_01585_),
    .B(_01656_),
    .C(_01681_),
    .D(_01682_),
    .X(_01683_));
 sg13g2_a21oi_1 _07145_ (.A1(_01673_),
    .A2(_01680_),
    .Y(_01684_),
    .B1(_01679_));
 sg13g2_a21o_1 _07146_ (.A2(_01672_),
    .A1(_01662_),
    .B1(_01671_),
    .X(_01685_));
 sg13g2_nand2b_1 _07147_ (.Y(_01686_),
    .B(_01685_),
    .A_N(_01684_));
 sg13g2_xnor2_1 _07148_ (.Y(_01687_),
    .A(_01684_),
    .B(_01685_));
 sg13g2_inv_1 _07149_ (.Y(_01688_),
    .A(_01687_));
 sg13g2_a22oi_1 _07150_ (.Y(_01689_),
    .B1(_01681_),
    .B2(_01682_),
    .A2(_01656_),
    .A1(_01585_));
 sg13g2_or3_1 _07151_ (.A(_01683_),
    .B(_01688_),
    .C(_01689_),
    .X(_01690_));
 sg13g2_nand2b_1 _07152_ (.Y(_01691_),
    .B(_01690_),
    .A_N(_01683_));
 sg13g2_a21o_1 _07153_ (.A2(_01589_),
    .A1(_01587_),
    .B1(_01588_),
    .X(_01692_));
 sg13g2_and3_1 _07154_ (.X(_01693_),
    .A(_01590_),
    .B(_01691_),
    .C(_01692_));
 sg13g2_a21oi_1 _07155_ (.A1(_01590_),
    .A2(_01692_),
    .Y(_01694_),
    .B1(_01691_));
 sg13g2_or3_1 _07156_ (.A(_01686_),
    .B(_01693_),
    .C(_01694_),
    .X(_01695_));
 sg13g2_nand2b_2 _07157_ (.Y(_01696_),
    .B(_01695_),
    .A_N(_01693_));
 sg13g2_nand2_1 _07158_ (.Y(_01697_),
    .A(_01655_),
    .B(_01696_));
 sg13g2_xnor2_1 _07159_ (.Y(_01698_),
    .A(_01655_),
    .B(_01696_));
 sg13g2_xor2_1 _07160_ (.B(_01682_),
    .A(_01681_),
    .X(_01699_));
 sg13g2_nor2_1 _07161_ (.A(_04807_),
    .B(_04826_),
    .Y(_01700_));
 sg13g2_nand2_2 _07162_ (.Y(_01701_),
    .A(net1399),
    .B(net1201));
 sg13g2_and4_1 _07163_ (.A(net1398),
    .B(net1390),
    .C(net1201),
    .D(net1197),
    .X(_01702_));
 sg13g2_a22oi_1 _07164_ (.Y(_01703_),
    .B1(net1197),
    .B2(net1398),
    .A2(net1201),
    .A1(net1390));
 sg13g2_nor2_1 _07165_ (.A(_01702_),
    .B(_01703_),
    .Y(_01704_));
 sg13g2_xor2_1 _07166_ (.B(_01704_),
    .A(_01700_),
    .X(_01705_));
 sg13g2_nand2b_1 _07167_ (.Y(_01706_),
    .B(_01705_),
    .A_N(_01471_));
 sg13g2_xor2_1 _07168_ (.B(_01676_),
    .A(_01674_),
    .X(_01707_));
 sg13g2_nor2b_1 _07169_ (.A(_01706_),
    .B_N(_01707_),
    .Y(_01708_));
 sg13g2_xnor2_1 _07170_ (.Y(_01709_),
    .A(_01706_),
    .B(_01707_));
 sg13g2_nand2_1 _07171_ (.Y(_01710_),
    .A(net1376),
    .B(net1210));
 sg13g2_nand2_1 _07172_ (.Y(_01711_),
    .A(net1355),
    .B(net1225));
 sg13g2_xor2_1 _07173_ (.B(_01710_),
    .A(_01657_),
    .X(_01712_));
 sg13g2_nand2b_1 _07174_ (.Y(_01713_),
    .B(_01712_),
    .A_N(_01711_));
 sg13g2_o21ai_1 _07175_ (.B1(_01713_),
    .Y(_01714_),
    .A1(_01657_),
    .A2(_01710_));
 sg13g2_a21oi_1 _07176_ (.A1(_01700_),
    .A2(_01704_),
    .Y(_01715_),
    .B1(_01702_));
 sg13g2_xnor2_1 _07177_ (.Y(_01716_),
    .A(_01659_),
    .B(_01660_));
 sg13g2_nor2b_1 _07178_ (.A(_01715_),
    .B_N(_01716_),
    .Y(_01717_));
 sg13g2_xnor2_1 _07179_ (.Y(_01718_),
    .A(_01715_),
    .B(_01716_));
 sg13g2_xnor2_1 _07180_ (.Y(_01719_),
    .A(_01714_),
    .B(_01718_));
 sg13g2_inv_1 _07181_ (.Y(_01720_),
    .A(_01719_));
 sg13g2_xnor2_1 _07182_ (.Y(_01721_),
    .A(_01709_),
    .B(_01719_));
 sg13g2_nand2_1 _07183_ (.Y(_01722_),
    .A(net1355),
    .B(net1221));
 sg13g2_and3_1 _07184_ (.X(_01723_),
    .A(net1355),
    .B(net1221),
    .C(_01721_));
 sg13g2_and2_1 _07185_ (.A(_01699_),
    .B(_01723_),
    .X(_01724_));
 sg13g2_a21oi_1 _07186_ (.A1(_01709_),
    .A2(_01720_),
    .Y(_01725_),
    .B1(_01708_));
 sg13g2_a21o_1 _07187_ (.A2(_01718_),
    .A1(_01714_),
    .B1(_01717_),
    .X(_01726_));
 sg13g2_nor2b_1 _07188_ (.A(_01725_),
    .B_N(_01726_),
    .Y(_01727_));
 sg13g2_xnor2_1 _07189_ (.Y(_01728_),
    .A(_01725_),
    .B(_01726_));
 sg13g2_xor2_1 _07190_ (.B(_01723_),
    .A(_01699_),
    .X(_01729_));
 sg13g2_a21o_1 _07191_ (.A2(_01729_),
    .A1(_01728_),
    .B1(_01724_),
    .X(_01730_));
 sg13g2_o21ai_1 _07192_ (.B1(_01688_),
    .Y(_01731_),
    .A1(_01683_),
    .A2(_01689_));
 sg13g2_nand3_1 _07193_ (.B(_01730_),
    .C(_01731_),
    .A(_01690_),
    .Y(_01732_));
 sg13g2_a21o_1 _07194_ (.A2(_01731_),
    .A1(_01690_),
    .B1(_01730_),
    .X(_01733_));
 sg13g2_nand3_1 _07195_ (.B(_01732_),
    .C(_01733_),
    .A(_01727_),
    .Y(_01734_));
 sg13g2_nand2_1 _07196_ (.Y(_01735_),
    .A(_01732_),
    .B(_01734_));
 sg13g2_o21ai_1 _07197_ (.B1(_01686_),
    .Y(_01736_),
    .A1(_01693_),
    .A2(_01694_));
 sg13g2_a21o_1 _07198_ (.A2(_01736_),
    .A1(_01695_),
    .B1(_01735_),
    .X(_01737_));
 sg13g2_and3_1 _07199_ (.X(_01738_),
    .A(_01695_),
    .B(_01735_),
    .C(_01736_));
 sg13g2_xor2_1 _07200_ (.B(_01722_),
    .A(_01721_),
    .X(_01739_));
 sg13g2_xnor2_1 _07201_ (.Y(_01740_),
    .A(_01471_),
    .B(_01705_));
 sg13g2_and4_1 _07202_ (.A(net1380),
    .B(net1374),
    .C(net1216),
    .D(net1210),
    .X(_01741_));
 sg13g2_nand2_1 _07203_ (.Y(_01742_),
    .A(net1360),
    .B(net1224));
 sg13g2_a22oi_1 _07204_ (.Y(_01743_),
    .B1(net1210),
    .B2(net1381),
    .A2(net1216),
    .A1(net1374));
 sg13g2_or3_1 _07205_ (.A(_01741_),
    .B(_01742_),
    .C(_01743_),
    .X(_01744_));
 sg13g2_nand2b_1 _07206_ (.Y(_01745_),
    .B(_01744_),
    .A_N(_01741_));
 sg13g2_nand2_1 _07207_ (.Y(_01746_),
    .A(net1403),
    .B(net1197));
 sg13g2_or2_1 _07208_ (.X(_01747_),
    .B(_01746_),
    .A(_01701_));
 sg13g2_nand2_1 _07209_ (.Y(_01748_),
    .A(net1387),
    .B(net1205));
 sg13g2_and2_1 _07210_ (.A(_01701_),
    .B(_01746_),
    .X(_01749_));
 sg13g2_xor2_1 _07211_ (.B(_01746_),
    .A(_01701_),
    .X(_01750_));
 sg13g2_o21ai_1 _07212_ (.B1(_01747_),
    .Y(_01751_),
    .A1(_01748_),
    .A2(_01749_));
 sg13g2_xnor2_1 _07213_ (.Y(_01752_),
    .A(_01711_),
    .B(_01712_));
 sg13g2_and2_1 _07214_ (.A(_01751_),
    .B(_01752_),
    .X(_01753_));
 sg13g2_xor2_1 _07215_ (.B(_01752_),
    .A(_01751_),
    .X(_01754_));
 sg13g2_xor2_1 _07216_ (.B(_01754_),
    .A(_01745_),
    .X(_01755_));
 sg13g2_nand2_1 _07217_ (.Y(_01756_),
    .A(_01740_),
    .B(_01755_));
 sg13g2_xnor2_1 _07218_ (.Y(_01757_),
    .A(_01740_),
    .B(_01755_));
 sg13g2_nand2_1 _07219_ (.Y(_01758_),
    .A(net1362),
    .B(net1220));
 sg13g2_nor2_1 _07220_ (.A(_01757_),
    .B(_01758_),
    .Y(_01759_));
 sg13g2_nand2b_1 _07221_ (.Y(_01760_),
    .B(_01759_),
    .A_N(_01739_));
 sg13g2_a21oi_1 _07222_ (.A1(_01745_),
    .A2(_01754_),
    .Y(_01761_),
    .B1(_01753_));
 sg13g2_or2_1 _07223_ (.X(_01762_),
    .B(_01761_),
    .A(_01756_));
 sg13g2_xnor2_1 _07224_ (.Y(_01763_),
    .A(_01756_),
    .B(_01761_));
 sg13g2_xnor2_1 _07225_ (.Y(_01764_),
    .A(_01739_),
    .B(_01759_));
 sg13g2_nand2b_1 _07226_ (.Y(_01765_),
    .B(_01764_),
    .A_N(_01763_));
 sg13g2_nand2_1 _07227_ (.Y(_01766_),
    .A(_01760_),
    .B(_01765_));
 sg13g2_xnor2_1 _07228_ (.Y(_01767_),
    .A(_01728_),
    .B(_01729_));
 sg13g2_nand2b_1 _07229_ (.Y(_01768_),
    .B(_01766_),
    .A_N(_01767_));
 sg13g2_xor2_1 _07230_ (.B(_01767_),
    .A(_01766_),
    .X(_01769_));
 sg13g2_o21ai_1 _07231_ (.B1(_01768_),
    .Y(_01770_),
    .A1(_01762_),
    .A2(_01769_));
 sg13g2_a21o_1 _07232_ (.A2(_01733_),
    .A1(_01732_),
    .B1(_01727_),
    .X(_01771_));
 sg13g2_a21oi_1 _07233_ (.A1(_01734_),
    .A2(_01771_),
    .Y(_01772_),
    .B1(_01770_));
 sg13g2_nand3_1 _07234_ (.B(_01770_),
    .C(_01771_),
    .A(_01734_),
    .Y(_01773_));
 sg13g2_xnor2_1 _07235_ (.Y(_01774_),
    .A(_01748_),
    .B(_01750_));
 sg13g2_and4_1 _07236_ (.A(net1389),
    .B(net1382),
    .C(net1216),
    .D(net1210),
    .X(_01775_));
 sg13g2_nand2_1 _07237_ (.Y(_01776_),
    .A(net1368),
    .B(net1224));
 sg13g2_a22oi_1 _07238_ (.Y(_01777_),
    .B1(net1210),
    .B2(net1389),
    .A2(net1216),
    .A1(net1382));
 sg13g2_or3_1 _07239_ (.A(_01775_),
    .B(_01776_),
    .C(_01777_),
    .X(_01778_));
 sg13g2_nand2b_1 _07240_ (.Y(_01779_),
    .B(_01778_),
    .A_N(_01775_));
 sg13g2_nor3_1 _07241_ (.A(_04804_),
    .B(_04826_),
    .C(_01701_),
    .Y(_01780_));
 sg13g2_o21ai_1 _07242_ (.B1(_01742_),
    .Y(_01781_),
    .A1(_01741_),
    .A2(_01743_));
 sg13g2_nand3_1 _07243_ (.B(_01780_),
    .C(_01781_),
    .A(_01744_),
    .Y(_01782_));
 sg13g2_a21o_1 _07244_ (.A2(_01781_),
    .A1(_01744_),
    .B1(_01780_),
    .X(_01783_));
 sg13g2_nand3_1 _07245_ (.B(_01782_),
    .C(_01783_),
    .A(_01779_),
    .Y(_01784_));
 sg13g2_a21o_1 _07246_ (.A2(_01783_),
    .A1(_01782_),
    .B1(_01779_),
    .X(_01785_));
 sg13g2_and3_1 _07247_ (.X(_01786_),
    .A(_01774_),
    .B(_01784_),
    .C(_01785_));
 sg13g2_nand3_1 _07248_ (.B(_01784_),
    .C(_01785_),
    .A(_01774_),
    .Y(_01787_));
 sg13g2_nand2_1 _07249_ (.Y(_01788_),
    .A(_01782_),
    .B(_01784_));
 sg13g2_nand2_1 _07250_ (.Y(_01789_),
    .A(_01786_),
    .B(_01788_));
 sg13g2_a21o_1 _07251_ (.A2(_01785_),
    .A1(_01784_),
    .B1(_01774_),
    .X(_01790_));
 sg13g2_and4_1 _07252_ (.A(net1366),
    .B(net1220),
    .C(_01787_),
    .D(_01790_),
    .X(_01791_));
 sg13g2_xor2_1 _07253_ (.B(_01758_),
    .A(_01757_),
    .X(_01792_));
 sg13g2_nand2_1 _07254_ (.Y(_01793_),
    .A(_01791_),
    .B(_01792_));
 sg13g2_xnor2_1 _07255_ (.Y(_01794_),
    .A(_01786_),
    .B(_01788_));
 sg13g2_xnor2_1 _07256_ (.Y(_01795_),
    .A(_01791_),
    .B(_01792_));
 sg13g2_o21ai_1 _07257_ (.B1(_01793_),
    .Y(_01796_),
    .A1(_01794_),
    .A2(_01795_));
 sg13g2_xnor2_1 _07258_ (.Y(_01797_),
    .A(_01763_),
    .B(_01764_));
 sg13g2_xnor2_1 _07259_ (.Y(_01798_),
    .A(_01796_),
    .B(_01797_));
 sg13g2_nor2_1 _07260_ (.A(_01789_),
    .B(_01798_),
    .Y(_01799_));
 sg13g2_xnor2_1 _07261_ (.Y(_01800_),
    .A(_01794_),
    .B(_01795_));
 sg13g2_a22oi_1 _07262_ (.Y(_01801_),
    .B1(_01787_),
    .B2(_01790_),
    .A2(net1220),
    .A1(net1367));
 sg13g2_nor2_1 _07263_ (.A(_04808_),
    .B(_04823_),
    .Y(_01802_));
 sg13g2_a22oi_1 _07264_ (.Y(_01803_),
    .B1(net1201),
    .B2(net1403),
    .A2(net1205),
    .A1(net1399));
 sg13g2_nor2_1 _07265_ (.A(_01780_),
    .B(_01803_),
    .Y(_01804_));
 sg13g2_and4_1 _07266_ (.A(net1400),
    .B(net1389),
    .C(net1214),
    .D(net1209),
    .X(_01805_));
 sg13g2_nand4_1 _07267_ (.B(net1389),
    .C(net1214),
    .A(net1400),
    .Y(_01806_),
    .D(net1209));
 sg13g2_nand2_1 _07268_ (.Y(_01807_),
    .A(net1375),
    .B(net1224));
 sg13g2_a22oi_1 _07269_ (.Y(_01808_),
    .B1(net1209),
    .B2(net1400),
    .A2(net1214),
    .A1(net1389));
 sg13g2_or3_1 _07270_ (.A(_01805_),
    .B(_01807_),
    .C(_01808_),
    .X(_01809_));
 sg13g2_o21ai_1 _07271_ (.B1(_01806_),
    .Y(_01810_),
    .A1(_01807_),
    .A2(_01808_));
 sg13g2_o21ai_1 _07272_ (.B1(_01776_),
    .Y(_01811_),
    .A1(_01775_),
    .A2(_01777_));
 sg13g2_nand3_1 _07273_ (.B(_01810_),
    .C(_01811_),
    .A(_01778_),
    .Y(_01812_));
 sg13g2_a21o_1 _07274_ (.A2(_01811_),
    .A1(_01778_),
    .B1(_01810_),
    .X(_01813_));
 sg13g2_nand3_1 _07275_ (.B(_01812_),
    .C(_01813_),
    .A(_01804_),
    .Y(_01814_));
 sg13g2_a21o_1 _07276_ (.A2(_01813_),
    .A1(_01812_),
    .B1(_01804_),
    .X(_01815_));
 sg13g2_nand3_1 _07277_ (.B(_01814_),
    .C(_01815_),
    .A(_01802_),
    .Y(_01816_));
 sg13g2_nor3_1 _07278_ (.A(_01791_),
    .B(_01801_),
    .C(_01816_),
    .Y(_01817_));
 sg13g2_nand2_1 _07279_ (.Y(_01818_),
    .A(_01812_),
    .B(_01814_));
 sg13g2_o21ai_1 _07280_ (.B1(_01816_),
    .Y(_01819_),
    .A1(_01791_),
    .A2(_01801_));
 sg13g2_nor2b_1 _07281_ (.A(_01817_),
    .B_N(_01819_),
    .Y(_01820_));
 sg13g2_a21oi_1 _07282_ (.A1(_01818_),
    .A2(_01819_),
    .Y(_01821_),
    .B1(_01817_));
 sg13g2_nand2_1 _07283_ (.Y(_01822_),
    .A(_01800_),
    .B(_01821_));
 sg13g2_xor2_1 _07284_ (.B(_01820_),
    .A(_01818_),
    .X(_01823_));
 sg13g2_and4_1 _07285_ (.A(net1403),
    .B(net1400),
    .C(net1214),
    .D(net1208),
    .X(_01824_));
 sg13g2_nand4_1 _07286_ (.B(net1400),
    .C(net1214),
    .A(net1403),
    .Y(_01825_),
    .D(net1208));
 sg13g2_nand2_1 _07287_ (.Y(_01826_),
    .A(net1382),
    .B(net1227));
 sg13g2_a22oi_1 _07288_ (.Y(_01827_),
    .B1(net1209),
    .B2(net1403),
    .A2(net1215),
    .A1(net1400));
 sg13g2_nor2_1 _07289_ (.A(_01824_),
    .B(_01827_),
    .Y(_01828_));
 sg13g2_o21ai_1 _07290_ (.B1(_01825_),
    .Y(_01829_),
    .A1(_01826_),
    .A2(_01827_));
 sg13g2_o21ai_1 _07291_ (.B1(_01807_),
    .Y(_01830_),
    .A1(_01805_),
    .A2(_01808_));
 sg13g2_and2_1 _07292_ (.A(_01809_),
    .B(_01830_),
    .X(_01831_));
 sg13g2_nand3_1 _07293_ (.B(_01829_),
    .C(_01830_),
    .A(_01809_),
    .Y(_01832_));
 sg13g2_a21o_1 _07294_ (.A2(_01830_),
    .A1(_01809_),
    .B1(_01829_),
    .X(_01833_));
 sg13g2_and4_1 _07295_ (.A(net1403),
    .B(net1207),
    .C(_01832_),
    .D(_01833_),
    .X(_01834_));
 sg13g2_a21oi_1 _07296_ (.A1(_01829_),
    .A2(_01831_),
    .Y(_01835_),
    .B1(_01834_));
 sg13g2_a22oi_1 _07297_ (.Y(_01836_),
    .B1(_01832_),
    .B2(_01833_),
    .A2(net1207),
    .A1(net1403));
 sg13g2_nand2_1 _07298_ (.Y(_01837_),
    .A(net1382),
    .B(net1219));
 sg13g2_nor3_1 _07299_ (.A(_01834_),
    .B(_01836_),
    .C(_01837_),
    .Y(_01838_));
 sg13g2_a21o_1 _07300_ (.A2(_01815_),
    .A1(_01814_),
    .B1(_01802_),
    .X(_01839_));
 sg13g2_and3_1 _07301_ (.X(_01840_),
    .A(_01816_),
    .B(_01838_),
    .C(_01839_));
 sg13g2_a21oi_1 _07302_ (.A1(_01816_),
    .A2(_01839_),
    .Y(_01841_),
    .B1(_01838_));
 sg13g2_or3_1 _07303_ (.A(_01835_),
    .B(_01840_),
    .C(_01841_),
    .X(_01842_));
 sg13g2_o21ai_1 _07304_ (.B1(_01835_),
    .Y(_01843_),
    .A1(_01840_),
    .A2(_01841_));
 sg13g2_xor2_1 _07305_ (.B(_01828_),
    .A(_01826_),
    .X(_01844_));
 sg13g2_nand2_1 _07306_ (.Y(_01845_),
    .A(net1406),
    .B(net1224));
 sg13g2_nor3_1 _07307_ (.A(_04806_),
    .B(_04824_),
    .C(_01845_),
    .Y(_01846_));
 sg13g2_nor2b_1 _07308_ (.A(_01844_),
    .B_N(_01846_),
    .Y(_01847_));
 sg13g2_o21ai_1 _07309_ (.B1(_01837_),
    .Y(_01848_),
    .A1(_01834_),
    .A2(_01836_));
 sg13g2_nand2b_1 _07310_ (.Y(_01849_),
    .B(_01848_),
    .A_N(_01838_));
 sg13g2_xnor2_1 _07311_ (.Y(_01850_),
    .A(_01844_),
    .B(_01846_));
 sg13g2_nand3_1 _07312_ (.B(net1220),
    .C(_01850_),
    .A(net1389),
    .Y(_01851_));
 sg13g2_o21ai_1 _07313_ (.B1(_01844_),
    .Y(_01852_),
    .A1(_04806_),
    .A2(_04823_));
 sg13g2_a22oi_1 _07314_ (.Y(_01853_),
    .B1(net1214),
    .B2(net1406),
    .A2(net1224),
    .A1(net1392));
 sg13g2_nor2_1 _07315_ (.A(_01846_),
    .B(_01853_),
    .Y(_01854_));
 sg13g2_nand3_1 _07316_ (.B(_01852_),
    .C(_01854_),
    .A(_01851_),
    .Y(_01855_));
 sg13g2_or3_1 _07317_ (.A(_01844_),
    .B(_01845_),
    .C(_01854_),
    .X(_01856_));
 sg13g2_nand2_1 _07318_ (.Y(_01857_),
    .A(net1400),
    .B(net1220));
 sg13g2_a21oi_1 _07319_ (.A1(_01855_),
    .A2(_01856_),
    .Y(_01858_),
    .B1(_01857_));
 sg13g2_xnor2_1 _07320_ (.Y(_01859_),
    .A(_01847_),
    .B(_01849_));
 sg13g2_nand4_1 _07321_ (.B(_01843_),
    .C(_01858_),
    .A(_01842_),
    .Y(_01860_),
    .D(_01859_));
 sg13g2_nor2b_1 _07322_ (.A(_01840_),
    .B_N(_01842_),
    .Y(_01861_));
 sg13g2_nor2_1 _07323_ (.A(_01860_),
    .B(_01861_),
    .Y(_01862_));
 sg13g2_nor2b_1 _07324_ (.A(_01847_),
    .B_N(_01851_),
    .Y(_01863_));
 sg13g2_nor2_1 _07325_ (.A(_01849_),
    .B(_01863_),
    .Y(_01864_));
 sg13g2_nand3_1 _07326_ (.B(_01843_),
    .C(_01864_),
    .A(_01842_),
    .Y(_01865_));
 sg13g2_nand3_1 _07327_ (.B(_01861_),
    .C(_01865_),
    .A(_01860_),
    .Y(_01866_));
 sg13g2_o21ai_1 _07328_ (.B1(_01866_),
    .Y(_01867_),
    .A1(_01823_),
    .A2(_01862_));
 sg13g2_or2_1 _07329_ (.X(_01868_),
    .B(_01821_),
    .A(_01800_));
 sg13g2_a22oi_1 _07330_ (.Y(_01869_),
    .B1(_01867_),
    .B2(_01868_),
    .A2(_01798_),
    .A1(_01789_));
 sg13g2_a221oi_1 _07331_ (.B2(_01869_),
    .C1(_01799_),
    .B1(_01822_),
    .A1(_01796_),
    .Y(_01870_),
    .A2(_01797_));
 sg13g2_xor2_1 _07332_ (.B(_01769_),
    .A(_01762_),
    .X(_01871_));
 sg13g2_nand2b_1 _07333_ (.Y(_01872_),
    .B(_01871_),
    .A_N(_01870_));
 sg13g2_a21oi_1 _07334_ (.A1(_01773_),
    .A2(_01872_),
    .Y(_01873_),
    .B1(_01772_));
 sg13g2_o21ai_1 _07335_ (.B1(_01737_),
    .Y(_01874_),
    .A1(_01738_),
    .A2(_01873_));
 sg13g2_xor2_1 _07336_ (.B(_01874_),
    .A(_01698_),
    .X(_01875_));
 sg13g2_o21ai_1 _07337_ (.B1(net1517),
    .Y(_01876_),
    .A1(net1143),
    .A2(_01875_));
 sg13g2_a21oi_1 _07338_ (.A1(net1143),
    .A2(_04781_),
    .Y(_00224_),
    .B1(_01876_));
 sg13g2_a21oi_1 _07339_ (.A1(_01592_),
    .A2(_01595_),
    .Y(_01877_),
    .B1(_01594_));
 sg13g2_a21o_1 _07340_ (.A2(_01648_),
    .A1(_01596_),
    .B1(_01646_),
    .X(_01878_));
 sg13g2_o21ai_1 _07341_ (.B1(_01613_),
    .Y(_01879_),
    .A1(_01605_),
    .A2(_01614_));
 sg13g2_nand2b_1 _07342_ (.Y(_01880_),
    .B(_01637_),
    .A_N(_01635_));
 sg13g2_nor2b_1 _07343_ (.A(_01642_),
    .B_N(_01880_),
    .Y(_01881_));
 sg13g2_xnor2_1 _07344_ (.Y(_01882_),
    .A(_01642_),
    .B(_01880_));
 sg13g2_xor2_1 _07345_ (.B(_01882_),
    .A(_01879_),
    .X(_01883_));
 sg13g2_nand2_1 _07346_ (.Y(_01884_),
    .A(net1454),
    .B(net1221));
 sg13g2_nand2_2 _07347_ (.Y(_01885_),
    .A(net1403),
    .B(net1159));
 sg13g2_or2_1 _07348_ (.X(_01886_),
    .B(_01885_),
    .A(_01884_));
 sg13g2_xnor2_1 _07349_ (.Y(_01887_),
    .A(_01884_),
    .B(_01885_));
 sg13g2_o21ai_1 _07350_ (.B1(_01610_),
    .Y(_01888_),
    .A1(_01607_),
    .A2(_01611_));
 sg13g2_inv_1 _07351_ (.Y(_01889_),
    .A(_01888_));
 sg13g2_o21ai_1 _07352_ (.B1(_01619_),
    .Y(_01890_),
    .A1(_01617_),
    .A2(_01620_));
 sg13g2_nand2_1 _07353_ (.Y(_01891_),
    .A(net1449),
    .B(net1226));
 sg13g2_nand2_1 _07354_ (.Y(_01892_),
    .A(net1458),
    .B(net1211));
 sg13g2_nand2_1 _07355_ (.Y(_01893_),
    .A(net1459),
    .B(net1217));
 sg13g2_or2_1 _07356_ (.X(_01894_),
    .B(_01892_),
    .A(_01609_));
 sg13g2_xnor2_1 _07357_ (.Y(_01895_),
    .A(_01608_),
    .B(_01893_));
 sg13g2_xor2_1 _07358_ (.B(_01895_),
    .A(_01891_),
    .X(_01896_));
 sg13g2_nand2_1 _07359_ (.Y(_01897_),
    .A(_01890_),
    .B(_01896_));
 sg13g2_xnor2_1 _07360_ (.Y(_01898_),
    .A(_01890_),
    .B(_01896_));
 sg13g2_xnor2_1 _07361_ (.Y(_01899_),
    .A(_01888_),
    .B(_01898_));
 sg13g2_xnor2_1 _07362_ (.Y(_01900_),
    .A(_01889_),
    .B(_01898_));
 sg13g2_o21ai_1 _07363_ (.B1(_01631_),
    .Y(_01901_),
    .A1(_01622_),
    .A2(_01632_));
 sg13g2_nand2_1 _07364_ (.Y(_01902_),
    .A(net1469),
    .B(net1206));
 sg13g2_nand2_1 _07365_ (.Y(_01903_),
    .A(net1473),
    .B(net1196));
 sg13g2_and4_1 _07366_ (.A(net1355),
    .B(net1473),
    .C(net1201),
    .D(net1196),
    .X(_01904_));
 sg13g2_a22oi_1 _07367_ (.Y(_01905_),
    .B1(net1197),
    .B2(net1355),
    .A2(net1202),
    .A1(net1473));
 sg13g2_nor3_1 _07368_ (.A(_01902_),
    .B(_01904_),
    .C(_01905_),
    .Y(_01906_));
 sg13g2_o21ai_1 _07369_ (.B1(_01902_),
    .Y(_01907_),
    .A1(_01904_),
    .A2(_01905_));
 sg13g2_nand2b_1 _07370_ (.Y(_01908_),
    .B(_01907_),
    .A_N(_01906_));
 sg13g2_o21ai_1 _07371_ (.B1(_01626_),
    .Y(_01909_),
    .A1(_01624_),
    .A2(_01627_));
 sg13g2_nand2_1 _07372_ (.Y(_01910_),
    .A(net1362),
    .B(net1192));
 sg13g2_and4_1 _07373_ (.A(net1376),
    .B(net1369),
    .C(net1185),
    .D(net1180),
    .X(_01911_));
 sg13g2_nand4_1 _07374_ (.B(net1369),
    .C(net1185),
    .A(net1377),
    .Y(_01912_),
    .D(net1180));
 sg13g2_a22oi_1 _07375_ (.Y(_01913_),
    .B1(net1180),
    .B2(net1377),
    .A2(net1185),
    .A1(net1369));
 sg13g2_or3_1 _07376_ (.A(_01910_),
    .B(_01911_),
    .C(_01913_),
    .X(_01914_));
 sg13g2_o21ai_1 _07377_ (.B1(_01910_),
    .Y(_01915_),
    .A1(_01911_),
    .A2(_01913_));
 sg13g2_and3_1 _07378_ (.X(_01916_),
    .A(_01909_),
    .B(_01914_),
    .C(_01915_));
 sg13g2_nand3_1 _07379_ (.B(_01914_),
    .C(_01915_),
    .A(_01909_),
    .Y(_01917_));
 sg13g2_a21oi_1 _07380_ (.A1(_01914_),
    .A2(_01915_),
    .Y(_01918_),
    .B1(_01909_));
 sg13g2_or3_1 _07381_ (.A(_01908_),
    .B(_01916_),
    .C(_01918_),
    .X(_01919_));
 sg13g2_o21ai_1 _07382_ (.B1(_01908_),
    .Y(_01920_),
    .A1(_01916_),
    .A2(_01918_));
 sg13g2_nand3_1 _07383_ (.B(_01919_),
    .C(_01920_),
    .A(_01901_),
    .Y(_01921_));
 sg13g2_a21oi_1 _07384_ (.A1(_01919_),
    .A2(_01920_),
    .Y(_01922_),
    .B1(_01901_));
 sg13g2_a21o_1 _07385_ (.A2(_01920_),
    .A1(_01919_),
    .B1(_01901_),
    .X(_01923_));
 sg13g2_and3_1 _07386_ (.X(_01924_),
    .A(_01899_),
    .B(_01921_),
    .C(_01923_));
 sg13g2_a21oi_1 _07387_ (.A1(_01921_),
    .A2(_01923_),
    .Y(_01925_),
    .B1(_01899_));
 sg13g2_nand2_1 _07388_ (.Y(_01926_),
    .A(net1383),
    .B(net1176));
 sg13g2_nand2_1 _07389_ (.Y(_01927_),
    .A(net1388),
    .B(net1165));
 sg13g2_and4_1 _07390_ (.A(net1399),
    .B(net1390),
    .C(net1172),
    .D(net1165),
    .X(_01928_));
 sg13g2_a22oi_1 _07391_ (.Y(_01929_),
    .B1(net1165),
    .B2(net1399),
    .A2(net1172),
    .A1(net1390));
 sg13g2_nor3_1 _07392_ (.A(_01926_),
    .B(_01928_),
    .C(_01929_),
    .Y(_01930_));
 sg13g2_o21ai_1 _07393_ (.B1(_01926_),
    .Y(_01931_),
    .A1(_01928_),
    .A2(_01929_));
 sg13g2_nor2b_1 _07394_ (.A(_01930_),
    .B_N(_01931_),
    .Y(_01932_));
 sg13g2_a21oi_1 _07395_ (.A1(_01597_),
    .A2(_01600_),
    .Y(_01933_),
    .B1(_01599_));
 sg13g2_nand2b_1 _07396_ (.Y(_01934_),
    .B(_01932_),
    .A_N(_01933_));
 sg13g2_xnor2_1 _07397_ (.Y(_01935_),
    .A(_01932_),
    .B(_01933_));
 sg13g2_nor2b_1 _07398_ (.A(_01602_),
    .B_N(_01935_),
    .Y(_01936_));
 sg13g2_xor2_1 _07399_ (.B(_01935_),
    .A(_01602_),
    .X(_01937_));
 sg13g2_o21ai_1 _07400_ (.B1(_01937_),
    .Y(_01938_),
    .A1(_01924_),
    .A2(_01925_));
 sg13g2_or3_1 _07401_ (.A(_01924_),
    .B(_01925_),
    .C(_01937_),
    .X(_01939_));
 sg13g2_and3_2 _07402_ (.X(_01940_),
    .A(_01640_),
    .B(_01938_),
    .C(_01939_));
 sg13g2_a21oi_1 _07403_ (.A1(_01938_),
    .A2(_01939_),
    .Y(_01941_),
    .B1(_01640_));
 sg13g2_or3_1 _07404_ (.A(_01887_),
    .B(_01940_),
    .C(_01941_),
    .X(_01942_));
 sg13g2_o21ai_1 _07405_ (.B1(_01887_),
    .Y(_01943_),
    .A1(_01940_),
    .A2(_01941_));
 sg13g2_nand3_1 _07406_ (.B(_01942_),
    .C(_01943_),
    .A(_01644_),
    .Y(_01944_));
 sg13g2_a21o_1 _07407_ (.A2(_01943_),
    .A1(_01942_),
    .B1(_01644_),
    .X(_01945_));
 sg13g2_nand3_1 _07408_ (.B(_01944_),
    .C(_01945_),
    .A(_01883_),
    .Y(_01946_));
 sg13g2_a21o_1 _07409_ (.A2(_01945_),
    .A1(_01944_),
    .B1(_01883_),
    .X(_01947_));
 sg13g2_and3_1 _07410_ (.X(_01948_),
    .A(_01878_),
    .B(_01946_),
    .C(_01947_));
 sg13g2_a21oi_1 _07411_ (.A1(_01946_),
    .A2(_01947_),
    .Y(_01949_),
    .B1(_01878_));
 sg13g2_or3_1 _07412_ (.A(_01877_),
    .B(_01948_),
    .C(_01949_),
    .X(_01950_));
 sg13g2_o21ai_1 _07413_ (.B1(_01877_),
    .Y(_01951_),
    .A1(_01948_),
    .A2(_01949_));
 sg13g2_and2_1 _07414_ (.A(_01950_),
    .B(_01951_),
    .X(_01952_));
 sg13g2_o21ai_1 _07415_ (.B1(_01652_),
    .Y(_01953_),
    .A1(_01532_),
    .A2(_01653_));
 sg13g2_or2_1 _07416_ (.X(_01954_),
    .B(_01953_),
    .A(_01952_));
 sg13g2_and3_1 _07417_ (.X(_01955_),
    .A(_01950_),
    .B(_01951_),
    .C(_01953_));
 sg13g2_xnor2_1 _07418_ (.Y(_01956_),
    .A(_01952_),
    .B(_01953_));
 sg13g2_o21ai_1 _07419_ (.B1(_01697_),
    .Y(_01957_),
    .A1(_01698_),
    .A2(_01874_));
 sg13g2_xor2_1 _07420_ (.B(_01957_),
    .A(_01956_),
    .X(_01958_));
 sg13g2_o21ai_1 _07421_ (.B1(net1517),
    .Y(_01959_),
    .A1(net1298),
    .A2(net283));
 sg13g2_a21oi_1 _07422_ (.A1(net1298),
    .A2(_01958_),
    .Y(_00225_),
    .B1(_01959_));
 sg13g2_nand2b_1 _07423_ (.Y(_01960_),
    .B(_01950_),
    .A_N(_01948_));
 sg13g2_a21oi_1 _07424_ (.A1(_01879_),
    .A2(_01882_),
    .Y(_01961_),
    .B1(_01881_));
 sg13g2_nand2_1 _07425_ (.Y(_01962_),
    .A(_01944_),
    .B(_01946_));
 sg13g2_o21ai_1 _07426_ (.B1(_01897_),
    .Y(_01963_),
    .A1(_01889_),
    .A2(_01898_));
 sg13g2_o21ai_1 _07427_ (.B1(_01921_),
    .Y(_01964_),
    .A1(_01900_),
    .A2(_01922_));
 sg13g2_and2_1 _07428_ (.A(_01940_),
    .B(_01964_),
    .X(_01965_));
 sg13g2_xor2_1 _07429_ (.B(_01964_),
    .A(_01940_),
    .X(_01966_));
 sg13g2_xnor2_1 _07430_ (.Y(_01967_),
    .A(_01963_),
    .B(_01966_));
 sg13g2_inv_1 _07431_ (.Y(_01968_),
    .A(_01967_));
 sg13g2_o21ai_1 _07432_ (.B1(_01894_),
    .Y(_01969_),
    .A1(_01891_),
    .A2(_01895_));
 sg13g2_inv_1 _07433_ (.Y(_01970_),
    .A(_01969_));
 sg13g2_or2_1 _07434_ (.X(_01971_),
    .B(_01906_),
    .A(_01904_));
 sg13g2_nand2_1 _07435_ (.Y(_01972_),
    .A(net1443),
    .B(net1225));
 sg13g2_nand2_1 _07436_ (.Y(_01973_),
    .A(net1454),
    .B(net1211));
 sg13g2_nand2_1 _07437_ (.Y(_01974_),
    .A(net1454),
    .B(net1218));
 sg13g2_or2_1 _07438_ (.X(_01975_),
    .B(_01973_),
    .A(_01893_));
 sg13g2_xnor2_1 _07439_ (.Y(_01976_),
    .A(_01892_),
    .B(_01974_));
 sg13g2_xor2_1 _07440_ (.B(_01976_),
    .A(_01972_),
    .X(_01977_));
 sg13g2_nand2_1 _07441_ (.Y(_01978_),
    .A(_01971_),
    .B(_01977_));
 sg13g2_xnor2_1 _07442_ (.Y(_01979_),
    .A(_01971_),
    .B(_01977_));
 sg13g2_xnor2_1 _07443_ (.Y(_01980_),
    .A(_01970_),
    .B(_01979_));
 sg13g2_o21ai_1 _07444_ (.B1(_01917_),
    .Y(_01981_),
    .A1(_01908_),
    .A2(_01918_));
 sg13g2_nand2_1 _07445_ (.Y(_01982_),
    .A(net1464),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ));
 sg13g2_nand2_1 _07446_ (.Y(_01983_),
    .A(net1469),
    .B(net1196));
 sg13g2_nand2_1 _07447_ (.Y(_01984_),
    .A(net1469),
    .B(net1202));
 sg13g2_xor2_1 _07448_ (.B(_01984_),
    .A(_01903_),
    .X(_01985_));
 sg13g2_nand2b_1 _07449_ (.Y(_01986_),
    .B(_01985_),
    .A_N(_01982_));
 sg13g2_xnor2_1 _07450_ (.Y(_01987_),
    .A(_01982_),
    .B(_01985_));
 sg13g2_o21ai_1 _07451_ (.B1(_01912_),
    .Y(_01988_),
    .A1(_01910_),
    .A2(_01913_));
 sg13g2_nand2_1 _07452_ (.Y(_01989_),
    .A(net1355),
    .B(net1191));
 sg13g2_and4_1 _07453_ (.A(net1369),
    .B(net1362),
    .C(net1185),
    .D(net1180),
    .X(_01990_));
 sg13g2_a22oi_1 _07454_ (.Y(_01991_),
    .B1(net1180),
    .B2(net1369),
    .A2(net1185),
    .A1(net1362));
 sg13g2_or3_1 _07455_ (.A(_01989_),
    .B(_01990_),
    .C(_01991_),
    .X(_01992_));
 sg13g2_o21ai_1 _07456_ (.B1(_01989_),
    .Y(_01993_),
    .A1(_01990_),
    .A2(_01991_));
 sg13g2_nand3_1 _07457_ (.B(_01992_),
    .C(_01993_),
    .A(_01988_),
    .Y(_01994_));
 sg13g2_a21o_1 _07458_ (.A2(_01993_),
    .A1(_01992_),
    .B1(_01988_),
    .X(_01995_));
 sg13g2_nand3_1 _07459_ (.B(_01994_),
    .C(_01995_),
    .A(_01987_),
    .Y(_01996_));
 sg13g2_a21o_1 _07460_ (.A2(_01995_),
    .A1(_01994_),
    .B1(_01987_),
    .X(_01997_));
 sg13g2_nand3_1 _07461_ (.B(_01996_),
    .C(_01997_),
    .A(_01981_),
    .Y(_01998_));
 sg13g2_a21o_1 _07462_ (.A2(_01997_),
    .A1(_01996_),
    .B1(_01981_),
    .X(_01999_));
 sg13g2_nand2_1 _07463_ (.Y(_02000_),
    .A(_01998_),
    .B(_01999_));
 sg13g2_xnor2_1 _07464_ (.Y(_02001_),
    .A(_01980_),
    .B(_02000_));
 sg13g2_nand2_1 _07465_ (.Y(_02002_),
    .A(net1374),
    .B(net1176));
 sg13g2_nand2_1 _07466_ (.Y(_02003_),
    .A(net1383),
    .B(net1172));
 sg13g2_or2_1 _07467_ (.X(_02004_),
    .B(_02003_),
    .A(_01927_));
 sg13g2_xor2_1 _07468_ (.B(_02003_),
    .A(_01927_),
    .X(_02005_));
 sg13g2_nand2b_1 _07469_ (.Y(_02006_),
    .B(_02005_),
    .A_N(_02002_));
 sg13g2_xnor2_1 _07470_ (.Y(_02007_),
    .A(_02002_),
    .B(_02005_));
 sg13g2_nor2_1 _07471_ (.A(_01928_),
    .B(_01930_),
    .Y(_02008_));
 sg13g2_nand2b_1 _07472_ (.Y(_02009_),
    .B(_02007_),
    .A_N(_02008_));
 sg13g2_xnor2_1 _07473_ (.Y(_02010_),
    .A(_02007_),
    .B(_02008_));
 sg13g2_nand2b_1 _07474_ (.Y(_02011_),
    .B(_02010_),
    .A_N(_01934_));
 sg13g2_xnor2_1 _07475_ (.Y(_02012_),
    .A(_01934_),
    .B(_02010_));
 sg13g2_nand2_1 _07476_ (.Y(_02013_),
    .A(_01936_),
    .B(_02010_));
 sg13g2_xnor2_1 _07477_ (.Y(_02014_),
    .A(_01936_),
    .B(_02012_));
 sg13g2_xor2_1 _07478_ (.B(_02014_),
    .A(_02001_),
    .X(_02015_));
 sg13g2_nand2b_1 _07479_ (.Y(_02016_),
    .B(_02015_),
    .A_N(_01939_));
 sg13g2_xnor2_1 _07480_ (.Y(_02017_),
    .A(_01939_),
    .B(_02015_));
 sg13g2_nand2_1 _07481_ (.Y(_02018_),
    .A(net1449),
    .B(net1219));
 sg13g2_nand2_2 _07482_ (.Y(_02019_),
    .A(net1399),
    .B(net1155));
 sg13g2_nor2_2 _07483_ (.A(_01885_),
    .B(_02019_),
    .Y(_02020_));
 sg13g2_a22oi_1 _07484_ (.Y(_02021_),
    .B1(net1155),
    .B2(net1404),
    .A2(net1160),
    .A1(net1399));
 sg13g2_nor3_2 _07485_ (.A(_02018_),
    .B(_02020_),
    .C(_02021_),
    .Y(_02022_));
 sg13g2_o21ai_1 _07486_ (.B1(_02018_),
    .Y(_02023_),
    .A1(_02020_),
    .A2(_02021_));
 sg13g2_nor2b_1 _07487_ (.A(_02022_),
    .B_N(_02023_),
    .Y(_02024_));
 sg13g2_nor2b_1 _07488_ (.A(_01886_),
    .B_N(_02024_),
    .Y(_02025_));
 sg13g2_xnor2_1 _07489_ (.Y(_02026_),
    .A(_01886_),
    .B(_02024_));
 sg13g2_xnor2_1 _07490_ (.Y(_02027_),
    .A(_02017_),
    .B(_02026_));
 sg13g2_nor2_1 _07491_ (.A(_01942_),
    .B(_02027_),
    .Y(_02028_));
 sg13g2_xor2_1 _07492_ (.B(_02027_),
    .A(_01942_),
    .X(_02029_));
 sg13g2_xnor2_1 _07493_ (.Y(_02030_),
    .A(_01967_),
    .B(_02029_));
 sg13g2_nand2_1 _07494_ (.Y(_02031_),
    .A(_01962_),
    .B(_02030_));
 sg13g2_xnor2_1 _07495_ (.Y(_02032_),
    .A(_01962_),
    .B(_02030_));
 sg13g2_or2_1 _07496_ (.X(_02033_),
    .B(_02032_),
    .A(_01961_));
 sg13g2_xnor2_1 _07497_ (.Y(_02034_),
    .A(_01961_),
    .B(_02032_));
 sg13g2_nor2b_1 _07498_ (.A(_02034_),
    .B_N(_01960_),
    .Y(_02035_));
 sg13g2_xnor2_1 _07499_ (.Y(_02036_),
    .A(_01960_),
    .B(_02034_));
 sg13g2_a21oi_1 _07500_ (.A1(_01655_),
    .A2(_01696_),
    .Y(_02037_),
    .B1(_01955_));
 sg13g2_a21o_1 _07501_ (.A2(_01696_),
    .A1(_01655_),
    .B1(_01955_),
    .X(_02038_));
 sg13g2_o21ai_1 _07502_ (.B1(_02037_),
    .Y(_02039_),
    .A1(_01698_),
    .A2(_01874_));
 sg13g2_or3_1 _07503_ (.A(_01698_),
    .B(_01874_),
    .C(_01956_),
    .X(_02040_));
 sg13g2_a21oi_1 _07504_ (.A1(_01954_),
    .A2(_02039_),
    .Y(_02041_),
    .B1(_02036_));
 sg13g2_nand3_1 _07505_ (.B(_02036_),
    .C(_02039_),
    .A(_01954_),
    .Y(_02042_));
 sg13g2_nand2b_2 _07506_ (.Y(_02043_),
    .B(_02042_),
    .A_N(_02041_));
 sg13g2_o21ai_1 _07507_ (.B1(net1519),
    .Y(_02044_),
    .A1(net1297),
    .A2(net310));
 sg13g2_a21oi_1 _07508_ (.A1(net1298),
    .A2(_02043_),
    .Y(_00226_),
    .B1(_02044_));
 sg13g2_a21oi_1 _07509_ (.A1(_01963_),
    .A2(_01966_),
    .Y(_02045_),
    .B1(_01965_));
 sg13g2_a21o_1 _07510_ (.A2(_02029_),
    .A1(_01968_),
    .B1(_02028_),
    .X(_02046_));
 sg13g2_o21ai_1 _07511_ (.B1(_01978_),
    .Y(_02047_),
    .A1(_01970_),
    .A2(_01979_));
 sg13g2_o21ai_1 _07512_ (.B1(_01998_),
    .Y(_02048_),
    .A1(_01980_),
    .A2(_02000_));
 sg13g2_nor2b_1 _07513_ (.A(_02016_),
    .B_N(_02048_),
    .Y(_02049_));
 sg13g2_xor2_1 _07514_ (.B(_02048_),
    .A(_02016_),
    .X(_02050_));
 sg13g2_nor2b_1 _07515_ (.A(_02050_),
    .B_N(_02047_),
    .Y(_02051_));
 sg13g2_xor2_1 _07516_ (.B(_02050_),
    .A(_02047_),
    .X(_02052_));
 sg13g2_a21o_1 _07517_ (.A2(_02026_),
    .A1(_02017_),
    .B1(_02025_),
    .X(_02053_));
 sg13g2_o21ai_1 _07518_ (.B1(_01975_),
    .Y(_02054_),
    .A1(_01972_),
    .A2(_01976_));
 sg13g2_o21ai_1 _07519_ (.B1(_01986_),
    .Y(_02055_),
    .A1(_01903_),
    .A2(_01984_));
 sg13g2_nand2_1 _07520_ (.Y(_02056_),
    .A(net1438),
    .B(net1225));
 sg13g2_nand2_1 _07521_ (.Y(_02057_),
    .A(net1449),
    .B(net1211));
 sg13g2_nand2_1 _07522_ (.Y(_02058_),
    .A(net1449),
    .B(net1216));
 sg13g2_xor2_1 _07523_ (.B(_02058_),
    .A(_01973_),
    .X(_02059_));
 sg13g2_nand2b_1 _07524_ (.Y(_02060_),
    .B(_02059_),
    .A_N(_02056_));
 sg13g2_xnor2_1 _07525_ (.Y(_02061_),
    .A(_02056_),
    .B(_02059_));
 sg13g2_xnor2_1 _07526_ (.Y(_02062_),
    .A(_02055_),
    .B(_02061_));
 sg13g2_nor2b_1 _07527_ (.A(_02062_),
    .B_N(_02054_),
    .Y(_02063_));
 sg13g2_xor2_1 _07528_ (.B(_02062_),
    .A(_02054_),
    .X(_02064_));
 sg13g2_nand2_1 _07529_ (.Y(_02065_),
    .A(_01994_),
    .B(_01996_));
 sg13g2_nand2_1 _07530_ (.Y(_02066_),
    .A(net1459),
    .B(net1205));
 sg13g2_nand2_1 _07531_ (.Y(_02067_),
    .A(net1462),
    .B(net1196));
 sg13g2_nand2_1 _07532_ (.Y(_02068_),
    .A(net1463),
    .B(net1202));
 sg13g2_xor2_1 _07533_ (.B(_02068_),
    .A(_01983_),
    .X(_02069_));
 sg13g2_nand2b_1 _07534_ (.Y(_02070_),
    .B(_02069_),
    .A_N(_02066_));
 sg13g2_xor2_1 _07535_ (.B(_02069_),
    .A(_02066_),
    .X(_02071_));
 sg13g2_nand2b_1 _07536_ (.Y(_02072_),
    .B(_01992_),
    .A_N(_01990_));
 sg13g2_nand2_1 _07537_ (.Y(_02073_),
    .A(net1472),
    .B(net1191));
 sg13g2_nand2_2 _07538_ (.Y(_02074_),
    .A(net1353),
    .B(net1182));
 sg13g2_and4_1 _07539_ (.A(net1360),
    .B(net1353),
    .C(net1188),
    .D(net1182),
    .X(_02075_));
 sg13g2_a22oi_1 _07540_ (.Y(_02076_),
    .B1(net1182),
    .B2(net1364),
    .A2(net1188),
    .A1(net1353));
 sg13g2_nor3_1 _07541_ (.A(_02073_),
    .B(_02075_),
    .C(_02076_),
    .Y(_02077_));
 sg13g2_o21ai_1 _07542_ (.B1(_02073_),
    .Y(_02078_),
    .A1(_02075_),
    .A2(_02076_));
 sg13g2_nor2b_2 _07543_ (.A(_02077_),
    .B_N(_02078_),
    .Y(_02079_));
 sg13g2_nand2_1 _07544_ (.Y(_02080_),
    .A(_02072_),
    .B(_02079_));
 sg13g2_xnor2_1 _07545_ (.Y(_02081_),
    .A(_02072_),
    .B(_02079_));
 sg13g2_xor2_1 _07546_ (.B(_02081_),
    .A(_02071_),
    .X(_02082_));
 sg13g2_nand2_1 _07547_ (.Y(_02083_),
    .A(_02065_),
    .B(_02082_));
 sg13g2_xnor2_1 _07548_ (.Y(_02084_),
    .A(_02065_),
    .B(_02082_));
 sg13g2_xnor2_1 _07549_ (.Y(_02085_),
    .A(_02064_),
    .B(_02084_));
 sg13g2_nand2_1 _07550_ (.Y(_02086_),
    .A(_02009_),
    .B(_02011_));
 sg13g2_and2_1 _07551_ (.A(_02004_),
    .B(_02006_),
    .X(_02087_));
 sg13g2_nand2_1 _07552_ (.Y(_02088_),
    .A(net1367),
    .B(net1176));
 sg13g2_and4_1 _07553_ (.A(net1381),
    .B(net1374),
    .C(net1170),
    .D(net1165),
    .X(_02089_));
 sg13g2_a22oi_1 _07554_ (.Y(_02090_),
    .B1(net1165),
    .B2(net1381),
    .A2(net1170),
    .A1(net1374));
 sg13g2_nor3_1 _07555_ (.A(_02088_),
    .B(_02089_),
    .C(_02090_),
    .Y(_02091_));
 sg13g2_o21ai_1 _07556_ (.B1(_02088_),
    .Y(_02092_),
    .A1(_02089_),
    .A2(_02090_));
 sg13g2_nor2b_2 _07557_ (.A(_02091_),
    .B_N(_02092_),
    .Y(_02093_));
 sg13g2_nand2_1 _07558_ (.Y(_02094_),
    .A(_02020_),
    .B(_02093_));
 sg13g2_nor2_1 _07559_ (.A(_02020_),
    .B(_02093_),
    .Y(_02095_));
 sg13g2_xor2_1 _07560_ (.B(_02093_),
    .A(_02020_),
    .X(_02096_));
 sg13g2_xnor2_1 _07561_ (.Y(_02097_),
    .A(_02087_),
    .B(_02096_));
 sg13g2_xnor2_1 _07562_ (.Y(_02098_),
    .A(_02086_),
    .B(_02097_));
 sg13g2_xnor2_1 _07563_ (.Y(_02099_),
    .A(_02085_),
    .B(_02098_));
 sg13g2_o21ai_1 _07564_ (.B1(_02013_),
    .Y(_02100_),
    .A1(_02001_),
    .A2(_02014_));
 sg13g2_nand2b_1 _07565_ (.Y(_02101_),
    .B(_02100_),
    .A_N(_02099_));
 sg13g2_xor2_1 _07566_ (.B(_02100_),
    .A(_02099_),
    .X(_02102_));
 sg13g2_nand2_1 _07567_ (.Y(_02103_),
    .A(net1443),
    .B(net1219));
 sg13g2_nand2_1 _07568_ (.Y(_02104_),
    .A(net1388),
    .B(net1159));
 sg13g2_nand2_1 _07569_ (.Y(_02105_),
    .A(net1404),
    .B(net1149));
 sg13g2_or2_1 _07570_ (.X(_02106_),
    .B(_02105_),
    .A(_02019_));
 sg13g2_and2_1 _07571_ (.A(_02019_),
    .B(_02105_),
    .X(_02107_));
 sg13g2_xor2_1 _07572_ (.B(_02105_),
    .A(_02019_),
    .X(_02108_));
 sg13g2_xnor2_1 _07573_ (.Y(_02109_),
    .A(_02104_),
    .B(_02108_));
 sg13g2_nand2b_1 _07574_ (.Y(_02110_),
    .B(_02109_),
    .A_N(_02103_));
 sg13g2_xnor2_1 _07575_ (.Y(_02111_),
    .A(_02103_),
    .B(_02109_));
 sg13g2_nand2_1 _07576_ (.Y(_02112_),
    .A(_02022_),
    .B(_02111_));
 sg13g2_xnor2_1 _07577_ (.Y(_02113_),
    .A(_02022_),
    .B(_02111_));
 sg13g2_xor2_1 _07578_ (.B(_02113_),
    .A(_02102_),
    .X(_02114_));
 sg13g2_nand2_1 _07579_ (.Y(_02115_),
    .A(_02053_),
    .B(_02114_));
 sg13g2_xnor2_1 _07580_ (.Y(_02116_),
    .A(_02053_),
    .B(_02114_));
 sg13g2_xor2_1 _07581_ (.B(_02116_),
    .A(_02052_),
    .X(_02117_));
 sg13g2_nand2_1 _07582_ (.Y(_02118_),
    .A(_02046_),
    .B(_02117_));
 sg13g2_xnor2_1 _07583_ (.Y(_02119_),
    .A(_02046_),
    .B(_02117_));
 sg13g2_xnor2_1 _07584_ (.Y(_02120_),
    .A(_02045_),
    .B(_02119_));
 sg13g2_nand3_1 _07585_ (.B(_02033_),
    .C(_02120_),
    .A(_02031_),
    .Y(_02121_));
 sg13g2_a21oi_1 _07586_ (.A1(_02031_),
    .A2(_02033_),
    .Y(_02122_),
    .B1(_02120_));
 sg13g2_inv_1 _07587_ (.Y(_02123_),
    .A(_02122_));
 sg13g2_nand2_1 _07588_ (.Y(_02124_),
    .A(_02121_),
    .B(_02123_));
 sg13g2_nor2b_1 _07589_ (.A(_02035_),
    .B_N(_02042_),
    .Y(_02125_));
 sg13g2_xnor2_1 _07590_ (.Y(_02126_),
    .A(_02124_),
    .B(_02125_));
 sg13g2_o21ai_1 _07591_ (.B1(net1519),
    .Y(_02127_),
    .A1(net1298),
    .A2(net300));
 sg13g2_a21oi_1 _07592_ (.A1(net1298),
    .A2(_02126_),
    .Y(_00227_),
    .B1(_02127_));
 sg13g2_nor2_1 _07593_ (.A(_02049_),
    .B(_02051_),
    .Y(_02128_));
 sg13g2_o21ai_1 _07594_ (.B1(_02115_),
    .Y(_02129_),
    .A1(_02052_),
    .A2(_02116_));
 sg13g2_a21o_1 _07595_ (.A2(_02061_),
    .A1(_02055_),
    .B1(_02063_),
    .X(_02130_));
 sg13g2_o21ai_1 _07596_ (.B1(_02083_),
    .Y(_02131_),
    .A1(_02064_),
    .A2(_02084_));
 sg13g2_inv_1 _07597_ (.Y(_02132_),
    .A(_02131_));
 sg13g2_xnor2_1 _07598_ (.Y(_02133_),
    .A(_02101_),
    .B(_02132_));
 sg13g2_nand2b_1 _07599_ (.Y(_02134_),
    .B(_02130_),
    .A_N(_02133_));
 sg13g2_xor2_1 _07600_ (.B(_02133_),
    .A(_02130_),
    .X(_02135_));
 sg13g2_o21ai_1 _07601_ (.B1(_02112_),
    .Y(_02136_),
    .A1(_02102_),
    .A2(_02113_));
 sg13g2_o21ai_1 _07602_ (.B1(_02060_),
    .Y(_02137_),
    .A1(_01973_),
    .A2(_02058_));
 sg13g2_o21ai_1 _07603_ (.B1(_02070_),
    .Y(_02138_),
    .A1(_01983_),
    .A2(_02068_));
 sg13g2_nand2_1 _07604_ (.Y(_02139_),
    .A(net1434),
    .B(net1225));
 sg13g2_nand2_1 _07605_ (.Y(_02140_),
    .A(net1444),
    .B(net1211));
 sg13g2_nand2_1 _07606_ (.Y(_02141_),
    .A(net1444),
    .B(net1216));
 sg13g2_xor2_1 _07607_ (.B(_02141_),
    .A(_02057_),
    .X(_02142_));
 sg13g2_nand2b_1 _07608_ (.Y(_02143_),
    .B(_02142_),
    .A_N(_02139_));
 sg13g2_xnor2_1 _07609_ (.Y(_02144_),
    .A(_02139_),
    .B(_02142_));
 sg13g2_xnor2_1 _07610_ (.Y(_02145_),
    .A(_02138_),
    .B(_02144_));
 sg13g2_nor2b_1 _07611_ (.A(_02145_),
    .B_N(_02137_),
    .Y(_02146_));
 sg13g2_xor2_1 _07612_ (.B(_02145_),
    .A(_02137_),
    .X(_02147_));
 sg13g2_o21ai_1 _07613_ (.B1(_02080_),
    .Y(_02148_),
    .A1(_02071_),
    .A2(_02081_));
 sg13g2_nand2_1 _07614_ (.Y(_02149_),
    .A(net1454),
    .B(net1206));
 sg13g2_nand2_1 _07615_ (.Y(_02150_),
    .A(net1457),
    .B(net1196));
 sg13g2_nand2_1 _07616_ (.Y(_02151_),
    .A(net1457),
    .B(net1202));
 sg13g2_xor2_1 _07617_ (.B(_02151_),
    .A(_02067_),
    .X(_02152_));
 sg13g2_nand2b_1 _07618_ (.Y(_02153_),
    .B(_02152_),
    .A_N(_02149_));
 sg13g2_xor2_1 _07619_ (.B(_02152_),
    .A(_02149_),
    .X(_02154_));
 sg13g2_or2_1 _07620_ (.X(_02155_),
    .B(_02077_),
    .A(_02075_));
 sg13g2_nand2_1 _07621_ (.Y(_02156_),
    .A(net1468),
    .B(net1192));
 sg13g2_nand2_1 _07622_ (.Y(_02157_),
    .A(net1471),
    .B(net1188));
 sg13g2_or2_1 _07623_ (.X(_02158_),
    .B(_02157_),
    .A(_02074_));
 sg13g2_and2_1 _07624_ (.A(_02074_),
    .B(_02157_),
    .X(_02159_));
 sg13g2_xor2_1 _07625_ (.B(_02157_),
    .A(_02074_),
    .X(_02160_));
 sg13g2_xnor2_1 _07626_ (.Y(_02161_),
    .A(_02156_),
    .B(_02160_));
 sg13g2_nand2_1 _07627_ (.Y(_02162_),
    .A(_02155_),
    .B(_02161_));
 sg13g2_xnor2_1 _07628_ (.Y(_02163_),
    .A(_02155_),
    .B(_02161_));
 sg13g2_xor2_1 _07629_ (.B(_02163_),
    .A(_02154_),
    .X(_02164_));
 sg13g2_nand2_1 _07630_ (.Y(_02165_),
    .A(_02148_),
    .B(_02164_));
 sg13g2_xnor2_1 _07631_ (.Y(_02166_),
    .A(_02148_),
    .B(_02164_));
 sg13g2_xor2_1 _07632_ (.B(_02166_),
    .A(_02147_),
    .X(_02167_));
 sg13g2_nor2b_2 _07633_ (.A(_02009_),
    .B_N(_02097_),
    .Y(_02168_));
 sg13g2_o21ai_1 _07634_ (.B1(_02094_),
    .Y(_02169_),
    .A1(_02087_),
    .A2(_02095_));
 sg13g2_or2_1 _07635_ (.X(_02170_),
    .B(_02091_),
    .A(_02089_));
 sg13g2_o21ai_1 _07636_ (.B1(_02106_),
    .Y(_02171_),
    .A1(_02104_),
    .A2(_02107_));
 sg13g2_nand2_1 _07637_ (.Y(_02172_),
    .A(net1360),
    .B(net1175));
 sg13g2_and4_1 _07638_ (.A(net1374),
    .B(net1366),
    .C(net1170),
    .D(net1163),
    .X(_02173_));
 sg13g2_a22oi_1 _07639_ (.Y(_02174_),
    .B1(net1164),
    .B2(net1374),
    .A2(net1170),
    .A1(net1367));
 sg13g2_nor3_1 _07640_ (.A(_02172_),
    .B(_02173_),
    .C(_02174_),
    .Y(_02175_));
 sg13g2_o21ai_1 _07641_ (.B1(_02172_),
    .Y(_02176_),
    .A1(_02173_),
    .A2(_02174_));
 sg13g2_nor2b_1 _07642_ (.A(_02175_),
    .B_N(_02176_),
    .Y(_02177_));
 sg13g2_and2_1 _07643_ (.A(_02171_),
    .B(_02177_),
    .X(_02178_));
 sg13g2_xor2_1 _07644_ (.B(_02177_),
    .A(_02171_),
    .X(_02179_));
 sg13g2_xnor2_1 _07645_ (.Y(_02180_),
    .A(_02170_),
    .B(_02179_));
 sg13g2_nand2b_1 _07646_ (.Y(_02181_),
    .B(_02169_),
    .A_N(_02180_));
 sg13g2_xnor2_1 _07647_ (.Y(_02182_),
    .A(_02169_),
    .B(_02180_));
 sg13g2_and2_1 _07648_ (.A(_02168_),
    .B(_02182_),
    .X(_02183_));
 sg13g2_or2_1 _07649_ (.X(_02184_),
    .B(_02182_),
    .A(_02168_));
 sg13g2_xor2_1 _07650_ (.B(_02182_),
    .A(_02168_),
    .X(_02185_));
 sg13g2_xnor2_1 _07651_ (.Y(_02186_),
    .A(_02167_),
    .B(_02185_));
 sg13g2_nand2b_1 _07652_ (.Y(_02187_),
    .B(_02097_),
    .A_N(_02011_));
 sg13g2_o21ai_1 _07653_ (.B1(_02187_),
    .Y(_02188_),
    .A1(_02085_),
    .A2(_02098_));
 sg13g2_nand2b_1 _07654_ (.Y(_02189_),
    .B(_02188_),
    .A_N(_02186_));
 sg13g2_xor2_1 _07655_ (.B(_02188_),
    .A(_02186_),
    .X(_02190_));
 sg13g2_nand2_1 _07656_ (.Y(_02191_),
    .A(net1438),
    .B(net1219));
 sg13g2_nand2_2 _07657_ (.Y(_02192_),
    .A(net1404),
    .B(net1350));
 sg13g2_nand2_1 _07658_ (.Y(_02193_),
    .A(net1381),
    .B(net1159));
 sg13g2_and4_1 _07659_ (.A(net1397),
    .B(net1388),
    .C(net1155),
    .D(net1149),
    .X(_02194_));
 sg13g2_nand4_1 _07660_ (.B(net1388),
    .C(net1155),
    .A(net1396),
    .Y(_02195_),
    .D(net1149));
 sg13g2_a22oi_1 _07661_ (.Y(_02196_),
    .B1(net1149),
    .B2(net1397),
    .A2(net1155),
    .A1(net1388));
 sg13g2_nor3_1 _07662_ (.A(_02193_),
    .B(_02194_),
    .C(_02196_),
    .Y(_02197_));
 sg13g2_o21ai_1 _07663_ (.B1(_02193_),
    .Y(_02198_),
    .A1(_02194_),
    .A2(_02196_));
 sg13g2_nor2b_1 _07664_ (.A(_02197_),
    .B_N(_02198_),
    .Y(_02199_));
 sg13g2_nor2b_2 _07665_ (.A(_02192_),
    .B_N(_02199_),
    .Y(_02200_));
 sg13g2_xnor2_1 _07666_ (.Y(_02201_),
    .A(_02192_),
    .B(_02199_));
 sg13g2_nor2b_1 _07667_ (.A(_02191_),
    .B_N(_02201_),
    .Y(_02202_));
 sg13g2_xnor2_1 _07668_ (.Y(_02203_),
    .A(_02191_),
    .B(_02201_));
 sg13g2_nand2b_1 _07669_ (.Y(_02204_),
    .B(_02203_),
    .A_N(_02110_));
 sg13g2_xnor2_1 _07670_ (.Y(_02205_),
    .A(_02110_),
    .B(_02203_));
 sg13g2_inv_1 _07671_ (.Y(_02206_),
    .A(_02205_));
 sg13g2_xnor2_1 _07672_ (.Y(_02207_),
    .A(_02190_),
    .B(_02205_));
 sg13g2_nand2_1 _07673_ (.Y(_02208_),
    .A(_02136_),
    .B(_02207_));
 sg13g2_xnor2_1 _07674_ (.Y(_02209_),
    .A(_02136_),
    .B(_02207_));
 sg13g2_xor2_1 _07675_ (.B(_02209_),
    .A(_02135_),
    .X(_02210_));
 sg13g2_nand2_1 _07676_ (.Y(_02211_),
    .A(_02129_),
    .B(_02210_));
 sg13g2_xnor2_1 _07677_ (.Y(_02212_),
    .A(_02129_),
    .B(_02210_));
 sg13g2_xor2_1 _07678_ (.B(_02212_),
    .A(_02128_),
    .X(_02213_));
 sg13g2_o21ai_1 _07679_ (.B1(_02118_),
    .Y(_02214_),
    .A1(_02045_),
    .A2(_02119_));
 sg13g2_and2_1 _07680_ (.A(_02213_),
    .B(_02214_),
    .X(_02215_));
 sg13g2_inv_1 _07681_ (.Y(_02216_),
    .A(_02215_));
 sg13g2_xor2_1 _07682_ (.B(_02214_),
    .A(_02213_),
    .X(_02217_));
 sg13g2_inv_1 _07683_ (.Y(_02218_),
    .A(_02217_));
 sg13g2_a21oi_1 _07684_ (.A1(_02035_),
    .A2(_02121_),
    .Y(_02219_),
    .B1(_02122_));
 sg13g2_nand3b_1 _07685_ (.B(_02036_),
    .C(_02121_),
    .Y(_02220_),
    .A_N(_02122_));
 sg13g2_a221oi_1 _07686_ (.B2(_02035_),
    .C1(_02122_),
    .B1(_02121_),
    .A1(_01954_),
    .Y(_02221_),
    .A2(_02038_));
 sg13g2_o21ai_1 _07687_ (.B1(_02219_),
    .Y(_02222_),
    .A1(_02042_),
    .A2(_02124_));
 sg13g2_a221oi_1 _07688_ (.B2(_02040_),
    .C1(_02218_),
    .B1(_02221_),
    .A1(_02219_),
    .Y(_02223_),
    .A2(_02220_));
 sg13g2_xnor2_1 _07689_ (.Y(_02224_),
    .A(_02218_),
    .B(_02222_));
 sg13g2_o21ai_1 _07690_ (.B1(net1517),
    .Y(_02225_),
    .A1(net1143),
    .A2(_02224_));
 sg13g2_a21oi_1 _07691_ (.A1(net1144),
    .A2(_04780_),
    .Y(_00228_),
    .B1(_02225_));
 sg13g2_o21ai_1 _07692_ (.B1(_02134_),
    .Y(_02226_),
    .A1(_02101_),
    .A2(_02132_));
 sg13g2_o21ai_1 _07693_ (.B1(_02208_),
    .Y(_02227_),
    .A1(_02135_),
    .A2(_02209_));
 sg13g2_a21o_1 _07694_ (.A2(_02144_),
    .A1(_02138_),
    .B1(_02146_),
    .X(_02228_));
 sg13g2_o21ai_1 _07695_ (.B1(_02165_),
    .Y(_02229_),
    .A1(_02147_),
    .A2(_02166_));
 sg13g2_inv_1 _07696_ (.Y(_02230_),
    .A(_02229_));
 sg13g2_xnor2_1 _07697_ (.Y(_02231_),
    .A(_02189_),
    .B(_02230_));
 sg13g2_nand2b_1 _07698_ (.Y(_02232_),
    .B(_02228_),
    .A_N(_02231_));
 sg13g2_xor2_1 _07699_ (.B(_02231_),
    .A(_02228_),
    .X(_02233_));
 sg13g2_o21ai_1 _07700_ (.B1(_02204_),
    .Y(_02234_),
    .A1(_02190_),
    .A2(_02206_));
 sg13g2_o21ai_1 _07701_ (.B1(_02143_),
    .Y(_02235_),
    .A1(_02057_),
    .A2(_02141_));
 sg13g2_o21ai_1 _07702_ (.B1(_02153_),
    .Y(_02236_),
    .A1(_02067_),
    .A2(_02151_));
 sg13g2_nand2_1 _07703_ (.Y(_02237_),
    .A(net1430),
    .B(net1225));
 sg13g2_nand2_1 _07704_ (.Y(_02238_),
    .A(net1439),
    .B(net1211));
 sg13g2_nand2_1 _07705_ (.Y(_02239_),
    .A(net1439),
    .B(net1218));
 sg13g2_or2_1 _07706_ (.X(_02240_),
    .B(_02238_),
    .A(_02141_));
 sg13g2_xnor2_1 _07707_ (.Y(_02241_),
    .A(_02140_),
    .B(_02239_));
 sg13g2_xor2_1 _07708_ (.B(_02241_),
    .A(_02237_),
    .X(_02242_));
 sg13g2_xnor2_1 _07709_ (.Y(_02243_),
    .A(_02236_),
    .B(_02242_));
 sg13g2_nor2b_1 _07710_ (.A(_02243_),
    .B_N(_02235_),
    .Y(_02244_));
 sg13g2_xor2_1 _07711_ (.B(_02243_),
    .A(_02235_),
    .X(_02245_));
 sg13g2_o21ai_1 _07712_ (.B1(_02162_),
    .Y(_02246_),
    .A1(_02154_),
    .A2(_02163_));
 sg13g2_nand2_1 _07713_ (.Y(_02247_),
    .A(net1449),
    .B(net1205));
 sg13g2_nand2_1 _07714_ (.Y(_02248_),
    .A(net1454),
    .B(net1196));
 sg13g2_nand2_1 _07715_ (.Y(_02249_),
    .A(net1454),
    .B(net1202));
 sg13g2_xor2_1 _07716_ (.B(_02249_),
    .A(_02150_),
    .X(_02250_));
 sg13g2_nand2b_1 _07717_ (.Y(_02251_),
    .B(_02250_),
    .A_N(_02247_));
 sg13g2_xor2_1 _07718_ (.B(_02250_),
    .A(_02247_),
    .X(_02252_));
 sg13g2_o21ai_1 _07719_ (.B1(_02158_),
    .Y(_02253_),
    .A1(_02156_),
    .A2(_02159_));
 sg13g2_nand2_1 _07720_ (.Y(_02254_),
    .A(net1462),
    .B(net1192));
 sg13g2_nand2_1 _07721_ (.Y(_02255_),
    .A(net1467),
    .B(net1182));
 sg13g2_and4_1 _07722_ (.A(net1471),
    .B(net1467),
    .C(net1188),
    .D(net1182),
    .X(_02256_));
 sg13g2_a22oi_1 _07723_ (.Y(_02257_),
    .B1(net1182),
    .B2(net1471),
    .A2(net1188),
    .A1(net1467));
 sg13g2_nor3_1 _07724_ (.A(_02254_),
    .B(_02256_),
    .C(_02257_),
    .Y(_02258_));
 sg13g2_o21ai_1 _07725_ (.B1(_02254_),
    .Y(_02259_),
    .A1(_02256_),
    .A2(_02257_));
 sg13g2_nor2b_1 _07726_ (.A(_02258_),
    .B_N(_02259_),
    .Y(_02260_));
 sg13g2_nand2_1 _07727_ (.Y(_02261_),
    .A(_02253_),
    .B(_02260_));
 sg13g2_xnor2_1 _07728_ (.Y(_02262_),
    .A(_02253_),
    .B(_02260_));
 sg13g2_xnor2_1 _07729_ (.Y(_02263_),
    .A(_02252_),
    .B(_02262_));
 sg13g2_nand2b_1 _07730_ (.Y(_02264_),
    .B(_02246_),
    .A_N(_02263_));
 sg13g2_xor2_1 _07731_ (.B(_02263_),
    .A(_02246_),
    .X(_02265_));
 sg13g2_xor2_1 _07732_ (.B(_02265_),
    .A(_02245_),
    .X(_02266_));
 sg13g2_a21oi_1 _07733_ (.A1(_02170_),
    .A2(_02179_),
    .Y(_02267_),
    .B1(_02178_));
 sg13g2_or2_1 _07734_ (.X(_02268_),
    .B(_02175_),
    .A(_02173_));
 sg13g2_o21ai_1 _07735_ (.B1(_02195_),
    .Y(_02269_),
    .A1(_02193_),
    .A2(_02196_));
 sg13g2_nand2_1 _07736_ (.Y(_02270_),
    .A(net1354),
    .B(net1175));
 sg13g2_and4_1 _07737_ (.A(net1367),
    .B(net1361),
    .C(net1170),
    .D(net1163),
    .X(_02271_));
 sg13g2_a22oi_1 _07738_ (.Y(_02272_),
    .B1(net1164),
    .B2(net1367),
    .A2(net1170),
    .A1(net1361));
 sg13g2_or3_1 _07739_ (.A(_02270_),
    .B(_02271_),
    .C(_02272_),
    .X(_02273_));
 sg13g2_o21ai_1 _07740_ (.B1(_02270_),
    .Y(_02274_),
    .A1(_02271_),
    .A2(_02272_));
 sg13g2_nand3_1 _07741_ (.B(_02273_),
    .C(_02274_),
    .A(_02269_),
    .Y(_02275_));
 sg13g2_a21o_1 _07742_ (.A2(_02274_),
    .A1(_02273_),
    .B1(_02269_),
    .X(_02276_));
 sg13g2_nand3_1 _07743_ (.B(_02275_),
    .C(_02276_),
    .A(_02268_),
    .Y(_02277_));
 sg13g2_a21o_2 _07744_ (.A2(_02276_),
    .A1(_02275_),
    .B1(_02268_),
    .X(_02278_));
 sg13g2_and3_1 _07745_ (.X(_02279_),
    .A(_02200_),
    .B(_02277_),
    .C(_02278_));
 sg13g2_nand3_1 _07746_ (.B(_02277_),
    .C(_02278_),
    .A(_02200_),
    .Y(_02280_));
 sg13g2_a21oi_1 _07747_ (.A1(_02277_),
    .A2(_02278_),
    .Y(_02281_),
    .B1(_02200_));
 sg13g2_a21o_1 _07748_ (.A2(_02278_),
    .A1(_02277_),
    .B1(_02200_),
    .X(_02282_));
 sg13g2_nor3_1 _07749_ (.A(_02267_),
    .B(_02279_),
    .C(_02281_),
    .Y(_02283_));
 sg13g2_a221oi_1 _07750_ (.B2(_02282_),
    .C1(_02178_),
    .B1(_02280_),
    .A1(_02170_),
    .Y(_02284_),
    .A2(_02179_));
 sg13g2_nor3_1 _07751_ (.A(_02181_),
    .B(_02283_),
    .C(_02284_),
    .Y(_02285_));
 sg13g2_or3_1 _07752_ (.A(_02181_),
    .B(_02283_),
    .C(_02284_),
    .X(_02286_));
 sg13g2_o21ai_1 _07753_ (.B1(_02181_),
    .Y(_02287_),
    .A1(_02283_),
    .A2(_02284_));
 sg13g2_nand3_1 _07754_ (.B(_02286_),
    .C(_02287_),
    .A(_02266_),
    .Y(_02288_));
 sg13g2_a21o_1 _07755_ (.A2(_02287_),
    .A1(_02286_),
    .B1(_02266_),
    .X(_02289_));
 sg13g2_a21o_1 _07756_ (.A2(_02184_),
    .A1(_02167_),
    .B1(_02183_),
    .X(_02290_));
 sg13g2_and3_2 _07757_ (.X(_02291_),
    .A(_02288_),
    .B(_02289_),
    .C(_02290_));
 sg13g2_a21oi_1 _07758_ (.A1(_02288_),
    .A2(_02289_),
    .Y(_02292_),
    .B1(_02290_));
 sg13g2_nand2_2 _07759_ (.Y(_02293_),
    .A(net1434),
    .B(net1222));
 sg13g2_a22oi_1 _07760_ (.Y(_02294_),
    .B1(net1345),
    .B2(net1404),
    .A2(net1349),
    .A1(net1396));
 sg13g2_nor3_2 _07761_ (.A(_04805_),
    .B(_04836_),
    .C(_02192_),
    .Y(_02295_));
 sg13g2_nor2_1 _07762_ (.A(_02294_),
    .B(_02295_),
    .Y(_02296_));
 sg13g2_nand2_1 _07763_ (.Y(_02297_),
    .A(net1373),
    .B(net1159));
 sg13g2_and4_1 _07764_ (.A(net1387),
    .B(net1380),
    .C(net1153),
    .D(net1147),
    .X(_02298_));
 sg13g2_nand4_1 _07765_ (.B(net1380),
    .C(net1154),
    .A(net1387),
    .Y(_02299_),
    .D(net1147));
 sg13g2_a22oi_1 _07766_ (.Y(_02300_),
    .B1(net1147),
    .B2(net1387),
    .A2(net1153),
    .A1(net1380));
 sg13g2_nor3_1 _07767_ (.A(_02297_),
    .B(_02298_),
    .C(_02300_),
    .Y(_02301_));
 sg13g2_o21ai_1 _07768_ (.B1(_02297_),
    .Y(_02302_),
    .A1(_02298_),
    .A2(_02300_));
 sg13g2_nor2b_1 _07769_ (.A(_02301_),
    .B_N(_02302_),
    .Y(_02303_));
 sg13g2_and2_1 _07770_ (.A(_02296_),
    .B(_02303_),
    .X(_02304_));
 sg13g2_xor2_1 _07771_ (.B(_02303_),
    .A(_02296_),
    .X(_02305_));
 sg13g2_nor2b_1 _07772_ (.A(_02293_),
    .B_N(_02305_),
    .Y(_02306_));
 sg13g2_xor2_1 _07773_ (.B(_02305_),
    .A(_02293_),
    .X(_02307_));
 sg13g2_inv_1 _07774_ (.Y(_02308_),
    .A(_02307_));
 sg13g2_nand2_1 _07775_ (.Y(_02309_),
    .A(_02202_),
    .B(_02308_));
 sg13g2_xor2_1 _07776_ (.B(_02307_),
    .A(_02202_),
    .X(_02310_));
 sg13g2_or3_1 _07777_ (.A(_02291_),
    .B(_02292_),
    .C(_02310_),
    .X(_02311_));
 sg13g2_o21ai_1 _07778_ (.B1(_02310_),
    .Y(_02312_),
    .A1(_02291_),
    .A2(_02292_));
 sg13g2_and3_1 _07779_ (.X(_02313_),
    .A(_02234_),
    .B(_02311_),
    .C(_02312_));
 sg13g2_a21oi_1 _07780_ (.A1(_02311_),
    .A2(_02312_),
    .Y(_02314_),
    .B1(_02234_));
 sg13g2_nor3_1 _07781_ (.A(_02233_),
    .B(_02313_),
    .C(_02314_),
    .Y(_02315_));
 sg13g2_o21ai_1 _07782_ (.B1(_02233_),
    .Y(_02316_),
    .A1(_02313_),
    .A2(_02314_));
 sg13g2_nor2b_1 _07783_ (.A(_02315_),
    .B_N(_02316_),
    .Y(_02317_));
 sg13g2_and2_1 _07784_ (.A(_02227_),
    .B(_02317_),
    .X(_02318_));
 sg13g2_or2_1 _07785_ (.X(_02319_),
    .B(_02317_),
    .A(_02227_));
 sg13g2_xor2_1 _07786_ (.B(_02317_),
    .A(_02227_),
    .X(_02320_));
 sg13g2_xnor2_1 _07787_ (.Y(_02321_),
    .A(_02226_),
    .B(_02320_));
 sg13g2_o21ai_1 _07788_ (.B1(_02211_),
    .Y(_02322_),
    .A1(_02128_),
    .A2(_02212_));
 sg13g2_nor2b_1 _07789_ (.A(_02322_),
    .B_N(_02321_),
    .Y(_02323_));
 sg13g2_nand2b_1 _07790_ (.Y(_02324_),
    .B(_02322_),
    .A_N(_02321_));
 sg13g2_nor2b_2 _07791_ (.A(_02323_),
    .B_N(_02324_),
    .Y(_02325_));
 sg13g2_nor2_1 _07792_ (.A(_02215_),
    .B(_02223_),
    .Y(_02326_));
 sg13g2_xnor2_1 _07793_ (.Y(_02327_),
    .A(_02325_),
    .B(_02326_));
 sg13g2_o21ai_1 _07794_ (.B1(net1518),
    .Y(_02328_),
    .A1(net1143),
    .A2(_02327_));
 sg13g2_a21oi_1 _07795_ (.A1(net1144),
    .A2(_04779_),
    .Y(_00229_),
    .B1(_02328_));
 sg13g2_o21ai_1 _07796_ (.B1(_02232_),
    .Y(_02329_),
    .A1(_02189_),
    .A2(_02230_));
 sg13g2_inv_1 _07797_ (.Y(_02330_),
    .A(_02329_));
 sg13g2_or2_1 _07798_ (.X(_02331_),
    .B(_02315_),
    .A(_02313_));
 sg13g2_a21o_1 _07799_ (.A2(_02242_),
    .A1(_02236_),
    .B1(_02244_),
    .X(_02332_));
 sg13g2_o21ai_1 _07800_ (.B1(_02264_),
    .Y(_02333_),
    .A1(_02245_),
    .A2(_02265_));
 sg13g2_xor2_1 _07801_ (.B(_02333_),
    .A(_02291_),
    .X(_02334_));
 sg13g2_and2_1 _07802_ (.A(_02332_),
    .B(_02334_),
    .X(_02335_));
 sg13g2_xor2_1 _07803_ (.B(_02334_),
    .A(_02332_),
    .X(_02336_));
 sg13g2_nand2_1 _07804_ (.Y(_02337_),
    .A(_02309_),
    .B(_02311_));
 sg13g2_o21ai_1 _07805_ (.B1(_02240_),
    .Y(_02338_),
    .A1(_02237_),
    .A2(_02241_));
 sg13g2_o21ai_1 _07806_ (.B1(_02251_),
    .Y(_02339_),
    .A1(_02150_),
    .A2(_02249_));
 sg13g2_nand2_1 _07807_ (.Y(_02340_),
    .A(net1426),
    .B(net1225));
 sg13g2_nand2_1 _07808_ (.Y(_02341_),
    .A(net1434),
    .B(net1211));
 sg13g2_nand2_1 _07809_ (.Y(_02342_),
    .A(net1435),
    .B(net1218));
 sg13g2_or2_1 _07810_ (.X(_02343_),
    .B(_02341_),
    .A(_02239_));
 sg13g2_xnor2_1 _07811_ (.Y(_02344_),
    .A(_02238_),
    .B(_02342_));
 sg13g2_xor2_1 _07812_ (.B(_02344_),
    .A(_02340_),
    .X(_02345_));
 sg13g2_xnor2_1 _07813_ (.Y(_02346_),
    .A(_02339_),
    .B(_02345_));
 sg13g2_nor2b_1 _07814_ (.A(_02346_),
    .B_N(_02338_),
    .Y(_02347_));
 sg13g2_xor2_1 _07815_ (.B(_02346_),
    .A(_02338_),
    .X(_02348_));
 sg13g2_o21ai_1 _07816_ (.B1(_02261_),
    .Y(_02349_),
    .A1(_02252_),
    .A2(_02262_));
 sg13g2_nand2_1 _07817_ (.Y(_02350_),
    .A(net1444),
    .B(net1205));
 sg13g2_nand2_1 _07818_ (.Y(_02351_),
    .A(net1449),
    .B(net1196));
 sg13g2_nand2_1 _07819_ (.Y(_02352_),
    .A(net1449),
    .B(net1202));
 sg13g2_xor2_1 _07820_ (.B(_02352_),
    .A(_02248_),
    .X(_02353_));
 sg13g2_nand2b_1 _07821_ (.Y(_02354_),
    .B(_02353_),
    .A_N(_02350_));
 sg13g2_xor2_1 _07822_ (.B(_02353_),
    .A(_02350_),
    .X(_02355_));
 sg13g2_or2_1 _07823_ (.X(_02356_),
    .B(_02258_),
    .A(_02256_));
 sg13g2_nand2_1 _07824_ (.Y(_02357_),
    .A(net1457),
    .B(net1191));
 sg13g2_nand2_1 _07825_ (.Y(_02358_),
    .A(net1462),
    .B(net1188));
 sg13g2_or2_1 _07826_ (.X(_02359_),
    .B(_02358_),
    .A(_02255_));
 sg13g2_and2_1 _07827_ (.A(_02255_),
    .B(_02358_),
    .X(_02360_));
 sg13g2_xor2_1 _07828_ (.B(_02358_),
    .A(_02255_),
    .X(_02361_));
 sg13g2_xnor2_1 _07829_ (.Y(_02362_),
    .A(_02357_),
    .B(_02361_));
 sg13g2_nand2_1 _07830_ (.Y(_02363_),
    .A(_02356_),
    .B(_02362_));
 sg13g2_xnor2_1 _07831_ (.Y(_02364_),
    .A(_02356_),
    .B(_02362_));
 sg13g2_xnor2_1 _07832_ (.Y(_02365_),
    .A(_02355_),
    .B(_02364_));
 sg13g2_nand2b_1 _07833_ (.Y(_02366_),
    .B(_02349_),
    .A_N(_02365_));
 sg13g2_xor2_1 _07834_ (.B(_02365_),
    .A(_02349_),
    .X(_02367_));
 sg13g2_xor2_1 _07835_ (.B(_02367_),
    .A(_02348_),
    .X(_02368_));
 sg13g2_o21ai_1 _07836_ (.B1(_02280_),
    .Y(_02369_),
    .A1(_02267_),
    .A2(_02281_));
 sg13g2_and2_1 _07837_ (.A(_02275_),
    .B(_02277_),
    .X(_02370_));
 sg13g2_nand2_1 _07838_ (.Y(_02371_),
    .A(_02275_),
    .B(_02277_));
 sg13g2_nand2b_1 _07839_ (.Y(_02372_),
    .B(_02273_),
    .A_N(_02271_));
 sg13g2_o21ai_1 _07840_ (.B1(_02299_),
    .Y(_02373_),
    .A1(_02297_),
    .A2(_02300_));
 sg13g2_nand2_1 _07841_ (.Y(_02374_),
    .A(net1471),
    .B(net1175));
 sg13g2_and4_1 _07842_ (.A(net1360),
    .B(net1353),
    .C(net1169),
    .D(net1163),
    .X(_02375_));
 sg13g2_a22oi_1 _07843_ (.Y(_02376_),
    .B1(net1163),
    .B2(net1360),
    .A2(net1169),
    .A1(net1353));
 sg13g2_or3_1 _07844_ (.A(_02374_),
    .B(_02375_),
    .C(_02376_),
    .X(_02377_));
 sg13g2_o21ai_1 _07845_ (.B1(_02374_),
    .Y(_02378_),
    .A1(_02375_),
    .A2(_02376_));
 sg13g2_nand3_1 _07846_ (.B(_02377_),
    .C(_02378_),
    .A(_02373_),
    .Y(_02379_));
 sg13g2_a21o_1 _07847_ (.A2(_02378_),
    .A1(_02377_),
    .B1(_02373_),
    .X(_02380_));
 sg13g2_nand3_1 _07848_ (.B(_02379_),
    .C(_02380_),
    .A(_02372_),
    .Y(_02381_));
 sg13g2_a21o_1 _07849_ (.A2(_02380_),
    .A1(_02379_),
    .B1(_02372_),
    .X(_02382_));
 sg13g2_nand3_1 _07850_ (.B(_02381_),
    .C(_02382_),
    .A(_02304_),
    .Y(_02383_));
 sg13g2_a21oi_1 _07851_ (.A1(_02381_),
    .A2(_02382_),
    .Y(_02384_),
    .B1(_02304_));
 sg13g2_a21o_1 _07852_ (.A2(_02382_),
    .A1(_02381_),
    .B1(_02304_),
    .X(_02385_));
 sg13g2_nand3_1 _07853_ (.B(_02383_),
    .C(_02385_),
    .A(_02371_),
    .Y(_02386_));
 sg13g2_a21o_1 _07854_ (.A2(_02385_),
    .A1(_02383_),
    .B1(_02371_),
    .X(_02387_));
 sg13g2_and3_1 _07855_ (.X(_02388_),
    .A(_02369_),
    .B(_02386_),
    .C(_02387_));
 sg13g2_nand3_1 _07856_ (.B(_02386_),
    .C(_02387_),
    .A(_02369_),
    .Y(_02389_));
 sg13g2_a21o_1 _07857_ (.A2(_02387_),
    .A1(_02386_),
    .B1(_02369_),
    .X(_02390_));
 sg13g2_and3_1 _07858_ (.X(_02391_),
    .A(_02368_),
    .B(_02389_),
    .C(_02390_));
 sg13g2_a21oi_1 _07859_ (.A1(_02389_),
    .A2(_02390_),
    .Y(_02392_),
    .B1(_02368_));
 sg13g2_a21oi_1 _07860_ (.A1(_02266_),
    .A2(_02287_),
    .Y(_02393_),
    .B1(_02285_));
 sg13g2_nor3_1 _07861_ (.A(_02391_),
    .B(_02392_),
    .C(_02393_),
    .Y(_02394_));
 sg13g2_o21ai_1 _07862_ (.B1(_02393_),
    .Y(_02395_),
    .A1(_02391_),
    .A2(_02392_));
 sg13g2_nand2b_1 _07863_ (.Y(_02396_),
    .B(_02395_),
    .A_N(_02394_));
 sg13g2_nand2_1 _07864_ (.Y(_02397_),
    .A(net1430),
    .B(net1219));
 sg13g2_nand2_1 _07865_ (.Y(_02398_),
    .A(net1366),
    .B(net1159));
 sg13g2_and4_1 _07866_ (.A(net1380),
    .B(net1373),
    .C(net1153),
    .D(net1147),
    .X(_02399_));
 sg13g2_nand4_1 _07867_ (.B(net1373),
    .C(net1153),
    .A(net1380),
    .Y(_02400_),
    .D(net1147));
 sg13g2_a22oi_1 _07868_ (.Y(_02401_),
    .B1(net1148),
    .B2(net1380),
    .A2(net1153),
    .A1(net1373));
 sg13g2_nor3_1 _07869_ (.A(_02398_),
    .B(_02399_),
    .C(_02401_),
    .Y(_02402_));
 sg13g2_o21ai_1 _07870_ (.B1(_02398_),
    .Y(_02403_),
    .A1(_02399_),
    .A2(_02401_));
 sg13g2_nor2b_1 _07871_ (.A(_02402_),
    .B_N(_02403_),
    .Y(_02404_));
 sg13g2_nand2_1 _07872_ (.Y(_02405_),
    .A(net1387),
    .B(net1349));
 sg13g2_and4_1 _07873_ (.A(net1404),
    .B(net1396),
    .C(net1344),
    .D(net1339),
    .X(_02406_));
 sg13g2_nand4_1 _07874_ (.B(net1396),
    .C(net1344),
    .A(net1404),
    .Y(_02407_),
    .D(net1339));
 sg13g2_a22oi_1 _07875_ (.Y(_02408_),
    .B1(net1339),
    .B2(net1404),
    .A2(net1344),
    .A1(net1396));
 sg13g2_or3_1 _07876_ (.A(_02405_),
    .B(_02406_),
    .C(_02408_),
    .X(_02409_));
 sg13g2_o21ai_1 _07877_ (.B1(_02405_),
    .Y(_02410_),
    .A1(_02406_),
    .A2(_02408_));
 sg13g2_and3_1 _07878_ (.X(_02411_),
    .A(_02295_),
    .B(_02409_),
    .C(_02410_));
 sg13g2_a21o_1 _07879_ (.A2(_02410_),
    .A1(_02409_),
    .B1(_02295_),
    .X(_02412_));
 sg13g2_nor2b_1 _07880_ (.A(_02411_),
    .B_N(_02412_),
    .Y(_02413_));
 sg13g2_xnor2_1 _07881_ (.Y(_02414_),
    .A(_02404_),
    .B(_02413_));
 sg13g2_nor2_1 _07882_ (.A(_02397_),
    .B(_02414_),
    .Y(_02415_));
 sg13g2_xor2_1 _07883_ (.B(_02414_),
    .A(_02397_),
    .X(_02416_));
 sg13g2_nand2_1 _07884_ (.Y(_02417_),
    .A(_02306_),
    .B(_02416_));
 sg13g2_xnor2_1 _07885_ (.Y(_02418_),
    .A(_02306_),
    .B(_02416_));
 sg13g2_xor2_1 _07886_ (.B(_02418_),
    .A(_02396_),
    .X(_02419_));
 sg13g2_and2_1 _07887_ (.A(_02337_),
    .B(_02419_),
    .X(_02420_));
 sg13g2_or2_1 _07888_ (.X(_02421_),
    .B(_02419_),
    .A(_02337_));
 sg13g2_xnor2_1 _07889_ (.Y(_02422_),
    .A(_02337_),
    .B(_02419_));
 sg13g2_xnor2_1 _07890_ (.Y(_02423_),
    .A(_02336_),
    .B(_02422_));
 sg13g2_nand2_1 _07891_ (.Y(_02424_),
    .A(_02331_),
    .B(_02423_));
 sg13g2_xnor2_1 _07892_ (.Y(_02425_),
    .A(_02331_),
    .B(_02423_));
 sg13g2_xnor2_1 _07893_ (.Y(_02426_),
    .A(_02330_),
    .B(_02425_));
 sg13g2_a21oi_1 _07894_ (.A1(_02226_),
    .A2(_02319_),
    .Y(_02427_),
    .B1(_02318_));
 sg13g2_or2_1 _07895_ (.X(_02428_),
    .B(_02427_),
    .A(_02426_));
 sg13g2_and2_1 _07896_ (.A(_02426_),
    .B(_02427_),
    .X(_02429_));
 sg13g2_xor2_1 _07897_ (.B(_02427_),
    .A(_02426_),
    .X(_02430_));
 sg13g2_a21oi_1 _07898_ (.A1(_02216_),
    .A2(_02324_),
    .Y(_02431_),
    .B1(_02323_));
 sg13g2_a21oi_1 _07899_ (.A1(_02223_),
    .A2(_02325_),
    .Y(_02432_),
    .B1(_02431_));
 sg13g2_xnor2_1 _07900_ (.Y(_02433_),
    .A(_02430_),
    .B(_02432_));
 sg13g2_o21ai_1 _07901_ (.B1(net1518),
    .Y(_02434_),
    .A1(net1143),
    .A2(_02433_));
 sg13g2_a21oi_1 _07902_ (.A1(net1143),
    .A2(_04778_),
    .Y(_00230_),
    .B1(_02434_));
 sg13g2_o21ai_1 _07903_ (.B1(_02428_),
    .Y(_02435_),
    .A1(_02429_),
    .A2(_02432_));
 sg13g2_o21ai_1 _07904_ (.B1(_02424_),
    .Y(_02436_),
    .A1(_02330_),
    .A2(_02425_));
 sg13g2_a21oi_1 _07905_ (.A1(_02291_),
    .A2(_02333_),
    .Y(_02437_),
    .B1(_02335_));
 sg13g2_a21oi_1 _07906_ (.A1(_02336_),
    .A2(_02421_),
    .Y(_02438_),
    .B1(_02420_));
 sg13g2_a21o_1 _07907_ (.A2(_02345_),
    .A1(_02339_),
    .B1(_02347_),
    .X(_02439_));
 sg13g2_o21ai_1 _07908_ (.B1(_02366_),
    .Y(_02440_),
    .A1(_02348_),
    .A2(_02367_));
 sg13g2_and2_1 _07909_ (.A(_02394_),
    .B(_02440_),
    .X(_02441_));
 sg13g2_xor2_1 _07910_ (.B(_02440_),
    .A(_02394_),
    .X(_02442_));
 sg13g2_xor2_1 _07911_ (.B(_02442_),
    .A(_02439_),
    .X(_02443_));
 sg13g2_o21ai_1 _07912_ (.B1(_02417_),
    .Y(_02444_),
    .A1(_02396_),
    .A2(_02418_));
 sg13g2_o21ai_1 _07913_ (.B1(_02343_),
    .Y(_02445_),
    .A1(_02340_),
    .A2(_02344_));
 sg13g2_o21ai_1 _07914_ (.B1(_02354_),
    .Y(_02446_),
    .A1(_02248_),
    .A2(_02352_));
 sg13g2_nand2_1 _07915_ (.Y(_02447_),
    .A(net1422),
    .B(net1224));
 sg13g2_nand2_1 _07916_ (.Y(_02448_),
    .A(net1430),
    .B(net1210));
 sg13g2_nand2_1 _07917_ (.Y(_02449_),
    .A(net1430),
    .B(net1216));
 sg13g2_or2_1 _07918_ (.X(_02450_),
    .B(_02448_),
    .A(_02342_));
 sg13g2_xnor2_1 _07919_ (.Y(_02451_),
    .A(_02341_),
    .B(_02449_));
 sg13g2_xor2_1 _07920_ (.B(_02451_),
    .A(_02447_),
    .X(_02452_));
 sg13g2_xnor2_1 _07921_ (.Y(_02453_),
    .A(_02446_),
    .B(_02452_));
 sg13g2_nor2b_1 _07922_ (.A(_02453_),
    .B_N(_02445_),
    .Y(_02454_));
 sg13g2_xor2_1 _07923_ (.B(_02453_),
    .A(_02445_),
    .X(_02455_));
 sg13g2_o21ai_1 _07924_ (.B1(_02363_),
    .Y(_02456_),
    .A1(_02355_),
    .A2(_02364_));
 sg13g2_nand2_1 _07925_ (.Y(_02457_),
    .A(net1439),
    .B(net1205));
 sg13g2_nand2_1 _07926_ (.Y(_02458_),
    .A(net1444),
    .B(net1196));
 sg13g2_nand2_1 _07927_ (.Y(_02459_),
    .A(net1444),
    .B(net1202));
 sg13g2_xor2_1 _07928_ (.B(_02459_),
    .A(_02351_),
    .X(_02460_));
 sg13g2_nand2b_1 _07929_ (.Y(_02461_),
    .B(_02460_),
    .A_N(_02457_));
 sg13g2_xor2_1 _07930_ (.B(_02460_),
    .A(_02457_),
    .X(_02462_));
 sg13g2_o21ai_1 _07931_ (.B1(_02359_),
    .Y(_02463_),
    .A1(_02357_),
    .A2(_02360_));
 sg13g2_nand2_1 _07932_ (.Y(_02464_),
    .A(net1454),
    .B(net1192));
 sg13g2_nand2_1 _07933_ (.Y(_02465_),
    .A(net1457),
    .B(net1183));
 sg13g2_and4_1 _07934_ (.A(net1462),
    .B(net1457),
    .C(net1188),
    .D(net1182),
    .X(_02466_));
 sg13g2_a22oi_1 _07935_ (.Y(_02467_),
    .B1(net1182),
    .B2(net1462),
    .A2(net1188),
    .A1(net1458));
 sg13g2_nor3_1 _07936_ (.A(_02464_),
    .B(_02466_),
    .C(_02467_),
    .Y(_02468_));
 sg13g2_o21ai_1 _07937_ (.B1(_02464_),
    .Y(_02469_),
    .A1(_02466_),
    .A2(_02467_));
 sg13g2_nor2b_1 _07938_ (.A(_02468_),
    .B_N(_02469_),
    .Y(_02470_));
 sg13g2_nand2_1 _07939_ (.Y(_02471_),
    .A(_02463_),
    .B(_02470_));
 sg13g2_xnor2_1 _07940_ (.Y(_02472_),
    .A(_02463_),
    .B(_02470_));
 sg13g2_xnor2_1 _07941_ (.Y(_02473_),
    .A(_02462_),
    .B(_02472_));
 sg13g2_nand2b_1 _07942_ (.Y(_02474_),
    .B(_02456_),
    .A_N(_02473_));
 sg13g2_xor2_1 _07943_ (.B(_02473_),
    .A(_02456_),
    .X(_02475_));
 sg13g2_xor2_1 _07944_ (.B(_02475_),
    .A(_02455_),
    .X(_02476_));
 sg13g2_o21ai_1 _07945_ (.B1(_02383_),
    .Y(_02477_),
    .A1(_02370_),
    .A2(_02384_));
 sg13g2_and2_1 _07946_ (.A(_02379_),
    .B(_02381_),
    .X(_02478_));
 sg13g2_a21o_1 _07947_ (.A2(_02412_),
    .A1(_02404_),
    .B1(_02411_),
    .X(_02479_));
 sg13g2_nand2b_1 _07948_ (.Y(_02480_),
    .B(_02377_),
    .A_N(_02375_));
 sg13g2_o21ai_1 _07949_ (.B1(_02400_),
    .Y(_02481_),
    .A1(_02398_),
    .A2(_02401_));
 sg13g2_nand2_1 _07950_ (.Y(_02482_),
    .A(net1467),
    .B(net1176));
 sg13g2_and4_1 _07951_ (.A(net1353),
    .B(net1471),
    .C(net1169),
    .D(net1163),
    .X(_02483_));
 sg13g2_a22oi_1 _07952_ (.Y(_02484_),
    .B1(net1163),
    .B2(net1353),
    .A2(net1169),
    .A1(net1471));
 sg13g2_or3_1 _07953_ (.A(_02482_),
    .B(_02483_),
    .C(_02484_),
    .X(_02485_));
 sg13g2_o21ai_1 _07954_ (.B1(_02482_),
    .Y(_02486_),
    .A1(_02483_),
    .A2(_02484_));
 sg13g2_nand3_1 _07955_ (.B(_02485_),
    .C(_02486_),
    .A(_02481_),
    .Y(_02487_));
 sg13g2_a21o_1 _07956_ (.A2(_02486_),
    .A1(_02485_),
    .B1(_02481_),
    .X(_02488_));
 sg13g2_nand3_1 _07957_ (.B(_02487_),
    .C(_02488_),
    .A(_02480_),
    .Y(_02489_));
 sg13g2_a21o_1 _07958_ (.A2(_02488_),
    .A1(_02487_),
    .B1(_02480_),
    .X(_02490_));
 sg13g2_and3_2 _07959_ (.X(_02491_),
    .A(_02479_),
    .B(_02489_),
    .C(_02490_));
 sg13g2_a21oi_1 _07960_ (.A1(_02489_),
    .A2(_02490_),
    .Y(_02492_),
    .B1(_02479_));
 sg13g2_or3_1 _07961_ (.A(_02478_),
    .B(_02491_),
    .C(_02492_),
    .X(_02493_));
 sg13g2_o21ai_1 _07962_ (.B1(_02478_),
    .Y(_02494_),
    .A1(_02491_),
    .A2(_02492_));
 sg13g2_nand3_1 _07963_ (.B(_02493_),
    .C(_02494_),
    .A(_02477_),
    .Y(_02495_));
 sg13g2_a21o_1 _07964_ (.A2(_02494_),
    .A1(_02493_),
    .B1(_02477_),
    .X(_02496_));
 sg13g2_and3_1 _07965_ (.X(_02497_),
    .A(_02476_),
    .B(_02495_),
    .C(_02496_));
 sg13g2_nand3_1 _07966_ (.B(_02495_),
    .C(_02496_),
    .A(_02476_),
    .Y(_02498_));
 sg13g2_a21oi_1 _07967_ (.A1(_02495_),
    .A2(_02496_),
    .Y(_02499_),
    .B1(_02476_));
 sg13g2_a21oi_1 _07968_ (.A1(_02368_),
    .A2(_02390_),
    .Y(_02500_),
    .B1(_02388_));
 sg13g2_nor3_1 _07969_ (.A(_02497_),
    .B(_02499_),
    .C(_02500_),
    .Y(_02501_));
 sg13g2_o21ai_1 _07970_ (.B1(_02500_),
    .Y(_02502_),
    .A1(_02497_),
    .A2(_02499_));
 sg13g2_nand2b_1 _07971_ (.Y(_02503_),
    .B(_02502_),
    .A_N(_02501_));
 sg13g2_nand2_1 _07972_ (.Y(_02504_),
    .A(net1426),
    .B(net1219));
 sg13g2_nand2_2 _07973_ (.Y(_02505_),
    .A(net1405),
    .B(net1336));
 sg13g2_nand2_1 _07974_ (.Y(_02506_),
    .A(net1360),
    .B(net1159));
 sg13g2_nand2_1 _07975_ (.Y(_02507_),
    .A(net1368),
    .B(net1148));
 sg13g2_and4_1 _07976_ (.A(net1373),
    .B(net1366),
    .C(net1153),
    .D(net1147),
    .X(_02508_));
 sg13g2_nand4_1 _07977_ (.B(net1366),
    .C(net1153),
    .A(net1373),
    .Y(_02509_),
    .D(net1147));
 sg13g2_a22oi_1 _07978_ (.Y(_02510_),
    .B1(net1147),
    .B2(net1373),
    .A2(net1153),
    .A1(net1366));
 sg13g2_nor3_1 _07979_ (.A(_02506_),
    .B(_02508_),
    .C(_02510_),
    .Y(_02511_));
 sg13g2_o21ai_1 _07980_ (.B1(_02506_),
    .Y(_02512_),
    .A1(_02508_),
    .A2(_02510_));
 sg13g2_nor2b_1 _07981_ (.A(_02511_),
    .B_N(_02512_),
    .Y(_02513_));
 sg13g2_o21ai_1 _07982_ (.B1(_02407_),
    .Y(_02514_),
    .A1(_02405_),
    .A2(_02408_));
 sg13g2_nand2_1 _07983_ (.Y(_02515_),
    .A(net1380),
    .B(net1349));
 sg13g2_and4_1 _07984_ (.A(net1396),
    .B(net1387),
    .C(net1344),
    .D(net1340),
    .X(_02516_));
 sg13g2_nand4_1 _07985_ (.B(net1387),
    .C(net1344),
    .A(net1396),
    .Y(_02517_),
    .D(net1339));
 sg13g2_a22oi_1 _07986_ (.Y(_02518_),
    .B1(net1339),
    .B2(net1396),
    .A2(net1344),
    .A1(net1387));
 sg13g2_or3_1 _07987_ (.A(_02515_),
    .B(_02516_),
    .C(_02518_),
    .X(_02519_));
 sg13g2_o21ai_1 _07988_ (.B1(_02515_),
    .Y(_02520_),
    .A1(_02516_),
    .A2(_02518_));
 sg13g2_and3_1 _07989_ (.X(_02521_),
    .A(_02514_),
    .B(_02519_),
    .C(_02520_));
 sg13g2_a21o_1 _07990_ (.A2(_02520_),
    .A1(_02519_),
    .B1(_02514_),
    .X(_02522_));
 sg13g2_nand2b_1 _07991_ (.Y(_02523_),
    .B(_02522_),
    .A_N(_02521_));
 sg13g2_xor2_1 _07992_ (.B(_02523_),
    .A(_02513_),
    .X(_02524_));
 sg13g2_nor2_1 _07993_ (.A(_02505_),
    .B(_02524_),
    .Y(_02525_));
 sg13g2_xor2_1 _07994_ (.B(_02524_),
    .A(_02505_),
    .X(_02526_));
 sg13g2_nor2b_1 _07995_ (.A(_02504_),
    .B_N(_02526_),
    .Y(_02527_));
 sg13g2_xnor2_1 _07996_ (.Y(_02528_),
    .A(_02504_),
    .B(_02526_));
 sg13g2_nand2_1 _07997_ (.Y(_02529_),
    .A(_02415_),
    .B(_02528_));
 sg13g2_xnor2_1 _07998_ (.Y(_02530_),
    .A(_02415_),
    .B(_02528_));
 sg13g2_xor2_1 _07999_ (.B(_02530_),
    .A(_02503_),
    .X(_02531_));
 sg13g2_and2_1 _08000_ (.A(_02444_),
    .B(_02531_),
    .X(_02532_));
 sg13g2_xor2_1 _08001_ (.B(_02531_),
    .A(_02444_),
    .X(_02533_));
 sg13g2_xor2_1 _08002_ (.B(_02533_),
    .A(_02443_),
    .X(_02534_));
 sg13g2_nand2b_1 _08003_ (.Y(_02535_),
    .B(_02534_),
    .A_N(_02438_));
 sg13g2_xnor2_1 _08004_ (.Y(_02536_),
    .A(_02438_),
    .B(_02534_));
 sg13g2_nand2b_1 _08005_ (.Y(_02537_),
    .B(_02536_),
    .A_N(_02437_));
 sg13g2_xnor2_1 _08006_ (.Y(_02538_),
    .A(_02437_),
    .B(_02536_));
 sg13g2_nor2_1 _08007_ (.A(_02436_),
    .B(_02538_),
    .Y(_02539_));
 sg13g2_xor2_1 _08008_ (.B(_02538_),
    .A(_02436_),
    .X(_02540_));
 sg13g2_xnor2_1 _08009_ (.Y(_02541_),
    .A(_02435_),
    .B(_02540_));
 sg13g2_o21ai_1 _08010_ (.B1(net1518),
    .Y(_02542_),
    .A1(net1297),
    .A2(net297));
 sg13g2_a21oi_1 _08011_ (.A1(net1297),
    .A2(_02541_),
    .Y(_00231_),
    .B1(_02542_));
 sg13g2_a21oi_1 _08012_ (.A1(_02439_),
    .A2(_02442_),
    .Y(_02543_),
    .B1(_02441_));
 sg13g2_a21oi_1 _08013_ (.A1(_02443_),
    .A2(_02533_),
    .Y(_02544_),
    .B1(_02532_));
 sg13g2_a21o_1 _08014_ (.A2(_02452_),
    .A1(_02446_),
    .B1(_02454_),
    .X(_02545_));
 sg13g2_o21ai_1 _08015_ (.B1(_02474_),
    .Y(_02546_),
    .A1(_02455_),
    .A2(_02475_));
 sg13g2_and2_1 _08016_ (.A(_02501_),
    .B(_02546_),
    .X(_02547_));
 sg13g2_xor2_1 _08017_ (.B(_02546_),
    .A(_02501_),
    .X(_02548_));
 sg13g2_xnor2_1 _08018_ (.Y(_02549_),
    .A(_02545_),
    .B(_02548_));
 sg13g2_o21ai_1 _08019_ (.B1(_02529_),
    .Y(_02550_),
    .A1(_02503_),
    .A2(_02530_));
 sg13g2_o21ai_1 _08020_ (.B1(_02450_),
    .Y(_02551_),
    .A1(_02447_),
    .A2(_02451_));
 sg13g2_o21ai_1 _08021_ (.B1(_02461_),
    .Y(_02552_),
    .A1(_02351_),
    .A2(_02459_));
 sg13g2_nand2_1 _08022_ (.Y(_02553_),
    .A(net1420),
    .B(net1224));
 sg13g2_nand2_1 _08023_ (.Y(_02554_),
    .A(net1426),
    .B(net1210));
 sg13g2_nand2_1 _08024_ (.Y(_02555_),
    .A(net1427),
    .B(net1216));
 sg13g2_or2_1 _08025_ (.X(_02556_),
    .B(_02554_),
    .A(_02449_));
 sg13g2_xnor2_1 _08026_ (.Y(_02557_),
    .A(_02448_),
    .B(_02555_));
 sg13g2_xor2_1 _08027_ (.B(_02557_),
    .A(_02553_),
    .X(_02558_));
 sg13g2_xnor2_1 _08028_ (.Y(_02559_),
    .A(_02552_),
    .B(_02558_));
 sg13g2_nor2b_1 _08029_ (.A(_02559_),
    .B_N(_02551_),
    .Y(_02560_));
 sg13g2_xor2_1 _08030_ (.B(_02559_),
    .A(_02551_),
    .X(_02561_));
 sg13g2_o21ai_1 _08031_ (.B1(_02471_),
    .Y(_02562_),
    .A1(_02462_),
    .A2(_02472_));
 sg13g2_nand2_1 _08032_ (.Y(_02563_),
    .A(net1435),
    .B(net1205));
 sg13g2_nand2_1 _08033_ (.Y(_02564_),
    .A(net1438),
    .B(net1198));
 sg13g2_nand2_1 _08034_ (.Y(_02565_),
    .A(net1439),
    .B(net1201));
 sg13g2_xor2_1 _08035_ (.B(_02565_),
    .A(_02458_),
    .X(_02566_));
 sg13g2_nand2b_1 _08036_ (.Y(_02567_),
    .B(_02566_),
    .A_N(_02563_));
 sg13g2_xor2_1 _08037_ (.B(_02566_),
    .A(_02563_),
    .X(_02568_));
 sg13g2_or2_1 _08038_ (.X(_02569_),
    .B(_02468_),
    .A(_02466_));
 sg13g2_nand2_1 _08039_ (.Y(_02570_),
    .A(net1448),
    .B(net1191));
 sg13g2_nand2_1 _08040_ (.Y(_02571_),
    .A(net1453),
    .B(net1189));
 sg13g2_or2_1 _08041_ (.X(_02572_),
    .B(_02571_),
    .A(_02465_));
 sg13g2_and2_1 _08042_ (.A(_02465_),
    .B(_02571_),
    .X(_02573_));
 sg13g2_xor2_1 _08043_ (.B(_02571_),
    .A(_02465_),
    .X(_02574_));
 sg13g2_xnor2_1 _08044_ (.Y(_02575_),
    .A(_02570_),
    .B(_02574_));
 sg13g2_nand2_1 _08045_ (.Y(_02576_),
    .A(_02569_),
    .B(_02575_));
 sg13g2_xnor2_1 _08046_ (.Y(_02577_),
    .A(_02569_),
    .B(_02575_));
 sg13g2_xnor2_1 _08047_ (.Y(_02578_),
    .A(_02568_),
    .B(_02577_));
 sg13g2_nand2b_1 _08048_ (.Y(_02579_),
    .B(_02562_),
    .A_N(_02578_));
 sg13g2_xor2_1 _08049_ (.B(_02578_),
    .A(_02562_),
    .X(_02580_));
 sg13g2_xor2_1 _08050_ (.B(_02580_),
    .A(_02561_),
    .X(_02581_));
 sg13g2_nor2b_2 _08051_ (.A(_02491_),
    .B_N(_02493_),
    .Y(_02582_));
 sg13g2_and2_1 _08052_ (.A(_02487_),
    .B(_02489_),
    .X(_02583_));
 sg13g2_a21o_1 _08053_ (.A2(_02522_),
    .A1(_02513_),
    .B1(_02521_),
    .X(_02584_));
 sg13g2_nand2b_1 _08054_ (.Y(_02585_),
    .B(_02485_),
    .A_N(_02483_));
 sg13g2_o21ai_1 _08055_ (.B1(_02509_),
    .Y(_02586_),
    .A1(_02506_),
    .A2(_02510_));
 sg13g2_nand2_1 _08056_ (.Y(_02587_),
    .A(net1462),
    .B(net1175));
 sg13g2_and4_1 _08057_ (.A(net1471),
    .B(net1467),
    .C(net1169),
    .D(net1163),
    .X(_02588_));
 sg13g2_a22oi_1 _08058_ (.Y(_02589_),
    .B1(net1163),
    .B2(net1471),
    .A2(net1169),
    .A1(net1467));
 sg13g2_or3_1 _08059_ (.A(_02587_),
    .B(_02588_),
    .C(_02589_),
    .X(_02590_));
 sg13g2_o21ai_1 _08060_ (.B1(_02587_),
    .Y(_02591_),
    .A1(_02588_),
    .A2(_02589_));
 sg13g2_nand3_1 _08061_ (.B(_02590_),
    .C(_02591_),
    .A(_02586_),
    .Y(_02592_));
 sg13g2_a21o_1 _08062_ (.A2(_02591_),
    .A1(_02590_),
    .B1(_02586_),
    .X(_02593_));
 sg13g2_nand3_1 _08063_ (.B(_02592_),
    .C(_02593_),
    .A(_02585_),
    .Y(_02594_));
 sg13g2_a21o_1 _08064_ (.A2(_02593_),
    .A1(_02592_),
    .B1(_02585_),
    .X(_02595_));
 sg13g2_and3_1 _08065_ (.X(_02596_),
    .A(_02584_),
    .B(_02594_),
    .C(_02595_));
 sg13g2_nand3_1 _08066_ (.B(_02594_),
    .C(_02595_),
    .A(_02584_),
    .Y(_02597_));
 sg13g2_a21oi_1 _08067_ (.A1(_02594_),
    .A2(_02595_),
    .Y(_02598_),
    .B1(_02584_));
 sg13g2_nor2_1 _08068_ (.A(_02596_),
    .B(_02598_),
    .Y(_02599_));
 sg13g2_xor2_1 _08069_ (.B(_02599_),
    .A(_02583_),
    .X(_02600_));
 sg13g2_nor2_1 _08070_ (.A(_02582_),
    .B(_02600_),
    .Y(_02601_));
 sg13g2_nand2_1 _08071_ (.Y(_02602_),
    .A(_02582_),
    .B(_02600_));
 sg13g2_xor2_1 _08072_ (.B(_02600_),
    .A(_02582_),
    .X(_02603_));
 sg13g2_xnor2_1 _08073_ (.Y(_02604_),
    .A(_02581_),
    .B(_02603_));
 sg13g2_and2_1 _08074_ (.A(_02495_),
    .B(_02498_),
    .X(_02605_));
 sg13g2_nor2_1 _08075_ (.A(_02604_),
    .B(_02605_),
    .Y(_02606_));
 sg13g2_xnor2_1 _08076_ (.Y(_02607_),
    .A(_02604_),
    .B(_02605_));
 sg13g2_nand2_2 _08077_ (.Y(_02608_),
    .A(net1422),
    .B(net1219));
 sg13g2_a22oi_1 _08078_ (.Y(_02609_),
    .B1(net1333),
    .B2(net1405),
    .A2(net1336),
    .A1(net1397));
 sg13g2_nand2_2 _08079_ (.Y(_02610_),
    .A(net1402),
    .B(net1333));
 sg13g2_or2_1 _08080_ (.X(_02611_),
    .B(_02610_),
    .A(_02505_));
 sg13g2_nand2b_2 _08081_ (.Y(_02612_),
    .B(_02611_),
    .A_N(_02609_));
 sg13g2_nand2_1 _08082_ (.Y(_02613_),
    .A(net1353),
    .B(net1159));
 sg13g2_nand2_1 _08083_ (.Y(_02614_),
    .A(net1361),
    .B(net1150));
 sg13g2_nand2_1 _08084_ (.Y(_02615_),
    .A(net1361),
    .B(net1154));
 sg13g2_nand4_1 _08085_ (.B(net1360),
    .C(net1154),
    .A(net1366),
    .Y(_02616_),
    .D(net1148));
 sg13g2_a22oi_1 _08086_ (.Y(_02617_),
    .B1(net1148),
    .B2(net1366),
    .A2(net1154),
    .A1(net1360));
 sg13g2_xor2_1 _08087_ (.B(_02615_),
    .A(_02507_),
    .X(_02618_));
 sg13g2_xnor2_1 _08088_ (.Y(_02619_),
    .A(_02613_),
    .B(_02618_));
 sg13g2_o21ai_1 _08089_ (.B1(_02517_),
    .Y(_02620_),
    .A1(_02515_),
    .A2(_02518_));
 sg13g2_nand2_1 _08090_ (.Y(_02621_),
    .A(net1373),
    .B(net1349));
 sg13g2_and4_1 _08091_ (.A(net1389),
    .B(net1382),
    .C(net1344),
    .D(net1339),
    .X(_02622_));
 sg13g2_a22oi_1 _08092_ (.Y(_02623_),
    .B1(net1340),
    .B2(net1389),
    .A2(net1344),
    .A1(net1382));
 sg13g2_or3_1 _08093_ (.A(_02621_),
    .B(_02622_),
    .C(_02623_),
    .X(_02624_));
 sg13g2_o21ai_1 _08094_ (.B1(_02621_),
    .Y(_02625_),
    .A1(_02622_),
    .A2(_02623_));
 sg13g2_and3_1 _08095_ (.X(_02626_),
    .A(_02620_),
    .B(_02624_),
    .C(_02625_));
 sg13g2_a21o_1 _08096_ (.A2(_02625_),
    .A1(_02624_),
    .B1(_02620_),
    .X(_02627_));
 sg13g2_nand2b_1 _08097_ (.Y(_02628_),
    .B(_02627_),
    .A_N(_02626_));
 sg13g2_xor2_1 _08098_ (.B(_02628_),
    .A(_02619_),
    .X(_02629_));
 sg13g2_or2_1 _08099_ (.X(_02630_),
    .B(_02629_),
    .A(_02612_));
 sg13g2_xor2_1 _08100_ (.B(_02629_),
    .A(_02612_),
    .X(_02631_));
 sg13g2_nand2_1 _08101_ (.Y(_02632_),
    .A(_02525_),
    .B(_02631_));
 sg13g2_xnor2_1 _08102_ (.Y(_02633_),
    .A(_02525_),
    .B(_02631_));
 sg13g2_nor2_1 _08103_ (.A(_02608_),
    .B(_02633_),
    .Y(_02634_));
 sg13g2_xnor2_1 _08104_ (.Y(_02635_),
    .A(_02608_),
    .B(_02633_));
 sg13g2_inv_1 _08105_ (.Y(_02636_),
    .A(_02635_));
 sg13g2_nand2_1 _08106_ (.Y(_02637_),
    .A(_02527_),
    .B(_02636_));
 sg13g2_xor2_1 _08107_ (.B(_02635_),
    .A(_02527_),
    .X(_02638_));
 sg13g2_xor2_1 _08108_ (.B(_02638_),
    .A(_02607_),
    .X(_02639_));
 sg13g2_nand2_1 _08109_ (.Y(_02640_),
    .A(_02550_),
    .B(_02639_));
 sg13g2_xnor2_1 _08110_ (.Y(_02641_),
    .A(_02550_),
    .B(_02639_));
 sg13g2_xor2_1 _08111_ (.B(_02641_),
    .A(_02549_),
    .X(_02642_));
 sg13g2_nand2b_1 _08112_ (.Y(_02643_),
    .B(_02642_),
    .A_N(_02544_));
 sg13g2_xnor2_1 _08113_ (.Y(_02644_),
    .A(_02544_),
    .B(_02642_));
 sg13g2_nand2b_1 _08114_ (.Y(_02645_),
    .B(_02644_),
    .A_N(_02543_));
 sg13g2_xor2_1 _08115_ (.B(_02644_),
    .A(_02543_),
    .X(_02646_));
 sg13g2_nand2_1 _08116_ (.Y(_02647_),
    .A(_02535_),
    .B(_02537_));
 sg13g2_nand2b_1 _08117_ (.Y(_02648_),
    .B(_02647_),
    .A_N(_02646_));
 sg13g2_inv_1 _08118_ (.Y(_02649_),
    .A(_02648_));
 sg13g2_xnor2_1 _08119_ (.Y(_02650_),
    .A(_02646_),
    .B(_02647_));
 sg13g2_and2_1 _08120_ (.A(_02430_),
    .B(_02540_),
    .X(_02651_));
 sg13g2_nand3_1 _08121_ (.B(_02325_),
    .C(_02651_),
    .A(_02223_),
    .Y(_02652_));
 sg13g2_nor2_1 _08122_ (.A(_02428_),
    .B(_02539_),
    .Y(_02653_));
 sg13g2_a221oi_1 _08123_ (.B2(_02431_),
    .C1(_02653_),
    .B1(_02651_),
    .A1(_02436_),
    .Y(_02654_),
    .A2(_02538_));
 sg13g2_nand2_1 _08124_ (.Y(_02655_),
    .A(_02652_),
    .B(_02654_));
 sg13g2_xnor2_1 _08125_ (.Y(_02656_),
    .A(_02650_),
    .B(_02655_));
 sg13g2_o21ai_1 _08126_ (.B1(net1518),
    .Y(_02657_),
    .A1(net1297),
    .A2(net304));
 sg13g2_a21oi_1 _08127_ (.A1(net1297),
    .A2(_02656_),
    .Y(_00232_),
    .B1(_02657_));
 sg13g2_nand2_1 _08128_ (.Y(_02658_),
    .A(_02643_),
    .B(_02645_));
 sg13g2_a21oi_1 _08129_ (.A1(_02545_),
    .A2(_02548_),
    .Y(_02659_),
    .B1(_02547_));
 sg13g2_o21ai_1 _08130_ (.B1(_02640_),
    .Y(_02660_),
    .A1(_02549_),
    .A2(_02641_));
 sg13g2_a21o_1 _08131_ (.A2(_02558_),
    .A1(_02552_),
    .B1(_02560_),
    .X(_02661_));
 sg13g2_o21ai_1 _08132_ (.B1(_02579_),
    .Y(_02662_),
    .A1(_02561_),
    .A2(_02580_));
 sg13g2_and2_1 _08133_ (.A(_02606_),
    .B(_02662_),
    .X(_02663_));
 sg13g2_xor2_1 _08134_ (.B(_02662_),
    .A(_02606_),
    .X(_02664_));
 sg13g2_xor2_1 _08135_ (.B(_02664_),
    .A(_02661_),
    .X(_02665_));
 sg13g2_o21ai_1 _08136_ (.B1(_02637_),
    .Y(_02666_),
    .A1(_02607_),
    .A2(_02638_));
 sg13g2_nand2_1 _08137_ (.Y(_02667_),
    .A(net1420),
    .B(net1219));
 sg13g2_nand2_1 _08138_ (.Y(_02668_),
    .A(net1394),
    .B(net1336));
 sg13g2_nand2_1 _08139_ (.Y(_02669_),
    .A(net1395),
    .B(net1330));
 sg13g2_nand2_1 _08140_ (.Y(_02670_),
    .A(net1405),
    .B(net1330));
 sg13g2_xor2_1 _08141_ (.B(_02670_),
    .A(_02610_),
    .X(_02671_));
 sg13g2_nand2b_1 _08142_ (.Y(_02672_),
    .B(_02671_),
    .A_N(_02668_));
 sg13g2_xnor2_1 _08143_ (.Y(_02673_),
    .A(_02668_),
    .B(_02671_));
 sg13g2_nand2b_1 _08144_ (.Y(_02674_),
    .B(_02673_),
    .A_N(_02611_));
 sg13g2_xnor2_1 _08145_ (.Y(_02675_),
    .A(_02611_),
    .B(_02673_));
 sg13g2_nand2_1 _08146_ (.Y(_02676_),
    .A(net1472),
    .B(net1159));
 sg13g2_nand2_1 _08147_ (.Y(_02677_),
    .A(net1354),
    .B(net1150));
 sg13g2_nand2_1 _08148_ (.Y(_02678_),
    .A(net1354),
    .B(net1156));
 sg13g2_or2_1 _08149_ (.X(_02679_),
    .B(_02677_),
    .A(_02615_));
 sg13g2_and2_1 _08150_ (.A(_02614_),
    .B(_02678_),
    .X(_02680_));
 sg13g2_xnor2_1 _08151_ (.Y(_02681_),
    .A(_02614_),
    .B(_02678_));
 sg13g2_xnor2_1 _08152_ (.Y(_02682_),
    .A(_02676_),
    .B(_02681_));
 sg13g2_nand2b_1 _08153_ (.Y(_02683_),
    .B(_02624_),
    .A_N(_02622_));
 sg13g2_and2_1 _08154_ (.A(net1368),
    .B(net1349),
    .X(_02684_));
 sg13g2_nand2_1 _08155_ (.Y(_02685_),
    .A(net1368),
    .B(net1349));
 sg13g2_nand2_1 _08156_ (.Y(_02686_),
    .A(net1375),
    .B(net1340));
 sg13g2_nand4_1 _08157_ (.B(net1375),
    .C(net1345),
    .A(net1382),
    .Y(_02687_),
    .D(net1339));
 sg13g2_inv_1 _08158_ (.Y(_02688_),
    .A(_02687_));
 sg13g2_a22oi_1 _08159_ (.Y(_02689_),
    .B1(net1339),
    .B2(net1382),
    .A2(net1345),
    .A1(net1375));
 sg13g2_nand3b_1 _08160_ (.B(_02684_),
    .C(_02687_),
    .Y(_02690_),
    .A_N(_02689_));
 sg13g2_o21ai_1 _08161_ (.B1(_02685_),
    .Y(_02691_),
    .A1(_02688_),
    .A2(_02689_));
 sg13g2_nand3_1 _08162_ (.B(_02690_),
    .C(_02691_),
    .A(_02683_),
    .Y(_02692_));
 sg13g2_a21oi_1 _08163_ (.A1(_02690_),
    .A2(_02691_),
    .Y(_02693_),
    .B1(_02683_));
 sg13g2_a21o_1 _08164_ (.A2(_02691_),
    .A1(_02690_),
    .B1(_02683_),
    .X(_02694_));
 sg13g2_nand2_1 _08165_ (.Y(_02695_),
    .A(_02692_),
    .B(_02694_));
 sg13g2_xor2_1 _08166_ (.B(_02695_),
    .A(_02682_),
    .X(_02696_));
 sg13g2_nand2_1 _08167_ (.Y(_02697_),
    .A(_02675_),
    .B(_02696_));
 sg13g2_xnor2_1 _08168_ (.Y(_02698_),
    .A(_02675_),
    .B(_02696_));
 sg13g2_nor2_1 _08169_ (.A(_02630_),
    .B(_02698_),
    .Y(_02699_));
 sg13g2_xnor2_1 _08170_ (.Y(_02700_),
    .A(_02630_),
    .B(_02698_));
 sg13g2_nor2_1 _08171_ (.A(_02667_),
    .B(_02700_),
    .Y(_02701_));
 sg13g2_xnor2_1 _08172_ (.Y(_02702_),
    .A(_02667_),
    .B(_02700_));
 sg13g2_or3_1 _08173_ (.A(_02608_),
    .B(_02633_),
    .C(_02702_),
    .X(_02703_));
 sg13g2_xnor2_1 _08174_ (.Y(_02704_),
    .A(_02634_),
    .B(_02702_));
 sg13g2_a21oi_1 _08175_ (.A1(_02581_),
    .A2(_02602_),
    .Y(_02705_),
    .B1(_02601_));
 sg13g2_o21ai_1 _08176_ (.B1(_02556_),
    .Y(_02706_),
    .A1(_02553_),
    .A2(_02557_));
 sg13g2_o21ai_1 _08177_ (.B1(_02567_),
    .Y(_02707_),
    .A1(_02458_),
    .A2(_02565_));
 sg13g2_nand2_1 _08178_ (.Y(_02708_),
    .A(net1416),
    .B(net1224));
 sg13g2_nand2_1 _08179_ (.Y(_02709_),
    .A(net1422),
    .B(net1210));
 sg13g2_nand2_1 _08180_ (.Y(_02710_),
    .A(net1423),
    .B(net1214));
 sg13g2_or2_1 _08181_ (.X(_02711_),
    .B(_02709_),
    .A(_02555_));
 sg13g2_xnor2_1 _08182_ (.Y(_02712_),
    .A(_02554_),
    .B(_02710_));
 sg13g2_xor2_1 _08183_ (.B(_02712_),
    .A(_02708_),
    .X(_02713_));
 sg13g2_xnor2_1 _08184_ (.Y(_02714_),
    .A(_02707_),
    .B(_02713_));
 sg13g2_nor2b_1 _08185_ (.A(_02714_),
    .B_N(_02706_),
    .Y(_02715_));
 sg13g2_xor2_1 _08186_ (.B(_02714_),
    .A(_02706_),
    .X(_02716_));
 sg13g2_o21ai_1 _08187_ (.B1(_02576_),
    .Y(_02717_),
    .A1(_02568_),
    .A2(_02577_));
 sg13g2_nand2_1 _08188_ (.Y(_02718_),
    .A(net1431),
    .B(net1205));
 sg13g2_nand2_1 _08189_ (.Y(_02719_),
    .A(net1434),
    .B(net1198));
 sg13g2_nand2_1 _08190_ (.Y(_02720_),
    .A(net1434),
    .B(net1201));
 sg13g2_xor2_1 _08191_ (.B(_02720_),
    .A(_02564_),
    .X(_02721_));
 sg13g2_nand2b_1 _08192_ (.Y(_02722_),
    .B(_02721_),
    .A_N(_02718_));
 sg13g2_xor2_1 _08193_ (.B(_02721_),
    .A(_02718_),
    .X(_02723_));
 sg13g2_o21ai_1 _08194_ (.B1(_02572_),
    .Y(_02724_),
    .A1(_02570_),
    .A2(_02573_));
 sg13g2_nand2_1 _08195_ (.Y(_02725_),
    .A(net1443),
    .B(net1191));
 sg13g2_nand2_1 _08196_ (.Y(_02726_),
    .A(net1448),
    .B(net1183));
 sg13g2_and4_1 _08197_ (.A(net1453),
    .B(net1448),
    .C(net1189),
    .D(net1183),
    .X(_02727_));
 sg13g2_a22oi_1 _08198_ (.Y(_02728_),
    .B1(net1183),
    .B2(net1453),
    .A2(net1189),
    .A1(net1448));
 sg13g2_nor3_1 _08199_ (.A(_02725_),
    .B(_02727_),
    .C(_02728_),
    .Y(_02729_));
 sg13g2_o21ai_1 _08200_ (.B1(_02725_),
    .Y(_02730_),
    .A1(_02727_),
    .A2(_02728_));
 sg13g2_nor2b_1 _08201_ (.A(_02729_),
    .B_N(_02730_),
    .Y(_02731_));
 sg13g2_nand2_1 _08202_ (.Y(_02732_),
    .A(_02724_),
    .B(_02731_));
 sg13g2_xnor2_1 _08203_ (.Y(_02733_),
    .A(_02724_),
    .B(_02731_));
 sg13g2_xor2_1 _08204_ (.B(_02733_),
    .A(_02723_),
    .X(_02734_));
 sg13g2_nand2_1 _08205_ (.Y(_02735_),
    .A(_02717_),
    .B(_02734_));
 sg13g2_xnor2_1 _08206_ (.Y(_02736_),
    .A(_02717_),
    .B(_02734_));
 sg13g2_xnor2_1 _08207_ (.Y(_02737_),
    .A(_02716_),
    .B(_02736_));
 sg13g2_o21ai_1 _08208_ (.B1(_02597_),
    .Y(_02738_),
    .A1(_02583_),
    .A2(_02598_));
 sg13g2_nand2_1 _08209_ (.Y(_02739_),
    .A(_02592_),
    .B(_02594_));
 sg13g2_a21o_1 _08210_ (.A2(_02627_),
    .A1(_02619_),
    .B1(_02626_),
    .X(_02740_));
 sg13g2_nand2b_1 _08211_ (.Y(_02741_),
    .B(_02590_),
    .A_N(_02588_));
 sg13g2_o21ai_1 _08212_ (.B1(_02616_),
    .Y(_02742_),
    .A1(_02613_),
    .A2(_02617_));
 sg13g2_nand2_1 _08213_ (.Y(_02743_),
    .A(net1458),
    .B(net1176));
 sg13g2_nand2_1 _08214_ (.Y(_02744_),
    .A(net1463),
    .B(net1166));
 sg13g2_and4_1 _08215_ (.A(net1467),
    .B(net1462),
    .C(net1169),
    .D(net1164),
    .X(_02745_));
 sg13g2_a22oi_1 _08216_ (.Y(_02746_),
    .B1(net1164),
    .B2(net1467),
    .A2(net1169),
    .A1(net1462));
 sg13g2_or3_1 _08217_ (.A(_02743_),
    .B(_02745_),
    .C(_02746_),
    .X(_02747_));
 sg13g2_o21ai_1 _08218_ (.B1(_02743_),
    .Y(_02748_),
    .A1(_02745_),
    .A2(_02746_));
 sg13g2_nand3_1 _08219_ (.B(_02747_),
    .C(_02748_),
    .A(_02742_),
    .Y(_02749_));
 sg13g2_a21o_1 _08220_ (.A2(_02748_),
    .A1(_02747_),
    .B1(_02742_),
    .X(_02750_));
 sg13g2_nand3_1 _08221_ (.B(_02749_),
    .C(_02750_),
    .A(_02741_),
    .Y(_02751_));
 sg13g2_a21o_1 _08222_ (.A2(_02750_),
    .A1(_02749_),
    .B1(_02741_),
    .X(_02752_));
 sg13g2_nand3_1 _08223_ (.B(_02751_),
    .C(_02752_),
    .A(_02740_),
    .Y(_02753_));
 sg13g2_a21o_1 _08224_ (.A2(_02752_),
    .A1(_02751_),
    .B1(_02740_),
    .X(_02754_));
 sg13g2_nand3_1 _08225_ (.B(_02753_),
    .C(_02754_),
    .A(_02739_),
    .Y(_02755_));
 sg13g2_a21o_1 _08226_ (.A2(_02754_),
    .A1(_02753_),
    .B1(_02739_),
    .X(_02756_));
 sg13g2_and3_1 _08227_ (.X(_02757_),
    .A(_02738_),
    .B(_02755_),
    .C(_02756_));
 sg13g2_nand3_1 _08228_ (.B(_02755_),
    .C(_02756_),
    .A(_02738_),
    .Y(_02758_));
 sg13g2_a21oi_1 _08229_ (.A1(_02755_),
    .A2(_02756_),
    .Y(_02759_),
    .B1(_02738_));
 sg13g2_a21o_1 _08230_ (.A2(_02756_),
    .A1(_02755_),
    .B1(_02738_),
    .X(_02760_));
 sg13g2_nor3_1 _08231_ (.A(_02737_),
    .B(_02757_),
    .C(_02759_),
    .Y(_02761_));
 sg13g2_nand3_1 _08232_ (.B(_02758_),
    .C(_02760_),
    .A(_02737_),
    .Y(_02762_));
 sg13g2_a21o_1 _08233_ (.A2(_02760_),
    .A1(_02758_),
    .B1(_02737_),
    .X(_02763_));
 sg13g2_a21oi_2 _08234_ (.B1(_02632_),
    .Y(_02764_),
    .A2(_02763_),
    .A1(_02762_));
 sg13g2_and3_1 _08235_ (.X(_02765_),
    .A(_02632_),
    .B(_02762_),
    .C(_02763_));
 sg13g2_nor3_1 _08236_ (.A(_02705_),
    .B(_02764_),
    .C(_02765_),
    .Y(_02766_));
 sg13g2_or3_1 _08237_ (.A(_02705_),
    .B(_02764_),
    .C(_02765_),
    .X(_02767_));
 sg13g2_o21ai_1 _08238_ (.B1(_02705_),
    .Y(_02768_),
    .A1(_02764_),
    .A2(_02765_));
 sg13g2_nand3_1 _08239_ (.B(_02767_),
    .C(_02768_),
    .A(_02704_),
    .Y(_02769_));
 sg13g2_a21o_1 _08240_ (.A2(_02768_),
    .A1(_02767_),
    .B1(_02704_),
    .X(_02770_));
 sg13g2_nand3_1 _08241_ (.B(_02769_),
    .C(_02770_),
    .A(_02666_),
    .Y(_02771_));
 sg13g2_a21o_1 _08242_ (.A2(_02770_),
    .A1(_02769_),
    .B1(_02666_),
    .X(_02772_));
 sg13g2_nand3_1 _08243_ (.B(_02771_),
    .C(_02772_),
    .A(_02665_),
    .Y(_02773_));
 sg13g2_a21o_1 _08244_ (.A2(_02772_),
    .A1(_02771_),
    .B1(_02665_),
    .X(_02774_));
 sg13g2_nand3_1 _08245_ (.B(_02773_),
    .C(_02774_),
    .A(_02660_),
    .Y(_02775_));
 sg13g2_a21o_1 _08246_ (.A2(_02774_),
    .A1(_02773_),
    .B1(_02660_),
    .X(_02776_));
 sg13g2_nand2_1 _08247_ (.Y(_02777_),
    .A(_02775_),
    .B(_02776_));
 sg13g2_xor2_1 _08248_ (.B(_02777_),
    .A(_02659_),
    .X(_02778_));
 sg13g2_nor2_1 _08249_ (.A(_02658_),
    .B(_02778_),
    .Y(_02779_));
 sg13g2_nand2_1 _08250_ (.Y(_02780_),
    .A(_02658_),
    .B(_02778_));
 sg13g2_xor2_1 _08251_ (.B(_02778_),
    .A(_02658_),
    .X(_02781_));
 sg13g2_a21oi_1 _08252_ (.A1(_02650_),
    .A2(_02655_),
    .Y(_02782_),
    .B1(_02649_));
 sg13g2_xor2_1 _08253_ (.B(_02782_),
    .A(_02781_),
    .X(_02783_));
 sg13g2_o21ai_1 _08254_ (.B1(net1518),
    .Y(_02784_),
    .A1(net1297),
    .A2(net256));
 sg13g2_a21oi_1 _08255_ (.A1(net1297),
    .A2(_02783_),
    .Y(_00233_),
    .B1(_02784_));
 sg13g2_a21oi_1 _08256_ (.A1(_02661_),
    .A2(_02664_),
    .Y(_02785_),
    .B1(_02663_));
 sg13g2_nand2_1 _08257_ (.Y(_02786_),
    .A(_02771_),
    .B(_02773_));
 sg13g2_a21o_1 _08258_ (.A2(_02713_),
    .A1(_02707_),
    .B1(_02715_),
    .X(_02787_));
 sg13g2_o21ai_1 _08259_ (.B1(_02735_),
    .Y(_02788_),
    .A1(_02716_),
    .A2(_02736_));
 sg13g2_o21ai_1 _08260_ (.B1(_02788_),
    .Y(_02789_),
    .A1(_02764_),
    .A2(_02766_));
 sg13g2_or3_1 _08261_ (.A(_02764_),
    .B(_02766_),
    .C(_02788_),
    .X(_02790_));
 sg13g2_nand2_1 _08262_ (.Y(_02791_),
    .A(_02789_),
    .B(_02790_));
 sg13g2_nand2b_1 _08263_ (.Y(_02792_),
    .B(_02787_),
    .A_N(_02791_));
 sg13g2_xnor2_1 _08264_ (.Y(_02793_),
    .A(_02787_),
    .B(_02791_));
 sg13g2_nand2_1 _08265_ (.Y(_02794_),
    .A(_02703_),
    .B(_02769_));
 sg13g2_a22oi_1 _08266_ (.Y(_02795_),
    .B1(net1328),
    .B2(net1405),
    .A2(net1223),
    .A1(net1416));
 sg13g2_nand4_1 _08267_ (.B(net1416),
    .C(net1223),
    .A(net1405),
    .Y(_02796_),
    .D(net1328));
 sg13g2_nand2b_2 _08268_ (.Y(_02797_),
    .B(_02796_),
    .A_N(_02795_));
 sg13g2_nand2_1 _08269_ (.Y(_02798_),
    .A(net1379),
    .B(net1336));
 sg13g2_nand2_1 _08270_ (.Y(_02799_),
    .A(net1394),
    .B(net1330));
 sg13g2_nand2_1 _08271_ (.Y(_02800_),
    .A(net1394),
    .B(net1333));
 sg13g2_or2_1 _08272_ (.X(_02801_),
    .B(_02799_),
    .A(_02610_));
 sg13g2_xor2_1 _08273_ (.B(_02800_),
    .A(_02669_),
    .X(_02802_));
 sg13g2_nand2b_1 _08274_ (.Y(_02803_),
    .B(_02802_),
    .A_N(_02798_));
 sg13g2_xnor2_1 _08275_ (.Y(_02804_),
    .A(_02798_),
    .B(_02802_));
 sg13g2_o21ai_1 _08276_ (.B1(_02672_),
    .Y(_02805_),
    .A1(_02610_),
    .A2(_02670_));
 sg13g2_nand2_1 _08277_ (.Y(_02806_),
    .A(_02804_),
    .B(_02805_));
 sg13g2_xor2_1 _08278_ (.B(_02805_),
    .A(_02804_),
    .X(_02807_));
 sg13g2_nor2b_1 _08279_ (.A(_02674_),
    .B_N(_02807_),
    .Y(_02808_));
 sg13g2_xnor2_1 _08280_ (.Y(_02809_),
    .A(_02674_),
    .B(_02807_));
 sg13g2_nand2_1 _08281_ (.Y(_02810_),
    .A(net1468),
    .B(net1160));
 sg13g2_nand2_1 _08282_ (.Y(_02811_),
    .A(net1472),
    .B(net1150));
 sg13g2_nand2_1 _08283_ (.Y(_02812_),
    .A(net1472),
    .B(net1156));
 sg13g2_or2_1 _08284_ (.X(_02813_),
    .B(_02811_),
    .A(_02678_));
 sg13g2_xnor2_1 _08285_ (.Y(_02814_),
    .A(_02677_),
    .B(_02812_));
 sg13g2_xor2_1 _08286_ (.B(_02814_),
    .A(_02810_),
    .X(_02815_));
 sg13g2_inv_1 _08287_ (.Y(_02816_),
    .A(_02815_));
 sg13g2_nand2_1 _08288_ (.Y(_02817_),
    .A(_02687_),
    .B(_02690_));
 sg13g2_nand2_1 _08289_ (.Y(_02818_),
    .A(net1361),
    .B(net1349));
 sg13g2_nand2_1 _08290_ (.Y(_02819_),
    .A(net1368),
    .B(net1346));
 sg13g2_or2_1 _08291_ (.X(_02820_),
    .B(_02819_),
    .A(_02686_));
 sg13g2_and2_1 _08292_ (.A(_02686_),
    .B(_02819_),
    .X(_02821_));
 sg13g2_xor2_1 _08293_ (.B(_02819_),
    .A(_02686_),
    .X(_02822_));
 sg13g2_xnor2_1 _08294_ (.Y(_02823_),
    .A(_02818_),
    .B(_02822_));
 sg13g2_nand2_1 _08295_ (.Y(_02824_),
    .A(_02817_),
    .B(_02823_));
 sg13g2_xnor2_1 _08296_ (.Y(_02825_),
    .A(_02817_),
    .B(_02823_));
 sg13g2_xnor2_1 _08297_ (.Y(_02826_),
    .A(_02815_),
    .B(_02825_));
 sg13g2_xnor2_1 _08298_ (.Y(_02827_),
    .A(_02809_),
    .B(_02826_));
 sg13g2_nor2_1 _08299_ (.A(_02697_),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_xor2_1 _08300_ (.B(_02827_),
    .A(_02697_),
    .X(_02829_));
 sg13g2_nand2b_1 _08301_ (.Y(_02830_),
    .B(_02829_),
    .A_N(_02797_));
 sg13g2_xnor2_1 _08302_ (.Y(_02831_),
    .A(_02797_),
    .B(_02829_));
 sg13g2_and2_1 _08303_ (.A(_02701_),
    .B(_02831_),
    .X(_02832_));
 sg13g2_xor2_1 _08304_ (.B(_02831_),
    .A(_02701_),
    .X(_02833_));
 sg13g2_nor2_1 _08305_ (.A(_02757_),
    .B(_02761_),
    .Y(_02834_));
 sg13g2_o21ai_1 _08306_ (.B1(_02711_),
    .Y(_02835_),
    .A1(_02708_),
    .A2(_02712_));
 sg13g2_o21ai_1 _08307_ (.B1(_02722_),
    .Y(_02836_),
    .A1(_02564_),
    .A2(_02720_));
 sg13g2_nand2_1 _08308_ (.Y(_02837_),
    .A(net1414),
    .B(net1227));
 sg13g2_nand2_2 _08309_ (.Y(_02838_),
    .A(net1420),
    .B(net1208));
 sg13g2_nand2_1 _08310_ (.Y(_02839_),
    .A(net1420),
    .B(net1214));
 sg13g2_or2_1 _08311_ (.X(_02840_),
    .B(_02838_),
    .A(_02710_));
 sg13g2_xnor2_1 _08312_ (.Y(_02841_),
    .A(_02709_),
    .B(_02839_));
 sg13g2_xor2_1 _08313_ (.B(_02841_),
    .A(_02837_),
    .X(_02842_));
 sg13g2_xnor2_1 _08314_ (.Y(_02843_),
    .A(_02836_),
    .B(_02842_));
 sg13g2_nor2b_1 _08315_ (.A(_02843_),
    .B_N(_02835_),
    .Y(_02844_));
 sg13g2_xor2_1 _08316_ (.B(_02843_),
    .A(_02835_),
    .X(_02845_));
 sg13g2_o21ai_1 _08317_ (.B1(_02732_),
    .Y(_02846_),
    .A1(_02723_),
    .A2(_02733_));
 sg13g2_nand2_1 _08318_ (.Y(_02847_),
    .A(net1426),
    .B(net1207));
 sg13g2_nand2_1 _08319_ (.Y(_02848_),
    .A(net1430),
    .B(net1198));
 sg13g2_nand2_1 _08320_ (.Y(_02849_),
    .A(net1430),
    .B(net1201));
 sg13g2_xor2_1 _08321_ (.B(_02849_),
    .A(_02719_),
    .X(_02850_));
 sg13g2_nand2b_1 _08322_ (.Y(_02851_),
    .B(_02850_),
    .A_N(_02847_));
 sg13g2_xor2_1 _08323_ (.B(_02850_),
    .A(_02847_),
    .X(_02852_));
 sg13g2_or2_1 _08324_ (.X(_02853_),
    .B(_02729_),
    .A(_02727_));
 sg13g2_nand2_1 _08325_ (.Y(_02854_),
    .A(net1438),
    .B(net1191));
 sg13g2_nand2_1 _08326_ (.Y(_02855_),
    .A(net1443),
    .B(net1183));
 sg13g2_nand2_1 _08327_ (.Y(_02856_),
    .A(net1443),
    .B(net1189));
 sg13g2_xor2_1 _08328_ (.B(_02856_),
    .A(_02726_),
    .X(_02857_));
 sg13g2_nand2b_1 _08329_ (.Y(_02858_),
    .B(_02857_),
    .A_N(_02854_));
 sg13g2_xnor2_1 _08330_ (.Y(_02859_),
    .A(_02854_),
    .B(_02857_));
 sg13g2_nand2_1 _08331_ (.Y(_02860_),
    .A(_02853_),
    .B(_02859_));
 sg13g2_xnor2_1 _08332_ (.Y(_02861_),
    .A(_02853_),
    .B(_02859_));
 sg13g2_xnor2_1 _08333_ (.Y(_02862_),
    .A(_02852_),
    .B(_02861_));
 sg13g2_nand2b_1 _08334_ (.Y(_02863_),
    .B(_02846_),
    .A_N(_02862_));
 sg13g2_xor2_1 _08335_ (.B(_02862_),
    .A(_02846_),
    .X(_02864_));
 sg13g2_xor2_1 _08336_ (.B(_02864_),
    .A(_02845_),
    .X(_02865_));
 sg13g2_nand2_1 _08337_ (.Y(_02866_),
    .A(_02753_),
    .B(_02755_));
 sg13g2_and2_1 _08338_ (.A(_02749_),
    .B(_02751_),
    .X(_02867_));
 sg13g2_o21ai_1 _08339_ (.B1(_02692_),
    .Y(_02868_),
    .A1(_02682_),
    .A2(_02693_));
 sg13g2_nand2b_1 _08340_ (.Y(_02869_),
    .B(_02747_),
    .A_N(_02745_));
 sg13g2_o21ai_1 _08341_ (.B1(_02679_),
    .Y(_02870_),
    .A1(_02676_),
    .A2(_02680_));
 sg13g2_nand2_1 _08342_ (.Y(_02871_),
    .A(net1453),
    .B(net1175));
 sg13g2_nand2_1 _08343_ (.Y(_02872_),
    .A(net1457),
    .B(net1166));
 sg13g2_nand2_1 _08344_ (.Y(_02873_),
    .A(net1457),
    .B(net1171));
 sg13g2_or2_1 _08345_ (.X(_02874_),
    .B(_02873_),
    .A(_02744_));
 sg13g2_xnor2_1 _08346_ (.Y(_02875_),
    .A(_02744_),
    .B(_02873_));
 sg13g2_xor2_1 _08347_ (.B(_02875_),
    .A(_02871_),
    .X(_02876_));
 sg13g2_xnor2_1 _08348_ (.Y(_02877_),
    .A(_02870_),
    .B(_02876_));
 sg13g2_nor2b_1 _08349_ (.A(_02877_),
    .B_N(_02869_),
    .Y(_02878_));
 sg13g2_xor2_1 _08350_ (.B(_02877_),
    .A(_02869_),
    .X(_02879_));
 sg13g2_nand2b_1 _08351_ (.Y(_02880_),
    .B(_02868_),
    .A_N(_02879_));
 sg13g2_xor2_1 _08352_ (.B(_02879_),
    .A(_02868_),
    .X(_02881_));
 sg13g2_xnor2_1 _08353_ (.Y(_02882_),
    .A(_02867_),
    .B(_02881_));
 sg13g2_nor2b_1 _08354_ (.A(_02882_),
    .B_N(_02866_),
    .Y(_02883_));
 sg13g2_nand2b_1 _08355_ (.Y(_02884_),
    .B(_02882_),
    .A_N(_02866_));
 sg13g2_xor2_1 _08356_ (.B(_02882_),
    .A(_02866_),
    .X(_02885_));
 sg13g2_xnor2_1 _08357_ (.Y(_02886_),
    .A(_02865_),
    .B(_02885_));
 sg13g2_nand2_1 _08358_ (.Y(_02887_),
    .A(_02699_),
    .B(_02886_));
 sg13g2_xnor2_1 _08359_ (.Y(_02888_),
    .A(_02699_),
    .B(_02886_));
 sg13g2_xor2_1 _08360_ (.B(_02888_),
    .A(_02834_),
    .X(_02889_));
 sg13g2_xor2_1 _08361_ (.B(_02889_),
    .A(_02833_),
    .X(_02890_));
 sg13g2_and2_1 _08362_ (.A(_02794_),
    .B(_02890_),
    .X(_02891_));
 sg13g2_xor2_1 _08363_ (.B(_02890_),
    .A(_02794_),
    .X(_02892_));
 sg13g2_xor2_1 _08364_ (.B(_02892_),
    .A(_02793_),
    .X(_02893_));
 sg13g2_nand2_1 _08365_ (.Y(_02894_),
    .A(_02786_),
    .B(_02893_));
 sg13g2_xnor2_1 _08366_ (.Y(_02895_),
    .A(_02786_),
    .B(_02893_));
 sg13g2_xor2_1 _08367_ (.B(_02895_),
    .A(_02785_),
    .X(_02896_));
 sg13g2_o21ai_1 _08368_ (.B1(_02775_),
    .Y(_02897_),
    .A1(_02659_),
    .A2(_02777_));
 sg13g2_nand2_1 _08369_ (.Y(_02898_),
    .A(_02896_),
    .B(_02897_));
 sg13g2_inv_1 _08370_ (.Y(_02899_),
    .A(_02898_));
 sg13g2_xor2_1 _08371_ (.B(_02897_),
    .A(_02896_),
    .X(_02900_));
 sg13g2_o21ai_1 _08372_ (.B1(_02780_),
    .Y(_02901_),
    .A1(_02648_),
    .A2(_02779_));
 sg13g2_and2_1 _08373_ (.A(_02650_),
    .B(_02781_),
    .X(_02902_));
 sg13g2_a21o_1 _08374_ (.A2(_02902_),
    .A1(_02655_),
    .B1(_02901_),
    .X(_02903_));
 sg13g2_xor2_1 _08375_ (.B(_02903_),
    .A(_02900_),
    .X(_02904_));
 sg13g2_o21ai_1 _08376_ (.B1(net1521),
    .Y(_02905_),
    .A1(net1143),
    .A2(_02904_));
 sg13g2_a21oi_1 _08377_ (.A1(net1143),
    .A2(_04777_),
    .Y(_00234_),
    .B1(_02905_));
 sg13g2_a21oi_1 _08378_ (.A1(_02900_),
    .A2(_02903_),
    .Y(_02906_),
    .B1(_02899_));
 sg13g2_o21ai_1 _08379_ (.B1(_02894_),
    .Y(_02907_),
    .A1(_02785_),
    .A2(_02895_));
 sg13g2_nand2_1 _08380_ (.Y(_02908_),
    .A(_02789_),
    .B(_02792_));
 sg13g2_a21oi_1 _08381_ (.A1(_02793_),
    .A2(_02892_),
    .Y(_02909_),
    .B1(_02891_));
 sg13g2_a21o_1 _08382_ (.A2(_02842_),
    .A1(_02836_),
    .B1(_02844_),
    .X(_02910_));
 sg13g2_o21ai_1 _08383_ (.B1(_02887_),
    .Y(_02911_),
    .A1(_02834_),
    .A2(_02888_));
 sg13g2_o21ai_1 _08384_ (.B1(_02863_),
    .Y(_02912_),
    .A1(_02845_),
    .A2(_02864_));
 sg13g2_and2_1 _08385_ (.A(_02911_),
    .B(_02912_),
    .X(_02913_));
 sg13g2_xor2_1 _08386_ (.B(_02912_),
    .A(_02911_),
    .X(_02914_));
 sg13g2_xor2_1 _08387_ (.B(_02914_),
    .A(_02910_),
    .X(_02915_));
 sg13g2_a21oi_1 _08388_ (.A1(_02833_),
    .A2(_02889_),
    .Y(_02916_),
    .B1(_02832_));
 sg13g2_nand2_1 _08389_ (.Y(_02917_),
    .A(net1372),
    .B(net1336));
 sg13g2_nand2_1 _08390_ (.Y(_02918_),
    .A(net1379),
    .B(net1330));
 sg13g2_nand2_1 _08391_ (.Y(_02919_),
    .A(net1379),
    .B(net1333));
 sg13g2_or2_1 _08392_ (.X(_02920_),
    .B(_02918_),
    .A(_02800_));
 sg13g2_xor2_1 _08393_ (.B(_02919_),
    .A(_02799_),
    .X(_02921_));
 sg13g2_nand2b_1 _08394_ (.Y(_02922_),
    .B(_02921_),
    .A_N(_02917_));
 sg13g2_xnor2_1 _08395_ (.Y(_02923_),
    .A(_02917_),
    .B(_02921_));
 sg13g2_and2_1 _08396_ (.A(_02801_),
    .B(_02803_),
    .X(_02924_));
 sg13g2_nand2b_1 _08397_ (.Y(_02925_),
    .B(_02923_),
    .A_N(_02924_));
 sg13g2_xnor2_1 _08398_ (.Y(_02926_),
    .A(_02923_),
    .B(_02924_));
 sg13g2_nor2b_1 _08399_ (.A(_02806_),
    .B_N(_02926_),
    .Y(_02927_));
 sg13g2_xnor2_1 _08400_ (.Y(_02928_),
    .A(_02806_),
    .B(_02926_));
 sg13g2_nand2_1 _08401_ (.Y(_02929_),
    .A(net1463),
    .B(net1160));
 sg13g2_nand2_1 _08402_ (.Y(_02930_),
    .A(net1468),
    .B(net1150));
 sg13g2_nand2_1 _08403_ (.Y(_02931_),
    .A(net1468),
    .B(net1156));
 sg13g2_or2_1 _08404_ (.X(_02932_),
    .B(_02930_),
    .A(_02812_));
 sg13g2_xnor2_1 _08405_ (.Y(_02933_),
    .A(_02811_),
    .B(_02931_));
 sg13g2_xnor2_1 _08406_ (.Y(_02934_),
    .A(_02929_),
    .B(_02933_));
 sg13g2_o21ai_1 _08407_ (.B1(_02820_),
    .Y(_02935_),
    .A1(_02818_),
    .A2(_02821_));
 sg13g2_nand2_1 _08408_ (.Y(_02936_),
    .A(net1354),
    .B(net1349));
 sg13g2_nand2_1 _08409_ (.Y(_02937_),
    .A(net1359),
    .B(net1341));
 sg13g2_and4_1 _08410_ (.A(net1368),
    .B(net1361),
    .C(net1346),
    .D(net1340),
    .X(_02938_));
 sg13g2_a22oi_1 _08411_ (.Y(_02939_),
    .B1(net1340),
    .B2(net1368),
    .A2(net1346),
    .A1(net1361));
 sg13g2_nor3_1 _08412_ (.A(_02936_),
    .B(_02938_),
    .C(_02939_),
    .Y(_02940_));
 sg13g2_o21ai_1 _08413_ (.B1(_02936_),
    .Y(_02941_),
    .A1(_02938_),
    .A2(_02939_));
 sg13g2_nor2b_1 _08414_ (.A(_02940_),
    .B_N(_02941_),
    .Y(_02942_));
 sg13g2_nand2_1 _08415_ (.Y(_02943_),
    .A(_02935_),
    .B(_02942_));
 sg13g2_xnor2_1 _08416_ (.Y(_02944_),
    .A(_02935_),
    .B(_02942_));
 sg13g2_xnor2_1 _08417_ (.Y(_02945_),
    .A(_02934_),
    .B(_02944_));
 sg13g2_inv_1 _08418_ (.Y(_02946_),
    .A(_02945_));
 sg13g2_xnor2_1 _08419_ (.Y(_02947_),
    .A(_02928_),
    .B(_02946_));
 sg13g2_a21oi_1 _08420_ (.A1(_02809_),
    .A2(_02826_),
    .Y(_02948_),
    .B1(_02808_));
 sg13g2_nor2_1 _08421_ (.A(_02947_),
    .B(_02948_),
    .Y(_02949_));
 sg13g2_inv_2 _08422_ (.Y(_02950_),
    .A(_02949_));
 sg13g2_xnor2_1 _08423_ (.Y(_02951_),
    .A(_02947_),
    .B(_02948_));
 sg13g2_nand2_1 _08424_ (.Y(_02952_),
    .A(net1414),
    .B(net1223));
 sg13g2_nand2_2 _08425_ (.Y(_02953_),
    .A(net1395),
    .B(net1324));
 sg13g2_and2_1 _08426_ (.A(net1405),
    .B(net1324),
    .X(_02954_));
 sg13g2_nand2_2 _08427_ (.Y(_02955_),
    .A(net1405),
    .B(net1324));
 sg13g2_nand2_1 _08428_ (.Y(_02956_),
    .A(net1395),
    .B(net1328));
 sg13g2_or2_1 _08429_ (.X(_02957_),
    .B(_02956_),
    .A(_02955_));
 sg13g2_xnor2_1 _08430_ (.Y(_02958_),
    .A(_02954_),
    .B(_02956_));
 sg13g2_nor2b_1 _08431_ (.A(_02952_),
    .B_N(_02958_),
    .Y(_02959_));
 sg13g2_xnor2_1 _08432_ (.Y(_02960_),
    .A(_02952_),
    .B(_02958_));
 sg13g2_inv_1 _08433_ (.Y(_02961_),
    .A(_02960_));
 sg13g2_xnor2_1 _08434_ (.Y(_02962_),
    .A(_02796_),
    .B(_02960_));
 sg13g2_nand2b_1 _08435_ (.Y(_02963_),
    .B(_02962_),
    .A_N(_02951_));
 sg13g2_xor2_1 _08436_ (.B(_02962_),
    .A(_02951_),
    .X(_02964_));
 sg13g2_nor2_1 _08437_ (.A(_02830_),
    .B(_02964_),
    .Y(_02965_));
 sg13g2_xor2_1 _08438_ (.B(_02964_),
    .A(_02830_),
    .X(_02966_));
 sg13g2_a21oi_1 _08439_ (.A1(_02865_),
    .A2(_02884_),
    .Y(_02967_),
    .B1(_02883_));
 sg13g2_o21ai_1 _08440_ (.B1(_02840_),
    .Y(_02968_),
    .A1(_02837_),
    .A2(_02841_));
 sg13g2_o21ai_1 _08441_ (.B1(_02851_),
    .Y(_02969_),
    .A1(_02719_),
    .A2(_02849_));
 sg13g2_nand2_2 _08442_ (.Y(_02970_),
    .A(net1411),
    .B(net1227));
 sg13g2_nand2_1 _08443_ (.Y(_02971_),
    .A(net1416),
    .B(net1215));
 sg13g2_xor2_1 _08444_ (.B(_02971_),
    .A(_02838_),
    .X(_02972_));
 sg13g2_nand2b_1 _08445_ (.Y(_02973_),
    .B(_02972_),
    .A_N(_02970_));
 sg13g2_xnor2_1 _08446_ (.Y(_02974_),
    .A(_02970_),
    .B(_02972_));
 sg13g2_xnor2_1 _08447_ (.Y(_02975_),
    .A(_02969_),
    .B(_02974_));
 sg13g2_nor2b_1 _08448_ (.A(_02975_),
    .B_N(_02968_),
    .Y(_02976_));
 sg13g2_xor2_1 _08449_ (.B(_02975_),
    .A(_02968_),
    .X(_02977_));
 sg13g2_o21ai_1 _08450_ (.B1(_02860_),
    .Y(_02978_),
    .A1(_02852_),
    .A2(_02861_));
 sg13g2_nand2_1 _08451_ (.Y(_02979_),
    .A(net1422),
    .B(net1207));
 sg13g2_nand2_1 _08452_ (.Y(_02980_),
    .A(net1426),
    .B(net1198));
 sg13g2_nand2_1 _08453_ (.Y(_02981_),
    .A(net1426),
    .B(net1200));
 sg13g2_xor2_1 _08454_ (.B(_02981_),
    .A(_02848_),
    .X(_02982_));
 sg13g2_nand2b_1 _08455_ (.Y(_02983_),
    .B(_02982_),
    .A_N(_02979_));
 sg13g2_xor2_1 _08456_ (.B(_02982_),
    .A(_02979_),
    .X(_02984_));
 sg13g2_o21ai_1 _08457_ (.B1(_02858_),
    .Y(_02985_),
    .A1(_02726_),
    .A2(_02856_));
 sg13g2_nand2_1 _08458_ (.Y(_02986_),
    .A(net1434),
    .B(net1191));
 sg13g2_nand2_1 _08459_ (.Y(_02987_),
    .A(net1438),
    .B(net1183));
 sg13g2_nand2_1 _08460_ (.Y(_02988_),
    .A(net1438),
    .B(net1189));
 sg13g2_xor2_1 _08461_ (.B(_02988_),
    .A(_02855_),
    .X(_02989_));
 sg13g2_nand2b_1 _08462_ (.Y(_02990_),
    .B(_02989_),
    .A_N(_02986_));
 sg13g2_xnor2_1 _08463_ (.Y(_02991_),
    .A(_02986_),
    .B(_02989_));
 sg13g2_nand2_1 _08464_ (.Y(_02992_),
    .A(_02985_),
    .B(_02991_));
 sg13g2_xnor2_1 _08465_ (.Y(_02993_),
    .A(_02985_),
    .B(_02991_));
 sg13g2_xnor2_1 _08466_ (.Y(_02994_),
    .A(_02984_),
    .B(_02993_));
 sg13g2_nor2b_1 _08467_ (.A(_02994_),
    .B_N(_02978_),
    .Y(_02995_));
 sg13g2_xor2_1 _08468_ (.B(_02994_),
    .A(_02978_),
    .X(_02996_));
 sg13g2_nor2_1 _08469_ (.A(_02977_),
    .B(_02996_),
    .Y(_02997_));
 sg13g2_xor2_1 _08470_ (.B(_02996_),
    .A(_02977_),
    .X(_02998_));
 sg13g2_inv_1 _08471_ (.Y(_02999_),
    .A(_02998_));
 sg13g2_o21ai_1 _08472_ (.B1(_02880_),
    .Y(_03000_),
    .A1(_02867_),
    .A2(_02881_));
 sg13g2_a21oi_1 _08473_ (.A1(_02870_),
    .A2(_02876_),
    .Y(_03001_),
    .B1(_02878_));
 sg13g2_o21ai_1 _08474_ (.B1(_02824_),
    .Y(_03002_),
    .A1(_02816_),
    .A2(_02825_));
 sg13g2_o21ai_1 _08475_ (.B1(_02874_),
    .Y(_03003_),
    .A1(_02871_),
    .A2(_02875_));
 sg13g2_o21ai_1 _08476_ (.B1(_02813_),
    .Y(_03004_),
    .A1(_02810_),
    .A2(_02814_));
 sg13g2_nand2_1 _08477_ (.Y(_03005_),
    .A(net1448),
    .B(net1175));
 sg13g2_nand2_1 _08478_ (.Y(_03006_),
    .A(net1453),
    .B(net1166));
 sg13g2_nand2_1 _08479_ (.Y(_03007_),
    .A(net1453),
    .B(net1171));
 sg13g2_xor2_1 _08480_ (.B(_03007_),
    .A(_02872_),
    .X(_03008_));
 sg13g2_nand2b_1 _08481_ (.Y(_03009_),
    .B(_03008_),
    .A_N(_03005_));
 sg13g2_xnor2_1 _08482_ (.Y(_03010_),
    .A(_03005_),
    .B(_03008_));
 sg13g2_xnor2_1 _08483_ (.Y(_03011_),
    .A(_03004_),
    .B(_03010_));
 sg13g2_nor2b_1 _08484_ (.A(_03011_),
    .B_N(_03003_),
    .Y(_03012_));
 sg13g2_xor2_1 _08485_ (.B(_03011_),
    .A(_03003_),
    .X(_03013_));
 sg13g2_nand2b_1 _08486_ (.Y(_03014_),
    .B(_03002_),
    .A_N(_03013_));
 sg13g2_xor2_1 _08487_ (.B(_03013_),
    .A(_03002_),
    .X(_03015_));
 sg13g2_xnor2_1 _08488_ (.Y(_03016_),
    .A(_03001_),
    .B(_03015_));
 sg13g2_nand2b_1 _08489_ (.Y(_03017_),
    .B(_03000_),
    .A_N(_03016_));
 sg13g2_xor2_1 _08490_ (.B(_03016_),
    .A(_03000_),
    .X(_03018_));
 sg13g2_xnor2_1 _08491_ (.Y(_03019_),
    .A(_02998_),
    .B(_03018_));
 sg13g2_nand2_1 _08492_ (.Y(_03020_),
    .A(_02828_),
    .B(_03019_));
 sg13g2_xnor2_1 _08493_ (.Y(_03021_),
    .A(_02828_),
    .B(_03019_));
 sg13g2_xor2_1 _08494_ (.B(_03021_),
    .A(_02967_),
    .X(_03022_));
 sg13g2_xnor2_1 _08495_ (.Y(_03023_),
    .A(_02966_),
    .B(_03022_));
 sg13g2_nor2_1 _08496_ (.A(_02916_),
    .B(_03023_),
    .Y(_03024_));
 sg13g2_xor2_1 _08497_ (.B(_03023_),
    .A(_02916_),
    .X(_03025_));
 sg13g2_xor2_1 _08498_ (.B(_03025_),
    .A(_02915_),
    .X(_03026_));
 sg13g2_nand2b_1 _08499_ (.Y(_03027_),
    .B(_03026_),
    .A_N(_02909_));
 sg13g2_xnor2_1 _08500_ (.Y(_03028_),
    .A(_02909_),
    .B(_03026_));
 sg13g2_nand2_1 _08501_ (.Y(_03029_),
    .A(_02908_),
    .B(_03028_));
 sg13g2_xnor2_1 _08502_ (.Y(_03030_),
    .A(_02908_),
    .B(_03028_));
 sg13g2_nand2b_1 _08503_ (.Y(_03031_),
    .B(_02907_),
    .A_N(_03030_));
 sg13g2_nor2b_1 _08504_ (.A(_02907_),
    .B_N(_03030_),
    .Y(_03032_));
 sg13g2_xnor2_1 _08505_ (.Y(_03033_),
    .A(_02907_),
    .B(_03030_));
 sg13g2_xor2_1 _08506_ (.B(_03033_),
    .A(_02906_),
    .X(_03034_));
 sg13g2_o21ai_1 _08507_ (.B1(net1518),
    .Y(_03035_),
    .A1(net1299),
    .A2(net367));
 sg13g2_a21oi_1 _08508_ (.A1(net1299),
    .A2(_03034_),
    .Y(_00235_),
    .B1(net368));
 sg13g2_a21o_1 _08509_ (.A2(_02914_),
    .A1(_02910_),
    .B1(_02913_),
    .X(_03036_));
 sg13g2_a21oi_1 _08510_ (.A1(_02915_),
    .A2(_03025_),
    .Y(_03037_),
    .B1(_03024_));
 sg13g2_a21o_1 _08511_ (.A2(_02974_),
    .A1(_02969_),
    .B1(_02976_),
    .X(_03038_));
 sg13g2_o21ai_1 _08512_ (.B1(_03020_),
    .Y(_03039_),
    .A1(_02967_),
    .A2(_03021_));
 sg13g2_nor2_1 _08513_ (.A(_02995_),
    .B(_02997_),
    .Y(_03040_));
 sg13g2_o21ai_1 _08514_ (.B1(_03039_),
    .Y(_03041_),
    .A1(_02995_),
    .A2(_02997_));
 sg13g2_xnor2_1 _08515_ (.Y(_03042_),
    .A(_03039_),
    .B(_03040_));
 sg13g2_nand2_1 _08516_ (.Y(_03043_),
    .A(_03038_),
    .B(_03042_));
 sg13g2_xor2_1 _08517_ (.B(_03042_),
    .A(_03038_),
    .X(_03044_));
 sg13g2_a21oi_1 _08518_ (.A1(_02966_),
    .A2(_03022_),
    .Y(_03045_),
    .B1(_02965_));
 sg13g2_o21ai_1 _08519_ (.B1(_02963_),
    .Y(_03046_),
    .A1(_02796_),
    .A2(_02961_));
 sg13g2_and2_1 _08520_ (.A(_02920_),
    .B(_02922_),
    .X(_03047_));
 sg13g2_nand2_1 _08521_ (.Y(_03048_),
    .A(net1365),
    .B(net1336));
 sg13g2_nand2_1 _08522_ (.Y(_03049_),
    .A(net1372),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ));
 sg13g2_nand2_1 _08523_ (.Y(_03050_),
    .A(net1372),
    .B(net1333));
 sg13g2_or2_1 _08524_ (.X(_03051_),
    .B(_03049_),
    .A(_02919_));
 sg13g2_xnor2_1 _08525_ (.Y(_03052_),
    .A(_02918_),
    .B(_03050_));
 sg13g2_xor2_1 _08526_ (.B(_03052_),
    .A(_03048_),
    .X(_03053_));
 sg13g2_nand2b_1 _08527_ (.Y(_03054_),
    .B(_03053_),
    .A_N(_02957_));
 sg13g2_xnor2_1 _08528_ (.Y(_03055_),
    .A(_02957_),
    .B(_03053_));
 sg13g2_nand2b_1 _08529_ (.Y(_03056_),
    .B(_03055_),
    .A_N(_03047_));
 sg13g2_xnor2_1 _08530_ (.Y(_03057_),
    .A(_03047_),
    .B(_03055_));
 sg13g2_nand2b_1 _08531_ (.Y(_03058_),
    .B(_03057_),
    .A_N(_02925_));
 sg13g2_xor2_1 _08532_ (.B(_03057_),
    .A(_02925_),
    .X(_03059_));
 sg13g2_nand2_1 _08533_ (.Y(_03060_),
    .A(net1457),
    .B(net1160));
 sg13g2_nand2_2 _08534_ (.Y(_03061_),
    .A(net1463),
    .B(net1150));
 sg13g2_nand2_2 _08535_ (.Y(_03062_),
    .A(net1463),
    .B(net1156));
 sg13g2_or2_1 _08536_ (.X(_03063_),
    .B(_03061_),
    .A(_02931_));
 sg13g2_xnor2_1 _08537_ (.Y(_03064_),
    .A(_02930_),
    .B(_03062_));
 sg13g2_xnor2_1 _08538_ (.Y(_03065_),
    .A(_03060_),
    .B(_03064_));
 sg13g2_or2_1 _08539_ (.X(_03066_),
    .B(_02940_),
    .A(_02938_));
 sg13g2_nand2_1 _08540_ (.Y(_03067_),
    .A(net1472),
    .B(net1350));
 sg13g2_nand2_1 _08541_ (.Y(_03068_),
    .A(net1352),
    .B(net1341));
 sg13g2_nand2_1 _08542_ (.Y(_03069_),
    .A(net1354),
    .B(net1347));
 sg13g2_xor2_1 _08543_ (.B(_03069_),
    .A(_02937_),
    .X(_03070_));
 sg13g2_nand2b_1 _08544_ (.Y(_03071_),
    .B(_03070_),
    .A_N(_03067_));
 sg13g2_xnor2_1 _08545_ (.Y(_03072_),
    .A(_03067_),
    .B(_03070_));
 sg13g2_nand2_1 _08546_ (.Y(_03073_),
    .A(_03066_),
    .B(_03072_));
 sg13g2_xnor2_1 _08547_ (.Y(_03074_),
    .A(_03066_),
    .B(_03072_));
 sg13g2_xnor2_1 _08548_ (.Y(_03075_),
    .A(_03065_),
    .B(_03074_));
 sg13g2_xnor2_1 _08549_ (.Y(_03076_),
    .A(_03059_),
    .B(_03075_));
 sg13g2_a21oi_1 _08550_ (.A1(_02928_),
    .A2(_02946_),
    .Y(_03077_),
    .B1(_02927_));
 sg13g2_nor2_1 _08551_ (.A(_03076_),
    .B(_03077_),
    .Y(_03078_));
 sg13g2_xnor2_1 _08552_ (.Y(_03079_),
    .A(_03076_),
    .B(_03077_));
 sg13g2_nor2_2 _08553_ (.A(_04822_),
    .B(_04823_),
    .Y(_03080_));
 sg13g2_nand2_2 _08554_ (.Y(_03081_),
    .A(net1411),
    .B(net1223));
 sg13g2_nor2_2 _08555_ (.A(_04805_),
    .B(_02955_),
    .Y(_03082_));
 sg13g2_nand2_2 _08556_ (.Y(_03083_),
    .A(net1395),
    .B(_02954_));
 sg13g2_a21oi_2 _08557_ (.B1(net1103),
    .Y(_03084_),
    .A2(_02955_),
    .A1(_02953_));
 sg13g2_a21o_2 _08558_ (.A2(_02955_),
    .A1(_02953_),
    .B1(net1103),
    .X(_03085_));
 sg13g2_and2_1 _08559_ (.A(net1394),
    .B(net1328),
    .X(_03086_));
 sg13g2_xnor2_1 _08560_ (.Y(_03087_),
    .A(_03085_),
    .B(_03086_));
 sg13g2_nor2_1 _08561_ (.A(net1118),
    .B(_03087_),
    .Y(_03088_));
 sg13g2_xnor2_1 _08562_ (.Y(_03089_),
    .A(net1118),
    .B(_03087_));
 sg13g2_xor2_1 _08563_ (.B(_03089_),
    .A(_02959_),
    .X(_03090_));
 sg13g2_nor2b_1 _08564_ (.A(_03079_),
    .B_N(_03090_),
    .Y(_03091_));
 sg13g2_xnor2_1 _08565_ (.Y(_03092_),
    .A(_03079_),
    .B(_03090_));
 sg13g2_and2_1 _08566_ (.A(_03046_),
    .B(_03092_),
    .X(_03093_));
 sg13g2_xor2_1 _08567_ (.B(_03092_),
    .A(_03046_),
    .X(_03094_));
 sg13g2_o21ai_1 _08568_ (.B1(_03017_),
    .Y(_03095_),
    .A1(_02999_),
    .A2(_03018_));
 sg13g2_o21ai_1 _08569_ (.B1(_02973_),
    .Y(_03096_),
    .A1(_02838_),
    .A2(_02971_));
 sg13g2_o21ai_1 _08570_ (.B1(_02983_),
    .Y(_03097_),
    .A1(_02848_),
    .A2(_02981_));
 sg13g2_nor3_1 _08571_ (.A(_04821_),
    .B(_04825_),
    .C(_02971_),
    .Y(_03098_));
 sg13g2_a22oi_1 _08572_ (.Y(_03099_),
    .B1(net1208),
    .B2(net1416),
    .A2(net1215),
    .A1(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ));
 sg13g2_nor3_1 _08573_ (.A(_02970_),
    .B(_03098_),
    .C(_03099_),
    .Y(_03100_));
 sg13g2_o21ai_1 _08574_ (.B1(_02970_),
    .Y(_03101_),
    .A1(_03098_),
    .A2(_03099_));
 sg13g2_nor2b_1 _08575_ (.A(_03100_),
    .B_N(_03101_),
    .Y(_03102_));
 sg13g2_xnor2_1 _08576_ (.Y(_03103_),
    .A(_03097_),
    .B(_03102_));
 sg13g2_nor2b_1 _08577_ (.A(_03103_),
    .B_N(_03096_),
    .Y(_03104_));
 sg13g2_xor2_1 _08578_ (.B(_03103_),
    .A(_03096_),
    .X(_03105_));
 sg13g2_o21ai_1 _08579_ (.B1(_02992_),
    .Y(_03106_),
    .A1(_02984_),
    .A2(_02993_));
 sg13g2_nand2_1 _08580_ (.Y(_03107_),
    .A(net1420),
    .B(net1207));
 sg13g2_nand2_1 _08581_ (.Y(_03108_),
    .A(net1422),
    .B(net1195));
 sg13g2_nand2_1 _08582_ (.Y(_03109_),
    .A(net1422),
    .B(net1200));
 sg13g2_xor2_1 _08583_ (.B(_03109_),
    .A(_02980_),
    .X(_03110_));
 sg13g2_nand2b_1 _08584_ (.Y(_03111_),
    .B(_03110_),
    .A_N(_03107_));
 sg13g2_xor2_1 _08585_ (.B(_03110_),
    .A(_03107_),
    .X(_03112_));
 sg13g2_o21ai_1 _08586_ (.B1(_02990_),
    .Y(_03113_),
    .A1(_02855_),
    .A2(_02988_));
 sg13g2_nand2_1 _08587_ (.Y(_03114_),
    .A(net1430),
    .B(net1191));
 sg13g2_nand2_1 _08588_ (.Y(_03115_),
    .A(net1433),
    .B(net1178));
 sg13g2_nand2_1 _08589_ (.Y(_03116_),
    .A(net1434),
    .B(net1190));
 sg13g2_xor2_1 _08590_ (.B(_03116_),
    .A(_02987_),
    .X(_03117_));
 sg13g2_nand2b_1 _08591_ (.Y(_03118_),
    .B(_03117_),
    .A_N(_03114_));
 sg13g2_xnor2_1 _08592_ (.Y(_03119_),
    .A(_03114_),
    .B(_03117_));
 sg13g2_nand2_1 _08593_ (.Y(_03120_),
    .A(_03113_),
    .B(_03119_));
 sg13g2_xnor2_1 _08594_ (.Y(_03121_),
    .A(_03113_),
    .B(_03119_));
 sg13g2_xor2_1 _08595_ (.B(_03121_),
    .A(_03112_),
    .X(_03122_));
 sg13g2_nand2_1 _08596_ (.Y(_03123_),
    .A(_03106_),
    .B(_03122_));
 sg13g2_xnor2_1 _08597_ (.Y(_03124_),
    .A(_03106_),
    .B(_03122_));
 sg13g2_xor2_1 _08598_ (.B(_03124_),
    .A(_03105_),
    .X(_03125_));
 sg13g2_inv_1 _08599_ (.Y(_03126_),
    .A(_03125_));
 sg13g2_o21ai_1 _08600_ (.B1(_03014_),
    .Y(_03127_),
    .A1(_03001_),
    .A2(_03015_));
 sg13g2_a21oi_1 _08601_ (.A1(_03004_),
    .A2(_03010_),
    .Y(_03128_),
    .B1(_03012_));
 sg13g2_o21ai_1 _08602_ (.B1(_02943_),
    .Y(_03129_),
    .A1(_02934_),
    .A2(_02944_));
 sg13g2_o21ai_1 _08603_ (.B1(_03009_),
    .Y(_03130_),
    .A1(_02872_),
    .A2(_03007_));
 sg13g2_o21ai_1 _08604_ (.B1(_02932_),
    .Y(_03131_),
    .A1(_02929_),
    .A2(_02933_));
 sg13g2_nand2_1 _08605_ (.Y(_03132_),
    .A(net1443),
    .B(net1175));
 sg13g2_nand2_1 _08606_ (.Y(_03133_),
    .A(net1448),
    .B(net1166));
 sg13g2_nand2_1 _08607_ (.Y(_03134_),
    .A(net1448),
    .B(net1171));
 sg13g2_xor2_1 _08608_ (.B(_03134_),
    .A(_03006_),
    .X(_03135_));
 sg13g2_nand2b_1 _08609_ (.Y(_03136_),
    .B(_03135_),
    .A_N(_03132_));
 sg13g2_xnor2_1 _08610_ (.Y(_03137_),
    .A(_03132_),
    .B(_03135_));
 sg13g2_xnor2_1 _08611_ (.Y(_03138_),
    .A(_03131_),
    .B(_03137_));
 sg13g2_nor2b_1 _08612_ (.A(_03138_),
    .B_N(_03130_),
    .Y(_03139_));
 sg13g2_xor2_1 _08613_ (.B(_03138_),
    .A(_03130_),
    .X(_03140_));
 sg13g2_nand2b_1 _08614_ (.Y(_03141_),
    .B(_03129_),
    .A_N(_03140_));
 sg13g2_xor2_1 _08615_ (.B(_03140_),
    .A(_03129_),
    .X(_03142_));
 sg13g2_xnor2_1 _08616_ (.Y(_03143_),
    .A(_03128_),
    .B(_03142_));
 sg13g2_nand2b_1 _08617_ (.Y(_03144_),
    .B(_03127_),
    .A_N(_03143_));
 sg13g2_xor2_1 _08618_ (.B(_03143_),
    .A(_03127_),
    .X(_03145_));
 sg13g2_xor2_1 _08619_ (.B(_03145_),
    .A(_03125_),
    .X(_03146_));
 sg13g2_nor2_1 _08620_ (.A(_02950_),
    .B(_03146_),
    .Y(_03147_));
 sg13g2_nand2_1 _08621_ (.Y(_03148_),
    .A(_02950_),
    .B(_03146_));
 sg13g2_xnor2_1 _08622_ (.Y(_03149_),
    .A(_02950_),
    .B(_03146_));
 sg13g2_xnor2_1 _08623_ (.Y(_03150_),
    .A(_03095_),
    .B(_03149_));
 sg13g2_xnor2_1 _08624_ (.Y(_03151_),
    .A(_03094_),
    .B(_03150_));
 sg13g2_nor2_1 _08625_ (.A(_03045_),
    .B(_03151_),
    .Y(_03152_));
 sg13g2_xor2_1 _08626_ (.B(_03151_),
    .A(_03045_),
    .X(_03153_));
 sg13g2_xor2_1 _08627_ (.B(_03153_),
    .A(_03044_),
    .X(_03154_));
 sg13g2_nand2b_1 _08628_ (.Y(_03155_),
    .B(_03154_),
    .A_N(_03037_));
 sg13g2_xnor2_1 _08629_ (.Y(_03156_),
    .A(_03037_),
    .B(_03154_));
 sg13g2_nand2_1 _08630_ (.Y(_03157_),
    .A(_03036_),
    .B(_03156_));
 sg13g2_xnor2_1 _08631_ (.Y(_03158_),
    .A(_03036_),
    .B(_03156_));
 sg13g2_a21o_1 _08632_ (.A2(_03029_),
    .A1(_03027_),
    .B1(_03158_),
    .X(_03159_));
 sg13g2_nand3_1 _08633_ (.B(_03029_),
    .C(_03158_),
    .A(_03027_),
    .Y(_03160_));
 sg13g2_and2_1 _08634_ (.A(_03159_),
    .B(_03160_),
    .X(_03161_));
 sg13g2_and2_1 _08635_ (.A(_02900_),
    .B(_03033_),
    .X(_03162_));
 sg13g2_a21oi_1 _08636_ (.A1(_02898_),
    .A2(_03031_),
    .Y(_03163_),
    .B1(_03032_));
 sg13g2_a21o_2 _08637_ (.A2(_03162_),
    .A1(_02901_),
    .B1(_03163_),
    .X(_03164_));
 sg13g2_nand4_1 _08638_ (.B(_02781_),
    .C(_02900_),
    .A(_02650_),
    .Y(_03165_),
    .D(_03033_));
 sg13g2_a21oi_2 _08639_ (.B1(_03165_),
    .Y(_03166_),
    .A2(_02654_),
    .A1(_02652_));
 sg13g2_or2_1 _08640_ (.X(_03167_),
    .B(_03166_),
    .A(_03164_));
 sg13g2_o21ai_1 _08641_ (.B1(_03161_),
    .Y(_03168_),
    .A1(_03164_),
    .A2(_03166_));
 sg13g2_xor2_1 _08642_ (.B(_03167_),
    .A(_03161_),
    .X(_03169_));
 sg13g2_o21ai_1 _08643_ (.B1(net1508),
    .Y(_03170_),
    .A1(net1141),
    .A2(_03169_));
 sg13g2_a21oi_1 _08644_ (.A1(net1142),
    .A2(_04776_),
    .Y(_00236_),
    .B1(_03170_));
 sg13g2_nand2_1 _08645_ (.Y(_03171_),
    .A(_03041_),
    .B(_03043_));
 sg13g2_a21oi_1 _08646_ (.A1(_03044_),
    .A2(_03153_),
    .Y(_03172_),
    .B1(_03152_));
 sg13g2_a21o_1 _08647_ (.A2(_03102_),
    .A1(_03097_),
    .B1(_03104_),
    .X(_03173_));
 sg13g2_a21oi_1 _08648_ (.A1(_03095_),
    .A2(_03148_),
    .Y(_03174_),
    .B1(_03147_));
 sg13g2_o21ai_1 _08649_ (.B1(_03123_),
    .Y(_03175_),
    .A1(_03105_),
    .A2(_03124_));
 sg13g2_nor2b_1 _08650_ (.A(_03174_),
    .B_N(_03175_),
    .Y(_03176_));
 sg13g2_xnor2_1 _08651_ (.Y(_03177_),
    .A(_03174_),
    .B(_03175_));
 sg13g2_xor2_1 _08652_ (.B(_03177_),
    .A(_03173_),
    .X(_03178_));
 sg13g2_a21oi_1 _08653_ (.A1(_03094_),
    .A2(_03150_),
    .Y(_03179_),
    .B1(_03093_));
 sg13g2_a21oi_1 _08654_ (.A1(_02959_),
    .A2(_03089_),
    .Y(_03180_),
    .B1(_03091_));
 sg13g2_nand2_1 _08655_ (.Y(_03181_),
    .A(_03054_),
    .B(_03056_));
 sg13g2_o21ai_1 _08656_ (.B1(_03051_),
    .Y(_03182_),
    .A1(_03048_),
    .A2(_03052_));
 sg13g2_a21oi_1 _08657_ (.A1(_03084_),
    .A2(_03086_),
    .Y(_03183_),
    .B1(_03082_));
 sg13g2_nand2_1 _08658_ (.Y(_03184_),
    .A(net1358),
    .B(net1336));
 sg13g2_nand2_1 _08659_ (.Y(_03185_),
    .A(net1365),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ));
 sg13g2_nand2_1 _08660_ (.Y(_03186_),
    .A(net1365),
    .B(net1333));
 sg13g2_or2_1 _08661_ (.X(_03187_),
    .B(_03185_),
    .A(_03050_));
 sg13g2_xnor2_1 _08662_ (.Y(_03188_),
    .A(_03049_),
    .B(_03186_));
 sg13g2_xor2_1 _08663_ (.B(_03188_),
    .A(_03184_),
    .X(_03189_));
 sg13g2_nor2b_1 _08664_ (.A(_03183_),
    .B_N(_03189_),
    .Y(_03190_));
 sg13g2_xnor2_1 _08665_ (.Y(_03191_),
    .A(_03183_),
    .B(_03189_));
 sg13g2_xnor2_1 _08666_ (.Y(_03192_),
    .A(_03182_),
    .B(_03191_));
 sg13g2_nand2b_1 _08667_ (.Y(_03193_),
    .B(_03181_),
    .A_N(_03192_));
 sg13g2_xor2_1 _08668_ (.B(_03192_),
    .A(_03181_),
    .X(_03194_));
 sg13g2_nand2_1 _08669_ (.Y(_03195_),
    .A(net1452),
    .B(net1160));
 sg13g2_nand2_2 _08670_ (.Y(_03196_),
    .A(net1456),
    .B(net1150));
 sg13g2_nand2_1 _08671_ (.Y(_03197_),
    .A(net1456),
    .B(net1156));
 sg13g2_or2_1 _08672_ (.X(_03198_),
    .B(_03196_),
    .A(_03062_));
 sg13g2_xnor2_1 _08673_ (.Y(_03199_),
    .A(_03061_),
    .B(_03197_));
 sg13g2_xnor2_1 _08674_ (.Y(_03200_),
    .A(_03195_),
    .B(_03199_));
 sg13g2_o21ai_1 _08675_ (.B1(_03071_),
    .Y(_03201_),
    .A1(_02937_),
    .A2(_03069_));
 sg13g2_nand2_1 _08676_ (.Y(_03202_),
    .A(net1466),
    .B(net1350));
 sg13g2_nand2_1 _08677_ (.Y(_03203_),
    .A(net1470),
    .B(net1338));
 sg13g2_nand2_1 _08678_ (.Y(_03204_),
    .A(net1474),
    .B(net1347));
 sg13g2_xor2_1 _08679_ (.B(_03204_),
    .A(_03068_),
    .X(_03205_));
 sg13g2_nand2b_1 _08680_ (.Y(_03206_),
    .B(_03205_),
    .A_N(_03202_));
 sg13g2_xnor2_1 _08681_ (.Y(_03207_),
    .A(_03202_),
    .B(_03205_));
 sg13g2_nand2_1 _08682_ (.Y(_03208_),
    .A(_03201_),
    .B(_03207_));
 sg13g2_xnor2_1 _08683_ (.Y(_03209_),
    .A(_03201_),
    .B(_03207_));
 sg13g2_xnor2_1 _08684_ (.Y(_03210_),
    .A(_03200_),
    .B(_03209_));
 sg13g2_xor2_1 _08685_ (.B(_03210_),
    .A(_03194_),
    .X(_03211_));
 sg13g2_o21ai_1 _08686_ (.B1(_03058_),
    .Y(_03212_),
    .A1(_03059_),
    .A2(_03075_));
 sg13g2_nand2_1 _08687_ (.Y(_03213_),
    .A(_03211_),
    .B(_03212_));
 sg13g2_xor2_1 _08688_ (.B(_03212_),
    .A(_03211_),
    .X(_03214_));
 sg13g2_and2_1 _08689_ (.A(net1394),
    .B(net1324),
    .X(_03215_));
 sg13g2_mux2_1 _08690_ (.A0(_02953_),
    .A1(net1395),
    .S(net1117),
    .X(_03216_));
 sg13g2_nand2_1 _08691_ (.Y(_03217_),
    .A(net1379),
    .B(net1327));
 sg13g2_nor2_1 _08692_ (.A(_03216_),
    .B(_03217_),
    .Y(_03218_));
 sg13g2_xor2_1 _08693_ (.B(_03217_),
    .A(_03216_),
    .X(_03219_));
 sg13g2_nand2_1 _08694_ (.Y(_03220_),
    .A(_02954_),
    .B(_03219_));
 sg13g2_xnor2_1 _08695_ (.Y(_03221_),
    .A(_02955_),
    .B(_03219_));
 sg13g2_xnor2_1 _08696_ (.Y(_03222_),
    .A(_03088_),
    .B(_03221_));
 sg13g2_inv_1 _08697_ (.Y(_03223_),
    .A(_03222_));
 sg13g2_xnor2_1 _08698_ (.Y(_03224_),
    .A(_03214_),
    .B(_03222_));
 sg13g2_nand2b_1 _08699_ (.Y(_03225_),
    .B(_03224_),
    .A_N(_03180_));
 sg13g2_xor2_1 _08700_ (.B(_03224_),
    .A(_03180_),
    .X(_03226_));
 sg13g2_o21ai_1 _08701_ (.B1(_03144_),
    .Y(_03227_),
    .A1(_03126_),
    .A2(_03145_));
 sg13g2_o21ai_1 _08702_ (.B1(_03141_),
    .Y(_03228_),
    .A1(_03128_),
    .A2(_03142_));
 sg13g2_inv_1 _08703_ (.Y(_03229_),
    .A(_03228_));
 sg13g2_a21o_1 _08704_ (.A2(_03137_),
    .A1(_03131_),
    .B1(_03139_),
    .X(_03230_));
 sg13g2_o21ai_1 _08705_ (.B1(_03073_),
    .Y(_03231_),
    .A1(_03065_),
    .A2(_03074_));
 sg13g2_o21ai_1 _08706_ (.B1(_03136_),
    .Y(_03232_),
    .A1(_03006_),
    .A2(_03134_));
 sg13g2_o21ai_1 _08707_ (.B1(_03063_),
    .Y(_03233_),
    .A1(_03060_),
    .A2(_03064_));
 sg13g2_nand2_1 _08708_ (.Y(_03234_),
    .A(net1438),
    .B(net1175));
 sg13g2_nand2_1 _08709_ (.Y(_03235_),
    .A(net1442),
    .B(net1162));
 sg13g2_nand2_1 _08710_ (.Y(_03236_),
    .A(net1443),
    .B(net1171));
 sg13g2_xor2_1 _08711_ (.B(_03236_),
    .A(_03133_),
    .X(_03237_));
 sg13g2_nand2b_1 _08712_ (.Y(_03238_),
    .B(_03237_),
    .A_N(_03234_));
 sg13g2_xnor2_1 _08713_ (.Y(_03239_),
    .A(_03234_),
    .B(_03237_));
 sg13g2_xnor2_1 _08714_ (.Y(_03240_),
    .A(_03233_),
    .B(_03239_));
 sg13g2_nor2b_1 _08715_ (.A(_03240_),
    .B_N(_03232_),
    .Y(_03241_));
 sg13g2_xnor2_1 _08716_ (.Y(_03242_),
    .A(_03232_),
    .B(_03240_));
 sg13g2_xnor2_1 _08717_ (.Y(_03243_),
    .A(_03231_),
    .B(_03242_));
 sg13g2_nor2b_1 _08718_ (.A(_03243_),
    .B_N(_03230_),
    .Y(_03244_));
 sg13g2_xor2_1 _08719_ (.B(_03243_),
    .A(_03230_),
    .X(_03245_));
 sg13g2_xor2_1 _08720_ (.B(_03245_),
    .A(_03228_),
    .X(_03246_));
 sg13g2_o21ai_1 _08721_ (.B1(_03120_),
    .Y(_03247_),
    .A1(_03112_),
    .A2(_03121_));
 sg13g2_nand2_1 _08722_ (.Y(_03248_),
    .A(net1416),
    .B(net1207));
 sg13g2_nand2_1 _08723_ (.Y(_03249_),
    .A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .B(net1195));
 sg13g2_nand2_1 _08724_ (.Y(_03250_),
    .A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .B(net1200));
 sg13g2_xor2_1 _08725_ (.B(_03250_),
    .A(_03108_),
    .X(_03251_));
 sg13g2_nand2b_1 _08726_ (.Y(_03252_),
    .B(_03251_),
    .A_N(_03248_));
 sg13g2_xor2_1 _08727_ (.B(_03251_),
    .A(_03248_),
    .X(_03253_));
 sg13g2_o21ai_1 _08728_ (.B1(_03118_),
    .Y(_03254_),
    .A1(_02987_),
    .A2(_03116_));
 sg13g2_nand2_1 _08729_ (.Y(_03255_),
    .A(net1426),
    .B(net1193));
 sg13g2_nand2_1 _08730_ (.Y(_03256_),
    .A(net1429),
    .B(net1178));
 sg13g2_nand2_1 _08731_ (.Y(_03257_),
    .A(net1429),
    .B(net1190));
 sg13g2_xor2_1 _08732_ (.B(_03257_),
    .A(_03115_),
    .X(_03258_));
 sg13g2_nand2b_1 _08733_ (.Y(_03259_),
    .B(_03258_),
    .A_N(_03255_));
 sg13g2_xnor2_1 _08734_ (.Y(_03260_),
    .A(_03255_),
    .B(_03258_));
 sg13g2_nand2_1 _08735_ (.Y(_03261_),
    .A(_03254_),
    .B(_03260_));
 sg13g2_xnor2_1 _08736_ (.Y(_03262_),
    .A(_03254_),
    .B(_03260_));
 sg13g2_xor2_1 _08737_ (.B(_03262_),
    .A(_03253_),
    .X(_03263_));
 sg13g2_nand2_1 _08738_ (.Y(_03264_),
    .A(_03247_),
    .B(_03263_));
 sg13g2_xnor2_1 _08739_ (.Y(_03265_),
    .A(_03247_),
    .B(_03263_));
 sg13g2_or2_1 _08740_ (.X(_03266_),
    .B(_03100_),
    .A(_03098_));
 sg13g2_o21ai_1 _08741_ (.B1(_03111_),
    .Y(_03267_),
    .A1(_02980_),
    .A2(_03109_));
 sg13g2_nand3_1 _08742_ (.B(net1215),
    .C(net1208),
    .A(net1411),
    .Y(_03268_));
 sg13g2_nor2_1 _08743_ (.A(_04821_),
    .B(_03268_),
    .Y(_03269_));
 sg13g2_a22oi_1 _08744_ (.Y(_03270_),
    .B1(net1208),
    .B2(net1414),
    .A2(net1215),
    .A1(net1411));
 sg13g2_nor3_1 _08745_ (.A(_02970_),
    .B(_03269_),
    .C(_03270_),
    .Y(_03271_));
 sg13g2_o21ai_1 _08746_ (.B1(_02970_),
    .Y(_03272_),
    .A1(_03269_),
    .A2(_03270_));
 sg13g2_nor2b_1 _08747_ (.A(_03271_),
    .B_N(_03272_),
    .Y(_03273_));
 sg13g2_xnor2_1 _08748_ (.Y(_03274_),
    .A(_03267_),
    .B(_03273_));
 sg13g2_nor2b_1 _08749_ (.A(_03274_),
    .B_N(_03266_),
    .Y(_03275_));
 sg13g2_xor2_1 _08750_ (.B(_03274_),
    .A(_03266_),
    .X(_03276_));
 sg13g2_xor2_1 _08751_ (.B(_03276_),
    .A(_03265_),
    .X(_03277_));
 sg13g2_nand2b_1 _08752_ (.Y(_03278_),
    .B(_03277_),
    .A_N(_03246_));
 sg13g2_xnor2_1 _08753_ (.Y(_03279_),
    .A(_03246_),
    .B(_03277_));
 sg13g2_xnor2_1 _08754_ (.Y(_03280_),
    .A(_03078_),
    .B(_03279_));
 sg13g2_nor2b_1 _08755_ (.A(_03280_),
    .B_N(_03227_),
    .Y(_03281_));
 sg13g2_xor2_1 _08756_ (.B(_03280_),
    .A(_03227_),
    .X(_03282_));
 sg13g2_xnor2_1 _08757_ (.Y(_03283_),
    .A(_03226_),
    .B(_03282_));
 sg13g2_nor2_1 _08758_ (.A(_03179_),
    .B(_03283_),
    .Y(_03284_));
 sg13g2_xor2_1 _08759_ (.B(_03283_),
    .A(_03179_),
    .X(_03285_));
 sg13g2_xor2_1 _08760_ (.B(_03285_),
    .A(_03178_),
    .X(_03286_));
 sg13g2_nor2b_1 _08761_ (.A(_03172_),
    .B_N(_03286_),
    .Y(_03287_));
 sg13g2_xnor2_1 _08762_ (.Y(_03288_),
    .A(_03172_),
    .B(_03286_));
 sg13g2_xnor2_1 _08763_ (.Y(_03289_),
    .A(_03171_),
    .B(_03288_));
 sg13g2_and3_1 _08764_ (.X(_03290_),
    .A(_03155_),
    .B(_03157_),
    .C(_03289_));
 sg13g2_a21o_1 _08765_ (.A2(_03157_),
    .A1(_03155_),
    .B1(_03289_),
    .X(_03291_));
 sg13g2_nor2b_2 _08766_ (.A(_03290_),
    .B_N(_03291_),
    .Y(_03292_));
 sg13g2_nand2_1 _08767_ (.Y(_03293_),
    .A(_03159_),
    .B(_03168_));
 sg13g2_xor2_1 _08768_ (.B(_03293_),
    .A(_03292_),
    .X(_03294_));
 sg13g2_o21ai_1 _08769_ (.B1(net1508),
    .Y(_03295_),
    .A1(net1142),
    .A2(_03294_));
 sg13g2_a21oi_1 _08770_ (.A1(net1141),
    .A2(_04775_),
    .Y(_00237_),
    .B1(_03295_));
 sg13g2_a21o_1 _08771_ (.A2(_03177_),
    .A1(_03173_),
    .B1(_03176_),
    .X(_03296_));
 sg13g2_a21oi_1 _08772_ (.A1(_03178_),
    .A2(_03285_),
    .Y(_03297_),
    .B1(_03284_));
 sg13g2_o21ai_1 _08773_ (.B1(_03225_),
    .Y(_03298_),
    .A1(_03226_),
    .A2(_03282_));
 sg13g2_nor2_1 _08774_ (.A(net1118),
    .B(_03221_),
    .Y(_03299_));
 sg13g2_a22oi_1 _08775_ (.Y(_03300_),
    .B1(_03299_),
    .B2(_03087_),
    .A2(_03223_),
    .A1(_03214_));
 sg13g2_a21o_1 _08776_ (.A2(_03191_),
    .A1(_03182_),
    .B1(_03190_),
    .X(_03301_));
 sg13g2_o21ai_1 _08777_ (.B1(_03187_),
    .Y(_03302_),
    .A1(_03184_),
    .A2(_03188_));
 sg13g2_a21oi_1 _08778_ (.A1(net1395),
    .A2(net1117),
    .Y(_03303_),
    .B1(_03218_));
 sg13g2_nand2_1 _08779_ (.Y(_03304_),
    .A(net1357),
    .B(net1336));
 sg13g2_nand2_1 _08780_ (.Y(_03305_),
    .A(net1358),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ));
 sg13g2_nand2_1 _08781_ (.Y(_03306_),
    .A(net1358),
    .B(net1333));
 sg13g2_or2_1 _08782_ (.X(_03307_),
    .B(_03305_),
    .A(_03186_));
 sg13g2_xnor2_1 _08783_ (.Y(_03308_),
    .A(_03185_),
    .B(_03306_));
 sg13g2_xor2_1 _08784_ (.B(_03308_),
    .A(_03304_),
    .X(_03309_));
 sg13g2_nor2b_1 _08785_ (.A(_03303_),
    .B_N(_03309_),
    .Y(_03310_));
 sg13g2_xnor2_1 _08786_ (.Y(_03311_),
    .A(_03303_),
    .B(_03309_));
 sg13g2_xnor2_1 _08787_ (.Y(_03312_),
    .A(_03302_),
    .B(_03311_));
 sg13g2_nand2b_1 _08788_ (.Y(_03313_),
    .B(_03301_),
    .A_N(_03312_));
 sg13g2_xor2_1 _08789_ (.B(_03312_),
    .A(_03301_),
    .X(_03314_));
 sg13g2_nand2_1 _08790_ (.Y(_03315_),
    .A(net1447),
    .B(net1158));
 sg13g2_nand2_2 _08791_ (.Y(_03316_),
    .A(net1452),
    .B(net1152));
 sg13g2_xor2_1 _08792_ (.B(_03316_),
    .A(_03196_),
    .X(_03317_));
 sg13g2_nand2b_1 _08793_ (.Y(_03318_),
    .B(_03317_),
    .A_N(_03315_));
 sg13g2_xor2_1 _08794_ (.B(_03317_),
    .A(_03315_),
    .X(_03319_));
 sg13g2_o21ai_1 _08795_ (.B1(_03206_),
    .Y(_03320_),
    .A1(_03068_),
    .A2(_03204_));
 sg13g2_nand2_1 _08796_ (.Y(_03321_),
    .A(net1461),
    .B(net1350));
 sg13g2_nand2_1 _08797_ (.Y(_03322_),
    .A(net1465),
    .B(net1338));
 sg13g2_nand2_1 _08798_ (.Y(_03323_),
    .A(net1466),
    .B(net1343));
 sg13g2_xor2_1 _08799_ (.B(_03323_),
    .A(_03203_),
    .X(_03324_));
 sg13g2_nand2b_1 _08800_ (.Y(_03325_),
    .B(_03324_),
    .A_N(_03321_));
 sg13g2_xnor2_1 _08801_ (.Y(_03326_),
    .A(_03321_),
    .B(_03324_));
 sg13g2_nand2_1 _08802_ (.Y(_03327_),
    .A(_03320_),
    .B(_03326_));
 sg13g2_xnor2_1 _08803_ (.Y(_03328_),
    .A(_03320_),
    .B(_03326_));
 sg13g2_xnor2_1 _08804_ (.Y(_03329_),
    .A(_03319_),
    .B(_03328_));
 sg13g2_xor2_1 _08805_ (.B(_03329_),
    .A(_03314_),
    .X(_03330_));
 sg13g2_o21ai_1 _08806_ (.B1(_03193_),
    .Y(_03331_),
    .A1(_03194_),
    .A2(_03210_));
 sg13g2_nand2_1 _08807_ (.Y(_03332_),
    .A(_03330_),
    .B(_03331_));
 sg13g2_xor2_1 _08808_ (.B(_03331_),
    .A(_03330_),
    .X(_03333_));
 sg13g2_and2_1 _08809_ (.A(net1379),
    .B(net1324),
    .X(_03334_));
 sg13g2_nand3_1 _08810_ (.B(net1379),
    .C(net1324),
    .A(net1394),
    .Y(_03335_));
 sg13g2_o21ai_1 _08811_ (.B1(_03335_),
    .Y(_03336_),
    .A1(net1117),
    .A2(_03334_));
 sg13g2_nand2_1 _08812_ (.Y(_03337_),
    .A(net1372),
    .B(net1327));
 sg13g2_nor2_1 _08813_ (.A(_03336_),
    .B(_03337_),
    .Y(_03338_));
 sg13g2_xor2_1 _08814_ (.B(_03337_),
    .A(_03336_),
    .X(_03339_));
 sg13g2_nand2_1 _08815_ (.Y(_03340_),
    .A(_03084_),
    .B(_03339_));
 sg13g2_xnor2_1 _08816_ (.Y(_03341_),
    .A(_03085_),
    .B(_03339_));
 sg13g2_nor2b_1 _08817_ (.A(_03220_),
    .B_N(_03341_),
    .Y(_03342_));
 sg13g2_xnor2_1 _08818_ (.Y(_03343_),
    .A(_03220_),
    .B(_03341_));
 sg13g2_inv_1 _08819_ (.Y(_03344_),
    .A(_03343_));
 sg13g2_xor2_1 _08820_ (.B(_03343_),
    .A(_03299_),
    .X(_03345_));
 sg13g2_xor2_1 _08821_ (.B(_03345_),
    .A(_03333_),
    .X(_03346_));
 sg13g2_nand2b_1 _08822_ (.Y(_03347_),
    .B(_03346_),
    .A_N(_03300_));
 sg13g2_xor2_1 _08823_ (.B(_03346_),
    .A(_03300_),
    .X(_03348_));
 sg13g2_o21ai_1 _08824_ (.B1(_03278_),
    .Y(_03349_),
    .A1(_03229_),
    .A2(_03245_));
 sg13g2_a21o_2 _08825_ (.A2(_03242_),
    .A1(_03231_),
    .B1(_03244_),
    .X(_03350_));
 sg13g2_a21o_2 _08826_ (.A2(_03239_),
    .A1(_03233_),
    .B1(_03241_),
    .X(_03351_));
 sg13g2_inv_1 _08827_ (.Y(_03352_),
    .A(_03351_));
 sg13g2_o21ai_1 _08828_ (.B1(_03208_),
    .Y(_03353_),
    .A1(_03200_),
    .A2(_03209_));
 sg13g2_o21ai_1 _08829_ (.B1(_03238_),
    .Y(_03354_),
    .A1(_03133_),
    .A2(_03236_));
 sg13g2_o21ai_1 _08830_ (.B1(_03198_),
    .Y(_03355_),
    .A1(_03195_),
    .A2(_03199_));
 sg13g2_nand2_1 _08831_ (.Y(_03356_),
    .A(net1433),
    .B(net1173));
 sg13g2_nand2_1 _08832_ (.Y(_03357_),
    .A(net1437),
    .B(net1162));
 sg13g2_nand2_1 _08833_ (.Y(_03358_),
    .A(net1437),
    .B(net1167));
 sg13g2_xor2_1 _08834_ (.B(_03358_),
    .A(_03235_),
    .X(_03359_));
 sg13g2_nand2b_1 _08835_ (.Y(_03360_),
    .B(_03359_),
    .A_N(_03356_));
 sg13g2_xnor2_1 _08836_ (.Y(_03361_),
    .A(_03356_),
    .B(_03359_));
 sg13g2_xnor2_1 _08837_ (.Y(_03362_),
    .A(_03355_),
    .B(_03361_));
 sg13g2_nor2b_1 _08838_ (.A(_03362_),
    .B_N(_03354_),
    .Y(_03363_));
 sg13g2_xor2_1 _08839_ (.B(_03362_),
    .A(_03354_),
    .X(_03364_));
 sg13g2_nand2b_1 _08840_ (.Y(_03365_),
    .B(_03353_),
    .A_N(_03364_));
 sg13g2_xor2_1 _08841_ (.B(_03364_),
    .A(_03353_),
    .X(_03366_));
 sg13g2_xnor2_1 _08842_ (.Y(_03367_),
    .A(_03351_),
    .B(_03366_));
 sg13g2_nand2_1 _08843_ (.Y(_03368_),
    .A(_03350_),
    .B(_03367_));
 sg13g2_xnor2_1 _08844_ (.Y(_03369_),
    .A(_03350_),
    .B(_03367_));
 sg13g2_or2_1 _08845_ (.X(_03370_),
    .B(_03271_),
    .A(_03269_));
 sg13g2_o21ai_1 _08846_ (.B1(_03252_),
    .Y(_03371_),
    .A1(_03108_),
    .A2(_03250_));
 sg13g2_o21ai_1 _08847_ (.B1(net1412),
    .Y(_03372_),
    .A1(net1215),
    .A2(net1208));
 sg13g2_nor2b_1 _08848_ (.A(_03372_),
    .B_N(_03268_),
    .Y(_03373_));
 sg13g2_xnor2_1 _08849_ (.Y(_03374_),
    .A(_02970_),
    .B(_03373_));
 sg13g2_xnor2_1 _08850_ (.Y(_03375_),
    .A(_03371_),
    .B(net1066));
 sg13g2_nor2b_1 _08851_ (.A(_03375_),
    .B_N(_03370_),
    .Y(_03376_));
 sg13g2_xor2_1 _08852_ (.B(_03375_),
    .A(_03370_),
    .X(_03377_));
 sg13g2_o21ai_1 _08853_ (.B1(_03261_),
    .Y(_03378_),
    .A1(_03253_),
    .A2(_03262_));
 sg13g2_nand2_1 _08854_ (.Y(_03379_),
    .A(net1414),
    .B(net1207));
 sg13g2_nand2_1 _08855_ (.Y(_03380_),
    .A(net1416),
    .B(net1200));
 sg13g2_xor2_1 _08856_ (.B(_03380_),
    .A(_03249_),
    .X(_03381_));
 sg13g2_nand2b_1 _08857_ (.Y(_03382_),
    .B(_03381_),
    .A_N(_03379_));
 sg13g2_xor2_1 _08858_ (.B(_03381_),
    .A(_03379_),
    .X(_03383_));
 sg13g2_o21ai_1 _08859_ (.B1(_03259_),
    .Y(_03384_),
    .A1(_03115_),
    .A2(_03257_));
 sg13g2_nand2_1 _08860_ (.Y(_03385_),
    .A(net1422),
    .B(net1193));
 sg13g2_nand2_1 _08861_ (.Y(_03386_),
    .A(net1425),
    .B(net1178));
 sg13g2_nand2_1 _08862_ (.Y(_03387_),
    .A(net1425),
    .B(net1190));
 sg13g2_xor2_1 _08863_ (.B(_03387_),
    .A(_03256_),
    .X(_03388_));
 sg13g2_nand2b_1 _08864_ (.Y(_03389_),
    .B(_03388_),
    .A_N(_03385_));
 sg13g2_xnor2_1 _08865_ (.Y(_03390_),
    .A(_03385_),
    .B(_03388_));
 sg13g2_nand2_1 _08866_ (.Y(_03391_),
    .A(_03384_),
    .B(_03390_));
 sg13g2_xnor2_1 _08867_ (.Y(_03392_),
    .A(_03384_),
    .B(_03390_));
 sg13g2_xor2_1 _08868_ (.B(_03392_),
    .A(_03383_),
    .X(_03393_));
 sg13g2_nand2_1 _08869_ (.Y(_03394_),
    .A(_03378_),
    .B(_03393_));
 sg13g2_xnor2_1 _08870_ (.Y(_03395_),
    .A(_03378_),
    .B(_03393_));
 sg13g2_xor2_1 _08871_ (.B(_03395_),
    .A(_03377_),
    .X(_03396_));
 sg13g2_inv_1 _08872_ (.Y(_03397_),
    .A(_03396_));
 sg13g2_xnor2_1 _08873_ (.Y(_03398_),
    .A(_03369_),
    .B(_03396_));
 sg13g2_nor2b_1 _08874_ (.A(_03213_),
    .B_N(_03398_),
    .Y(_03399_));
 sg13g2_xnor2_1 _08875_ (.Y(_03400_),
    .A(_03213_),
    .B(_03398_));
 sg13g2_xnor2_1 _08876_ (.Y(_03401_),
    .A(_03349_),
    .B(_03400_));
 sg13g2_xnor2_1 _08877_ (.Y(_03402_),
    .A(_03348_),
    .B(_03401_));
 sg13g2_nor2b_1 _08878_ (.A(_03402_),
    .B_N(_03298_),
    .Y(_03403_));
 sg13g2_nand2b_1 _08879_ (.Y(_03404_),
    .B(_03402_),
    .A_N(_03298_));
 sg13g2_xor2_1 _08880_ (.B(_03402_),
    .A(_03298_),
    .X(_03405_));
 sg13g2_a21o_1 _08881_ (.A2(_03273_),
    .A1(_03267_),
    .B1(_03275_),
    .X(_03406_));
 sg13g2_a21oi_1 _08882_ (.A1(_03078_),
    .A2(_03279_),
    .Y(_03407_),
    .B1(_03281_));
 sg13g2_o21ai_1 _08883_ (.B1(_03264_),
    .Y(_03408_),
    .A1(_03265_),
    .A2(_03276_));
 sg13g2_nand2b_1 _08884_ (.Y(_03409_),
    .B(_03408_),
    .A_N(_03407_));
 sg13g2_xor2_1 _08885_ (.B(_03408_),
    .A(_03407_),
    .X(_03410_));
 sg13g2_nand2b_1 _08886_ (.Y(_03411_),
    .B(_03406_),
    .A_N(_03410_));
 sg13g2_xnor2_1 _08887_ (.Y(_03412_),
    .A(_03406_),
    .B(_03410_));
 sg13g2_xnor2_1 _08888_ (.Y(_03413_),
    .A(_03405_),
    .B(_03412_));
 sg13g2_nor2b_1 _08889_ (.A(_03297_),
    .B_N(_03413_),
    .Y(_03414_));
 sg13g2_xnor2_1 _08890_ (.Y(_03415_),
    .A(_03297_),
    .B(_03413_));
 sg13g2_xnor2_1 _08891_ (.Y(_03416_),
    .A(_03296_),
    .B(_03415_));
 sg13g2_a21o_1 _08892_ (.A2(_03288_),
    .A1(_03171_),
    .B1(_03287_),
    .X(_03417_));
 sg13g2_nand2b_1 _08893_ (.Y(_03418_),
    .B(_03417_),
    .A_N(_03416_));
 sg13g2_xnor2_1 _08894_ (.Y(_03419_),
    .A(_03416_),
    .B(_03417_));
 sg13g2_inv_1 _08895_ (.Y(_03420_),
    .A(_03419_));
 sg13g2_and2_1 _08896_ (.A(_03161_),
    .B(_03292_),
    .X(_03421_));
 sg13g2_o21ai_1 _08897_ (.B1(_03291_),
    .Y(_03422_),
    .A1(_03159_),
    .A2(_03290_));
 sg13g2_a21oi_1 _08898_ (.A1(_03167_),
    .A2(_03421_),
    .Y(_03423_),
    .B1(_03422_));
 sg13g2_xnor2_1 _08899_ (.Y(_03424_),
    .A(_03419_),
    .B(_03423_));
 sg13g2_o21ai_1 _08900_ (.B1(net1509),
    .Y(_03425_),
    .A1(net1142),
    .A2(_03424_));
 sg13g2_a21oi_1 _08901_ (.A1(net1142),
    .A2(_04774_),
    .Y(_00238_),
    .B1(_03425_));
 sg13g2_a21o_1 _08902_ (.A2(_03415_),
    .A1(_03296_),
    .B1(_03414_),
    .X(_03426_));
 sg13g2_nand2_1 _08903_ (.Y(_03427_),
    .A(_03409_),
    .B(_03411_));
 sg13g2_a21oi_1 _08904_ (.A1(_03404_),
    .A2(_03412_),
    .Y(_03428_),
    .B1(_03403_));
 sg13g2_o21ai_1 _08905_ (.B1(_03347_),
    .Y(_03429_),
    .A1(_03348_),
    .A2(_03401_));
 sg13g2_nor2_1 _08906_ (.A(_03081_),
    .B(_03343_),
    .Y(_03430_));
 sg13g2_a22oi_1 _08907_ (.Y(_03431_),
    .B1(_03430_),
    .B2(_03221_),
    .A2(_03345_),
    .A1(_03333_));
 sg13g2_o21ai_1 _08908_ (.B1(_03313_),
    .Y(_03432_),
    .A1(_03314_),
    .A2(_03329_));
 sg13g2_a21o_1 _08909_ (.A2(_03311_),
    .A1(_03302_),
    .B1(_03310_),
    .X(_03433_));
 sg13g2_o21ai_1 _08910_ (.B1(_03307_),
    .Y(_03434_),
    .A1(_03304_),
    .A2(_03308_));
 sg13g2_a21oi_1 _08911_ (.A1(net1379),
    .A2(_03215_),
    .Y(_03435_),
    .B1(_03338_));
 sg13g2_nand2_1 _08912_ (.Y(_03436_),
    .A(net1470),
    .B(net1334));
 sg13g2_nand2_1 _08913_ (.Y(_03437_),
    .A(net1352),
    .B(net1329));
 sg13g2_nand2_1 _08914_ (.Y(_03438_),
    .A(net1352),
    .B(net1331));
 sg13g2_or2_1 _08915_ (.X(_03439_),
    .B(_03437_),
    .A(_03306_));
 sg13g2_xnor2_1 _08916_ (.Y(_03440_),
    .A(_03305_),
    .B(_03438_));
 sg13g2_xor2_1 _08917_ (.B(_03440_),
    .A(_03436_),
    .X(_03441_));
 sg13g2_nor2b_1 _08918_ (.A(_03435_),
    .B_N(_03441_),
    .Y(_03442_));
 sg13g2_xnor2_1 _08919_ (.Y(_03443_),
    .A(_03435_),
    .B(_03441_));
 sg13g2_xor2_1 _08920_ (.B(_03443_),
    .A(_03434_),
    .X(_03444_));
 sg13g2_nand2_1 _08921_ (.Y(_03445_),
    .A(_03433_),
    .B(_03444_));
 sg13g2_xnor2_1 _08922_ (.Y(_03446_),
    .A(_03433_),
    .B(_03444_));
 sg13g2_nand2_1 _08923_ (.Y(_03447_),
    .A(net1442),
    .B(net1158));
 sg13g2_nand2_2 _08924_ (.Y(_03448_),
    .A(net1447),
    .B(net1146));
 sg13g2_nor2_1 _08925_ (.A(_03316_),
    .B(_03448_),
    .Y(_03449_));
 sg13g2_or2_1 _08926_ (.X(_03450_),
    .B(_03448_),
    .A(_03316_));
 sg13g2_a22oi_1 _08927_ (.Y(_03451_),
    .B1(net1146),
    .B2(net1452),
    .A2(net1152),
    .A1(net1447));
 sg13g2_or2_1 _08928_ (.X(_03452_),
    .B(_03451_),
    .A(_03449_));
 sg13g2_xnor2_1 _08929_ (.Y(_03453_),
    .A(_03447_),
    .B(_03452_));
 sg13g2_o21ai_1 _08930_ (.B1(_03325_),
    .Y(_03454_),
    .A1(_03203_),
    .A2(_03323_));
 sg13g2_nand2_1 _08931_ (.Y(_03455_),
    .A(net1456),
    .B(net1351));
 sg13g2_nand2_1 _08932_ (.Y(_03456_),
    .A(net1461),
    .B(net1338));
 sg13g2_nand2_1 _08933_ (.Y(_03457_),
    .A(net1460),
    .B(net1343));
 sg13g2_xor2_1 _08934_ (.B(_03457_),
    .A(_03322_),
    .X(_03458_));
 sg13g2_nand2b_1 _08935_ (.Y(_03459_),
    .B(_03458_),
    .A_N(_03455_));
 sg13g2_xnor2_1 _08936_ (.Y(_03460_),
    .A(_03455_),
    .B(_03458_));
 sg13g2_nand2_1 _08937_ (.Y(_03461_),
    .A(_03454_),
    .B(_03460_));
 sg13g2_xnor2_1 _08938_ (.Y(_03462_),
    .A(_03454_),
    .B(_03460_));
 sg13g2_xnor2_1 _08939_ (.Y(_03463_),
    .A(_03453_),
    .B(_03462_));
 sg13g2_xor2_1 _08940_ (.B(_03463_),
    .A(_03446_),
    .X(_03464_));
 sg13g2_xnor2_1 _08941_ (.Y(_03465_),
    .A(_03342_),
    .B(_03464_));
 sg13g2_nor2b_1 _08942_ (.A(_03465_),
    .B_N(_03432_),
    .Y(_03466_));
 sg13g2_xor2_1 _08943_ (.B(_03465_),
    .A(_03432_),
    .X(_03467_));
 sg13g2_nand2_1 _08944_ (.Y(_03468_),
    .A(net1103),
    .B(net1117));
 sg13g2_inv_2 _08945_ (.Y(_03469_),
    .A(_03468_));
 sg13g2_and2_1 _08946_ (.A(_03084_),
    .B(net1117),
    .X(_03470_));
 sg13g2_xnor2_1 _08947_ (.Y(_03471_),
    .A(_03084_),
    .B(net1117));
 sg13g2_a21oi_2 _08948_ (.B1(_03469_),
    .Y(_03472_),
    .A2(_03471_),
    .A1(_03083_));
 sg13g2_and2_1 _08949_ (.A(net1372),
    .B(net1324),
    .X(_03473_));
 sg13g2_nand2_1 _08950_ (.Y(_03474_),
    .A(net1372),
    .B(net1325));
 sg13g2_nand2_1 _08951_ (.Y(_03475_),
    .A(net1372),
    .B(_03334_));
 sg13g2_o21ai_1 _08952_ (.B1(_03475_),
    .Y(_03476_),
    .A1(_03334_),
    .A2(_03473_));
 sg13g2_nand2_1 _08953_ (.Y(_03477_),
    .A(net1365),
    .B(net1326));
 sg13g2_nor2_1 _08954_ (.A(_03476_),
    .B(_03477_),
    .Y(_03478_));
 sg13g2_xor2_1 _08955_ (.B(_03477_),
    .A(_03476_),
    .X(_03479_));
 sg13g2_xnor2_1 _08956_ (.Y(_03480_),
    .A(_03472_),
    .B(_03479_));
 sg13g2_nor2_1 _08957_ (.A(_03340_),
    .B(_03480_),
    .Y(_03481_));
 sg13g2_xor2_1 _08958_ (.B(_03480_),
    .A(_03340_),
    .X(_03482_));
 sg13g2_xnor2_1 _08959_ (.Y(_03483_),
    .A(_03430_),
    .B(_03482_));
 sg13g2_nor2_1 _08960_ (.A(_03467_),
    .B(_03483_),
    .Y(_03484_));
 sg13g2_xnor2_1 _08961_ (.Y(_03485_),
    .A(_03467_),
    .B(_03483_));
 sg13g2_nor2_1 _08962_ (.A(_03431_),
    .B(_03485_),
    .Y(_03486_));
 sg13g2_xor2_1 _08963_ (.B(_03485_),
    .A(_03431_),
    .X(_03487_));
 sg13g2_o21ai_1 _08964_ (.B1(_03368_),
    .Y(_03488_),
    .A1(_03369_),
    .A2(_03397_));
 sg13g2_o21ai_1 _08965_ (.B1(_03268_),
    .Y(_03489_),
    .A1(_02970_),
    .A2(_03372_));
 sg13g2_o21ai_1 _08966_ (.B1(_03382_),
    .Y(_03490_),
    .A1(_03249_),
    .A2(_03380_));
 sg13g2_and2_1 _08967_ (.A(net1066),
    .B(_03490_),
    .X(_03491_));
 sg13g2_xor2_1 _08968_ (.B(_03490_),
    .A(_03374_),
    .X(_03492_));
 sg13g2_xnor2_1 _08969_ (.Y(_03493_),
    .A(_03489_),
    .B(_03492_));
 sg13g2_o21ai_1 _08970_ (.B1(_03391_),
    .Y(_03494_),
    .A1(_03383_),
    .A2(_03392_));
 sg13g2_nand2_2 _08971_ (.Y(_03495_),
    .A(net1412),
    .B(net1207));
 sg13g2_nor3_1 _08972_ (.A(_04821_),
    .B(_04828_),
    .C(_03380_),
    .Y(_03496_));
 sg13g2_a22oi_1 _08973_ (.Y(_03497_),
    .B1(net1195),
    .B2(net1416),
    .A2(net1200),
    .A1(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ));
 sg13g2_nor3_1 _08974_ (.A(_03495_),
    .B(_03496_),
    .C(_03497_),
    .Y(_03498_));
 sg13g2_o21ai_1 _08975_ (.B1(_03495_),
    .Y(_03499_),
    .A1(_03496_),
    .A2(_03497_));
 sg13g2_nor2b_1 _08976_ (.A(_03498_),
    .B_N(_03499_),
    .Y(_03500_));
 sg13g2_inv_1 _08977_ (.Y(_03501_),
    .A(_03500_));
 sg13g2_o21ai_1 _08978_ (.B1(_03389_),
    .Y(_03502_),
    .A1(_03256_),
    .A2(_03387_));
 sg13g2_nand2_1 _08979_ (.Y(_03503_),
    .A(net1419),
    .B(net1193));
 sg13g2_nand2_1 _08980_ (.Y(_03504_),
    .A(net1423),
    .B(net1178));
 sg13g2_nand2_1 _08981_ (.Y(_03505_),
    .A(net1423),
    .B(net1184));
 sg13g2_xor2_1 _08982_ (.B(_03505_),
    .A(_03386_),
    .X(_03506_));
 sg13g2_nand2b_1 _08983_ (.Y(_03507_),
    .B(_03506_),
    .A_N(_03503_));
 sg13g2_xnor2_1 _08984_ (.Y(_03508_),
    .A(_03503_),
    .B(_03506_));
 sg13g2_nand2_1 _08985_ (.Y(_03509_),
    .A(_03502_),
    .B(_03508_));
 sg13g2_xnor2_1 _08986_ (.Y(_03510_),
    .A(_03502_),
    .B(_03508_));
 sg13g2_xnor2_1 _08987_ (.Y(_03511_),
    .A(_03501_),
    .B(_03510_));
 sg13g2_nand2b_1 _08988_ (.Y(_03512_),
    .B(_03494_),
    .A_N(_03511_));
 sg13g2_xor2_1 _08989_ (.B(_03511_),
    .A(_03494_),
    .X(_03513_));
 sg13g2_xor2_1 _08990_ (.B(_03513_),
    .A(_03493_),
    .X(_03514_));
 sg13g2_inv_1 _08991_ (.Y(_03515_),
    .A(_03514_));
 sg13g2_o21ai_1 _08992_ (.B1(_03365_),
    .Y(_03516_),
    .A1(_03352_),
    .A2(_03366_));
 sg13g2_a21o_1 _08993_ (.A2(_03361_),
    .A1(_03355_),
    .B1(_03363_),
    .X(_03517_));
 sg13g2_o21ai_1 _08994_ (.B1(_03327_),
    .Y(_03518_),
    .A1(_03319_),
    .A2(_03328_));
 sg13g2_inv_1 _08995_ (.Y(_03519_),
    .A(_03518_));
 sg13g2_o21ai_1 _08996_ (.B1(_03360_),
    .Y(_03520_),
    .A1(_03235_),
    .A2(_03358_));
 sg13g2_o21ai_1 _08997_ (.B1(_03318_),
    .Y(_03521_),
    .A1(_03196_),
    .A2(_03316_));
 sg13g2_nand2_1 _08998_ (.Y(_03522_),
    .A(net1429),
    .B(net1173));
 sg13g2_nand2_1 _08999_ (.Y(_03523_),
    .A(net1433),
    .B(net1162));
 sg13g2_nand2_1 _09000_ (.Y(_03524_),
    .A(net1433),
    .B(net1168));
 sg13g2_xor2_1 _09001_ (.B(_03524_),
    .A(_03357_),
    .X(_03525_));
 sg13g2_nand2b_1 _09002_ (.Y(_03526_),
    .B(_03525_),
    .A_N(_03522_));
 sg13g2_xnor2_1 _09003_ (.Y(_03527_),
    .A(_03522_),
    .B(_03525_));
 sg13g2_xnor2_1 _09004_ (.Y(_03528_),
    .A(_03521_),
    .B(_03527_));
 sg13g2_nor2b_1 _09005_ (.A(_03528_),
    .B_N(_03520_),
    .Y(_03529_));
 sg13g2_xor2_1 _09006_ (.B(_03528_),
    .A(_03520_),
    .X(_03530_));
 sg13g2_xor2_1 _09007_ (.B(_03530_),
    .A(_03518_),
    .X(_03531_));
 sg13g2_nand2b_1 _09008_ (.Y(_03532_),
    .B(_03517_),
    .A_N(_03531_));
 sg13g2_xor2_1 _09009_ (.B(_03531_),
    .A(_03517_),
    .X(_03533_));
 sg13g2_nor2b_1 _09010_ (.A(_03533_),
    .B_N(_03516_),
    .Y(_03534_));
 sg13g2_xor2_1 _09011_ (.B(_03533_),
    .A(_03516_),
    .X(_03535_));
 sg13g2_nor2_1 _09012_ (.A(_03515_),
    .B(_03535_),
    .Y(_03536_));
 sg13g2_xnor2_1 _09013_ (.Y(_03537_),
    .A(_03515_),
    .B(_03535_));
 sg13g2_xor2_1 _09014_ (.B(_03537_),
    .A(_03332_),
    .X(_03538_));
 sg13g2_nand2_1 _09015_ (.Y(_03539_),
    .A(_03488_),
    .B(_03538_));
 sg13g2_xor2_1 _09016_ (.B(_03538_),
    .A(_03488_),
    .X(_03540_));
 sg13g2_xnor2_1 _09017_ (.Y(_03541_),
    .A(_03487_),
    .B(_03540_));
 sg13g2_nor2b_1 _09018_ (.A(_03541_),
    .B_N(_03429_),
    .Y(_03542_));
 sg13g2_nand2b_1 _09019_ (.Y(_03543_),
    .B(_03541_),
    .A_N(_03429_));
 sg13g2_xor2_1 _09020_ (.B(_03541_),
    .A(_03429_),
    .X(_03544_));
 sg13g2_a21o_1 _09021_ (.A2(_03374_),
    .A1(_03371_),
    .B1(_03376_),
    .X(_03545_));
 sg13g2_a21oi_1 _09022_ (.A1(_03349_),
    .A2(_03400_),
    .Y(_03546_),
    .B1(_03399_));
 sg13g2_o21ai_1 _09023_ (.B1(_03394_),
    .Y(_03547_),
    .A1(_03377_),
    .A2(_03395_));
 sg13g2_nand2b_1 _09024_ (.Y(_03548_),
    .B(_03547_),
    .A_N(_03546_));
 sg13g2_xor2_1 _09025_ (.B(_03547_),
    .A(_03546_),
    .X(_03549_));
 sg13g2_nand2b_1 _09026_ (.Y(_03550_),
    .B(_03545_),
    .A_N(_03549_));
 sg13g2_xnor2_1 _09027_ (.Y(_03551_),
    .A(_03545_),
    .B(_03549_));
 sg13g2_xnor2_1 _09028_ (.Y(_03552_),
    .A(_03544_),
    .B(_03551_));
 sg13g2_nor2b_1 _09029_ (.A(_03428_),
    .B_N(_03552_),
    .Y(_03553_));
 sg13g2_xnor2_1 _09030_ (.Y(_03554_),
    .A(_03428_),
    .B(_03552_));
 sg13g2_xnor2_1 _09031_ (.Y(_03555_),
    .A(_03427_),
    .B(_03554_));
 sg13g2_nand2b_1 _09032_ (.Y(_03556_),
    .B(_03426_),
    .A_N(_03555_));
 sg13g2_nand2b_1 _09033_ (.Y(_03557_),
    .B(_03555_),
    .A_N(_03426_));
 sg13g2_xnor2_1 _09034_ (.Y(_03558_),
    .A(_03426_),
    .B(_03555_));
 sg13g2_o21ai_1 _09035_ (.B1(_03418_),
    .Y(_03559_),
    .A1(_03420_),
    .A2(_03423_));
 sg13g2_xor2_1 _09036_ (.B(_03559_),
    .A(_03558_),
    .X(_03560_));
 sg13g2_o21ai_1 _09037_ (.B1(net1509),
    .Y(_03561_),
    .A1(net1142),
    .A2(_03560_));
 sg13g2_a21oi_1 _09038_ (.A1(net1142),
    .A2(_04773_),
    .Y(_00239_),
    .B1(_03561_));
 sg13g2_and2_1 _09039_ (.A(_03419_),
    .B(_03558_),
    .X(_03562_));
 sg13g2_and4_1 _09040_ (.A(_03161_),
    .B(_03292_),
    .C(_03419_),
    .D(_03558_),
    .X(_03563_));
 sg13g2_o21ai_1 _09041_ (.B1(_03563_),
    .Y(_03564_),
    .A1(_03164_),
    .A2(_03166_));
 sg13g2_nand2_1 _09042_ (.Y(_03565_),
    .A(_03418_),
    .B(_03556_));
 sg13g2_a22oi_1 _09043_ (.Y(_03566_),
    .B1(_03565_),
    .B2(_03557_),
    .A2(_03562_),
    .A1(_03422_));
 sg13g2_nand2_1 _09044_ (.Y(_03567_),
    .A(_03564_),
    .B(_03566_));
 sg13g2_nand2_1 _09045_ (.Y(_03568_),
    .A(_03548_),
    .B(_03550_));
 sg13g2_a21oi_1 _09046_ (.A1(_03543_),
    .A2(_03551_),
    .Y(_03569_),
    .B1(_03542_));
 sg13g2_a21oi_1 _09047_ (.A1(_03487_),
    .A2(_03540_),
    .Y(_03570_),
    .B1(_03486_));
 sg13g2_nor3_1 _09048_ (.A(_03081_),
    .B(_03344_),
    .C(_03482_),
    .Y(_03571_));
 sg13g2_nor2_1 _09049_ (.A(_03484_),
    .B(_03571_),
    .Y(_03572_));
 sg13g2_nand2_1 _09050_ (.Y(_03573_),
    .A(_03080_),
    .B(_03482_));
 sg13g2_nand2_1 _09051_ (.Y(_03574_),
    .A(_02955_),
    .B(net1118));
 sg13g2_xnor2_1 _09052_ (.Y(_03575_),
    .A(_02954_),
    .B(net1118));
 sg13g2_inv_1 _09053_ (.Y(_03576_),
    .A(_03575_));
 sg13g2_nor2_2 _09054_ (.A(net1103),
    .B(_03470_),
    .Y(_03577_));
 sg13g2_nor2b_1 _09055_ (.A(_03216_),
    .B_N(_03334_),
    .Y(_03578_));
 sg13g2_xnor2_1 _09056_ (.Y(_03579_),
    .A(_03216_),
    .B(_03334_));
 sg13g2_o21ai_1 _09057_ (.B1(_03579_),
    .Y(_03580_),
    .A1(net1103),
    .A2(_03470_));
 sg13g2_xnor2_1 _09058_ (.Y(_03581_),
    .A(_03577_),
    .B(_03579_));
 sg13g2_and2_1 _09059_ (.A(net1365),
    .B(net1323),
    .X(_03582_));
 sg13g2_nand2_1 _09060_ (.Y(_03583_),
    .A(net1365),
    .B(net1323));
 sg13g2_nand2_1 _09061_ (.Y(_03584_),
    .A(net1365),
    .B(_03473_));
 sg13g2_o21ai_1 _09062_ (.B1(_03584_),
    .Y(_03585_),
    .A1(_03473_),
    .A2(_03582_));
 sg13g2_nand2_1 _09063_ (.Y(_03586_),
    .A(net1358),
    .B(net1327));
 sg13g2_nor2_1 _09064_ (.A(_03585_),
    .B(_03586_),
    .Y(_03587_));
 sg13g2_xor2_1 _09065_ (.B(_03586_),
    .A(_03585_),
    .X(_03588_));
 sg13g2_nand2_1 _09066_ (.Y(_03589_),
    .A(_03581_),
    .B(_03588_));
 sg13g2_xnor2_1 _09067_ (.Y(_03590_),
    .A(_03581_),
    .B(_03588_));
 sg13g2_a21o_1 _09068_ (.A2(_03479_),
    .A1(_03472_),
    .B1(_03469_),
    .X(_03591_));
 sg13g2_nand2b_1 _09069_ (.Y(_03592_),
    .B(_03591_),
    .A_N(_03590_));
 sg13g2_xor2_1 _09070_ (.B(_03591_),
    .A(_03590_),
    .X(_03593_));
 sg13g2_nor2_1 _09071_ (.A(_03576_),
    .B(_03593_),
    .Y(_03594_));
 sg13g2_xnor2_1 _09072_ (.Y(_03595_),
    .A(_03576_),
    .B(_03593_));
 sg13g2_or2_1 _09073_ (.X(_03596_),
    .B(_03595_),
    .A(_03573_));
 sg13g2_xnor2_1 _09074_ (.Y(_03597_),
    .A(_03573_),
    .B(_03595_));
 sg13g2_o21ai_1 _09075_ (.B1(_03445_),
    .Y(_03598_),
    .A1(_03446_),
    .A2(_03463_));
 sg13g2_a21o_1 _09076_ (.A2(_03443_),
    .A1(_03434_),
    .B1(_03442_),
    .X(_03599_));
 sg13g2_o21ai_1 _09077_ (.B1(_03439_),
    .Y(_03600_),
    .A1(_03436_),
    .A2(_03440_));
 sg13g2_a21oi_1 _09078_ (.A1(net1379),
    .A2(_03473_),
    .Y(_03601_),
    .B1(_03478_));
 sg13g2_nand2_1 _09079_ (.Y(_03602_),
    .A(net1465),
    .B(net1334));
 sg13g2_nand2_1 _09080_ (.Y(_03603_),
    .A(net1470),
    .B(net1329));
 sg13g2_nand2_1 _09081_ (.Y(_03604_),
    .A(net1470),
    .B(net1332));
 sg13g2_or2_1 _09082_ (.X(_03605_),
    .B(_03603_),
    .A(_03438_));
 sg13g2_xnor2_1 _09083_ (.Y(_03606_),
    .A(_03437_),
    .B(_03604_));
 sg13g2_xor2_1 _09084_ (.B(_03606_),
    .A(_03602_),
    .X(_03607_));
 sg13g2_nor2b_1 _09085_ (.A(_03601_),
    .B_N(_03607_),
    .Y(_03608_));
 sg13g2_xnor2_1 _09086_ (.Y(_03609_),
    .A(_03601_),
    .B(_03607_));
 sg13g2_xnor2_1 _09087_ (.Y(_03610_),
    .A(_03600_),
    .B(_03609_));
 sg13g2_nand2b_1 _09088_ (.Y(_03611_),
    .B(_03599_),
    .A_N(_03610_));
 sg13g2_xor2_1 _09089_ (.B(_03610_),
    .A(_03599_),
    .X(_03612_));
 sg13g2_nand2_1 _09090_ (.Y(_03613_),
    .A(net1437),
    .B(net1158));
 sg13g2_nand2_1 _09091_ (.Y(_03614_),
    .A(net1441),
    .B(net1145));
 sg13g2_nand2_1 _09092_ (.Y(_03615_),
    .A(net1442),
    .B(net1152));
 sg13g2_xor2_1 _09093_ (.B(_03615_),
    .A(_03448_),
    .X(_03616_));
 sg13g2_nand2b_1 _09094_ (.Y(_03617_),
    .B(_03616_),
    .A_N(_03613_));
 sg13g2_xor2_1 _09095_ (.B(_03616_),
    .A(_03613_),
    .X(_03618_));
 sg13g2_o21ai_1 _09096_ (.B1(_03459_),
    .Y(_03619_),
    .A1(_03322_),
    .A2(_03457_));
 sg13g2_nand2_1 _09097_ (.Y(_03620_),
    .A(net1452),
    .B(net1351));
 sg13g2_nand2_1 _09098_ (.Y(_03621_),
    .A(net1456),
    .B(net1337));
 sg13g2_nand2_1 _09099_ (.Y(_03622_),
    .A(net1456),
    .B(net1343));
 sg13g2_xor2_1 _09100_ (.B(_03622_),
    .A(_03456_),
    .X(_03623_));
 sg13g2_nand2b_1 _09101_ (.Y(_03624_),
    .B(_03623_),
    .A_N(_03620_));
 sg13g2_xnor2_1 _09102_ (.Y(_03625_),
    .A(_03620_),
    .B(_03623_));
 sg13g2_nand2_1 _09103_ (.Y(_03626_),
    .A(_03619_),
    .B(_03625_));
 sg13g2_xnor2_1 _09104_ (.Y(_03627_),
    .A(_03619_),
    .B(_03625_));
 sg13g2_xnor2_1 _09105_ (.Y(_03628_),
    .A(_03618_),
    .B(_03627_));
 sg13g2_xor2_1 _09106_ (.B(_03628_),
    .A(_03612_),
    .X(_03629_));
 sg13g2_and2_1 _09107_ (.A(_03481_),
    .B(_03629_),
    .X(_03630_));
 sg13g2_xor2_1 _09108_ (.B(_03629_),
    .A(_03481_),
    .X(_03631_));
 sg13g2_xnor2_1 _09109_ (.Y(_03632_),
    .A(_03598_),
    .B(_03631_));
 sg13g2_xnor2_1 _09110_ (.Y(_03633_),
    .A(_03597_),
    .B(_03632_));
 sg13g2_or2_1 _09111_ (.X(_03634_),
    .B(_03633_),
    .A(_03572_));
 sg13g2_xnor2_1 _09112_ (.Y(_03635_),
    .A(_03572_),
    .B(_03633_));
 sg13g2_nor2_1 _09113_ (.A(_03534_),
    .B(_03536_),
    .Y(_03636_));
 sg13g2_a21o_1 _09114_ (.A2(_03464_),
    .A1(_03342_),
    .B1(_03466_),
    .X(_03637_));
 sg13g2_or2_1 _09115_ (.X(_03638_),
    .B(_03498_),
    .A(_03496_));
 sg13g2_and2_1 _09116_ (.A(net1066),
    .B(_03638_),
    .X(_03639_));
 sg13g2_xor2_1 _09117_ (.B(_03638_),
    .A(net1066),
    .X(_03640_));
 sg13g2_xnor2_1 _09118_ (.Y(_03641_),
    .A(_03489_),
    .B(_03640_));
 sg13g2_o21ai_1 _09119_ (.B1(_03509_),
    .Y(_03642_),
    .A1(_03501_),
    .A2(_03510_));
 sg13g2_nand3_1 _09120_ (.B(net1200),
    .C(net1195),
    .A(net1412),
    .Y(_03643_));
 sg13g2_nor2_1 _09121_ (.A(_04821_),
    .B(_03643_),
    .Y(_03644_));
 sg13g2_a22oi_1 _09122_ (.Y(_03645_),
    .B1(net1195),
    .B2(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ),
    .A2(net1200),
    .A1(net1412));
 sg13g2_nor3_1 _09123_ (.A(_03495_),
    .B(_03644_),
    .C(_03645_),
    .Y(_03646_));
 sg13g2_o21ai_1 _09124_ (.B1(_03495_),
    .Y(_03647_),
    .A1(_03644_),
    .A2(_03645_));
 sg13g2_nor2b_1 _09125_ (.A(_03646_),
    .B_N(_03647_),
    .Y(_03648_));
 sg13g2_inv_1 _09126_ (.Y(_03649_),
    .A(_03648_));
 sg13g2_o21ai_1 _09127_ (.B1(_03507_),
    .Y(_03650_),
    .A1(_03386_),
    .A2(_03505_));
 sg13g2_nand2_1 _09128_ (.Y(_03651_),
    .A(net1415),
    .B(net1193));
 sg13g2_nand2_1 _09129_ (.Y(_03652_),
    .A(net1419),
    .B(net1177));
 sg13g2_nand2_1 _09130_ (.Y(_03653_),
    .A(net1419),
    .B(net1184));
 sg13g2_xor2_1 _09131_ (.B(_03653_),
    .A(_03504_),
    .X(_03654_));
 sg13g2_nand2b_1 _09132_ (.Y(_03655_),
    .B(_03654_),
    .A_N(_03651_));
 sg13g2_xnor2_1 _09133_ (.Y(_03656_),
    .A(_03651_),
    .B(_03654_));
 sg13g2_nand2_1 _09134_ (.Y(_03657_),
    .A(_03650_),
    .B(_03656_));
 sg13g2_xnor2_1 _09135_ (.Y(_03658_),
    .A(_03650_),
    .B(_03656_));
 sg13g2_xnor2_1 _09136_ (.Y(_03659_),
    .A(_03648_),
    .B(_03658_));
 sg13g2_nand2_1 _09137_ (.Y(_03660_),
    .A(_03642_),
    .B(_03659_));
 sg13g2_xnor2_1 _09138_ (.Y(_03661_),
    .A(_03642_),
    .B(_03659_));
 sg13g2_xor2_1 _09139_ (.B(_03661_),
    .A(_03641_),
    .X(_03662_));
 sg13g2_inv_1 _09140_ (.Y(_03663_),
    .A(_03662_));
 sg13g2_o21ai_1 _09141_ (.B1(_03532_),
    .Y(_03664_),
    .A1(_03519_),
    .A2(_03530_));
 sg13g2_a21o_1 _09142_ (.A2(_03527_),
    .A1(_03521_),
    .B1(_03529_),
    .X(_03665_));
 sg13g2_o21ai_1 _09143_ (.B1(_03461_),
    .Y(_03666_),
    .A1(_03453_),
    .A2(_03462_));
 sg13g2_o21ai_1 _09144_ (.B1(_03526_),
    .Y(_03667_),
    .A1(_03357_),
    .A2(_03524_));
 sg13g2_o21ai_1 _09145_ (.B1(_03450_),
    .Y(_03668_),
    .A1(_03447_),
    .A2(_03452_));
 sg13g2_nand2_1 _09146_ (.Y(_03669_),
    .A(net1425),
    .B(net1173));
 sg13g2_nand2_1 _09147_ (.Y(_03670_),
    .A(net1428),
    .B(net1161));
 sg13g2_nand2_1 _09148_ (.Y(_03671_),
    .A(net1429),
    .B(net1167));
 sg13g2_xor2_1 _09149_ (.B(_03671_),
    .A(_03523_),
    .X(_03672_));
 sg13g2_nand2b_1 _09150_ (.Y(_03673_),
    .B(_03672_),
    .A_N(_03669_));
 sg13g2_xnor2_1 _09151_ (.Y(_03674_),
    .A(_03669_),
    .B(_03672_));
 sg13g2_xnor2_1 _09152_ (.Y(_03675_),
    .A(_03668_),
    .B(_03674_));
 sg13g2_nor2b_1 _09153_ (.A(_03675_),
    .B_N(_03667_),
    .Y(_03676_));
 sg13g2_xor2_1 _09154_ (.B(_03675_),
    .A(_03667_),
    .X(_03677_));
 sg13g2_nand2b_1 _09155_ (.Y(_03678_),
    .B(_03666_),
    .A_N(_03677_));
 sg13g2_xor2_1 _09156_ (.B(_03677_),
    .A(_03666_),
    .X(_03679_));
 sg13g2_nand2b_1 _09157_ (.Y(_03680_),
    .B(_03665_),
    .A_N(_03679_));
 sg13g2_xor2_1 _09158_ (.B(_03679_),
    .A(_03665_),
    .X(_03681_));
 sg13g2_nand2b_1 _09159_ (.Y(_03682_),
    .B(_03664_),
    .A_N(_03681_));
 sg13g2_xor2_1 _09160_ (.B(_03681_),
    .A(_03664_),
    .X(_03683_));
 sg13g2_xnor2_1 _09161_ (.Y(_03684_),
    .A(_03663_),
    .B(_03683_));
 sg13g2_nand2b_1 _09162_ (.Y(_03685_),
    .B(_03637_),
    .A_N(_03684_));
 sg13g2_xor2_1 _09163_ (.B(_03684_),
    .A(_03637_),
    .X(_03686_));
 sg13g2_xnor2_1 _09164_ (.Y(_03687_),
    .A(_03636_),
    .B(_03686_));
 sg13g2_xnor2_1 _09165_ (.Y(_03688_),
    .A(_03635_),
    .B(_03687_));
 sg13g2_nor2_1 _09166_ (.A(_03570_),
    .B(_03688_),
    .Y(_03689_));
 sg13g2_xor2_1 _09167_ (.B(_03688_),
    .A(_03570_),
    .X(_03690_));
 sg13g2_a21o_1 _09168_ (.A2(_03492_),
    .A1(_03489_),
    .B1(_03491_),
    .X(_03691_));
 sg13g2_o21ai_1 _09169_ (.B1(_03539_),
    .Y(_03692_),
    .A1(_03332_),
    .A2(_03537_));
 sg13g2_o21ai_1 _09170_ (.B1(_03512_),
    .Y(_03693_),
    .A1(_03493_),
    .A2(_03513_));
 sg13g2_xnor2_1 _09171_ (.Y(_03694_),
    .A(_03692_),
    .B(_03693_));
 sg13g2_nor2b_1 _09172_ (.A(_03694_),
    .B_N(_03691_),
    .Y(_03695_));
 sg13g2_xnor2_1 _09173_ (.Y(_03696_),
    .A(_03691_),
    .B(_03694_));
 sg13g2_xnor2_1 _09174_ (.Y(_03697_),
    .A(_03690_),
    .B(_03696_));
 sg13g2_nor2_1 _09175_ (.A(_03569_),
    .B(_03697_),
    .Y(_03698_));
 sg13g2_xor2_1 _09176_ (.B(_03697_),
    .A(_03569_),
    .X(_03699_));
 sg13g2_xnor2_1 _09177_ (.Y(_03700_),
    .A(_03568_),
    .B(_03699_));
 sg13g2_a21o_1 _09178_ (.A2(_03554_),
    .A1(_03427_),
    .B1(_03553_),
    .X(_03701_));
 sg13g2_nor2b_1 _09179_ (.A(_03700_),
    .B_N(_03701_),
    .Y(_03702_));
 sg13g2_xnor2_1 _09180_ (.Y(_03703_),
    .A(_03700_),
    .B(_03701_));
 sg13g2_xnor2_1 _09181_ (.Y(_03704_),
    .A(_03567_),
    .B(_03703_));
 sg13g2_o21ai_1 _09182_ (.B1(net1498),
    .Y(_03705_),
    .A1(net1296),
    .A2(net288));
 sg13g2_a21oi_1 _09183_ (.A1(net1296),
    .A2(_03704_),
    .Y(_00240_),
    .B1(net289));
 sg13g2_a21o_1 _09184_ (.A2(_03699_),
    .A1(_03568_),
    .B1(_03698_),
    .X(_03706_));
 sg13g2_a21oi_1 _09185_ (.A1(_03692_),
    .A2(_03693_),
    .Y(_03707_),
    .B1(_03695_));
 sg13g2_a21oi_1 _09186_ (.A1(_03690_),
    .A2(_03696_),
    .Y(_03708_),
    .B1(_03689_));
 sg13g2_o21ai_1 _09187_ (.B1(_03634_),
    .Y(_03709_),
    .A1(_03635_),
    .A2(_03687_));
 sg13g2_o21ai_1 _09188_ (.B1(_03596_),
    .Y(_03710_),
    .A1(_03597_),
    .A2(_03632_));
 sg13g2_a21oi_2 _09189_ (.B1(_03578_),
    .Y(_03711_),
    .A2(net1117),
    .A1(net1395));
 sg13g2_xnor2_1 _09190_ (.Y(_03712_),
    .A(_03336_),
    .B(_03473_));
 sg13g2_nand2b_2 _09191_ (.Y(_03713_),
    .B(_03712_),
    .A_N(_03711_));
 sg13g2_xnor2_1 _09192_ (.Y(_03714_),
    .A(_03711_),
    .B(_03712_));
 sg13g2_and2_1 _09193_ (.A(net1358),
    .B(net1322),
    .X(_03715_));
 sg13g2_nand2_1 _09194_ (.Y(_03716_),
    .A(net1358),
    .B(net1323));
 sg13g2_nand2_1 _09195_ (.Y(_03717_),
    .A(net1358),
    .B(_03582_));
 sg13g2_o21ai_1 _09196_ (.B1(_03717_),
    .Y(_03718_),
    .A1(_03582_),
    .A2(_03715_));
 sg13g2_nand2_1 _09197_ (.Y(_03719_),
    .A(net1352),
    .B(net1326));
 sg13g2_nor2_1 _09198_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sg13g2_xor2_1 _09199_ (.B(_03719_),
    .A(_03718_),
    .X(_03721_));
 sg13g2_nand2_1 _09200_ (.Y(_03722_),
    .A(_03714_),
    .B(_03721_));
 sg13g2_xnor2_1 _09201_ (.Y(_03723_),
    .A(_03714_),
    .B(_03721_));
 sg13g2_nand2_1 _09202_ (.Y(_03724_),
    .A(_03580_),
    .B(_03589_));
 sg13g2_nand2b_1 _09203_ (.Y(_03725_),
    .B(_03724_),
    .A_N(_03723_));
 sg13g2_xor2_1 _09204_ (.B(_03724_),
    .A(_03723_),
    .X(_03726_));
 sg13g2_xor2_1 _09205_ (.B(_03574_),
    .A(_02953_),
    .X(_03727_));
 sg13g2_inv_1 _09206_ (.Y(_03728_),
    .A(_03727_));
 sg13g2_nor2_1 _09207_ (.A(_03726_),
    .B(_03727_),
    .Y(_03729_));
 sg13g2_xnor2_1 _09208_ (.Y(_03730_),
    .A(_03726_),
    .B(_03728_));
 sg13g2_nand2_1 _09209_ (.Y(_03731_),
    .A(_03594_),
    .B(_03730_));
 sg13g2_xnor2_1 _09210_ (.Y(_03732_),
    .A(_03594_),
    .B(_03730_));
 sg13g2_o21ai_1 _09211_ (.B1(_03611_),
    .Y(_03733_),
    .A1(_03612_),
    .A2(_03628_));
 sg13g2_a21o_1 _09212_ (.A2(_03609_),
    .A1(_03600_),
    .B1(_03608_),
    .X(_03734_));
 sg13g2_o21ai_1 _09213_ (.B1(_03605_),
    .Y(_03735_),
    .A1(_03602_),
    .A2(_03606_));
 sg13g2_a21oi_1 _09214_ (.A1(net1372),
    .A2(_03582_),
    .Y(_03736_),
    .B1(_03587_));
 sg13g2_nand2_1 _09215_ (.Y(_03737_),
    .A(net1460),
    .B(net1335));
 sg13g2_nand2_1 _09216_ (.Y(_03738_),
    .A(net1465),
    .B(net1329));
 sg13g2_nand2_1 _09217_ (.Y(_03739_),
    .A(net1465),
    .B(net1331));
 sg13g2_or2_1 _09218_ (.X(_03740_),
    .B(_03738_),
    .A(_03604_));
 sg13g2_xnor2_1 _09219_ (.Y(_03741_),
    .A(_03603_),
    .B(_03739_));
 sg13g2_xor2_1 _09220_ (.B(_03741_),
    .A(_03737_),
    .X(_03742_));
 sg13g2_nor2b_1 _09221_ (.A(_03736_),
    .B_N(_03742_),
    .Y(_03743_));
 sg13g2_xnor2_1 _09222_ (.Y(_03744_),
    .A(_03736_),
    .B(_03742_));
 sg13g2_xnor2_1 _09223_ (.Y(_03745_),
    .A(_03735_),
    .B(_03744_));
 sg13g2_nand2b_1 _09224_ (.Y(_03746_),
    .B(_03734_),
    .A_N(_03745_));
 sg13g2_xor2_1 _09225_ (.B(_03745_),
    .A(_03734_),
    .X(_03747_));
 sg13g2_nand2_1 _09226_ (.Y(_03748_),
    .A(net1432),
    .B(net1157));
 sg13g2_nand2_1 _09227_ (.Y(_03749_),
    .A(net1436),
    .B(net1145));
 sg13g2_nand2_1 _09228_ (.Y(_03750_),
    .A(net1436),
    .B(net1151));
 sg13g2_xor2_1 _09229_ (.B(_03750_),
    .A(_03614_),
    .X(_03751_));
 sg13g2_nand2b_1 _09230_ (.Y(_03752_),
    .B(_03751_),
    .A_N(_03748_));
 sg13g2_xnor2_1 _09231_ (.Y(_03753_),
    .A(_03748_),
    .B(_03751_));
 sg13g2_inv_1 _09232_ (.Y(_03754_),
    .A(_03753_));
 sg13g2_o21ai_1 _09233_ (.B1(_03624_),
    .Y(_03755_),
    .A1(_03456_),
    .A2(_03622_));
 sg13g2_nand2_1 _09234_ (.Y(_03756_),
    .A(net1446),
    .B(net1348));
 sg13g2_nand2_1 _09235_ (.Y(_03757_),
    .A(net1451),
    .B(net1337));
 sg13g2_nand2_1 _09236_ (.Y(_03758_),
    .A(net1451),
    .B(net1342));
 sg13g2_xor2_1 _09237_ (.B(_03758_),
    .A(_03621_),
    .X(_03759_));
 sg13g2_nand2b_1 _09238_ (.Y(_03760_),
    .B(_03759_),
    .A_N(_03756_));
 sg13g2_xnor2_1 _09239_ (.Y(_03761_),
    .A(_03756_),
    .B(_03759_));
 sg13g2_nand2_1 _09240_ (.Y(_03762_),
    .A(_03755_),
    .B(_03761_));
 sg13g2_xnor2_1 _09241_ (.Y(_03763_),
    .A(_03755_),
    .B(_03761_));
 sg13g2_xnor2_1 _09242_ (.Y(_03764_),
    .A(_03754_),
    .B(_03763_));
 sg13g2_xor2_1 _09243_ (.B(_03764_),
    .A(_03747_),
    .X(_03765_));
 sg13g2_nor2b_1 _09244_ (.A(_03592_),
    .B_N(_03765_),
    .Y(_03766_));
 sg13g2_xnor2_1 _09245_ (.Y(_03767_),
    .A(_03592_),
    .B(_03765_));
 sg13g2_xnor2_1 _09246_ (.Y(_03768_),
    .A(_03733_),
    .B(_03767_));
 sg13g2_xor2_1 _09247_ (.B(_03768_),
    .A(_03732_),
    .X(_03769_));
 sg13g2_nand2_1 _09248_ (.Y(_03770_),
    .A(_03710_),
    .B(_03769_));
 sg13g2_xnor2_1 _09249_ (.Y(_03771_),
    .A(_03710_),
    .B(_03769_));
 sg13g2_o21ai_1 _09250_ (.B1(_03682_),
    .Y(_03772_),
    .A1(_03663_),
    .A2(_03683_));
 sg13g2_a21oi_1 _09251_ (.A1(_03598_),
    .A2(_03631_),
    .Y(_03773_),
    .B1(_03630_));
 sg13g2_or2_1 _09252_ (.X(_03774_),
    .B(_03646_),
    .A(_03644_));
 sg13g2_and2_1 _09253_ (.A(net1066),
    .B(_03774_),
    .X(_03775_));
 sg13g2_xor2_1 _09254_ (.B(_03774_),
    .A(net1066),
    .X(_03776_));
 sg13g2_xnor2_1 _09255_ (.Y(_03777_),
    .A(_03489_),
    .B(_03776_));
 sg13g2_o21ai_1 _09256_ (.B1(_03657_),
    .Y(_03778_),
    .A1(_03649_),
    .A2(_03658_));
 sg13g2_o21ai_1 _09257_ (.B1(net1411),
    .Y(_03779_),
    .A1(net1200),
    .A2(net1195));
 sg13g2_nand2b_2 _09258_ (.Y(_03780_),
    .B(_03643_),
    .A_N(_03779_));
 sg13g2_xor2_1 _09259_ (.B(_03780_),
    .A(_03495_),
    .X(_03781_));
 sg13g2_xnor2_1 _09260_ (.Y(_03782_),
    .A(_03495_),
    .B(_03780_));
 sg13g2_o21ai_1 _09261_ (.B1(_03655_),
    .Y(_03783_),
    .A1(_03504_),
    .A2(_03653_));
 sg13g2_nand2_1 _09262_ (.Y(_03784_),
    .A(net1413),
    .B(net1193));
 sg13g2_nand2_1 _09263_ (.Y(_03785_),
    .A(net1417),
    .B(net1177));
 sg13g2_nand2_1 _09264_ (.Y(_03786_),
    .A(net1417),
    .B(net1184));
 sg13g2_xor2_1 _09265_ (.B(_03786_),
    .A(_03652_),
    .X(_03787_));
 sg13g2_nand2b_1 _09266_ (.Y(_03788_),
    .B(_03787_),
    .A_N(_03784_));
 sg13g2_xnor2_1 _09267_ (.Y(_03789_),
    .A(_03784_),
    .B(_03787_));
 sg13g2_nand2_1 _09268_ (.Y(_03790_),
    .A(_03783_),
    .B(_03789_));
 sg13g2_xnor2_1 _09269_ (.Y(_03791_),
    .A(_03783_),
    .B(_03789_));
 sg13g2_xnor2_1 _09270_ (.Y(_03792_),
    .A(_03781_),
    .B(_03791_));
 sg13g2_nand2_1 _09271_ (.Y(_03793_),
    .A(_03778_),
    .B(_03792_));
 sg13g2_xnor2_1 _09272_ (.Y(_03794_),
    .A(_03778_),
    .B(_03792_));
 sg13g2_xor2_1 _09273_ (.B(_03794_),
    .A(_03777_),
    .X(_03795_));
 sg13g2_inv_1 _09274_ (.Y(_03796_),
    .A(_03795_));
 sg13g2_nand2_1 _09275_ (.Y(_03797_),
    .A(_03678_),
    .B(_03680_));
 sg13g2_a21o_1 _09276_ (.A2(_03674_),
    .A1(_03668_),
    .B1(_03676_),
    .X(_03798_));
 sg13g2_o21ai_1 _09277_ (.B1(_03626_),
    .Y(_03799_),
    .A1(_03618_),
    .A2(_03627_));
 sg13g2_inv_1 _09278_ (.Y(_03800_),
    .A(_03799_));
 sg13g2_o21ai_1 _09279_ (.B1(_03673_),
    .Y(_03801_),
    .A1(_03523_),
    .A2(_03671_));
 sg13g2_o21ai_1 _09280_ (.B1(_03617_),
    .Y(_03802_),
    .A1(_03448_),
    .A2(_03615_));
 sg13g2_nand2_1 _09281_ (.Y(_03803_),
    .A(net1423),
    .B(net1173));
 sg13g2_nand2_1 _09282_ (.Y(_03804_),
    .A(net1424),
    .B(net1161));
 sg13g2_nand2_1 _09283_ (.Y(_03805_),
    .A(net1425),
    .B(net1168));
 sg13g2_xor2_1 _09284_ (.B(_03805_),
    .A(_03670_),
    .X(_03806_));
 sg13g2_nand2b_1 _09285_ (.Y(_03807_),
    .B(_03806_),
    .A_N(_03803_));
 sg13g2_xnor2_1 _09286_ (.Y(_03808_),
    .A(_03803_),
    .B(_03806_));
 sg13g2_xnor2_1 _09287_ (.Y(_03809_),
    .A(_03802_),
    .B(_03808_));
 sg13g2_nor2b_1 _09288_ (.A(_03809_),
    .B_N(_03801_),
    .Y(_03810_));
 sg13g2_xor2_1 _09289_ (.B(_03809_),
    .A(_03801_),
    .X(_03811_));
 sg13g2_xor2_1 _09290_ (.B(_03811_),
    .A(_03799_),
    .X(_03812_));
 sg13g2_nand2b_1 _09291_ (.Y(_03813_),
    .B(_03798_),
    .A_N(_03812_));
 sg13g2_xor2_1 _09292_ (.B(_03812_),
    .A(_03798_),
    .X(_03814_));
 sg13g2_nand2b_1 _09293_ (.Y(_03815_),
    .B(_03797_),
    .A_N(_03814_));
 sg13g2_xor2_1 _09294_ (.B(_03814_),
    .A(_03797_),
    .X(_03816_));
 sg13g2_xnor2_1 _09295_ (.Y(_03817_),
    .A(_03796_),
    .B(_03816_));
 sg13g2_nor2_1 _09296_ (.A(_03773_),
    .B(_03817_),
    .Y(_03818_));
 sg13g2_xor2_1 _09297_ (.B(_03817_),
    .A(_03773_),
    .X(_03819_));
 sg13g2_xnor2_1 _09298_ (.Y(_03820_),
    .A(_03772_),
    .B(_03819_));
 sg13g2_xor2_1 _09299_ (.B(_03820_),
    .A(_03771_),
    .X(_03821_));
 sg13g2_and2_1 _09300_ (.A(_03709_),
    .B(_03821_),
    .X(_03822_));
 sg13g2_or2_1 _09301_ (.X(_03823_),
    .B(_03821_),
    .A(_03709_));
 sg13g2_xnor2_1 _09302_ (.Y(_03824_),
    .A(_03709_),
    .B(_03821_));
 sg13g2_a21o_1 _09303_ (.A2(_03640_),
    .A1(_03489_),
    .B1(_03639_),
    .X(_03825_));
 sg13g2_o21ai_1 _09304_ (.B1(_03685_),
    .Y(_03826_),
    .A1(_03636_),
    .A2(_03686_));
 sg13g2_o21ai_1 _09305_ (.B1(_03660_),
    .Y(_03827_),
    .A1(_03641_),
    .A2(_03661_));
 sg13g2_and2_1 _09306_ (.A(_03826_),
    .B(_03827_),
    .X(_03828_));
 sg13g2_xor2_1 _09307_ (.B(_03827_),
    .A(_03826_),
    .X(_03829_));
 sg13g2_xor2_1 _09308_ (.B(_03829_),
    .A(_03825_),
    .X(_03830_));
 sg13g2_xnor2_1 _09309_ (.Y(_03831_),
    .A(_03824_),
    .B(_03830_));
 sg13g2_nand2b_1 _09310_ (.Y(_03832_),
    .B(_03831_),
    .A_N(_03708_));
 sg13g2_xnor2_1 _09311_ (.Y(_03833_),
    .A(_03708_),
    .B(_03831_));
 sg13g2_nand2b_1 _09312_ (.Y(_03834_),
    .B(_03833_),
    .A_N(_03707_));
 sg13g2_xnor2_1 _09313_ (.Y(_03835_),
    .A(_03707_),
    .B(_03833_));
 sg13g2_and2_1 _09314_ (.A(_03706_),
    .B(_03835_),
    .X(_03836_));
 sg13g2_xor2_1 _09315_ (.B(_03835_),
    .A(_03706_),
    .X(_03837_));
 sg13g2_a21oi_1 _09316_ (.A1(_03567_),
    .A2(_03703_),
    .Y(_03838_),
    .B1(_03702_));
 sg13g2_xnor2_1 _09317_ (.Y(_03839_),
    .A(_03837_),
    .B(_03838_));
 sg13g2_o21ai_1 _09318_ (.B1(net1507),
    .Y(_03840_),
    .A1(net1141),
    .A2(_03839_));
 sg13g2_a21oi_1 _09319_ (.A1(net1141),
    .A2(_04772_),
    .Y(_00241_),
    .B1(_03840_));
 sg13g2_nand2_1 _09320_ (.Y(_03841_),
    .A(_03703_),
    .B(_03837_));
 sg13g2_a21o_1 _09321_ (.A2(_03566_),
    .A1(_03564_),
    .B1(_03841_),
    .X(_03842_));
 sg13g2_a21oi_1 _09322_ (.A1(_03702_),
    .A2(_03837_),
    .Y(_03843_),
    .B1(_03836_));
 sg13g2_nand2_1 _09323_ (.Y(_03844_),
    .A(_03832_),
    .B(_03834_));
 sg13g2_a21oi_1 _09324_ (.A1(_03825_),
    .A2(_03829_),
    .Y(_03845_),
    .B1(_03828_));
 sg13g2_a21oi_1 _09325_ (.A1(_03823_),
    .A2(_03830_),
    .Y(_03846_),
    .B1(_03822_));
 sg13g2_o21ai_1 _09326_ (.B1(_03770_),
    .Y(_03847_),
    .A1(_03771_),
    .A2(_03820_));
 sg13g2_o21ai_1 _09327_ (.B1(_03731_),
    .Y(_03848_),
    .A1(_03732_),
    .A2(_03768_));
 sg13g2_a21oi_1 _09328_ (.A1(_03080_),
    .A2(net1103),
    .Y(_03849_),
    .B1(_03729_));
 sg13g2_o21ai_1 _09329_ (.B1(_03335_),
    .Y(_03850_),
    .A1(_03336_),
    .A2(_03474_));
 sg13g2_xnor2_1 _09330_ (.Y(_03851_),
    .A(_03476_),
    .B(_03582_));
 sg13g2_nand2_1 _09331_ (.Y(_03852_),
    .A(_03850_),
    .B(_03851_));
 sg13g2_xnor2_1 _09332_ (.Y(_03853_),
    .A(_03850_),
    .B(_03851_));
 sg13g2_and2_1 _09333_ (.A(net1352),
    .B(net1322),
    .X(_03854_));
 sg13g2_nand2_1 _09334_ (.Y(_03855_),
    .A(net1352),
    .B(net1323));
 sg13g2_nand2_1 _09335_ (.Y(_03856_),
    .A(net1352),
    .B(_03715_));
 sg13g2_o21ai_1 _09336_ (.B1(_03856_),
    .Y(_03857_),
    .A1(_03715_),
    .A2(_03854_));
 sg13g2_nand2_1 _09337_ (.Y(_03858_),
    .A(net1470),
    .B(net1326));
 sg13g2_nor2_1 _09338_ (.A(_03857_),
    .B(_03858_),
    .Y(_03859_));
 sg13g2_xor2_1 _09339_ (.B(_03858_),
    .A(_03857_),
    .X(_03860_));
 sg13g2_inv_1 _09340_ (.Y(_03861_),
    .A(_03860_));
 sg13g2_xnor2_1 _09341_ (.Y(_03862_),
    .A(_03853_),
    .B(_03860_));
 sg13g2_nand2_1 _09342_ (.Y(_03863_),
    .A(_03713_),
    .B(_03722_));
 sg13g2_nand2_1 _09343_ (.Y(_03864_),
    .A(_03862_),
    .B(_03863_));
 sg13g2_xor2_1 _09344_ (.B(_03863_),
    .A(_03862_),
    .X(_03865_));
 sg13g2_nand2_1 _09345_ (.Y(_03866_),
    .A(_03080_),
    .B(_03085_));
 sg13g2_xor2_1 _09346_ (.B(_03866_),
    .A(_03472_),
    .X(_03867_));
 sg13g2_inv_1 _09347_ (.Y(_03868_),
    .A(_03867_));
 sg13g2_xnor2_1 _09348_ (.Y(_03869_),
    .A(_03865_),
    .B(_03868_));
 sg13g2_xor2_1 _09349_ (.B(_03869_),
    .A(_03849_),
    .X(_03870_));
 sg13g2_o21ai_1 _09350_ (.B1(_03746_),
    .Y(_03871_),
    .A1(_03747_),
    .A2(_03764_));
 sg13g2_a21o_1 _09351_ (.A2(_03744_),
    .A1(_03735_),
    .B1(_03743_),
    .X(_03872_));
 sg13g2_o21ai_1 _09352_ (.B1(_03740_),
    .Y(_03873_),
    .A1(_03737_),
    .A2(_03741_));
 sg13g2_a21oi_1 _09353_ (.A1(net1365),
    .A2(_03715_),
    .Y(_03874_),
    .B1(_03720_));
 sg13g2_nand2_1 _09354_ (.Y(_03875_),
    .A(net1455),
    .B(net1334));
 sg13g2_nand2_1 _09355_ (.Y(_03876_),
    .A(net1460),
    .B(net1329));
 sg13g2_nand2_1 _09356_ (.Y(_03877_),
    .A(net1460),
    .B(net1331));
 sg13g2_or2_1 _09357_ (.X(_03878_),
    .B(_03876_),
    .A(_03739_));
 sg13g2_xnor2_1 _09358_ (.Y(_03879_),
    .A(_03738_),
    .B(_03877_));
 sg13g2_xor2_1 _09359_ (.B(_03879_),
    .A(_03875_),
    .X(_03880_));
 sg13g2_nor2b_1 _09360_ (.A(_03874_),
    .B_N(_03880_),
    .Y(_03881_));
 sg13g2_xnor2_1 _09361_ (.Y(_03882_),
    .A(_03874_),
    .B(_03880_));
 sg13g2_xor2_1 _09362_ (.B(_03882_),
    .A(_03873_),
    .X(_03883_));
 sg13g2_nand2_1 _09363_ (.Y(_03884_),
    .A(_03872_),
    .B(_03883_));
 sg13g2_xnor2_1 _09364_ (.Y(_03885_),
    .A(_03872_),
    .B(_03883_));
 sg13g2_nand2_1 _09365_ (.Y(_03886_),
    .A(net1428),
    .B(net1157));
 sg13g2_nand2_1 _09366_ (.Y(_03887_),
    .A(net1432),
    .B(net1145));
 sg13g2_nand2_1 _09367_ (.Y(_03888_),
    .A(net1432),
    .B(net1151));
 sg13g2_or2_1 _09368_ (.X(_03889_),
    .B(_03887_),
    .A(_03750_));
 sg13g2_xnor2_1 _09369_ (.Y(_03890_),
    .A(_03749_),
    .B(_03888_));
 sg13g2_xnor2_1 _09370_ (.Y(_03891_),
    .A(_03886_),
    .B(_03890_));
 sg13g2_o21ai_1 _09371_ (.B1(_03760_),
    .Y(_03892_),
    .A1(_03621_),
    .A2(_03758_));
 sg13g2_nand2_1 _09372_ (.Y(_03893_),
    .A(net1441),
    .B(net1348));
 sg13g2_nand2_1 _09373_ (.Y(_03894_),
    .A(net1446),
    .B(net1337));
 sg13g2_nand2_1 _09374_ (.Y(_03895_),
    .A(net1446),
    .B(net1342));
 sg13g2_xor2_1 _09375_ (.B(_03895_),
    .A(_03757_),
    .X(_03896_));
 sg13g2_nand2b_1 _09376_ (.Y(_03897_),
    .B(_03896_),
    .A_N(_03893_));
 sg13g2_xnor2_1 _09377_ (.Y(_03898_),
    .A(_03893_),
    .B(_03896_));
 sg13g2_nand2_1 _09378_ (.Y(_03899_),
    .A(_03892_),
    .B(_03898_));
 sg13g2_xnor2_1 _09379_ (.Y(_03900_),
    .A(_03892_),
    .B(_03898_));
 sg13g2_xnor2_1 _09380_ (.Y(_03901_),
    .A(_03891_),
    .B(_03900_));
 sg13g2_xor2_1 _09381_ (.B(_03901_),
    .A(_03885_),
    .X(_03902_));
 sg13g2_nor2b_1 _09382_ (.A(_03725_),
    .B_N(_03902_),
    .Y(_03903_));
 sg13g2_xnor2_1 _09383_ (.Y(_03904_),
    .A(_03725_),
    .B(_03902_));
 sg13g2_xnor2_1 _09384_ (.Y(_03905_),
    .A(_03871_),
    .B(_03904_));
 sg13g2_inv_1 _09385_ (.Y(_03906_),
    .A(_03905_));
 sg13g2_nand2_1 _09386_ (.Y(_03907_),
    .A(_03870_),
    .B(_03906_));
 sg13g2_xnor2_1 _09387_ (.Y(_03908_),
    .A(_03870_),
    .B(_03905_));
 sg13g2_nand2_1 _09388_ (.Y(_03909_),
    .A(_03848_),
    .B(_03908_));
 sg13g2_xnor2_1 _09389_ (.Y(_03910_),
    .A(_03848_),
    .B(_03908_));
 sg13g2_o21ai_1 _09390_ (.B1(_03815_),
    .Y(_03911_),
    .A1(_03796_),
    .A2(_03816_));
 sg13g2_a21oi_1 _09391_ (.A1(_03733_),
    .A2(_03767_),
    .Y(_03912_),
    .B1(_03766_));
 sg13g2_o21ai_1 _09392_ (.B1(_03813_),
    .Y(_03913_),
    .A1(_03800_),
    .A2(_03811_));
 sg13g2_a21o_2 _09393_ (.A2(_03808_),
    .A1(_03802_),
    .B1(_03810_),
    .X(_03914_));
 sg13g2_o21ai_1 _09394_ (.B1(_03762_),
    .Y(_03915_),
    .A1(_03754_),
    .A2(_03763_));
 sg13g2_inv_1 _09395_ (.Y(_03916_),
    .A(_03915_));
 sg13g2_o21ai_1 _09396_ (.B1(_03807_),
    .Y(_03917_),
    .A1(_03670_),
    .A2(_03805_));
 sg13g2_o21ai_1 _09397_ (.B1(_03752_),
    .Y(_03918_),
    .A1(_03614_),
    .A2(_03750_));
 sg13g2_nand2_1 _09398_ (.Y(_03919_),
    .A(net1418),
    .B(net1173));
 sg13g2_nand2_1 _09399_ (.Y(_03920_),
    .A(net1421),
    .B(net1161));
 sg13g2_nand2_1 _09400_ (.Y(_03921_),
    .A(net1421),
    .B(net1167));
 sg13g2_xor2_1 _09401_ (.B(_03921_),
    .A(_03804_),
    .X(_03922_));
 sg13g2_nand2b_1 _09402_ (.Y(_03923_),
    .B(_03922_),
    .A_N(_03919_));
 sg13g2_xnor2_1 _09403_ (.Y(_03924_),
    .A(_03919_),
    .B(_03922_));
 sg13g2_xnor2_1 _09404_ (.Y(_03925_),
    .A(_03918_),
    .B(_03924_));
 sg13g2_nor2b_1 _09405_ (.A(_03925_),
    .B_N(_03917_),
    .Y(_03926_));
 sg13g2_xor2_1 _09406_ (.B(_03925_),
    .A(_03917_),
    .X(_03927_));
 sg13g2_xor2_1 _09407_ (.B(_03927_),
    .A(_03915_),
    .X(_03928_));
 sg13g2_nand2b_1 _09408_ (.Y(_03929_),
    .B(_03914_),
    .A_N(_03928_));
 sg13g2_xor2_1 _09409_ (.B(_03928_),
    .A(_03914_),
    .X(_03930_));
 sg13g2_nand2b_1 _09410_ (.Y(_03931_),
    .B(_03913_),
    .A_N(_03930_));
 sg13g2_xor2_1 _09411_ (.B(_03930_),
    .A(_03913_),
    .X(_03932_));
 sg13g2_o21ai_1 _09412_ (.B1(_03643_),
    .Y(_03933_),
    .A1(_03495_),
    .A2(_03779_));
 sg13g2_and2_1 _09413_ (.A(net1066),
    .B(_03933_),
    .X(_03934_));
 sg13g2_xor2_1 _09414_ (.B(_03933_),
    .A(net1066),
    .X(_03935_));
 sg13g2_xnor2_1 _09415_ (.Y(_03936_),
    .A(_03489_),
    .B(_03935_));
 sg13g2_o21ai_1 _09416_ (.B1(_03790_),
    .Y(_03937_),
    .A1(_03782_),
    .A2(_03791_));
 sg13g2_o21ai_1 _09417_ (.B1(_03788_),
    .Y(_03938_),
    .A1(_03652_),
    .A2(_03786_));
 sg13g2_nand2_2 _09418_ (.Y(_03939_),
    .A(net1410),
    .B(net1193));
 sg13g2_nand2_1 _09419_ (.Y(_03940_),
    .A(net1414),
    .B(net1184));
 sg13g2_xor2_1 _09420_ (.B(_03940_),
    .A(_03785_),
    .X(_03941_));
 sg13g2_nand2b_1 _09421_ (.Y(_03942_),
    .B(_03941_),
    .A_N(_03939_));
 sg13g2_xnor2_1 _09422_ (.Y(_03943_),
    .A(_03939_),
    .B(_03941_));
 sg13g2_nand2_1 _09423_ (.Y(_03944_),
    .A(_03938_),
    .B(_03943_));
 sg13g2_xnor2_1 _09424_ (.Y(_03945_),
    .A(_03938_),
    .B(_03943_));
 sg13g2_xnor2_1 _09425_ (.Y(_03946_),
    .A(_03782_),
    .B(_03945_));
 sg13g2_nand2b_1 _09426_ (.Y(_03947_),
    .B(_03937_),
    .A_N(_03946_));
 sg13g2_xor2_1 _09427_ (.B(_03946_),
    .A(_03937_),
    .X(_03948_));
 sg13g2_xor2_1 _09428_ (.B(_03948_),
    .A(net1030),
    .X(_03949_));
 sg13g2_inv_1 _09429_ (.Y(_03950_),
    .A(_03949_));
 sg13g2_xnor2_1 _09430_ (.Y(_03951_),
    .A(_03932_),
    .B(_03949_));
 sg13g2_nor2b_1 _09431_ (.A(_03912_),
    .B_N(_03951_),
    .Y(_03952_));
 sg13g2_xnor2_1 _09432_ (.Y(_03953_),
    .A(_03912_),
    .B(_03951_));
 sg13g2_xnor2_1 _09433_ (.Y(_03954_),
    .A(_03911_),
    .B(_03953_));
 sg13g2_xor2_1 _09434_ (.B(_03954_),
    .A(_03910_),
    .X(_03955_));
 sg13g2_xnor2_1 _09435_ (.Y(_03956_),
    .A(_03847_),
    .B(_03955_));
 sg13g2_a21o_1 _09436_ (.A2(_03776_),
    .A1(_03489_),
    .B1(_03775_),
    .X(_03957_));
 sg13g2_a21oi_1 _09437_ (.A1(_03772_),
    .A2(_03819_),
    .Y(_03958_),
    .B1(_03818_));
 sg13g2_o21ai_1 _09438_ (.B1(_03793_),
    .Y(_03959_),
    .A1(_03777_),
    .A2(_03794_));
 sg13g2_nand2b_1 _09439_ (.Y(_03960_),
    .B(_03959_),
    .A_N(_03958_));
 sg13g2_xor2_1 _09440_ (.B(_03959_),
    .A(_03958_),
    .X(_03961_));
 sg13g2_nand2b_1 _09441_ (.Y(_03962_),
    .B(_03957_),
    .A_N(_03961_));
 sg13g2_xor2_1 _09442_ (.B(_03961_),
    .A(_03957_),
    .X(_03963_));
 sg13g2_nor2_1 _09443_ (.A(_03956_),
    .B(_03963_),
    .Y(_03964_));
 sg13g2_xor2_1 _09444_ (.B(_03963_),
    .A(_03956_),
    .X(_03965_));
 sg13g2_nand2b_1 _09445_ (.Y(_03966_),
    .B(_03965_),
    .A_N(_03846_));
 sg13g2_xnor2_1 _09446_ (.Y(_03967_),
    .A(_03846_),
    .B(_03965_));
 sg13g2_nand2b_1 _09447_ (.Y(_03968_),
    .B(_03967_),
    .A_N(_03845_));
 sg13g2_xnor2_1 _09448_ (.Y(_03969_),
    .A(_03845_),
    .B(_03967_));
 sg13g2_nand2_1 _09449_ (.Y(_03970_),
    .A(_03844_),
    .B(_03969_));
 sg13g2_inv_1 _09450_ (.Y(_03971_),
    .A(_03970_));
 sg13g2_xnor2_1 _09451_ (.Y(_03972_),
    .A(_03844_),
    .B(_03969_));
 sg13g2_a21oi_1 _09452_ (.A1(_03842_),
    .A2(_03843_),
    .Y(_03973_),
    .B1(_03972_));
 sg13g2_nand3_1 _09453_ (.B(_03843_),
    .C(_03972_),
    .A(_03842_),
    .Y(_03974_));
 sg13g2_nor2b_2 _09454_ (.A(_03973_),
    .B_N(_03974_),
    .Y(_03975_));
 sg13g2_o21ai_1 _09455_ (.B1(net1507),
    .Y(_03976_),
    .A1(net1141),
    .A2(_03975_));
 sg13g2_a21oi_1 _09456_ (.A1(net1141),
    .A2(_04771_),
    .Y(_00242_),
    .B1(_03976_));
 sg13g2_nand2_1 _09457_ (.Y(_03977_),
    .A(_03966_),
    .B(_03968_));
 sg13g2_nand2_1 _09458_ (.Y(_03978_),
    .A(_03960_),
    .B(_03962_));
 sg13g2_a21oi_1 _09459_ (.A1(_03847_),
    .A2(_03955_),
    .Y(_03979_),
    .B1(_03964_));
 sg13g2_o21ai_1 _09460_ (.B1(_03909_),
    .Y(_03980_),
    .A1(_03910_),
    .A2(_03954_));
 sg13g2_o21ai_1 _09461_ (.B1(_03907_),
    .Y(_03981_),
    .A1(_03849_),
    .A2(_03869_));
 sg13g2_a22oi_1 _09462_ (.Y(_03982_),
    .B1(_03865_),
    .B2(_03868_),
    .A2(_03470_),
    .A1(_03080_));
 sg13g2_nand2_1 _09463_ (.Y(_03983_),
    .A(_03080_),
    .B(_03472_));
 sg13g2_xnor2_1 _09464_ (.Y(_03984_),
    .A(_03575_),
    .B(_03581_));
 sg13g2_xnor2_1 _09465_ (.Y(_03985_),
    .A(_03983_),
    .B(_03984_));
 sg13g2_o21ai_1 _09466_ (.B1(_03852_),
    .Y(_03986_),
    .A1(_03853_),
    .A2(_03861_));
 sg13g2_o21ai_1 _09467_ (.B1(_03475_),
    .Y(_03987_),
    .A1(_03476_),
    .A2(_03583_));
 sg13g2_xnor2_1 _09468_ (.Y(_03988_),
    .A(_03585_),
    .B(_03715_));
 sg13g2_xnor2_1 _09469_ (.Y(_03989_),
    .A(_03987_),
    .B(_03988_));
 sg13g2_and2_1 _09470_ (.A(net1470),
    .B(net1322),
    .X(_03990_));
 sg13g2_nand2_1 _09471_ (.Y(_03991_),
    .A(net1470),
    .B(net1322));
 sg13g2_nand2_1 _09472_ (.Y(_03992_),
    .A(net1470),
    .B(_03854_));
 sg13g2_o21ai_1 _09473_ (.B1(_03992_),
    .Y(_03993_),
    .A1(_03854_),
    .A2(_03990_));
 sg13g2_nand2_1 _09474_ (.Y(_03994_),
    .A(net1465),
    .B(net1326));
 sg13g2_nor2_1 _09475_ (.A(_03993_),
    .B(_03994_),
    .Y(_03995_));
 sg13g2_xor2_1 _09476_ (.B(_03994_),
    .A(_03993_),
    .X(_03996_));
 sg13g2_nor2b_1 _09477_ (.A(_03989_),
    .B_N(_03996_),
    .Y(_03997_));
 sg13g2_xnor2_1 _09478_ (.Y(_03998_),
    .A(_03989_),
    .B(_03996_));
 sg13g2_xnor2_1 _09479_ (.Y(_03999_),
    .A(_03468_),
    .B(_03998_));
 sg13g2_and2_1 _09480_ (.A(_03986_),
    .B(_03999_),
    .X(_04000_));
 sg13g2_xnor2_1 _09481_ (.Y(_04001_),
    .A(_03986_),
    .B(_03999_));
 sg13g2_or2_1 _09482_ (.X(_04002_),
    .B(_04001_),
    .A(_03985_));
 sg13g2_xor2_1 _09483_ (.B(_04001_),
    .A(_03985_),
    .X(_04003_));
 sg13g2_nor2b_1 _09484_ (.A(_03982_),
    .B_N(_04003_),
    .Y(_04004_));
 sg13g2_xnor2_1 _09485_ (.Y(_04005_),
    .A(_03982_),
    .B(_04003_));
 sg13g2_o21ai_1 _09486_ (.B1(_03884_),
    .Y(_04006_),
    .A1(_03885_),
    .A2(_03901_));
 sg13g2_a21o_2 _09487_ (.A2(_03882_),
    .A1(_03873_),
    .B1(_03881_),
    .X(_04007_));
 sg13g2_o21ai_1 _09488_ (.B1(_03878_),
    .Y(_04008_),
    .A1(_03875_),
    .A2(_03879_));
 sg13g2_a21oi_1 _09489_ (.A1(net1358),
    .A2(_03854_),
    .Y(_04009_),
    .B1(_03859_));
 sg13g2_nand2_1 _09490_ (.Y(_04010_),
    .A(net1451),
    .B(net1334));
 sg13g2_nand2_1 _09491_ (.Y(_04011_),
    .A(net1455),
    .B(net1329));
 sg13g2_nand2_1 _09492_ (.Y(_04012_),
    .A(net1455),
    .B(net1331));
 sg13g2_or2_1 _09493_ (.X(_04013_),
    .B(_04011_),
    .A(_03877_));
 sg13g2_xnor2_1 _09494_ (.Y(_04014_),
    .A(_03876_),
    .B(_04012_));
 sg13g2_xor2_1 _09495_ (.B(_04014_),
    .A(_04010_),
    .X(_04015_));
 sg13g2_nor2b_1 _09496_ (.A(_04009_),
    .B_N(_04015_),
    .Y(_04016_));
 sg13g2_xnor2_1 _09497_ (.Y(_04017_),
    .A(_04009_),
    .B(_04015_));
 sg13g2_xor2_1 _09498_ (.B(_04017_),
    .A(_04008_),
    .X(_04018_));
 sg13g2_nand2_1 _09499_ (.Y(_04019_),
    .A(_04007_),
    .B(_04018_));
 sg13g2_xnor2_1 _09500_ (.Y(_04020_),
    .A(_04007_),
    .B(_04018_));
 sg13g2_nand2_1 _09501_ (.Y(_04021_),
    .A(net1424),
    .B(net1157));
 sg13g2_nand2_1 _09502_ (.Y(_04022_),
    .A(net1428),
    .B(net1145));
 sg13g2_nand2_1 _09503_ (.Y(_04023_),
    .A(net1428),
    .B(net1151));
 sg13g2_or2_1 _09504_ (.X(_04024_),
    .B(_04022_),
    .A(_03888_));
 sg13g2_xnor2_1 _09505_ (.Y(_04025_),
    .A(_03887_),
    .B(_04023_));
 sg13g2_xnor2_1 _09506_ (.Y(_04026_),
    .A(_04021_),
    .B(_04025_));
 sg13g2_o21ai_1 _09507_ (.B1(_03897_),
    .Y(_04027_),
    .A1(_03757_),
    .A2(_03895_));
 sg13g2_nand2_1 _09508_ (.Y(_04028_),
    .A(net1436),
    .B(net1348));
 sg13g2_nand2_1 _09509_ (.Y(_04029_),
    .A(net1441),
    .B(net1337));
 sg13g2_nand2_1 _09510_ (.Y(_04030_),
    .A(net1441),
    .B(net1342));
 sg13g2_xor2_1 _09511_ (.B(_04030_),
    .A(_03894_),
    .X(_04031_));
 sg13g2_nand2b_1 _09512_ (.Y(_04032_),
    .B(_04031_),
    .A_N(_04028_));
 sg13g2_xnor2_1 _09513_ (.Y(_04033_),
    .A(_04028_),
    .B(_04031_));
 sg13g2_nand2_1 _09514_ (.Y(_04034_),
    .A(_04027_),
    .B(_04033_));
 sg13g2_xnor2_1 _09515_ (.Y(_04035_),
    .A(_04027_),
    .B(_04033_));
 sg13g2_xnor2_1 _09516_ (.Y(_04036_),
    .A(_04026_),
    .B(_04035_));
 sg13g2_xnor2_1 _09517_ (.Y(_04037_),
    .A(_04020_),
    .B(_04036_));
 sg13g2_nor2_1 _09518_ (.A(_03864_),
    .B(_04037_),
    .Y(_04038_));
 sg13g2_xor2_1 _09519_ (.B(_04037_),
    .A(_03864_),
    .X(_04039_));
 sg13g2_xnor2_1 _09520_ (.Y(_04040_),
    .A(_04006_),
    .B(_04039_));
 sg13g2_inv_1 _09521_ (.Y(_04041_),
    .A(_04040_));
 sg13g2_xnor2_1 _09522_ (.Y(_04042_),
    .A(_04005_),
    .B(_04040_));
 sg13g2_nand2_1 _09523_ (.Y(_04043_),
    .A(_03981_),
    .B(_04042_));
 sg13g2_xnor2_1 _09524_ (.Y(_04044_),
    .A(_03981_),
    .B(_04042_));
 sg13g2_o21ai_1 _09525_ (.B1(_03931_),
    .Y(_04045_),
    .A1(_03932_),
    .A2(_03950_));
 sg13g2_a21oi_1 _09526_ (.A1(_03871_),
    .A2(_03904_),
    .Y(_04046_),
    .B1(_03903_));
 sg13g2_o21ai_1 _09527_ (.B1(_03929_),
    .Y(_04047_),
    .A1(_03916_),
    .A2(_03927_));
 sg13g2_a21o_1 _09528_ (.A2(_03924_),
    .A1(_03918_),
    .B1(_03926_),
    .X(_04048_));
 sg13g2_o21ai_1 _09529_ (.B1(_03899_),
    .Y(_04049_),
    .A1(_03891_),
    .A2(_03900_));
 sg13g2_o21ai_1 _09530_ (.B1(_03923_),
    .Y(_04050_),
    .A1(_03804_),
    .A2(_03921_));
 sg13g2_o21ai_1 _09531_ (.B1(_03889_),
    .Y(_04051_),
    .A1(_03886_),
    .A2(_03890_));
 sg13g2_nand2_1 _09532_ (.Y(_04052_),
    .A(net1415),
    .B(net1173));
 sg13g2_nand2_1 _09533_ (.Y(_04053_),
    .A(net1418),
    .B(net1161));
 sg13g2_nand2_1 _09534_ (.Y(_04054_),
    .A(net1418),
    .B(net1167));
 sg13g2_xor2_1 _09535_ (.B(_04054_),
    .A(_03920_),
    .X(_04055_));
 sg13g2_nand2b_1 _09536_ (.Y(_04056_),
    .B(_04055_),
    .A_N(_04052_));
 sg13g2_xnor2_1 _09537_ (.Y(_04057_),
    .A(_04052_),
    .B(_04055_));
 sg13g2_xnor2_1 _09538_ (.Y(_04058_),
    .A(_04051_),
    .B(_04057_));
 sg13g2_nor2b_1 _09539_ (.A(_04058_),
    .B_N(_04050_),
    .Y(_04059_));
 sg13g2_xnor2_1 _09540_ (.Y(_04060_),
    .A(_04050_),
    .B(_04058_));
 sg13g2_xnor2_1 _09541_ (.Y(_04061_),
    .A(_04049_),
    .B(_04060_));
 sg13g2_nor2b_1 _09542_ (.A(_04061_),
    .B_N(_04048_),
    .Y(_04062_));
 sg13g2_xor2_1 _09543_ (.B(_04061_),
    .A(_04048_),
    .X(_04063_));
 sg13g2_nand2b_1 _09544_ (.Y(_04064_),
    .B(_04047_),
    .A_N(_04063_));
 sg13g2_xor2_1 _09545_ (.B(_04063_),
    .A(_04047_),
    .X(_04065_));
 sg13g2_o21ai_1 _09546_ (.B1(_03944_),
    .Y(_04066_),
    .A1(_03782_),
    .A2(_03945_));
 sg13g2_o21ai_1 _09547_ (.B1(_03942_),
    .Y(_04067_),
    .A1(_03785_),
    .A2(_03940_));
 sg13g2_nor3_1 _09548_ (.A(_04822_),
    .B(_04831_),
    .C(_03940_),
    .Y(_04068_));
 sg13g2_a22oi_1 _09549_ (.Y(_04069_),
    .B1(net1177),
    .B2(net1414),
    .A2(net1184),
    .A1(net1410));
 sg13g2_nor3_1 _09550_ (.A(_03939_),
    .B(_04068_),
    .C(_04069_),
    .Y(_04070_));
 sg13g2_o21ai_1 _09551_ (.B1(_03939_),
    .Y(_04071_),
    .A1(_04068_),
    .A2(_04069_));
 sg13g2_nor2b_1 _09552_ (.A(_04070_),
    .B_N(_04071_),
    .Y(_04072_));
 sg13g2_nand2_1 _09553_ (.Y(_04073_),
    .A(_04067_),
    .B(_04072_));
 sg13g2_xnor2_1 _09554_ (.Y(_04074_),
    .A(_04067_),
    .B(_04072_));
 sg13g2_xnor2_1 _09555_ (.Y(_04075_),
    .A(_03782_),
    .B(_04074_));
 sg13g2_nand2b_1 _09556_ (.Y(_04076_),
    .B(_04066_),
    .A_N(_04075_));
 sg13g2_xor2_1 _09557_ (.B(_04075_),
    .A(_04066_),
    .X(_04077_));
 sg13g2_xor2_1 _09558_ (.B(_04077_),
    .A(_03936_),
    .X(_04078_));
 sg13g2_inv_1 _09559_ (.Y(_04079_),
    .A(_04078_));
 sg13g2_xnor2_1 _09560_ (.Y(_04080_),
    .A(_04065_),
    .B(_04078_));
 sg13g2_nor2b_1 _09561_ (.A(_04046_),
    .B_N(_04080_),
    .Y(_04081_));
 sg13g2_xnor2_1 _09562_ (.Y(_04082_),
    .A(_04046_),
    .B(_04080_));
 sg13g2_xnor2_1 _09563_ (.Y(_04083_),
    .A(_04045_),
    .B(_04082_));
 sg13g2_xor2_1 _09564_ (.B(_04083_),
    .A(_04044_),
    .X(_04084_));
 sg13g2_xnor2_1 _09565_ (.Y(_04085_),
    .A(_03980_),
    .B(_04084_));
 sg13g2_a21o_2 _09566_ (.A2(_03935_),
    .A1(_03489_),
    .B1(_03934_),
    .X(_04086_));
 sg13g2_inv_4 _09567_ (.A(_04086_),
    .Y(_04087_));
 sg13g2_a21oi_1 _09568_ (.A1(_03911_),
    .A2(_03953_),
    .Y(_04088_),
    .B1(_03952_));
 sg13g2_o21ai_1 _09569_ (.B1(_03947_),
    .Y(_04089_),
    .A1(net1030),
    .A2(_03948_));
 sg13g2_nand2b_1 _09570_ (.Y(_04090_),
    .B(_04089_),
    .A_N(_04088_));
 sg13g2_xor2_1 _09571_ (.B(_04089_),
    .A(_04088_),
    .X(_04091_));
 sg13g2_xnor2_1 _09572_ (.Y(_04092_),
    .A(_04087_),
    .B(_04091_));
 sg13g2_nor2_1 _09573_ (.A(_04085_),
    .B(_04092_),
    .Y(_04093_));
 sg13g2_xor2_1 _09574_ (.B(_04092_),
    .A(_04085_),
    .X(_04094_));
 sg13g2_nor2b_1 _09575_ (.A(_03979_),
    .B_N(_04094_),
    .Y(_04095_));
 sg13g2_xnor2_1 _09576_ (.Y(_04096_),
    .A(_03979_),
    .B(_04094_));
 sg13g2_xor2_1 _09577_ (.B(_04096_),
    .A(_03978_),
    .X(_04097_));
 sg13g2_nand2_1 _09578_ (.Y(_04098_),
    .A(_03977_),
    .B(_04097_));
 sg13g2_xnor2_1 _09579_ (.Y(_04099_),
    .A(_03977_),
    .B(_04097_));
 sg13g2_inv_1 _09580_ (.Y(_04100_),
    .A(_04099_));
 sg13g2_o21ai_1 _09581_ (.B1(_04100_),
    .Y(_04101_),
    .A1(_03971_),
    .A2(_03973_));
 sg13g2_or3_1 _09582_ (.A(_03971_),
    .B(_03973_),
    .C(_04100_),
    .X(_04102_));
 sg13g2_nand2_1 _09583_ (.Y(_04103_),
    .A(_04101_),
    .B(_04102_));
 sg13g2_o21ai_1 _09584_ (.B1(net1507),
    .Y(_04104_),
    .A1(net1300),
    .A2(net285));
 sg13g2_a21oi_1 _09585_ (.A1(net1300),
    .A2(_04103_),
    .Y(_00243_),
    .B1(net286));
 sg13g2_a21o_1 _09586_ (.A2(_04096_),
    .A1(_03978_),
    .B1(_04095_),
    .X(_04105_));
 sg13g2_o21ai_1 _09587_ (.B1(_04090_),
    .Y(_04106_),
    .A1(_04087_),
    .A2(_04091_));
 sg13g2_a21oi_1 _09588_ (.A1(_03980_),
    .A2(_04084_),
    .Y(_04107_),
    .B1(_04093_));
 sg13g2_o21ai_1 _09589_ (.B1(_04043_),
    .Y(_04108_),
    .A1(_04044_),
    .A2(_04083_));
 sg13g2_a21oi_1 _09590_ (.A1(_04005_),
    .A2(_04041_),
    .Y(_04109_),
    .B1(_04004_));
 sg13g2_o21ai_1 _09591_ (.B1(_04002_),
    .Y(_04110_),
    .A1(_03983_),
    .A2(_03984_));
 sg13g2_xnor2_1 _09592_ (.Y(_04111_),
    .A(_03714_),
    .B(_03727_));
 sg13g2_nand3_1 _09593_ (.B(_03581_),
    .C(_04111_),
    .A(_03575_),
    .Y(_04112_));
 sg13g2_a21o_1 _09594_ (.A2(_03581_),
    .A1(_03575_),
    .B1(_04111_),
    .X(_04113_));
 sg13g2_nand2_1 _09595_ (.Y(_04114_),
    .A(_04112_),
    .B(_04113_));
 sg13g2_a21o_1 _09596_ (.A2(_03988_),
    .A1(_03987_),
    .B1(_03997_),
    .X(_04115_));
 sg13g2_and2_1 _09597_ (.A(net1465),
    .B(net1322),
    .X(_04116_));
 sg13g2_nand2_1 _09598_ (.Y(_04117_),
    .A(net1465),
    .B(net1322));
 sg13g2_nand2_1 _09599_ (.Y(_04118_),
    .A(net1465),
    .B(_03990_));
 sg13g2_o21ai_1 _09600_ (.B1(_04118_),
    .Y(_04119_),
    .A1(_03990_),
    .A2(_04116_));
 sg13g2_nand2_1 _09601_ (.Y(_04120_),
    .A(net1460),
    .B(net1326));
 sg13g2_xnor2_1 _09602_ (.Y(_04121_),
    .A(_04119_),
    .B(_04120_));
 sg13g2_o21ai_1 _09603_ (.B1(_03584_),
    .Y(_04122_),
    .A1(_03585_),
    .A2(_03716_));
 sg13g2_xnor2_1 _09604_ (.Y(_04123_),
    .A(_03718_),
    .B(_03854_));
 sg13g2_nand2_1 _09605_ (.Y(_04124_),
    .A(_04122_),
    .B(_04123_));
 sg13g2_xnor2_1 _09606_ (.Y(_04125_),
    .A(_04122_),
    .B(_04123_));
 sg13g2_xnor2_1 _09607_ (.Y(_04126_),
    .A(_04121_),
    .B(_04125_));
 sg13g2_xor2_1 _09608_ (.B(_04126_),
    .A(_03580_),
    .X(_04127_));
 sg13g2_nand2_1 _09609_ (.Y(_04128_),
    .A(_04115_),
    .B(_04127_));
 sg13g2_xnor2_1 _09610_ (.Y(_04129_),
    .A(_04115_),
    .B(_04127_));
 sg13g2_xor2_1 _09611_ (.B(_04129_),
    .A(_04114_),
    .X(_04130_));
 sg13g2_nand2_1 _09612_ (.Y(_04131_),
    .A(_04110_),
    .B(_04130_));
 sg13g2_xnor2_1 _09613_ (.Y(_04132_),
    .A(_04110_),
    .B(_04130_));
 sg13g2_o21ai_1 _09614_ (.B1(_04019_),
    .Y(_04133_),
    .A1(_04020_),
    .A2(_04036_));
 sg13g2_a21o_2 _09615_ (.A2(_03998_),
    .A1(_03469_),
    .B1(_04000_),
    .X(_04134_));
 sg13g2_a21o_1 _09616_ (.A2(_04017_),
    .A1(_04008_),
    .B1(_04016_),
    .X(_04135_));
 sg13g2_o21ai_1 _09617_ (.B1(_04013_),
    .Y(_04136_),
    .A1(_04010_),
    .A2(_04014_));
 sg13g2_a21oi_1 _09618_ (.A1(net1352),
    .A2(_03990_),
    .Y(_04137_),
    .B1(_03995_));
 sg13g2_nand2_1 _09619_ (.Y(_04138_),
    .A(net1446),
    .B(net1334));
 sg13g2_nand2_1 _09620_ (.Y(_04139_),
    .A(net1451),
    .B(net1329));
 sg13g2_nand2_1 _09621_ (.Y(_04140_),
    .A(net1451),
    .B(net1331));
 sg13g2_or2_1 _09622_ (.X(_04141_),
    .B(_04139_),
    .A(_04012_));
 sg13g2_xnor2_1 _09623_ (.Y(_04142_),
    .A(_04011_),
    .B(_04140_));
 sg13g2_xor2_1 _09624_ (.B(_04142_),
    .A(_04138_),
    .X(_04143_));
 sg13g2_nor2b_1 _09625_ (.A(_04137_),
    .B_N(_04143_),
    .Y(_04144_));
 sg13g2_xnor2_1 _09626_ (.Y(_04145_),
    .A(_04137_),
    .B(_04143_));
 sg13g2_xor2_1 _09627_ (.B(_04145_),
    .A(_04136_),
    .X(_04146_));
 sg13g2_nand2_1 _09628_ (.Y(_04147_),
    .A(_04135_),
    .B(_04146_));
 sg13g2_xnor2_1 _09629_ (.Y(_04148_),
    .A(_04135_),
    .B(_04146_));
 sg13g2_nand2_1 _09630_ (.Y(_04149_),
    .A(net1421),
    .B(net1157));
 sg13g2_nand2_1 _09631_ (.Y(_04150_),
    .A(net1424),
    .B(net1145));
 sg13g2_nand2_1 _09632_ (.Y(_04151_),
    .A(net1424),
    .B(net1151));
 sg13g2_or2_1 _09633_ (.X(_04152_),
    .B(_04150_),
    .A(_04023_));
 sg13g2_xnor2_1 _09634_ (.Y(_04153_),
    .A(_04022_),
    .B(_04151_));
 sg13g2_xnor2_1 _09635_ (.Y(_04154_),
    .A(_04149_),
    .B(_04153_));
 sg13g2_o21ai_1 _09636_ (.B1(_04032_),
    .Y(_04155_),
    .A1(_03894_),
    .A2(_04030_));
 sg13g2_nand2_1 _09637_ (.Y(_04156_),
    .A(net1432),
    .B(net1348));
 sg13g2_nand2_1 _09638_ (.Y(_04157_),
    .A(net1436),
    .B(net1337));
 sg13g2_nand2_1 _09639_ (.Y(_04158_),
    .A(net1436),
    .B(net1342));
 sg13g2_xor2_1 _09640_ (.B(_04158_),
    .A(_04029_),
    .X(_04159_));
 sg13g2_nand2b_1 _09641_ (.Y(_04160_),
    .B(_04159_),
    .A_N(_04156_));
 sg13g2_xnor2_1 _09642_ (.Y(_04161_),
    .A(_04156_),
    .B(_04159_));
 sg13g2_nand2_1 _09643_ (.Y(_04162_),
    .A(_04155_),
    .B(_04161_));
 sg13g2_xnor2_1 _09644_ (.Y(_04163_),
    .A(_04155_),
    .B(_04161_));
 sg13g2_xnor2_1 _09645_ (.Y(_04164_),
    .A(_04154_),
    .B(_04163_));
 sg13g2_xor2_1 _09646_ (.B(_04164_),
    .A(_04148_),
    .X(_04165_));
 sg13g2_xor2_1 _09647_ (.B(_04165_),
    .A(_04134_),
    .X(_04166_));
 sg13g2_and2_1 _09648_ (.A(_04133_),
    .B(_04166_),
    .X(_04167_));
 sg13g2_xnor2_1 _09649_ (.Y(_04168_),
    .A(_04133_),
    .B(_04166_));
 sg13g2_xor2_1 _09650_ (.B(_04168_),
    .A(_04132_),
    .X(_04169_));
 sg13g2_nand2b_1 _09651_ (.Y(_04170_),
    .B(_04169_),
    .A_N(_04109_));
 sg13g2_xor2_1 _09652_ (.B(_04169_),
    .A(_04109_),
    .X(_04171_));
 sg13g2_o21ai_1 _09653_ (.B1(_04064_),
    .Y(_04172_),
    .A1(_04065_),
    .A2(_04079_));
 sg13g2_a21oi_1 _09654_ (.A1(_04006_),
    .A2(_04039_),
    .Y(_04173_),
    .B1(_04038_));
 sg13g2_a21o_1 _09655_ (.A2(_04060_),
    .A1(_04049_),
    .B1(_04062_),
    .X(_04174_));
 sg13g2_a21o_1 _09656_ (.A2(_04057_),
    .A1(_04051_),
    .B1(_04059_),
    .X(_04175_));
 sg13g2_o21ai_1 _09657_ (.B1(_04034_),
    .Y(_04176_),
    .A1(_04026_),
    .A2(_04035_));
 sg13g2_o21ai_1 _09658_ (.B1(_04056_),
    .Y(_04177_),
    .A1(_03920_),
    .A2(_04054_));
 sg13g2_o21ai_1 _09659_ (.B1(_04024_),
    .Y(_04178_),
    .A1(_04021_),
    .A2(_04025_));
 sg13g2_nand2_1 _09660_ (.Y(_04179_),
    .A(net1413),
    .B(net1174));
 sg13g2_nand2_1 _09661_ (.Y(_04180_),
    .A(net1415),
    .B(net1167));
 sg13g2_xor2_1 _09662_ (.B(_04180_),
    .A(_04053_),
    .X(_04181_));
 sg13g2_nand2b_1 _09663_ (.Y(_04182_),
    .B(_04181_),
    .A_N(_04179_));
 sg13g2_xnor2_1 _09664_ (.Y(_04183_),
    .A(_04179_),
    .B(_04181_));
 sg13g2_xnor2_1 _09665_ (.Y(_04184_),
    .A(_04178_),
    .B(_04183_));
 sg13g2_nor2b_1 _09666_ (.A(_04184_),
    .B_N(_04177_),
    .Y(_04185_));
 sg13g2_xnor2_1 _09667_ (.Y(_04186_),
    .A(_04177_),
    .B(_04184_));
 sg13g2_xnor2_1 _09668_ (.Y(_04187_),
    .A(_04176_),
    .B(_04186_));
 sg13g2_nor2b_1 _09669_ (.A(_04187_),
    .B_N(_04175_),
    .Y(_04188_));
 sg13g2_xnor2_1 _09670_ (.Y(_04189_),
    .A(_04175_),
    .B(_04187_));
 sg13g2_nand2_1 _09671_ (.Y(_04190_),
    .A(_04174_),
    .B(_04189_));
 sg13g2_xnor2_1 _09672_ (.Y(_04191_),
    .A(_04174_),
    .B(_04189_));
 sg13g2_o21ai_1 _09673_ (.B1(_04073_),
    .Y(_04192_),
    .A1(_03782_),
    .A2(_04074_));
 sg13g2_inv_1 _09674_ (.Y(_04193_),
    .A(_04192_));
 sg13g2_or2_1 _09675_ (.X(_04194_),
    .B(_04070_),
    .A(_04068_));
 sg13g2_o21ai_1 _09676_ (.B1(net1411),
    .Y(_04195_),
    .A1(net1184),
    .A2(net1177));
 sg13g2_nand3_1 _09677_ (.B(net1184),
    .C(net1177),
    .A(net1411),
    .Y(_04196_));
 sg13g2_nand2b_1 _09678_ (.Y(_04197_),
    .B(_04196_),
    .A_N(_04195_));
 sg13g2_xnor2_1 _09679_ (.Y(_04198_),
    .A(_03939_),
    .B(_04197_));
 sg13g2_nand2b_1 _09680_ (.Y(_04199_),
    .B(_04194_),
    .A_N(_04198_));
 sg13g2_xnor2_1 _09681_ (.Y(_04200_),
    .A(_04194_),
    .B(_04198_));
 sg13g2_xnor2_1 _09682_ (.Y(_04201_),
    .A(_03781_),
    .B(_04200_));
 sg13g2_xnor2_1 _09683_ (.Y(_04202_),
    .A(_04192_),
    .B(_04201_));
 sg13g2_nand2b_1 _09684_ (.Y(_04203_),
    .B(_04202_),
    .A_N(net1030));
 sg13g2_xnor2_1 _09685_ (.Y(_04204_),
    .A(net1030),
    .B(_04202_));
 sg13g2_inv_1 _09686_ (.Y(_04205_),
    .A(_04204_));
 sg13g2_xnor2_1 _09687_ (.Y(_04206_),
    .A(_04191_),
    .B(_04204_));
 sg13g2_nor2b_1 _09688_ (.A(_04173_),
    .B_N(_04206_),
    .Y(_04207_));
 sg13g2_xnor2_1 _09689_ (.Y(_04208_),
    .A(_04173_),
    .B(_04206_));
 sg13g2_xnor2_1 _09690_ (.Y(_04209_),
    .A(_04172_),
    .B(_04208_));
 sg13g2_xnor2_1 _09691_ (.Y(_04210_),
    .A(_04171_),
    .B(_04209_));
 sg13g2_nor2b_1 _09692_ (.A(_04210_),
    .B_N(_04108_),
    .Y(_04211_));
 sg13g2_xor2_1 _09693_ (.B(_04210_),
    .A(_04108_),
    .X(_04212_));
 sg13g2_a21oi_1 _09694_ (.A1(_04045_),
    .A2(_04082_),
    .Y(_04213_),
    .B1(_04081_));
 sg13g2_o21ai_1 _09695_ (.B1(_04076_),
    .Y(_04214_),
    .A1(_03936_),
    .A2(_04077_));
 sg13g2_nand2b_1 _09696_ (.Y(_04215_),
    .B(_04214_),
    .A_N(_04213_));
 sg13g2_xor2_1 _09697_ (.B(_04214_),
    .A(_04213_),
    .X(_04216_));
 sg13g2_xnor2_1 _09698_ (.Y(_04217_),
    .A(_04087_),
    .B(_04216_));
 sg13g2_nor2_1 _09699_ (.A(_04212_),
    .B(_04217_),
    .Y(_04218_));
 sg13g2_xor2_1 _09700_ (.B(_04217_),
    .A(_04212_),
    .X(_04219_));
 sg13g2_nor2b_1 _09701_ (.A(_04107_),
    .B_N(_04219_),
    .Y(_04220_));
 sg13g2_xnor2_1 _09702_ (.Y(_04221_),
    .A(_04107_),
    .B(_04219_));
 sg13g2_xor2_1 _09703_ (.B(_04221_),
    .A(_04106_),
    .X(_04222_));
 sg13g2_and2_1 _09704_ (.A(_04105_),
    .B(_04222_),
    .X(_04223_));
 sg13g2_xnor2_1 _09705_ (.Y(_04224_),
    .A(_04105_),
    .B(_04222_));
 sg13g2_a21oi_1 _09706_ (.A1(_04098_),
    .A2(_04101_),
    .Y(_04225_),
    .B1(_04224_));
 sg13g2_nand3_1 _09707_ (.B(_04101_),
    .C(_04224_),
    .A(_04098_),
    .Y(_04226_));
 sg13g2_nand2b_2 _09708_ (.Y(_04227_),
    .B(_04226_),
    .A_N(_04225_));
 sg13g2_o21ai_1 _09709_ (.B1(net1499),
    .Y(_04228_),
    .A1(net1296),
    .A2(net271));
 sg13g2_a21oi_1 _09710_ (.A1(net1296),
    .A2(_04227_),
    .Y(_00244_),
    .B1(net272));
 sg13g2_a21o_1 _09711_ (.A2(_04221_),
    .A1(_04106_),
    .B1(_04220_),
    .X(_04229_));
 sg13g2_o21ai_1 _09712_ (.B1(_04215_),
    .Y(_04230_),
    .A1(_04087_),
    .A2(_04216_));
 sg13g2_nor2_1 _09713_ (.A(_04211_),
    .B(_04218_),
    .Y(_04231_));
 sg13g2_o21ai_1 _09714_ (.B1(_04170_),
    .Y(_04232_),
    .A1(_04171_),
    .A2(_04209_));
 sg13g2_o21ai_1 _09715_ (.B1(_04131_),
    .Y(_04233_),
    .A1(_04132_),
    .A2(_04168_));
 sg13g2_o21ai_1 _09716_ (.B1(_04112_),
    .Y(_04234_),
    .A1(_04114_),
    .A2(_04129_));
 sg13g2_a22oi_1 _09717_ (.Y(_04235_),
    .B1(_03714_),
    .B2(_03728_),
    .A2(net1103),
    .A1(_03080_));
 sg13g2_and2_1 _09718_ (.A(net1103),
    .B(_03851_),
    .X(_04236_));
 sg13g2_xnor2_1 _09719_ (.Y(_04237_),
    .A(_03083_),
    .B(_03851_));
 sg13g2_xnor2_1 _09720_ (.Y(_04238_),
    .A(_03850_),
    .B(_04237_));
 sg13g2_inv_1 _09721_ (.Y(_04239_),
    .A(_04238_));
 sg13g2_or2_1 _09722_ (.X(_04240_),
    .B(net1117),
    .A(net1118));
 sg13g2_o21ai_1 _09723_ (.B1(_04240_),
    .Y(_04241_),
    .A1(_03080_),
    .A2(_03471_));
 sg13g2_xnor2_1 _09724_ (.Y(_04242_),
    .A(_04239_),
    .B(_04241_));
 sg13g2_nor2_1 _09725_ (.A(_04235_),
    .B(_04242_),
    .Y(_04243_));
 sg13g2_xor2_1 _09726_ (.B(_04242_),
    .A(_04235_),
    .X(_04244_));
 sg13g2_o21ai_1 _09727_ (.B1(_04124_),
    .Y(_04245_),
    .A1(_04121_),
    .A2(_04125_));
 sg13g2_and2_1 _09728_ (.A(net1460),
    .B(net1322),
    .X(_04246_));
 sg13g2_nand2_1 _09729_ (.Y(_04247_),
    .A(net1460),
    .B(_04116_));
 sg13g2_o21ai_1 _09730_ (.B1(_04247_),
    .Y(_04248_),
    .A1(_04116_),
    .A2(_04246_));
 sg13g2_nand2_1 _09731_ (.Y(_04249_),
    .A(net1455),
    .B(net1326));
 sg13g2_xor2_1 _09732_ (.B(_04249_),
    .A(_04248_),
    .X(_04250_));
 sg13g2_inv_1 _09733_ (.Y(_04251_),
    .A(_04250_));
 sg13g2_o21ai_1 _09734_ (.B1(_03717_),
    .Y(_04252_),
    .A1(_03718_),
    .A2(_03855_));
 sg13g2_xnor2_1 _09735_ (.Y(_04253_),
    .A(_03857_),
    .B(_03990_));
 sg13g2_nand2_1 _09736_ (.Y(_04254_),
    .A(_04252_),
    .B(_04253_));
 sg13g2_xnor2_1 _09737_ (.Y(_04255_),
    .A(_04252_),
    .B(_04253_));
 sg13g2_xnor2_1 _09738_ (.Y(_04256_),
    .A(_04251_),
    .B(_04255_));
 sg13g2_nor2_1 _09739_ (.A(_03713_),
    .B(_04256_),
    .Y(_04257_));
 sg13g2_xor2_1 _09740_ (.B(_04256_),
    .A(_03713_),
    .X(_04258_));
 sg13g2_xnor2_1 _09741_ (.Y(_04259_),
    .A(_04245_),
    .B(_04258_));
 sg13g2_inv_1 _09742_ (.Y(_04260_),
    .A(_04259_));
 sg13g2_xnor2_1 _09743_ (.Y(_04261_),
    .A(_04244_),
    .B(_04259_));
 sg13g2_nand2_1 _09744_ (.Y(_04262_),
    .A(_04234_),
    .B(_04261_));
 sg13g2_xnor2_1 _09745_ (.Y(_04263_),
    .A(_04234_),
    .B(_04261_));
 sg13g2_o21ai_1 _09746_ (.B1(_04147_),
    .Y(_04264_),
    .A1(_04148_),
    .A2(_04164_));
 sg13g2_o21ai_1 _09747_ (.B1(_04128_),
    .Y(_04265_),
    .A1(_03580_),
    .A2(_04126_));
 sg13g2_a21o_1 _09748_ (.A2(_04145_),
    .A1(_04136_),
    .B1(_04144_),
    .X(_04266_));
 sg13g2_o21ai_1 _09749_ (.B1(_04141_),
    .Y(_04267_),
    .A1(_04138_),
    .A2(_04142_));
 sg13g2_o21ai_1 _09750_ (.B1(_04118_),
    .Y(_04268_),
    .A1(_04119_),
    .A2(_04120_));
 sg13g2_nand2_1 _09751_ (.Y(_04269_),
    .A(net1441),
    .B(net1334));
 sg13g2_nand2_2 _09752_ (.Y(_04270_),
    .A(net1446),
    .B(net1331));
 sg13g2_or2_1 _09753_ (.X(_04271_),
    .B(_04270_),
    .A(_04139_));
 sg13g2_xnor2_1 _09754_ (.Y(_04272_),
    .A(_04139_),
    .B(_04270_));
 sg13g2_xor2_1 _09755_ (.B(_04272_),
    .A(_04269_),
    .X(_04273_));
 sg13g2_xnor2_1 _09756_ (.Y(_04274_),
    .A(_04268_),
    .B(_04273_));
 sg13g2_nor2b_1 _09757_ (.A(_04274_),
    .B_N(_04267_),
    .Y(_04275_));
 sg13g2_xnor2_1 _09758_ (.Y(_04276_),
    .A(_04267_),
    .B(_04274_));
 sg13g2_nand2_1 _09759_ (.Y(_04277_),
    .A(_04266_),
    .B(_04276_));
 sg13g2_xnor2_1 _09760_ (.Y(_04278_),
    .A(_04266_),
    .B(_04276_));
 sg13g2_nand2_1 _09761_ (.Y(_04279_),
    .A(net1418),
    .B(net1157));
 sg13g2_nand2_1 _09762_ (.Y(_04280_),
    .A(net1421),
    .B(net1145));
 sg13g2_nand2_1 _09763_ (.Y(_04281_),
    .A(net1421),
    .B(net1151));
 sg13g2_xor2_1 _09764_ (.B(_04281_),
    .A(_04150_),
    .X(_04282_));
 sg13g2_nand2b_1 _09765_ (.Y(_04283_),
    .B(_04282_),
    .A_N(_04279_));
 sg13g2_xor2_1 _09766_ (.B(_04282_),
    .A(_04279_),
    .X(_04284_));
 sg13g2_o21ai_1 _09767_ (.B1(_04160_),
    .Y(_04285_),
    .A1(_04029_),
    .A2(_04158_));
 sg13g2_nand2_1 _09768_ (.Y(_04286_),
    .A(net1428),
    .B(net1348));
 sg13g2_nand2_2 _09769_ (.Y(_04287_),
    .A(net1432),
    .B(net1342));
 sg13g2_xor2_1 _09770_ (.B(_04287_),
    .A(_04157_),
    .X(_04288_));
 sg13g2_nand2b_1 _09771_ (.Y(_04289_),
    .B(_04288_),
    .A_N(_04286_));
 sg13g2_xnor2_1 _09772_ (.Y(_04290_),
    .A(_04286_),
    .B(_04288_));
 sg13g2_nand2_1 _09773_ (.Y(_04291_),
    .A(_04285_),
    .B(_04290_));
 sg13g2_xnor2_1 _09774_ (.Y(_04292_),
    .A(_04285_),
    .B(_04290_));
 sg13g2_xnor2_1 _09775_ (.Y(_04293_),
    .A(_04284_),
    .B(_04292_));
 sg13g2_xor2_1 _09776_ (.B(_04293_),
    .A(_04278_),
    .X(_04294_));
 sg13g2_xor2_1 _09777_ (.B(_04294_),
    .A(_04265_),
    .X(_04295_));
 sg13g2_and2_1 _09778_ (.A(_04264_),
    .B(_04295_),
    .X(_04296_));
 sg13g2_xnor2_1 _09779_ (.Y(_04297_),
    .A(_04264_),
    .B(_04295_));
 sg13g2_xor2_1 _09780_ (.B(_04297_),
    .A(_04263_),
    .X(_04298_));
 sg13g2_nand2_1 _09781_ (.Y(_04299_),
    .A(_04233_),
    .B(_04298_));
 sg13g2_xnor2_1 _09782_ (.Y(_04300_),
    .A(_04233_),
    .B(_04298_));
 sg13g2_o21ai_1 _09783_ (.B1(_04190_),
    .Y(_04301_),
    .A1(_04191_),
    .A2(_04205_));
 sg13g2_a21oi_1 _09784_ (.A1(_04134_),
    .A2(_04165_),
    .Y(_04302_),
    .B1(_04167_));
 sg13g2_nand2_1 _09785_ (.Y(_04303_),
    .A(_03939_),
    .B(_04195_));
 sg13g2_nand3b_1 _09786_ (.B(_04303_),
    .C(_03781_),
    .Y(_04304_),
    .A_N(_04200_));
 sg13g2_nor2_1 _09787_ (.A(_03781_),
    .B(_04303_),
    .Y(_04305_));
 sg13g2_nor2_1 _09788_ (.A(_03782_),
    .B(_04199_),
    .Y(_04306_));
 sg13g2_inv_1 _09789_ (.Y(_04307_),
    .A(_04306_));
 sg13g2_o21ai_1 _09790_ (.B1(_04304_),
    .Y(_04308_),
    .A1(_03781_),
    .A2(_04303_));
 sg13g2_nor2_1 _09791_ (.A(net1030),
    .B(_04308_),
    .Y(_04309_));
 sg13g2_xnor2_1 _09792_ (.Y(_04310_),
    .A(net1030),
    .B(_04308_));
 sg13g2_a21o_1 _09793_ (.A2(_04186_),
    .A1(_04176_),
    .B1(_04188_),
    .X(_04311_));
 sg13g2_a21o_1 _09794_ (.A2(_04183_),
    .A1(_04178_),
    .B1(_04185_),
    .X(_04312_));
 sg13g2_o21ai_1 _09795_ (.B1(_04162_),
    .Y(_04313_),
    .A1(_04154_),
    .A2(_04163_));
 sg13g2_o21ai_1 _09796_ (.B1(_04182_),
    .Y(_04314_),
    .A1(_04053_),
    .A2(_04180_));
 sg13g2_o21ai_1 _09797_ (.B1(_04152_),
    .Y(_04315_),
    .A1(_04149_),
    .A2(_04153_));
 sg13g2_nand2_2 _09798_ (.Y(_04316_),
    .A(net1410),
    .B(net1174));
 sg13g2_nor3_1 _09799_ (.A(_04821_),
    .B(_04833_),
    .C(_04180_),
    .Y(_04317_));
 sg13g2_a22oi_1 _09800_ (.Y(_04318_),
    .B1(net1161),
    .B2(net1415),
    .A2(net1167),
    .A1(net1413));
 sg13g2_nor3_1 _09801_ (.A(_04316_),
    .B(_04317_),
    .C(_04318_),
    .Y(_04319_));
 sg13g2_o21ai_1 _09802_ (.B1(_04316_),
    .Y(_04320_),
    .A1(_04317_),
    .A2(_04318_));
 sg13g2_nor2b_1 _09803_ (.A(_04319_),
    .B_N(_04320_),
    .Y(_04321_));
 sg13g2_xnor2_1 _09804_ (.Y(_04322_),
    .A(_04315_),
    .B(_04321_));
 sg13g2_nor2b_1 _09805_ (.A(_04322_),
    .B_N(_04314_),
    .Y(_04323_));
 sg13g2_xnor2_1 _09806_ (.Y(_04324_),
    .A(_04314_),
    .B(_04322_));
 sg13g2_xnor2_1 _09807_ (.Y(_04325_),
    .A(_04313_),
    .B(_04324_));
 sg13g2_nor2b_1 _09808_ (.A(_04325_),
    .B_N(_04312_),
    .Y(_04326_));
 sg13g2_xnor2_1 _09809_ (.Y(_04327_),
    .A(_04312_),
    .B(_04325_));
 sg13g2_nand2_1 _09810_ (.Y(_04328_),
    .A(_04311_),
    .B(_04327_));
 sg13g2_xnor2_1 _09811_ (.Y(_04329_),
    .A(_04311_),
    .B(_04327_));
 sg13g2_xnor2_1 _09812_ (.Y(_04330_),
    .A(_04310_),
    .B(_04329_));
 sg13g2_nor2_1 _09813_ (.A(_04302_),
    .B(_04330_),
    .Y(_04331_));
 sg13g2_xor2_1 _09814_ (.B(_04330_),
    .A(_04302_),
    .X(_04332_));
 sg13g2_xnor2_1 _09815_ (.Y(_04333_),
    .A(_04301_),
    .B(_04332_));
 sg13g2_xor2_1 _09816_ (.B(_04333_),
    .A(_04300_),
    .X(_04334_));
 sg13g2_nand2_1 _09817_ (.Y(_04335_),
    .A(_04232_),
    .B(_04334_));
 sg13g2_xnor2_1 _09818_ (.Y(_04336_),
    .A(_04232_),
    .B(_04334_));
 sg13g2_a21oi_1 _09819_ (.A1(_04172_),
    .A2(_04208_),
    .Y(_04337_),
    .B1(_04207_));
 sg13g2_o21ai_1 _09820_ (.B1(_04203_),
    .Y(_04338_),
    .A1(_04193_),
    .A2(_04201_));
 sg13g2_nand2b_1 _09821_ (.Y(_04339_),
    .B(_04338_),
    .A_N(_04337_));
 sg13g2_xor2_1 _09822_ (.B(_04338_),
    .A(_04337_),
    .X(_04340_));
 sg13g2_xnor2_1 _09823_ (.Y(_04341_),
    .A(_04086_),
    .B(_04340_));
 sg13g2_nand2b_1 _09824_ (.Y(_04342_),
    .B(_04341_),
    .A_N(_04336_));
 sg13g2_xnor2_1 _09825_ (.Y(_04343_),
    .A(_04336_),
    .B(_04341_));
 sg13g2_nor2b_1 _09826_ (.A(_04231_),
    .B_N(_04343_),
    .Y(_04344_));
 sg13g2_xnor2_1 _09827_ (.Y(_04345_),
    .A(_04231_),
    .B(_04343_));
 sg13g2_xor2_1 _09828_ (.B(_04345_),
    .A(_04230_),
    .X(_04346_));
 sg13g2_nand2_1 _09829_ (.Y(_04347_),
    .A(_04229_),
    .B(_04346_));
 sg13g2_xnor2_1 _09830_ (.Y(_04348_),
    .A(_04229_),
    .B(_04346_));
 sg13g2_inv_1 _09831_ (.Y(_04349_),
    .A(_04348_));
 sg13g2_o21ai_1 _09832_ (.B1(_04349_),
    .Y(_04350_),
    .A1(_04223_),
    .A2(_04225_));
 sg13g2_or3_1 _09833_ (.A(_04223_),
    .B(_04225_),
    .C(_04349_),
    .X(_04351_));
 sg13g2_nand2_1 _09834_ (.Y(_04352_),
    .A(_04350_),
    .B(_04351_));
 sg13g2_o21ai_1 _09835_ (.B1(net1498),
    .Y(_04353_),
    .A1(net1296),
    .A2(net276));
 sg13g2_a21oi_1 _09836_ (.A1(net1296),
    .A2(_04352_),
    .Y(_00245_),
    .B1(net277));
 sg13g2_a21o_1 _09837_ (.A2(_04345_),
    .A1(_04230_),
    .B1(_04344_),
    .X(_04354_));
 sg13g2_o21ai_1 _09838_ (.B1(_04339_),
    .Y(_04355_),
    .A1(_04087_),
    .A2(_04340_));
 sg13g2_and2_1 _09839_ (.A(_04335_),
    .B(_04342_),
    .X(_04356_));
 sg13g2_a21oi_1 _09840_ (.A1(_04301_),
    .A2(_04332_),
    .Y(_04357_),
    .B1(_04331_));
 sg13g2_nor2_1 _09841_ (.A(_04306_),
    .B(_04309_),
    .Y(_04358_));
 sg13g2_or2_1 _09842_ (.X(_04359_),
    .B(_04358_),
    .A(_04357_));
 sg13g2_xnor2_1 _09843_ (.Y(_04360_),
    .A(_04357_),
    .B(_04358_));
 sg13g2_xnor2_1 _09844_ (.Y(_04361_),
    .A(_04086_),
    .B(_04360_));
 sg13g2_o21ai_1 _09845_ (.B1(_04299_),
    .Y(_04362_),
    .A1(_04300_),
    .A2(_04333_));
 sg13g2_o21ai_1 _09846_ (.B1(_04328_),
    .Y(_04363_),
    .A1(_04310_),
    .A2(_04329_));
 sg13g2_a21oi_1 _09847_ (.A1(_04265_),
    .A2(_04294_),
    .Y(_04364_),
    .B1(_04296_));
 sg13g2_nor2_1 _09848_ (.A(_04305_),
    .B(_04306_),
    .Y(_04365_));
 sg13g2_xnor2_1 _09849_ (.Y(_04366_),
    .A(net1030),
    .B(_04365_));
 sg13g2_inv_1 _09850_ (.Y(_04367_),
    .A(_04366_));
 sg13g2_a21o_1 _09851_ (.A2(_04324_),
    .A1(_04313_),
    .B1(_04326_),
    .X(_04368_));
 sg13g2_a21o_1 _09852_ (.A2(_04321_),
    .A1(_04315_),
    .B1(_04323_),
    .X(_04369_));
 sg13g2_o21ai_1 _09853_ (.B1(_04291_),
    .Y(_04370_),
    .A1(_04284_),
    .A2(_04292_));
 sg13g2_or2_1 _09854_ (.X(_04371_),
    .B(_04319_),
    .A(_04317_));
 sg13g2_o21ai_1 _09855_ (.B1(_04283_),
    .Y(_04372_),
    .A1(_04150_),
    .A2(_04281_));
 sg13g2_and4_1 _09856_ (.A(net1413),
    .B(net1410),
    .C(net1167),
    .D(net1161),
    .X(_04373_));
 sg13g2_a22oi_1 _09857_ (.Y(_04374_),
    .B1(net1161),
    .B2(net1413),
    .A2(net1167),
    .A1(net1410));
 sg13g2_nor3_1 _09858_ (.A(_04316_),
    .B(_04373_),
    .C(_04374_),
    .Y(_04375_));
 sg13g2_o21ai_1 _09859_ (.B1(_04316_),
    .Y(_04376_),
    .A1(_04373_),
    .A2(_04374_));
 sg13g2_nor2b_1 _09860_ (.A(_04375_),
    .B_N(_04376_),
    .Y(_04377_));
 sg13g2_xnor2_1 _09861_ (.Y(_04378_),
    .A(_04372_),
    .B(_04377_));
 sg13g2_nor2b_1 _09862_ (.A(_04378_),
    .B_N(_04371_),
    .Y(_04379_));
 sg13g2_xnor2_1 _09863_ (.Y(_04380_),
    .A(_04371_),
    .B(_04378_));
 sg13g2_xnor2_1 _09864_ (.Y(_04381_),
    .A(_04370_),
    .B(_04380_));
 sg13g2_nor2b_1 _09865_ (.A(_04381_),
    .B_N(_04369_),
    .Y(_04382_));
 sg13g2_xnor2_1 _09866_ (.Y(_04383_),
    .A(_04369_),
    .B(_04381_));
 sg13g2_xnor2_1 _09867_ (.Y(_04384_),
    .A(_04368_),
    .B(_04383_));
 sg13g2_nor2_1 _09868_ (.A(_04367_),
    .B(_04384_),
    .Y(_04385_));
 sg13g2_xnor2_1 _09869_ (.Y(_04386_),
    .A(_04367_),
    .B(_04384_));
 sg13g2_xor2_1 _09870_ (.B(_04386_),
    .A(_04364_),
    .X(_04387_));
 sg13g2_nand2_1 _09871_ (.Y(_04388_),
    .A(_04363_),
    .B(_04387_));
 sg13g2_xnor2_1 _09872_ (.Y(_04389_),
    .A(_04363_),
    .B(_04387_));
 sg13g2_o21ai_1 _09873_ (.B1(_04262_),
    .Y(_04390_),
    .A1(_04263_),
    .A2(_04297_));
 sg13g2_o21ai_1 _09874_ (.B1(_04277_),
    .Y(_04391_),
    .A1(_04278_),
    .A2(_04293_));
 sg13g2_a21oi_1 _09875_ (.A1(_04245_),
    .A2(_04258_),
    .Y(_04392_),
    .B1(_04257_));
 sg13g2_a21o_1 _09876_ (.A2(_04273_),
    .A1(_04268_),
    .B1(_04275_),
    .X(_04393_));
 sg13g2_o21ai_1 _09877_ (.B1(_04271_),
    .Y(_04394_),
    .A1(_04269_),
    .A2(_04272_));
 sg13g2_o21ai_1 _09878_ (.B1(_04247_),
    .Y(_04395_),
    .A1(_04248_),
    .A2(_04249_));
 sg13g2_nand2_1 _09879_ (.Y(_04396_),
    .A(net1436),
    .B(net1334));
 sg13g2_nand2_1 _09880_ (.Y(_04397_),
    .A(net1441),
    .B(net1329));
 sg13g2_nor2_1 _09881_ (.A(_04270_),
    .B(_04397_),
    .Y(_04398_));
 sg13g2_or2_1 _09882_ (.X(_04399_),
    .B(_04397_),
    .A(_04270_));
 sg13g2_a22oi_1 _09883_ (.Y(_04400_),
    .B1(net1329),
    .B2(net1446),
    .A2(net1331),
    .A1(net1441));
 sg13g2_nor2_1 _09884_ (.A(_04398_),
    .B(_04400_),
    .Y(_04401_));
 sg13g2_xnor2_1 _09885_ (.Y(_04402_),
    .A(_04396_),
    .B(_04401_));
 sg13g2_xnor2_1 _09886_ (.Y(_04403_),
    .A(_04395_),
    .B(_04402_));
 sg13g2_nor2b_1 _09887_ (.A(_04403_),
    .B_N(_04394_),
    .Y(_04404_));
 sg13g2_xnor2_1 _09888_ (.Y(_04405_),
    .A(_04394_),
    .B(_04403_));
 sg13g2_xnor2_1 _09889_ (.Y(_04406_),
    .A(_04393_),
    .B(_04405_));
 sg13g2_nand2_1 _09890_ (.Y(_04407_),
    .A(net1415),
    .B(net1157));
 sg13g2_nand2_1 _09891_ (.Y(_04408_),
    .A(net1418),
    .B(net1145));
 sg13g2_nand2_1 _09892_ (.Y(_04409_),
    .A(net1418),
    .B(net1151));
 sg13g2_xor2_1 _09893_ (.B(_04409_),
    .A(_04280_),
    .X(_04410_));
 sg13g2_nand2b_1 _09894_ (.Y(_04411_),
    .B(_04410_),
    .A_N(_04407_));
 sg13g2_xor2_1 _09895_ (.B(_04410_),
    .A(_04407_),
    .X(_04412_));
 sg13g2_o21ai_1 _09896_ (.B1(_04289_),
    .Y(_04413_),
    .A1(_04157_),
    .A2(_04287_));
 sg13g2_nand2_1 _09897_ (.Y(_04414_),
    .A(net1424),
    .B(net1348));
 sg13g2_nand2_1 _09898_ (.Y(_04415_),
    .A(net1428),
    .B(net1337));
 sg13g2_nor2_1 _09899_ (.A(_04287_),
    .B(_04415_),
    .Y(_04416_));
 sg13g2_or2_1 _09900_ (.X(_04417_),
    .B(_04415_),
    .A(_04287_));
 sg13g2_a22oi_1 _09901_ (.Y(_04418_),
    .B1(net1337),
    .B2(net1432),
    .A2(net1342),
    .A1(net1428));
 sg13g2_nor2_1 _09902_ (.A(_04416_),
    .B(_04418_),
    .Y(_04419_));
 sg13g2_xnor2_1 _09903_ (.Y(_04420_),
    .A(_04414_),
    .B(_04419_));
 sg13g2_xnor2_1 _09904_ (.Y(_04421_),
    .A(_04413_),
    .B(_04420_));
 sg13g2_nor2_1 _09905_ (.A(_04412_),
    .B(_04421_),
    .Y(_04422_));
 sg13g2_xnor2_1 _09906_ (.Y(_04423_),
    .A(_04412_),
    .B(_04421_));
 sg13g2_nor2_1 _09907_ (.A(_04406_),
    .B(_04423_),
    .Y(_04424_));
 sg13g2_xnor2_1 _09908_ (.Y(_04425_),
    .A(_04406_),
    .B(_04423_));
 sg13g2_nor2_1 _09909_ (.A(_04392_),
    .B(_04425_),
    .Y(_04426_));
 sg13g2_xor2_1 _09910_ (.B(_04425_),
    .A(_04392_),
    .X(_04427_));
 sg13g2_xnor2_1 _09911_ (.Y(_04428_),
    .A(_04391_),
    .B(_04427_));
 sg13g2_a21oi_1 _09912_ (.A1(_04244_),
    .A2(_04260_),
    .Y(_04429_),
    .B1(_04243_));
 sg13g2_o21ai_1 _09913_ (.B1(_04254_),
    .Y(_04430_),
    .A1(_04251_),
    .A2(_04255_));
 sg13g2_a21o_2 _09914_ (.A2(_04237_),
    .A1(_03850_),
    .B1(_04236_),
    .X(_04431_));
 sg13g2_nand2_1 _09915_ (.Y(_04432_),
    .A(net1455),
    .B(_04246_));
 sg13g2_o21ai_1 _09916_ (.B1(net1322),
    .Y(_04433_),
    .A1(net1460),
    .A2(net1455));
 sg13g2_a21oi_1 _09917_ (.A1(net1456),
    .A2(_04246_),
    .Y(_04434_),
    .B1(_04433_));
 sg13g2_nand2_1 _09918_ (.Y(_04435_),
    .A(net1451),
    .B(net1326));
 sg13g2_xor2_1 _09919_ (.B(_04435_),
    .A(_04434_),
    .X(_04436_));
 sg13g2_o21ai_1 _09920_ (.B1(_03856_),
    .Y(_04437_),
    .A1(_03857_),
    .A2(_03991_));
 sg13g2_xnor2_1 _09921_ (.Y(_04438_),
    .A(_03993_),
    .B(_04116_));
 sg13g2_nand2_1 _09922_ (.Y(_04439_),
    .A(_04437_),
    .B(_04438_));
 sg13g2_xnor2_1 _09923_ (.Y(_04440_),
    .A(_04437_),
    .B(_04438_));
 sg13g2_xor2_1 _09924_ (.B(_04440_),
    .A(_04436_),
    .X(_04441_));
 sg13g2_xnor2_1 _09925_ (.Y(_04442_),
    .A(_04431_),
    .B(_04441_));
 sg13g2_nor2b_1 _09926_ (.A(_04442_),
    .B_N(_04430_),
    .Y(_04443_));
 sg13g2_xor2_1 _09927_ (.B(_04442_),
    .A(_04430_),
    .X(_04444_));
 sg13g2_a22oi_1 _09928_ (.Y(_04445_),
    .B1(_04239_),
    .B2(_04241_),
    .A2(_03470_),
    .A1(_03080_));
 sg13g2_nor2b_1 _09929_ (.A(_03577_),
    .B_N(_03988_),
    .Y(_04446_));
 sg13g2_xnor2_1 _09930_ (.Y(_04447_),
    .A(_03577_),
    .B(_03988_));
 sg13g2_xor2_1 _09931_ (.B(_04447_),
    .A(_03987_),
    .X(_04448_));
 sg13g2_nand2_1 _09932_ (.Y(_04449_),
    .A(_03575_),
    .B(_03579_));
 sg13g2_xnor2_1 _09933_ (.Y(_04450_),
    .A(_03575_),
    .B(_03579_));
 sg13g2_nor3_1 _09934_ (.A(net1118),
    .B(_03471_),
    .C(_04450_),
    .Y(_04451_));
 sg13g2_o21ai_1 _09935_ (.B1(_04450_),
    .Y(_04452_),
    .A1(net1118),
    .A2(_03471_));
 sg13g2_nor2b_1 _09936_ (.A(_04451_),
    .B_N(_04452_),
    .Y(_04453_));
 sg13g2_xor2_1 _09937_ (.B(_04453_),
    .A(_04448_),
    .X(_04454_));
 sg13g2_nand2b_1 _09938_ (.Y(_04455_),
    .B(_04454_),
    .A_N(_04445_));
 sg13g2_xnor2_1 _09939_ (.Y(_04456_),
    .A(_04445_),
    .B(_04454_));
 sg13g2_nand2b_1 _09940_ (.Y(_04457_),
    .B(_04456_),
    .A_N(_04444_));
 sg13g2_xnor2_1 _09941_ (.Y(_04458_),
    .A(_04444_),
    .B(_04456_));
 sg13g2_nand2b_1 _09942_ (.Y(_04459_),
    .B(_04458_),
    .A_N(_04429_));
 sg13g2_xnor2_1 _09943_ (.Y(_04460_),
    .A(_04429_),
    .B(_04458_));
 sg13g2_nand2b_1 _09944_ (.Y(_04461_),
    .B(_04460_),
    .A_N(_04428_));
 sg13g2_xnor2_1 _09945_ (.Y(_04462_),
    .A(_04428_),
    .B(_04460_));
 sg13g2_nand2_1 _09946_ (.Y(_04463_),
    .A(_04390_),
    .B(_04462_));
 sg13g2_xnor2_1 _09947_ (.Y(_04464_),
    .A(_04390_),
    .B(_04462_));
 sg13g2_xor2_1 _09948_ (.B(_04464_),
    .A(_04389_),
    .X(_04465_));
 sg13g2_and2_1 _09949_ (.A(_04362_),
    .B(_04465_),
    .X(_04466_));
 sg13g2_xor2_1 _09950_ (.B(_04465_),
    .A(_04362_),
    .X(_04467_));
 sg13g2_xor2_1 _09951_ (.B(_04467_),
    .A(_04361_),
    .X(_04468_));
 sg13g2_nor2b_1 _09952_ (.A(_04356_),
    .B_N(_04468_),
    .Y(_04469_));
 sg13g2_xnor2_1 _09953_ (.Y(_04470_),
    .A(_04356_),
    .B(_04468_));
 sg13g2_xor2_1 _09954_ (.B(_04470_),
    .A(_04355_),
    .X(_04471_));
 sg13g2_xnor2_1 _09955_ (.Y(_04472_),
    .A(_04354_),
    .B(_04471_));
 sg13g2_a21oi_1 _09956_ (.A1(_04347_),
    .A2(_04350_),
    .Y(_04473_),
    .B1(_04472_));
 sg13g2_nand3_1 _09957_ (.B(_04350_),
    .C(_04472_),
    .A(_04347_),
    .Y(_04474_));
 sg13g2_nand2b_2 _09958_ (.Y(_04475_),
    .B(_04474_),
    .A_N(_04473_));
 sg13g2_o21ai_1 _09959_ (.B1(net1499),
    .Y(_04476_),
    .A1(net1296),
    .A2(net260));
 sg13g2_a21oi_1 _09960_ (.A1(net1296),
    .A2(_04475_),
    .Y(_00246_),
    .B1(net261));
 sg13g2_a21oi_1 _09961_ (.A1(_04354_),
    .A2(_04471_),
    .Y(_04477_),
    .B1(_04473_));
 sg13g2_a21oi_1 _09962_ (.A1(_04355_),
    .A2(_04470_),
    .Y(_04478_),
    .B1(_04469_));
 sg13g2_o21ai_1 _09963_ (.B1(_04359_),
    .Y(_04479_),
    .A1(_04087_),
    .A2(_04360_));
 sg13g2_a21oi_1 _09964_ (.A1(_04361_),
    .A2(_04467_),
    .Y(_04480_),
    .B1(_04466_));
 sg13g2_o21ai_1 _09965_ (.B1(_04463_),
    .Y(_04481_),
    .A1(_04389_),
    .A2(_04464_));
 sg13g2_o21ai_1 _09966_ (.B1(_04388_),
    .Y(_04482_),
    .A1(_04364_),
    .A2(_04386_));
 sg13g2_xnor2_1 _09967_ (.Y(_04483_),
    .A(_04481_),
    .B(_04482_));
 sg13g2_o21ai_1 _09968_ (.B1(_04307_),
    .Y(_04484_),
    .A1(net1030),
    .A2(_04305_));
 sg13g2_xnor2_1 _09969_ (.Y(_04485_),
    .A(_04087_),
    .B(_04484_));
 sg13g2_a21oi_1 _09970_ (.A1(_04368_),
    .A2(_04383_),
    .Y(_04486_),
    .B1(_04385_));
 sg13g2_nand2_1 _09971_ (.Y(_04487_),
    .A(_04459_),
    .B(_04461_));
 sg13g2_xnor2_1 _09972_ (.Y(_04488_),
    .A(_04486_),
    .B(_04487_));
 sg13g2_nand2_1 _09973_ (.Y(_04489_),
    .A(_04455_),
    .B(_04457_));
 sg13g2_a21oi_1 _09974_ (.A1(_04393_),
    .A2(_04405_),
    .Y(_04490_),
    .B1(_04424_));
 sg13g2_xnor2_1 _09975_ (.Y(_04491_),
    .A(_04489_),
    .B(_04490_));
 sg13g2_a21oi_1 _09976_ (.A1(_04372_),
    .A2(_04377_),
    .Y(_04492_),
    .B1(_04379_));
 sg13g2_xor2_1 _09977_ (.B(net1162),
    .A(net1168),
    .X(_04493_));
 sg13g2_a21oi_1 _09978_ (.A1(net1174),
    .A2(_04493_),
    .Y(_04494_),
    .B1(_04822_));
 sg13g2_o21ai_1 _09979_ (.B1(_04494_),
    .Y(_04495_),
    .A1(net1174),
    .A2(_04493_));
 sg13g2_nor2_1 _09980_ (.A(_04373_),
    .B(_04375_),
    .Y(_04496_));
 sg13g2_o21ai_1 _09981_ (.B1(_04411_),
    .Y(_04497_),
    .A1(_04280_),
    .A2(_04409_));
 sg13g2_xnor2_1 _09982_ (.Y(_04498_),
    .A(_04496_),
    .B(_04497_));
 sg13g2_xnor2_1 _09983_ (.Y(_04499_),
    .A(_04495_),
    .B(_04498_));
 sg13g2_xnor2_1 _09984_ (.Y(_04500_),
    .A(_04492_),
    .B(_04499_));
 sg13g2_a21oi_1 _09985_ (.A1(_04413_),
    .A2(_04420_),
    .Y(_04501_),
    .B1(_04422_));
 sg13g2_a21oi_1 _09986_ (.A1(_04370_),
    .A2(_04380_),
    .Y(_04502_),
    .B1(_04382_));
 sg13g2_xnor2_1 _09987_ (.Y(_04503_),
    .A(_04366_),
    .B(_04501_));
 sg13g2_xnor2_1 _09988_ (.Y(_04504_),
    .A(_04502_),
    .B(_04503_));
 sg13g2_xnor2_1 _09989_ (.Y(_04505_),
    .A(_04500_),
    .B(_04504_));
 sg13g2_xnor2_1 _09990_ (.Y(_04506_),
    .A(_04491_),
    .B(_04505_));
 sg13g2_xor2_1 _09991_ (.B(_03727_),
    .A(_03712_),
    .X(_04507_));
 sg13g2_xnor2_1 _09992_ (.Y(_04508_),
    .A(_04449_),
    .B(_04507_));
 sg13g2_xor2_1 _09993_ (.B(_04125_),
    .A(_03711_),
    .X(_04509_));
 sg13g2_o21ai_1 _09994_ (.B1(_03992_),
    .Y(_04510_),
    .A1(_03993_),
    .A2(_04117_));
 sg13g2_o21ai_1 _09995_ (.B1(net1323),
    .Y(_04511_),
    .A1(net1455),
    .A2(net1451));
 sg13g2_a21oi_1 _09996_ (.A1(net1455),
    .A2(net1451),
    .Y(_04512_),
    .B1(_04511_));
 sg13g2_nand2_1 _09997_ (.Y(_04513_),
    .A(net1446),
    .B(net1326));
 sg13g2_xnor2_1 _09998_ (.Y(_04514_),
    .A(_04512_),
    .B(_04513_));
 sg13g2_xor2_1 _09999_ (.B(_04246_),
    .A(_04119_),
    .X(_04515_));
 sg13g2_xnor2_1 _10000_ (.Y(_04516_),
    .A(_04510_),
    .B(_04515_));
 sg13g2_xnor2_1 _10001_ (.Y(_04517_),
    .A(_04514_),
    .B(_04516_));
 sg13g2_o21ai_1 _10002_ (.B1(_04439_),
    .Y(_04518_),
    .A1(_04436_),
    .A2(_04440_));
 sg13g2_xnor2_1 _10003_ (.Y(_04519_),
    .A(_04508_),
    .B(_04517_));
 sg13g2_xnor2_1 _10004_ (.Y(_04520_),
    .A(_04509_),
    .B(_04518_));
 sg13g2_xnor2_1 _10005_ (.Y(_04521_),
    .A(_04519_),
    .B(_04520_));
 sg13g2_nand2_1 _10006_ (.Y(_04522_),
    .A(net1413),
    .B(net1157));
 sg13g2_o21ai_1 _10007_ (.B1(_04417_),
    .Y(_04523_),
    .A1(_04414_),
    .A2(_04418_));
 sg13g2_xnor2_1 _10008_ (.Y(_04524_),
    .A(_04522_),
    .B(_04523_));
 sg13g2_nand2_1 _10009_ (.Y(_04525_),
    .A(net1436),
    .B(net1331));
 sg13g2_xnor2_1 _10010_ (.Y(_04526_),
    .A(_04397_),
    .B(_04525_));
 sg13g2_nand2_1 _10011_ (.Y(_04527_),
    .A(net1421),
    .B(net1348));
 sg13g2_nand2_1 _10012_ (.Y(_04528_),
    .A(net1432),
    .B(net1334));
 sg13g2_xor2_1 _10013_ (.B(_04528_),
    .A(_04527_),
    .X(_04529_));
 sg13g2_xnor2_1 _10014_ (.Y(_04530_),
    .A(_04526_),
    .B(_04529_));
 sg13g2_nand2_1 _10015_ (.Y(_04531_),
    .A(net1415),
    .B(net1151));
 sg13g2_xor2_1 _10016_ (.B(_04531_),
    .A(_04408_),
    .X(_04532_));
 sg13g2_nand2_1 _10017_ (.Y(_04533_),
    .A(net1424),
    .B(net1342));
 sg13g2_xor2_1 _10018_ (.B(_04533_),
    .A(_04415_),
    .X(_04534_));
 sg13g2_xnor2_1 _10019_ (.Y(_04535_),
    .A(_04532_),
    .B(_04534_));
 sg13g2_o21ai_1 _10020_ (.B1(_04399_),
    .Y(_04536_),
    .A1(_04396_),
    .A2(_04400_));
 sg13g2_xnor2_1 _10021_ (.Y(_04537_),
    .A(_04535_),
    .B(_04536_));
 sg13g2_xnor2_1 _10022_ (.Y(_04538_),
    .A(_04530_),
    .B(_04537_));
 sg13g2_xnor2_1 _10023_ (.Y(_04539_),
    .A(_04524_),
    .B(_04538_));
 sg13g2_a21oi_1 _10024_ (.A1(_04395_),
    .A2(_04402_),
    .Y(_04540_),
    .B1(_04404_));
 sg13g2_o21ai_1 _10025_ (.B1(_04432_),
    .Y(_04541_),
    .A1(_04433_),
    .A2(_04435_));
 sg13g2_xnor2_1 _10026_ (.Y(_04542_),
    .A(_04540_),
    .B(_04541_));
 sg13g2_xnor2_1 _10027_ (.Y(_04543_),
    .A(_04539_),
    .B(_04542_));
 sg13g2_xnor2_1 _10028_ (.Y(_04544_),
    .A(_04521_),
    .B(_04543_));
 sg13g2_a21oi_1 _10029_ (.A1(_04448_),
    .A2(_04453_),
    .Y(_04545_),
    .B1(_04451_));
 sg13g2_a21oi_1 _10030_ (.A1(_03987_),
    .A2(_04447_),
    .Y(_04546_),
    .B1(_04446_));
 sg13g2_xnor2_1 _10031_ (.Y(_04547_),
    .A(_04545_),
    .B(_04546_));
 sg13g2_a21oi_1 _10032_ (.A1(_04431_),
    .A2(_04441_),
    .Y(_04548_),
    .B1(_04443_));
 sg13g2_xnor2_1 _10033_ (.Y(_04549_),
    .A(_04547_),
    .B(_04548_));
 sg13g2_xnor2_1 _10034_ (.Y(_04550_),
    .A(_04544_),
    .B(_04549_));
 sg13g2_a21oi_1 _10035_ (.A1(_04391_),
    .A2(_04427_),
    .Y(_04551_),
    .B1(_04426_));
 sg13g2_xnor2_1 _10036_ (.Y(_04552_),
    .A(_04550_),
    .B(_04551_));
 sg13g2_xnor2_1 _10037_ (.Y(_04553_),
    .A(_04506_),
    .B(_04552_));
 sg13g2_xnor2_1 _10038_ (.Y(_04554_),
    .A(_04488_),
    .B(_04553_));
 sg13g2_xnor2_1 _10039_ (.Y(_04555_),
    .A(_04485_),
    .B(_04554_));
 sg13g2_xnor2_1 _10040_ (.Y(_04556_),
    .A(_04483_),
    .B(_04555_));
 sg13g2_xnor2_1 _10041_ (.Y(_04557_),
    .A(_04480_),
    .B(_04556_));
 sg13g2_xor2_1 _10042_ (.B(_04557_),
    .A(_04479_),
    .X(_04558_));
 sg13g2_xnor2_1 _10043_ (.Y(_04559_),
    .A(_04478_),
    .B(_04558_));
 sg13g2_xnor2_1 _10044_ (.Y(_04560_),
    .A(_04477_),
    .B(_04559_));
 sg13g2_o21ai_1 _10045_ (.B1(net1507),
    .Y(_04561_),
    .A1(net1141),
    .A2(_04560_));
 sg13g2_a21oi_1 _10046_ (.A1(_04769_),
    .A2(net1141),
    .Y(_00247_),
    .B1(_04561_));
 sg13g2_nor2_1 _10047_ (.A(net1295),
    .B(mac_en_clear),
    .Y(_04562_));
 sg13g2_nand2_2 _10048_ (.Y(_04563_),
    .A(net397),
    .B(_01875_));
 sg13g2_inv_1 _10049_ (.Y(_04564_),
    .A(_04563_));
 sg13g2_o21ai_1 _10050_ (.B1(net1294),
    .Y(_04565_),
    .A1(net397),
    .A2(_01875_));
 sg13g2_inv_1 _10051_ (.Y(_04566_),
    .A(_04565_));
 sg13g2_a22oi_1 _10052_ (.Y(_04567_),
    .B1(_04563_),
    .B2(_04566_),
    .A2(net1115),
    .A1(net397));
 sg13g2_nor2_1 _10053_ (.A(net1485),
    .B(_04567_),
    .Y(_00248_));
 sg13g2_nor2b_1 _10054_ (.A(_01958_),
    .B_N(\mac_inst.accumulator[1] ),
    .Y(_04568_));
 sg13g2_nand2b_1 _10055_ (.Y(_04569_),
    .B(_01958_),
    .A_N(net281));
 sg13g2_nand2b_1 _10056_ (.Y(_04570_),
    .B(_04569_),
    .A_N(_04568_));
 sg13g2_o21ai_1 _10057_ (.B1(net1294),
    .Y(_04571_),
    .A1(_04563_),
    .A2(_04570_));
 sg13g2_a21oi_1 _10058_ (.A1(_04563_),
    .A2(_04570_),
    .Y(_04572_),
    .B1(_04571_));
 sg13g2_a21oi_1 _10059_ (.A1(net281),
    .A2(net1115),
    .Y(_04573_),
    .B1(_04572_));
 sg13g2_nor2_1 _10060_ (.A(net1485),
    .B(net282),
    .Y(_00249_));
 sg13g2_a21oi_1 _10061_ (.A1(_04564_),
    .A2(_04569_),
    .Y(_04574_),
    .B1(_04568_));
 sg13g2_or2_1 _10062_ (.X(_04575_),
    .B(_02043_),
    .A(_04768_));
 sg13g2_xnor2_1 _10063_ (.Y(_04576_),
    .A(_04768_),
    .B(_02043_));
 sg13g2_o21ai_1 _10064_ (.B1(net1294),
    .Y(_04577_),
    .A1(_04574_),
    .A2(_04576_));
 sg13g2_a21oi_1 _10065_ (.A1(_04574_),
    .A2(_04576_),
    .Y(_04578_),
    .B1(_04577_));
 sg13g2_a21oi_1 _10066_ (.A1(net315),
    .A2(net1115),
    .Y(_04579_),
    .B1(_04578_));
 sg13g2_nor2_1 _10067_ (.A(net1486),
    .B(net316),
    .Y(_00250_));
 sg13g2_o21ai_1 _10068_ (.B1(_04575_),
    .Y(_04580_),
    .A1(_04574_),
    .A2(_04576_));
 sg13g2_nor2b_1 _10069_ (.A(_02126_),
    .B_N(\mac_inst.accumulator[3] ),
    .Y(_04581_));
 sg13g2_xnor2_1 _10070_ (.Y(_04582_),
    .A(net393),
    .B(_02126_));
 sg13g2_or2_1 _10071_ (.X(_04583_),
    .B(_04582_),
    .A(_04580_));
 sg13g2_a21oi_1 _10072_ (.A1(_04580_),
    .A2(_04582_),
    .Y(_04584_),
    .B1(_04803_));
 sg13g2_a22oi_1 _10073_ (.Y(_04585_),
    .B1(_04583_),
    .B2(_04584_),
    .A2(net1115),
    .A1(net393));
 sg13g2_nor2_1 _10074_ (.A(net1486),
    .B(net394),
    .Y(_00251_));
 sg13g2_nand2_1 _10075_ (.Y(_04586_),
    .A(net559),
    .B(_02224_));
 sg13g2_xnor2_1 _10076_ (.Y(_04587_),
    .A(net385),
    .B(_02224_));
 sg13g2_a21oi_1 _10077_ (.A1(_04580_),
    .A2(_04582_),
    .Y(_04588_),
    .B1(_04581_));
 sg13g2_nor2_1 _10078_ (.A(_04587_),
    .B(_04588_),
    .Y(_04589_));
 sg13g2_nand2_1 _10079_ (.Y(_04590_),
    .A(_04587_),
    .B(_04588_));
 sg13g2_nor2_1 _10080_ (.A(_04803_),
    .B(_04589_),
    .Y(_04591_));
 sg13g2_a22oi_1 _10081_ (.Y(_04592_),
    .B1(_04590_),
    .B2(_04591_),
    .A2(net1114),
    .A1(net385));
 sg13g2_nor2_1 _10082_ (.A(net1486),
    .B(net386),
    .Y(_00252_));
 sg13g2_nand2_1 _10083_ (.Y(_04593_),
    .A(net267),
    .B(net1114));
 sg13g2_xnor2_1 _10084_ (.Y(_04594_),
    .A(\mac_inst.accumulator[5] ),
    .B(_02327_));
 sg13g2_nand2_1 _10085_ (.Y(_04595_),
    .A(_04586_),
    .B(_04594_));
 sg13g2_or2_1 _10086_ (.X(_04596_),
    .B(_04595_),
    .A(_04589_));
 sg13g2_or3_1 _10087_ (.A(_04587_),
    .B(_04588_),
    .C(_04594_),
    .X(_04597_));
 sg13g2_nor2_1 _10088_ (.A(_04586_),
    .B(_04594_),
    .Y(_04598_));
 sg13g2_o21ai_1 _10089_ (.B1(net1294),
    .Y(_04599_),
    .A1(_04586_),
    .A2(_04594_));
 sg13g2_nand3b_1 _10090_ (.B(_04597_),
    .C(_04596_),
    .Y(_04600_),
    .A_N(_04599_));
 sg13g2_a21oi_1 _10091_ (.A1(net268),
    .A2(_04600_),
    .Y(_00253_),
    .B1(net1486));
 sg13g2_a21oi_1 _10092_ (.A1(\mac_inst.accumulator[5] ),
    .A2(_02327_),
    .Y(_04601_),
    .B1(_04598_));
 sg13g2_and2_1 _10093_ (.A(_04597_),
    .B(_04601_),
    .X(_04602_));
 sg13g2_nand2_1 _10094_ (.Y(_04603_),
    .A(\mac_inst.accumulator[6] ),
    .B(_02433_));
 sg13g2_xnor2_1 _10095_ (.Y(_04604_),
    .A(net387),
    .B(_02433_));
 sg13g2_or2_1 _10096_ (.X(_04605_),
    .B(_04604_),
    .A(_04602_));
 sg13g2_a21oi_1 _10097_ (.A1(_04602_),
    .A2(_04604_),
    .Y(_04606_),
    .B1(_04803_));
 sg13g2_a22oi_1 _10098_ (.Y(_04607_),
    .B1(_04605_),
    .B2(_04606_),
    .A2(net1114),
    .A1(net387));
 sg13g2_nor2_1 _10099_ (.A(net1485),
    .B(net388),
    .Y(_00254_));
 sg13g2_nand2_1 _10100_ (.Y(_04608_),
    .A(_04603_),
    .B(_04605_));
 sg13g2_nand2b_1 _10101_ (.Y(_04609_),
    .B(\mac_inst.accumulator[7] ),
    .A_N(_02541_));
 sg13g2_nor2b_1 _10102_ (.A(\mac_inst.accumulator[7] ),
    .B_N(_02541_),
    .Y(_04610_));
 sg13g2_xnor2_1 _10103_ (.Y(_04611_),
    .A(net347),
    .B(_02541_));
 sg13g2_o21ai_1 _10104_ (.B1(net1294),
    .Y(_04612_),
    .A1(_04608_),
    .A2(_04611_));
 sg13g2_a21oi_1 _10105_ (.A1(_04608_),
    .A2(_04611_),
    .Y(_04613_),
    .B1(_04612_));
 sg13g2_a21oi_1 _10106_ (.A1(net347),
    .A2(net1114),
    .Y(_04614_),
    .B1(_04613_));
 sg13g2_nor2_1 _10107_ (.A(net1485),
    .B(net348),
    .Y(_00255_));
 sg13g2_nor2_1 _10108_ (.A(_04767_),
    .B(_02656_),
    .Y(_04615_));
 sg13g2_xnor2_1 _10109_ (.Y(_04616_),
    .A(_04767_),
    .B(_02656_));
 sg13g2_inv_1 _10110_ (.Y(_04617_),
    .A(_04616_));
 sg13g2_nand2b_1 _10111_ (.Y(_04618_),
    .B(_04611_),
    .A_N(_04604_));
 sg13g2_a21oi_1 _10112_ (.A1(_04597_),
    .A2(_04601_),
    .Y(_04619_),
    .B1(_04618_));
 sg13g2_a21oi_1 _10113_ (.A1(_04603_),
    .A2(_04609_),
    .Y(_04620_),
    .B1(_04610_));
 sg13g2_or2_1 _10114_ (.X(_04621_),
    .B(_04620_),
    .A(_04619_));
 sg13g2_and2_1 _10115_ (.A(_04617_),
    .B(_04621_),
    .X(_04622_));
 sg13g2_o21ai_1 _10116_ (.B1(net1294),
    .Y(_04623_),
    .A1(_04617_),
    .A2(_04621_));
 sg13g2_nor2_1 _10117_ (.A(_04622_),
    .B(_04623_),
    .Y(_04624_));
 sg13g2_a21oi_1 _10118_ (.A1(net254),
    .A2(net1114),
    .Y(_04625_),
    .B1(_04624_));
 sg13g2_nor2_1 _10119_ (.A(net1485),
    .B(net255),
    .Y(_00256_));
 sg13g2_nand2b_1 _10120_ (.Y(_04626_),
    .B(_02783_),
    .A_N(\mac_inst.accumulator[9] ));
 sg13g2_nor2b_1 _10121_ (.A(_02783_),
    .B_N(\mac_inst.accumulator[9] ),
    .Y(_04627_));
 sg13g2_xnor2_1 _10122_ (.Y(_04628_),
    .A(net411),
    .B(_02783_));
 sg13g2_o21ai_1 _10123_ (.B1(_04628_),
    .Y(_04629_),
    .A1(_04615_),
    .A2(_04622_));
 sg13g2_nor3_1 _10124_ (.A(_04615_),
    .B(_04622_),
    .C(_04628_),
    .Y(_04630_));
 sg13g2_nor2_1 _10125_ (.A(_04803_),
    .B(_04630_),
    .Y(_04631_));
 sg13g2_a22oi_1 _10126_ (.Y(_04632_),
    .B1(_04629_),
    .B2(_04631_),
    .A2(net1114),
    .A1(net411));
 sg13g2_nor2_1 _10127_ (.A(net1485),
    .B(net412),
    .Y(_00257_));
 sg13g2_nand2_1 _10128_ (.Y(_04633_),
    .A(\mac_inst.accumulator[10] ),
    .B(_02904_));
 sg13g2_inv_1 _10129_ (.Y(_04634_),
    .A(_04633_));
 sg13g2_xor2_1 _10130_ (.B(_02904_),
    .A(net381),
    .X(_04635_));
 sg13g2_and2_1 _10131_ (.A(_04617_),
    .B(_04628_),
    .X(_04636_));
 sg13g2_o21ai_1 _10132_ (.B1(_04636_),
    .Y(_04637_),
    .A1(_04619_),
    .A2(_04620_));
 sg13g2_o21ai_1 _10133_ (.B1(_04626_),
    .Y(_04638_),
    .A1(_04615_),
    .A2(_04627_));
 sg13g2_nand2_1 _10134_ (.Y(_04639_),
    .A(_04637_),
    .B(_04638_));
 sg13g2_and2_1 _10135_ (.A(_04635_),
    .B(_04639_),
    .X(_04640_));
 sg13g2_o21ai_1 _10136_ (.B1(net1294),
    .Y(_04641_),
    .A1(_04635_),
    .A2(_04639_));
 sg13g2_nor2_1 _10137_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sg13g2_a21oi_1 _10138_ (.A1(net381),
    .A2(net1114),
    .Y(_04643_),
    .B1(_04642_));
 sg13g2_nor2_1 _10139_ (.A(net1485),
    .B(net382),
    .Y(_00258_));
 sg13g2_nand2_1 _10140_ (.Y(_04644_),
    .A(net204),
    .B(net1114));
 sg13g2_nand2_1 _10141_ (.Y(_04645_),
    .A(_04766_),
    .B(_03034_));
 sg13g2_or2_1 _10142_ (.X(_04646_),
    .B(_03034_),
    .A(_04766_));
 sg13g2_and2_1 _10143_ (.A(_04645_),
    .B(_04646_),
    .X(_04647_));
 sg13g2_o21ai_1 _10144_ (.B1(_04647_),
    .Y(_04648_),
    .A1(_04634_),
    .A2(_04640_));
 sg13g2_or3_1 _10145_ (.A(_04634_),
    .B(_04640_),
    .C(_04647_),
    .X(_04649_));
 sg13g2_nand3_1 _10146_ (.B(_04648_),
    .C(_04649_),
    .A(net1294),
    .Y(_04650_));
 sg13g2_a21oi_1 _10147_ (.A1(net205),
    .A2(_04650_),
    .Y(_00259_),
    .B1(net1485));
 sg13g2_nand2_1 _10148_ (.Y(_04651_),
    .A(net249),
    .B(net1116));
 sg13g2_a21o_1 _10149_ (.A2(_03034_),
    .A1(_04766_),
    .B1(_04633_),
    .X(_04652_));
 sg13g2_and3_1 _10150_ (.X(_04653_),
    .A(_04638_),
    .B(_04646_),
    .C(_04652_));
 sg13g2_o21ai_1 _10151_ (.B1(_04645_),
    .Y(_04654_),
    .A1(\mac_inst.accumulator[10] ),
    .A2(_02904_));
 sg13g2_a22oi_1 _10152_ (.Y(_04655_),
    .B1(_04654_),
    .B2(_04646_),
    .A2(_04653_),
    .A1(_04637_));
 sg13g2_and2_1 _10153_ (.A(\mac_inst.accumulator[12] ),
    .B(_03169_),
    .X(_04656_));
 sg13g2_inv_1 _10154_ (.Y(_04657_),
    .A(_04656_));
 sg13g2_xnor2_1 _10155_ (.Y(_04658_),
    .A(net249),
    .B(_03169_));
 sg13g2_inv_1 _10156_ (.Y(_04659_),
    .A(_04658_));
 sg13g2_a21oi_1 _10157_ (.A1(_04655_),
    .A2(_04659_),
    .Y(_04660_),
    .B1(_04803_));
 sg13g2_o21ai_1 _10158_ (.B1(_04660_),
    .Y(_04661_),
    .A1(_04655_),
    .A2(_04659_));
 sg13g2_a21oi_1 _10159_ (.A1(net250),
    .A2(_04661_),
    .Y(_00260_),
    .B1(net1483));
 sg13g2_nand2_1 _10160_ (.Y(_04662_),
    .A(net234),
    .B(net1113));
 sg13g2_nand2_1 _10161_ (.Y(_04663_),
    .A(\mac_inst.accumulator[13] ),
    .B(_03294_));
 sg13g2_xnor2_1 _10162_ (.Y(_04664_),
    .A(\mac_inst.accumulator[13] ),
    .B(_03294_));
 sg13g2_a21oi_1 _10163_ (.A1(_04655_),
    .A2(_04659_),
    .Y(_04665_),
    .B1(_04656_));
 sg13g2_a21oi_1 _10164_ (.A1(_04664_),
    .A2(_04665_),
    .Y(_04666_),
    .B1(_04803_));
 sg13g2_o21ai_1 _10165_ (.B1(_04666_),
    .Y(_04667_),
    .A1(_04664_),
    .A2(_04665_));
 sg13g2_a21oi_1 _10166_ (.A1(_04662_),
    .A2(_04667_),
    .Y(_00261_),
    .B1(net1483));
 sg13g2_nand2_1 _10167_ (.Y(_04668_),
    .A(net240),
    .B(net1113));
 sg13g2_nand2_1 _10168_ (.Y(_04669_),
    .A(net240),
    .B(_03424_));
 sg13g2_xnor2_1 _10169_ (.Y(_04670_),
    .A(net240),
    .B(_03424_));
 sg13g2_inv_1 _10170_ (.Y(_04671_),
    .A(_04670_));
 sg13g2_o21ai_1 _10171_ (.B1(_04663_),
    .Y(_04672_),
    .A1(_04664_),
    .A2(_04665_));
 sg13g2_nand2_1 _10172_ (.Y(_04673_),
    .A(_04671_),
    .B(_04672_));
 sg13g2_o21ai_1 _10173_ (.B1(net1293),
    .Y(_04674_),
    .A1(_04671_),
    .A2(_04672_));
 sg13g2_nand2b_1 _10174_ (.Y(_04675_),
    .B(_04673_),
    .A_N(_04674_));
 sg13g2_a21oi_1 _10175_ (.A1(_04668_),
    .A2(_04675_),
    .Y(_00262_),
    .B1(net1483));
 sg13g2_nand2_1 _10176_ (.Y(_04676_),
    .A(net301),
    .B(net1113));
 sg13g2_and2_1 _10177_ (.A(_04669_),
    .B(_04673_),
    .X(_04677_));
 sg13g2_nor2_1 _10178_ (.A(\mac_inst.accumulator[15] ),
    .B(_03560_),
    .Y(_04678_));
 sg13g2_nand2_1 _10179_ (.Y(_04679_),
    .A(\mac_inst.accumulator[15] ),
    .B(_03560_));
 sg13g2_xor2_1 _10180_ (.B(_03560_),
    .A(\mac_inst.accumulator[15] ),
    .X(_04680_));
 sg13g2_nand2b_1 _10181_ (.Y(_04681_),
    .B(_04680_),
    .A_N(_04677_));
 sg13g2_nand2b_1 _10182_ (.Y(_04682_),
    .B(_04677_),
    .A_N(_04680_));
 sg13g2_nand3_1 _10183_ (.B(_04681_),
    .C(_04682_),
    .A(net1293),
    .Y(_04683_));
 sg13g2_a21oi_1 _10184_ (.A1(_04676_),
    .A2(_04683_),
    .Y(_00263_),
    .B1(net1483));
 sg13g2_and2_1 _10185_ (.A(_04671_),
    .B(_04680_),
    .X(_04684_));
 sg13g2_nor2_1 _10186_ (.A(_04658_),
    .B(_04664_),
    .Y(_04685_));
 sg13g2_and3_1 _10187_ (.X(_04686_),
    .A(_04671_),
    .B(_04680_),
    .C(_04685_));
 sg13g2_o21ai_1 _10188_ (.B1(_04663_),
    .Y(_04687_),
    .A1(_04657_),
    .A2(_04664_));
 sg13g2_a21oi_1 _10189_ (.A1(_04669_),
    .A2(_04679_),
    .Y(_04688_),
    .B1(_04678_));
 sg13g2_a221oi_1 _10190_ (.B2(_04684_),
    .C1(_04688_),
    .B1(_04687_),
    .A1(_04655_),
    .Y(_04689_),
    .A2(_04686_));
 sg13g2_or2_1 _10191_ (.X(_04690_),
    .B(_03704_),
    .A(_04765_));
 sg13g2_xnor2_1 _10192_ (.Y(_04691_),
    .A(_04765_),
    .B(_03704_));
 sg13g2_nor2_1 _10193_ (.A(_04689_),
    .B(_04691_),
    .Y(_04692_));
 sg13g2_nand2_1 _10194_ (.Y(_04693_),
    .A(_04689_),
    .B(_04691_));
 sg13g2_nor2_1 _10195_ (.A(_04803_),
    .B(_04692_),
    .Y(_04694_));
 sg13g2_a22oi_1 _10196_ (.Y(_04695_),
    .B1(_04693_),
    .B2(_04694_),
    .A2(net1112),
    .A1(net293));
 sg13g2_nor2_1 _10197_ (.A(net1482),
    .B(net294),
    .Y(_00264_));
 sg13g2_nand2_1 _10198_ (.Y(_04696_),
    .A(\mac_inst.accumulator[17] ),
    .B(_03839_));
 sg13g2_inv_1 _10199_ (.Y(_04697_),
    .A(_04696_));
 sg13g2_xnor2_1 _10200_ (.Y(_04698_),
    .A(\mac_inst.accumulator[17] ),
    .B(_03839_));
 sg13g2_inv_1 _10201_ (.Y(_04699_),
    .A(_04698_));
 sg13g2_o21ai_1 _10202_ (.B1(_04690_),
    .Y(_04700_),
    .A1(_04689_),
    .A2(_04691_));
 sg13g2_and2_1 _10203_ (.A(_04699_),
    .B(_04700_),
    .X(_04701_));
 sg13g2_o21ai_1 _10204_ (.B1(net1293),
    .Y(_04702_),
    .A1(_04699_),
    .A2(_04700_));
 sg13g2_nor2_1 _10205_ (.A(_04701_),
    .B(_04702_),
    .Y(_04703_));
 sg13g2_a21oi_1 _10206_ (.A1(net284),
    .A2(net1112),
    .Y(_04704_),
    .B1(_04703_));
 sg13g2_nor2_1 _10207_ (.A(net1482),
    .B(_04704_),
    .Y(_00265_));
 sg13g2_nand2_1 _10208_ (.Y(_04705_),
    .A(net224),
    .B(net1112));
 sg13g2_nand2_1 _10209_ (.Y(_04706_),
    .A(\mac_inst.accumulator[18] ),
    .B(_03975_));
 sg13g2_xnor2_1 _10210_ (.Y(_04707_),
    .A(\mac_inst.accumulator[18] ),
    .B(_03975_));
 sg13g2_inv_1 _10211_ (.Y(_04708_),
    .A(_04707_));
 sg13g2_o21ai_1 _10212_ (.B1(_04708_),
    .Y(_04709_),
    .A1(_04697_),
    .A2(_04701_));
 sg13g2_or3_1 _10213_ (.A(_04697_),
    .B(_04701_),
    .C(_04708_),
    .X(_04710_));
 sg13g2_nand3_1 _10214_ (.B(_04709_),
    .C(_04710_),
    .A(net1293),
    .Y(_04711_));
 sg13g2_a21oi_1 _10215_ (.A1(_04705_),
    .A2(_04711_),
    .Y(_00266_),
    .B1(net1482));
 sg13g2_nand2_1 _10216_ (.Y(_04712_),
    .A(net216),
    .B(net1112));
 sg13g2_a21oi_1 _10217_ (.A1(_04101_),
    .A2(_04102_),
    .Y(_04713_),
    .B1(\mac_inst.accumulator[19] ));
 sg13g2_and3_1 _10218_ (.X(_04714_),
    .A(\mac_inst.accumulator[19] ),
    .B(_04101_),
    .C(_04102_));
 sg13g2_nand3_1 _10219_ (.B(_04101_),
    .C(_04102_),
    .A(\mac_inst.accumulator[19] ),
    .Y(_04715_));
 sg13g2_nand2b_1 _10220_ (.Y(_04716_),
    .B(_04715_),
    .A_N(_04713_));
 sg13g2_a21o_1 _10221_ (.A2(_04709_),
    .A1(_04706_),
    .B1(_04716_),
    .X(_04717_));
 sg13g2_nand3_1 _10222_ (.B(_04709_),
    .C(_04716_),
    .A(_04706_),
    .Y(_04718_));
 sg13g2_nand3_1 _10223_ (.B(_04717_),
    .C(_04718_),
    .A(net1293),
    .Y(_04719_));
 sg13g2_a21oi_1 _10224_ (.A1(_04712_),
    .A2(_04719_),
    .Y(_00267_),
    .B1(net1482));
 sg13g2_nand2_1 _10225_ (.Y(_04720_),
    .A(net197),
    .B(net1112));
 sg13g2_nor3_1 _10226_ (.A(_04707_),
    .B(_04713_),
    .C(_04714_),
    .Y(_04721_));
 sg13g2_nand3b_1 _10227_ (.B(_04699_),
    .C(_04721_),
    .Y(_04722_),
    .A_N(_04691_));
 sg13g2_nor2_1 _10228_ (.A(_04689_),
    .B(_04722_),
    .Y(_04723_));
 sg13g2_o21ai_1 _10229_ (.B1(_04696_),
    .Y(_04724_),
    .A1(_04690_),
    .A2(_04698_));
 sg13g2_o21ai_1 _10230_ (.B1(_04715_),
    .Y(_04725_),
    .A1(_04706_),
    .A2(_04713_));
 sg13g2_a21oi_1 _10231_ (.A1(_04721_),
    .A2(_04724_),
    .Y(_04726_),
    .B1(_04725_));
 sg13g2_nor2b_1 _10232_ (.A(_04723_),
    .B_N(_04726_),
    .Y(_04727_));
 sg13g2_o21ai_1 _10233_ (.B1(_04726_),
    .Y(_04728_),
    .A1(_04689_),
    .A2(_04722_));
 sg13g2_or2_1 _10234_ (.X(_04729_),
    .B(_04227_),
    .A(_04764_));
 sg13g2_xnor2_1 _10235_ (.Y(_04730_),
    .A(_04764_),
    .B(_04227_));
 sg13g2_o21ai_1 _10236_ (.B1(net1293),
    .Y(_04731_),
    .A1(_04727_),
    .A2(_04730_));
 sg13g2_a21o_1 _10237_ (.A2(_04730_),
    .A1(_04727_),
    .B1(_04731_),
    .X(_04732_));
 sg13g2_a21oi_1 _10238_ (.A1(_04720_),
    .A2(_04732_),
    .Y(_00268_),
    .B1(net1478));
 sg13g2_nand2_1 _10239_ (.Y(_04733_),
    .A(net236),
    .B(net1112));
 sg13g2_a21oi_1 _10240_ (.A1(_04350_),
    .A2(_04351_),
    .Y(_04734_),
    .B1(net236));
 sg13g2_and3_1 _10241_ (.X(_04735_),
    .A(\mac_inst.accumulator[21] ),
    .B(_04350_),
    .C(_04351_));
 sg13g2_nand3_1 _10242_ (.B(_04350_),
    .C(_04351_),
    .A(\mac_inst.accumulator[21] ),
    .Y(_04736_));
 sg13g2_nor2_1 _10243_ (.A(_04734_),
    .B(_04735_),
    .Y(_04737_));
 sg13g2_o21ai_1 _10244_ (.B1(_04729_),
    .Y(_04738_),
    .A1(_04727_),
    .A2(_04730_));
 sg13g2_a21oi_1 _10245_ (.A1(_04737_),
    .A2(_04738_),
    .Y(_04739_),
    .B1(_04803_));
 sg13g2_o21ai_1 _10246_ (.B1(_04739_),
    .Y(_04740_),
    .A1(_04737_),
    .A2(_04738_));
 sg13g2_a21oi_1 _10247_ (.A1(_04733_),
    .A2(_04740_),
    .Y(_00269_),
    .B1(net1478));
 sg13g2_nor3_1 _10248_ (.A(_04730_),
    .B(_04734_),
    .C(_04735_),
    .Y(_04741_));
 sg13g2_o21ai_1 _10249_ (.B1(_04736_),
    .Y(_04742_),
    .A1(_04729_),
    .A2(_04734_));
 sg13g2_a21oi_1 _10250_ (.A1(_04728_),
    .A2(_04741_),
    .Y(_04743_),
    .B1(_04742_));
 sg13g2_or2_1 _10251_ (.X(_04744_),
    .B(_04475_),
    .A(_04763_));
 sg13g2_xnor2_1 _10252_ (.Y(_04745_),
    .A(_04763_),
    .B(_04475_));
 sg13g2_o21ai_1 _10253_ (.B1(net1293),
    .Y(_04746_),
    .A1(_04743_),
    .A2(_04745_));
 sg13g2_a21oi_1 _10254_ (.A1(_04743_),
    .A2(_04745_),
    .Y(_04747_),
    .B1(_04746_));
 sg13g2_a21oi_1 _10255_ (.A1(net263),
    .A2(net1112),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_nor2_1 _10256_ (.A(net1478),
    .B(net264),
    .Y(_00270_));
 sg13g2_nand2_1 _10257_ (.Y(_04749_),
    .A(net242),
    .B(net1112));
 sg13g2_o21ai_1 _10258_ (.B1(_04744_),
    .Y(_04750_),
    .A1(_04743_),
    .A2(_04745_));
 sg13g2_xor2_1 _10259_ (.B(_04560_),
    .A(net242),
    .X(_04751_));
 sg13g2_o21ai_1 _10260_ (.B1(net1293),
    .Y(_04752_),
    .A1(_04750_),
    .A2(_04751_));
 sg13g2_a21o_1 _10261_ (.A2(_04751_),
    .A1(_04750_),
    .B1(_04752_),
    .X(_04753_));
 sg13g2_a21oi_1 _10262_ (.A1(_04749_),
    .A2(_04753_),
    .Y(_00271_),
    .B1(net1478));
 sg13g2_o21ai_1 _10263_ (.B1(net1516),
    .Y(_04754_),
    .A1(\mac_inst.RDY_get_multiply ),
    .A2(net1299));
 sg13g2_nor2_1 _10264_ (.A(net177),
    .B(_04754_),
    .Y(_00272_));
 sg13g2_o21ai_1 _10265_ (.B1(net1516),
    .Y(_04755_),
    .A1(\mac_inst.RDY_get_mac ),
    .A2(net1295));
 sg13g2_nor2_1 _10266_ (.A(net175),
    .B(_04755_),
    .Y(_00273_));
 sg13g2_nor2b_2 _10267_ (.A(_04865_),
    .B_N(net1104),
    .Y(_04756_));
 sg13g2_nand2_1 _10268_ (.Y(_04757_),
    .A(net1),
    .B(net1064));
 sg13g2_o21ai_1 _10269_ (.B1(_04757_),
    .Y(_00274_),
    .A1(_04830_),
    .A2(net1064));
 sg13g2_nand2_1 _10270_ (.Y(_04758_),
    .A(net2),
    .B(net1064));
 sg13g2_o21ai_1 _10271_ (.B1(_04758_),
    .Y(_00275_),
    .A1(_04831_),
    .A2(net1065));
 sg13g2_nand2_1 _10272_ (.Y(_04759_),
    .A(net3),
    .B(net1064));
 sg13g2_o21ai_1 _10273_ (.B1(_04759_),
    .Y(_00276_),
    .A1(_04832_),
    .A2(net1065));
 sg13g2_mux2_1 _10274_ (.A0(net1168),
    .A1(net4),
    .S(net1065),
    .X(_00277_));
 sg13g2_nand2_1 _10275_ (.Y(_04760_),
    .A(net5),
    .B(net1064));
 sg13g2_o21ai_1 _10276_ (.B1(_04760_),
    .Y(_00278_),
    .A1(_04833_),
    .A2(net1064));
 sg13g2_mux2_1 _10277_ (.A0(net1158),
    .A1(net6),
    .S(net1065),
    .X(_00279_));
 sg13g2_nand2_1 _10278_ (.Y(_04761_),
    .A(net7),
    .B(net1064));
 sg13g2_o21ai_1 _10279_ (.B1(_04761_),
    .Y(_00280_),
    .A1(_04834_),
    .A2(net1064));
 sg13g2_mux2_1 _10280_ (.A0(net1146),
    .A1(net8),
    .S(net1065),
    .X(_00281_));
 sg13g2_dfrbpq_1 _10281_ (.RESET_B(net33),
    .D(_00025_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _10282_ (.RESET_B(net1502),
    .D(net453),
    .Q(\byte_counter[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _10283_ (.RESET_B(net1502),
    .D(net451),
    .Q(\byte_counter[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _10284_ (.RESET_B(net1502),
    .D(net202),
    .Q(\byte_counter[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _10285_ (.RESET_B(net1500),
    .D(_00029_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _10286_ (.RESET_B(net1521),
    .D(_00030_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _10287_ (.RESET_B(net1499),
    .D(_00031_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _10288_ (.RESET_B(net1507),
    .D(_00032_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10289_ (.RESET_B(net1499),
    .D(_00033_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _10290_ (.RESET_B(net1521),
    .D(_00034_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10291_ (.RESET_B(net1499),
    .D(_00035_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _10292_ (.RESET_B(net1508),
    .D(_00036_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10293_ (.RESET_B(net34),
    .D(_00018_),
    .Q(\cordic_inst.current_op[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10294_ (.RESET_B(net36),
    .D(_00019_),
    .Q(\cordic_inst.current_op[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10295_ (.RESET_B(net41),
    .D(_00020_),
    .Q(\cordic_inst.current_op[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _10296_ (.RESET_B(net1497),
    .D(_00037_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _10297_ (.RESET_B(net1508),
    .D(_00038_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10298_ (.RESET_B(net1497),
    .D(_00039_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _10299_ (.RESET_B(net1506),
    .D(_00040_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _10300_ (.RESET_B(net1497),
    .D(_00041_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _10301_ (.RESET_B(net1508),
    .D(_00042_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10302_ (.RESET_B(net1497),
    .D(_00043_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _10303_ (.RESET_B(net1506),
    .D(_00044_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _10304_ (.RESET_B(net37),
    .D(_00001_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _10305_ (.RESET_B(net38),
    .D(_00002_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _10306_ (.RESET_B(net39),
    .D(_00003_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _10307_ (.RESET_B(net40),
    .D(_00004_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _10308_ (.RESET_B(net122),
    .D(_00005_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _10309_ (.RESET_B(net35),
    .D(_00000_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _10310_ (.RESET_B(net32),
    .D(_00045_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _10311_ (.RESET_B(net31),
    .D(_00046_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10312_ (.RESET_B(net30),
    .D(_00047_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _10313_ (.RESET_B(net29),
    .D(_00048_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _10314_ (.RESET_B(net28),
    .D(_00049_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _10315_ (.RESET_B(net27),
    .D(_00050_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _10316_ (.RESET_B(net1517),
    .D(_00051_),
    .Q(\result_reg[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _10317_ (.RESET_B(net1501),
    .D(net244),
    .Q(\result_reg[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _10318_ (.RESET_B(net1517),
    .D(net408),
    .Q(\result_reg[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _10319_ (.RESET_B(net1516),
    .D(net371),
    .Q(\result_reg[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10320_ (.RESET_B(net1501),
    .D(_00055_),
    .Q(\result_reg[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _10321_ (.RESET_B(net1517),
    .D(net446),
    .Q(\result_reg[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _10322_ (.RESET_B(net1516),
    .D(net392),
    .Q(\result_reg[6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _10323_ (.RESET_B(net1518),
    .D(_00058_),
    .Q(\result_reg[7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _10324_ (.RESET_B(net1503),
    .D(net259),
    .Q(\result_reg[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _10325_ (.RESET_B(net1517),
    .D(_00060_),
    .Q(\result_reg[9] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _10326_ (.RESET_B(net1517),
    .D(_00061_),
    .Q(\result_reg[10] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _10327_ (.RESET_B(net1503),
    .D(net229),
    .Q(\result_reg[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _10328_ (.RESET_B(net1510),
    .D(net346),
    .Q(\result_reg[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10329_ (.RESET_B(net1510),
    .D(net215),
    .Q(\result_reg[13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10330_ (.RESET_B(net1514),
    .D(net309),
    .Q(\result_reg[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _10331_ (.RESET_B(net1501),
    .D(net213),
    .Q(\result_reg[15] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _10332_ (.RESET_B(net1502),
    .D(net192),
    .Q(\result_reg[16] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _10333_ (.RESET_B(net1503),
    .D(net248),
    .Q(\result_reg[17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10334_ (.RESET_B(net1501),
    .D(net210),
    .Q(\result_reg[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _10335_ (.RESET_B(net1512),
    .D(net208),
    .Q(\result_reg[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10336_ (.RESET_B(net1504),
    .D(net199),
    .Q(\result_reg[20] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10337_ (.RESET_B(net1510),
    .D(net231),
    .Q(\result_reg[21] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10338_ (.RESET_B(net1501),
    .D(net307),
    .Q(\result_reg[22] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _10339_ (.RESET_B(net1510),
    .D(net375),
    .Q(\result_reg[23] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _10340_ (.RESET_B(net1501),
    .D(_00075_),
    .Q(uo_out[0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _10341_ (.RESET_B(net1501),
    .D(_00076_),
    .Q(uo_out[1]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10342_ (.RESET_B(net1494),
    .D(_00077_),
    .Q(uo_out[2]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10343_ (.RESET_B(net1494),
    .D(_00078_),
    .Q(uo_out[3]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10344_ (.RESET_B(net1495),
    .D(_00079_),
    .Q(uo_out[4]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10345_ (.RESET_B(net1495),
    .D(_00080_),
    .Q(uo_out[5]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _10346_ (.RESET_B(net1494),
    .D(_00081_),
    .Q(uo_out[6]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10347_ (.RESET_B(net1495),
    .D(net443),
    .Q(uo_out[7]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _10348_ (.RESET_B(net1503),
    .D(_00083_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _10349_ (.RESET_B(net1503),
    .D(_00084_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _10350_ (.RESET_B(net1503),
    .D(_00085_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _10351_ (.RESET_B(net1511),
    .D(_00086_),
    .Q(\cmd_reg[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _10352_ (.RESET_B(net1512),
    .D(_00087_),
    .Q(\cmd_reg[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10353_ (.RESET_B(net1511),
    .D(_00088_),
    .Q(\cmd_reg[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10354_ (.RESET_B(net1512),
    .D(_00089_),
    .Q(\cmd_reg[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10355_ (.RESET_B(net1514),
    .D(_00090_),
    .Q(\cmd_reg[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10356_ (.RESET_B(net1515),
    .D(_00091_),
    .Q(\cmd_reg[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10357_ (.RESET_B(net1514),
    .D(_00092_),
    .Q(\cmd_reg[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10358_ (.RESET_B(net1515),
    .D(_00093_),
    .Q(\cmd_reg[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10359_ (.RESET_B(net1506),
    .D(_00094_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _10360_ (.RESET_B(net1521),
    .D(_00095_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _10361_ (.RESET_B(net1506),
    .D(_00096_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _10362_ (.RESET_B(net1521),
    .D(_00097_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10363_ (.RESET_B(net1508),
    .D(_00098_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _10364_ (.RESET_B(net1520),
    .D(_00099_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _10365_ (.RESET_B(net1508),
    .D(_00100_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _10366_ (.RESET_B(net1513),
    .D(_00101_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _10367_ (.RESET_B(net1489),
    .D(_00102_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _10368_ (.RESET_B(net1500),
    .D(_00103_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _10369_ (.RESET_B(net1497),
    .D(_00104_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _10370_ (.RESET_B(net1497),
    .D(_00105_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _10371_ (.RESET_B(net1490),
    .D(_00106_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _10372_ (.RESET_B(net1498),
    .D(_00107_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _10373_ (.RESET_B(net1489),
    .D(_00108_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _10374_ (.RESET_B(net1500),
    .D(_00109_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _10375_ (.RESET_B(net1502),
    .D(net219),
    .Q(\result_reg[24] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10376_ (.RESET_B(net1501),
    .D(net223),
    .Q(\result_reg[25] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _10377_ (.RESET_B(net1495),
    .D(net180),
    .Q(\result_reg[26] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10378_ (.RESET_B(net1494),
    .D(net227),
    .Q(\result_reg[27] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10379_ (.RESET_B(net1494),
    .D(net233),
    .Q(\result_reg[28] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _10380_ (.RESET_B(net1494),
    .D(net246),
    .Q(\result_reg[29] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10381_ (.RESET_B(net1494),
    .D(net239),
    .Q(\result_reg[30] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _10382_ (.RESET_B(net1491),
    .D(net335),
    .Q(\result_reg[31] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _10383_ (.RESET_B(net1491),
    .D(net344),
    .Q(\result_reg[32] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _10384_ (.RESET_B(net1491),
    .D(net275),
    .Q(\result_reg[33] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _10385_ (.RESET_B(net1491),
    .D(net337),
    .Q(\result_reg[34] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _10386_ (.RESET_B(net1492),
    .D(net324),
    .Q(\result_reg[35] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _10387_ (.RESET_B(net1491),
    .D(net384),
    .Q(\result_reg[36] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _10388_ (.RESET_B(net1492),
    .D(net318),
    .Q(\result_reg[37] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _10389_ (.RESET_B(net1491),
    .D(net339),
    .Q(\result_reg[38] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _10390_ (.RESET_B(net1492),
    .D(net292),
    .Q(\result_reg[39] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _10391_ (.RESET_B(net1491),
    .D(net360),
    .Q(\result_reg[40] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _10392_ (.RESET_B(net1491),
    .D(net358),
    .Q(\result_reg[41] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10393_ (.RESET_B(net1492),
    .D(net296),
    .Q(\result_reg[42] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10394_ (.RESET_B(net1492),
    .D(net314),
    .Q(\result_reg[43] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10395_ (.RESET_B(net1493),
    .D(net270),
    .Q(\result_reg[44] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _10396_ (.RESET_B(net1492),
    .D(net356),
    .Q(\result_reg[45] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10397_ (.RESET_B(net1492),
    .D(net266),
    .Q(\result_reg[46] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10398_ (.RESET_B(net1494),
    .D(net253),
    .Q(\result_reg[47] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _10399_ (.RESET_B(net1503),
    .D(net9),
    .Q(wr_prev),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _10400_ (.RESET_B(net1502),
    .D(net10),
    .Q(rd_prev),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _10401_ (.RESET_B(net1514),
    .D(_00011_),
    .Q(cordic_en_sin_cos),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _10402_ (.RESET_B(net1511),
    .D(_00007_),
    .Q(cordic_en_atan2),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10403_ (.RESET_B(net1504),
    .D(_00012_),
    .Q(cordic_en_sqrt),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _10404_ (.RESET_B(net1511),
    .D(_00009_),
    .Q(cordic_en_get_sin_cos),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10405_ (.RESET_B(net1511),
    .D(_00008_),
    .Q(cordic_en_get_atan2),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10406_ (.RESET_B(net1511),
    .D(_00010_),
    .Q(cordic_en_get_sqrt),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10407_ (.RESET_B(net1514),
    .D(_00017_),
    .Q(mac_en_multiply),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _10408_ (.RESET_B(net1515),
    .D(_00015_),
    .Q(mac_en_get_multiply),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10409_ (.RESET_B(net1514),
    .D(net331),
    .Q(mac_en_mac),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _10410_ (.RESET_B(net1514),
    .D(net379),
    .Q(mac_en_get_mac),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _10411_ (.RESET_B(net1514),
    .D(_00013_),
    .Q(mac_en_clear),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _10412_ (.RESET_B(net174),
    .D(net441),
    .Q(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _10413_ (.RESET_B(net172),
    .D(_00135_),
    .Q(cordic_busy),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10414_ (.RESET_B(net170),
    .D(_00136_),
    .Q(\cordic_inst.cordic_state[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _10415_ (.RESET_B(net168),
    .D(_00137_),
    .Q(\cordic_inst.cordic_state[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _10416_ (.RESET_B(net166),
    .D(_00138_),
    .Q(\cordic_inst.cordic_state[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _10417_ (.RESET_B(net164),
    .D(_00139_),
    .Q(\cordic_inst.cordic_state[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _10418_ (.RESET_B(net163),
    .D(_00140_),
    .Q(\cordic_inst.cordic_state[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _10419_ (.RESET_B(net161),
    .D(_00141_),
    .Q(\cordic_inst.cordic_state[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _10420_ (.RESET_B(net159),
    .D(_00142_),
    .Q(\cordic_atan2_result[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _10421_ (.RESET_B(net157),
    .D(_00143_),
    .Q(\cordic_atan2_result[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _10422_ (.RESET_B(net155),
    .D(_00144_),
    .Q(\cordic_atan2_result[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10423_ (.RESET_B(net153),
    .D(_00145_),
    .Q(\cordic_atan2_result[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10424_ (.RESET_B(net151),
    .D(_00146_),
    .Q(\cordic_atan2_result[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10425_ (.RESET_B(net149),
    .D(_00147_),
    .Q(\cordic_atan2_result[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _10426_ (.RESET_B(net148),
    .D(_00148_),
    .Q(\cordic_atan2_result[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _10427_ (.RESET_B(net147),
    .D(_00149_),
    .Q(\cordic_atan2_result[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10428_ (.RESET_B(net145),
    .D(_00150_),
    .Q(\cordic_atan2_result[8] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10429_ (.RESET_B(net144),
    .D(_00151_),
    .Q(\cordic_atan2_result[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10430_ (.RESET_B(net143),
    .D(_00152_),
    .Q(\cordic_atan2_result[10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _10431_ (.RESET_B(net142),
    .D(_00153_),
    .Q(\cordic_atan2_result[11] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _10432_ (.RESET_B(net141),
    .D(_00154_),
    .Q(\cordic_atan2_result[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10433_ (.RESET_B(net140),
    .D(net402),
    .Q(\cordic_atan2_result[13] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _10434_ (.RESET_B(net139),
    .D(_00156_),
    .Q(\cordic_atan2_result[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _10435_ (.RESET_B(net138),
    .D(_00157_),
    .Q(\cordic_atan2_result[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10436_ (.RESET_B(net137),
    .D(_00158_),
    .Q(\cordic_atan2_result[16] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _10437_ (.RESET_B(net135),
    .D(_00159_),
    .Q(\cordic_atan2_result[17] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _10438_ (.RESET_B(net133),
    .D(_00160_),
    .Q(\cordic_atan2_result[18] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _10439_ (.RESET_B(net131),
    .D(_00161_),
    .Q(\cordic_atan2_result[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10440_ (.RESET_B(net129),
    .D(_00162_),
    .Q(\cordic_atan2_result[20] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10441_ (.RESET_B(net127),
    .D(_00163_),
    .Q(\cordic_atan2_result[21] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10442_ (.RESET_B(net126),
    .D(_00164_),
    .Q(\cordic_atan2_result[22] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _10443_ (.RESET_B(net124),
    .D(net459),
    .Q(\cordic_atan2_result[23] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10444_ (.RESET_B(net121),
    .D(_00166_),
    .Q(\cordic_inst.cordic_state[32] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _10445_ (.RESET_B(net119),
    .D(_00167_),
    .Q(\cordic_inst.cordic_state[33] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _10446_ (.RESET_B(net117),
    .D(_00168_),
    .Q(\cordic_inst.cordic_state[34] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _10447_ (.RESET_B(net115),
    .D(_00169_),
    .Q(\cordic_inst.cordic_state[35] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _10448_ (.RESET_B(net113),
    .D(_00170_),
    .Q(\cordic_inst.cordic_state[36] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _10449_ (.RESET_B(net111),
    .D(net475),
    .Q(\cordic_inst.cordic_state[37] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _10450_ (.RESET_B(net110),
    .D(net468),
    .Q(\cordic_inst.cordic_state[38] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _10451_ (.RESET_B(net108),
    .D(_00173_),
    .Q(\cordic_inst.cordic_state[39] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _10452_ (.RESET_B(net106),
    .D(_00174_),
    .Q(\cordic_inst.cordic_state[40] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _10453_ (.RESET_B(net104),
    .D(_00175_),
    .Q(\cordic_inst.cordic_state[41] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _10454_ (.RESET_B(net102),
    .D(_00176_),
    .Q(\cordic_inst.cordic_state[42] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _10455_ (.RESET_B(net100),
    .D(_00177_),
    .Q(\cordic_inst.cordic_state[43] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _10456_ (.RESET_B(net98),
    .D(_00178_),
    .Q(\cordic_inst.cordic_state[44] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _10457_ (.RESET_B(net96),
    .D(_00179_),
    .Q(\cordic_inst.cordic_state[45] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _10458_ (.RESET_B(net95),
    .D(_00180_),
    .Q(\cordic_inst.cordic_state[46] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _10459_ (.RESET_B(net93),
    .D(_00181_),
    .Q(\cordic_inst.cordic_state[47] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _10460_ (.RESET_B(net91),
    .D(_00182_),
    .Q(\cordic_inst.cordic_state[48] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _10461_ (.RESET_B(net89),
    .D(_00183_),
    .Q(\cordic_inst.cordic_state[49] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _10462_ (.RESET_B(net87),
    .D(_00184_),
    .Q(\cordic_inst.cordic_state[50] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _10463_ (.RESET_B(net85),
    .D(_00185_),
    .Q(\cordic_inst.cordic_state[51] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _10464_ (.RESET_B(net83),
    .D(_00186_),
    .Q(\cordic_inst.cordic_state[52] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _10465_ (.RESET_B(net81),
    .D(net489),
    .Q(\cordic_inst.cordic_state[53] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _10466_ (.RESET_B(net80),
    .D(_00188_),
    .Q(\cordic_inst.cordic_state[54] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _10467_ (.RESET_B(net78),
    .D(_00189_),
    .Q(\cordic_inst.cordic_state[55] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _10468_ (.RESET_B(net76),
    .D(net416),
    .Q(\cordic_inst.cordic_state[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10469_ (.RESET_B(net74),
    .D(net484),
    .Q(\cordic_inst.cordic_state[57] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _10470_ (.RESET_B(net72),
    .D(_00192_),
    .Q(\cordic_inst.cordic_state[58] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _10471_ (.RESET_B(net70),
    .D(net486),
    .Q(\cordic_inst.cordic_state[59] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10472_ (.RESET_B(net68),
    .D(_00194_),
    .Q(\cordic_inst.cordic_state[60] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10473_ (.RESET_B(net66),
    .D(net491),
    .Q(\cordic_inst.cordic_state[61] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10474_ (.RESET_B(net65),
    .D(net461),
    .Q(\cordic_inst.cordic_state[62] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10475_ (.RESET_B(net63),
    .D(_00197_),
    .Q(\cordic_inst.cordic_state[63] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10476_ (.RESET_B(net61),
    .D(_00198_),
    .Q(\cordic_inst.cordic_state[64] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10477_ (.RESET_B(net59),
    .D(_00199_),
    .Q(\cordic_inst.cordic_state[65] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _10478_ (.RESET_B(net57),
    .D(_00200_),
    .Q(\cordic_inst.cordic_state[66] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _10479_ (.RESET_B(net55),
    .D(_00201_),
    .Q(\cordic_inst.cordic_state[67] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _10480_ (.RESET_B(net53),
    .D(_00202_),
    .Q(\cordic_inst.cordic_state[68] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10481_ (.RESET_B(net51),
    .D(_00203_),
    .Q(\cordic_inst.cordic_state[69] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _10482_ (.RESET_B(net50),
    .D(_00204_),
    .Q(\cordic_inst.cordic_state[70] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _10483_ (.RESET_B(net48),
    .D(_00205_),
    .Q(\cordic_inst.cordic_state[71] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _10484_ (.RESET_B(net46),
    .D(_00206_),
    .Q(\cordic_inst.cordic_state[72] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _10485_ (.RESET_B(net44),
    .D(_00207_),
    .Q(\cordic_inst.cordic_state[73] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _10486_ (.RESET_B(net43),
    .D(_00208_),
    .Q(\cordic_inst.cordic_state[74] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _10487_ (.RESET_B(net173),
    .D(_00209_),
    .Q(\cordic_inst.cordic_state[75] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _10488_ (.RESET_B(net169),
    .D(_00210_),
    .Q(\cordic_inst.cordic_state[76] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _10489_ (.RESET_B(net165),
    .D(_00211_),
    .Q(\cordic_inst.cordic_state[77] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _10490_ (.RESET_B(net162),
    .D(_00212_),
    .Q(\cordic_inst.cordic_state[78] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _10491_ (.RESET_B(net158),
    .D(_00213_),
    .Q(\cordic_inst.cordic_state[79] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _10492_ (.RESET_B(net154),
    .D(_00214_),
    .Q(\cordic_inst.operation_pending ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _10493_ (.RESET_B(net150),
    .D(_00215_),
    .Q(\cordic_inst.result_ready ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _10494_ (.RESET_B(net1503),
    .D(_00024_),
    .Q(_00023_),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _10495_ (.RESET_B(net1511),
    .D(net354),
    .Q(\exec_phase[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _10496_ (.RESET_B(net1511),
    .D(_00022_),
    .Q(\exec_phase[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _10497_ (.RESET_B(net1498),
    .D(_00216_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10498_ (.RESET_B(net1498),
    .D(_00217_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10499_ (.RESET_B(net1506),
    .D(_00218_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _10500_ (.RESET_B(net1506),
    .D(_00219_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10501_ (.RESET_B(net1498),
    .D(_00220_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _10502_ (.RESET_B(net1510),
    .D(_00221_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _10503_ (.RESET_B(net1506),
    .D(_00222_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _10504_ (.RESET_B(net1510),
    .D(_00223_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10505_ (.RESET_B(net136),
    .D(_00224_),
    .Q(\mac_inst.get_multiply[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _10506_ (.RESET_B(net132),
    .D(_00225_),
    .Q(\mac_inst.get_multiply[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _10507_ (.RESET_B(net128),
    .D(_00226_),
    .Q(\mac_inst.get_multiply[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _10508_ (.RESET_B(net125),
    .D(_00227_),
    .Q(\mac_inst.get_multiply[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _10509_ (.RESET_B(net120),
    .D(_00228_),
    .Q(\mac_inst.get_multiply[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _10510_ (.RESET_B(net116),
    .D(_00229_),
    .Q(\mac_inst.get_multiply[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _10511_ (.RESET_B(net112),
    .D(_00230_),
    .Q(\mac_inst.get_multiply[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _10512_ (.RESET_B(net109),
    .D(net298),
    .Q(\mac_inst.get_multiply[7] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _10513_ (.RESET_B(net105),
    .D(net305),
    .Q(\mac_inst.get_multiply[8] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _10514_ (.RESET_B(net101),
    .D(net257),
    .Q(\mac_inst.get_multiply[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _10515_ (.RESET_B(net97),
    .D(_00234_),
    .Q(\mac_inst.get_multiply[10] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10516_ (.RESET_B(net94),
    .D(net369),
    .Q(\mac_inst.get_multiply[11] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _10517_ (.RESET_B(net90),
    .D(_00236_),
    .Q(\mac_inst.get_multiply[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10518_ (.RESET_B(net86),
    .D(_00237_),
    .Q(\mac_inst.get_multiply[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10519_ (.RESET_B(net82),
    .D(_00238_),
    .Q(\mac_inst.get_multiply[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _10520_ (.RESET_B(net79),
    .D(_00239_),
    .Q(\mac_inst.get_multiply[15] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _10521_ (.RESET_B(net75),
    .D(net290),
    .Q(\mac_inst.get_multiply[16] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _10522_ (.RESET_B(net71),
    .D(_00241_),
    .Q(\mac_inst.get_multiply[17] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _10523_ (.RESET_B(net67),
    .D(_00242_),
    .Q(\mac_inst.get_multiply[18] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _10524_ (.RESET_B(net64),
    .D(net287),
    .Q(\mac_inst.get_multiply[19] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _10525_ (.RESET_B(net60),
    .D(net273),
    .Q(\mac_inst.get_multiply[20] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _10526_ (.RESET_B(net56),
    .D(net278),
    .Q(\mac_inst.get_multiply[21] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _10527_ (.RESET_B(net52),
    .D(net262),
    .Q(\mac_inst.get_multiply[22] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _10528_ (.RESET_B(net49),
    .D(_00247_),
    .Q(\mac_inst.get_multiply[23] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _10529_ (.RESET_B(net45),
    .D(_00248_),
    .Q(\mac_inst.accumulator[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _10530_ (.RESET_B(net42),
    .D(_00249_),
    .Q(\mac_inst.accumulator[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _10531_ (.RESET_B(net167),
    .D(_00250_),
    .Q(\mac_inst.accumulator[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10532_ (.RESET_B(net160),
    .D(_00251_),
    .Q(\mac_inst.accumulator[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10533_ (.RESET_B(net152),
    .D(_00252_),
    .Q(\mac_inst.accumulator[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _10534_ (.RESET_B(net146),
    .D(_00253_),
    .Q(\mac_inst.accumulator[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _10535_ (.RESET_B(net130),
    .D(_00254_),
    .Q(\mac_inst.accumulator[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _10536_ (.RESET_B(net123),
    .D(_00255_),
    .Q(\mac_inst.accumulator[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10537_ (.RESET_B(net114),
    .D(_00256_),
    .Q(\mac_inst.accumulator[8] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10538_ (.RESET_B(net107),
    .D(_00257_),
    .Q(\mac_inst.accumulator[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _10539_ (.RESET_B(net99),
    .D(_00258_),
    .Q(\mac_inst.accumulator[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _10540_ (.RESET_B(net92),
    .D(net206),
    .Q(\mac_inst.accumulator[11] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _10541_ (.RESET_B(net84),
    .D(net251),
    .Q(\mac_inst.accumulator[12] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _10542_ (.RESET_B(net77),
    .D(net235),
    .Q(\mac_inst.accumulator[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _10543_ (.RESET_B(net69),
    .D(net241),
    .Q(\mac_inst.accumulator[14] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _10544_ (.RESET_B(net62),
    .D(net302),
    .Q(\mac_inst.accumulator[15] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _10545_ (.RESET_B(net54),
    .D(_00264_),
    .Q(\mac_inst.accumulator[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _10546_ (.RESET_B(net47),
    .D(_00265_),
    .Q(\mac_inst.accumulator[17] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _10547_ (.RESET_B(net171),
    .D(net225),
    .Q(\mac_inst.accumulator[18] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _10548_ (.RESET_B(net156),
    .D(net217),
    .Q(\mac_inst.accumulator[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _10549_ (.RESET_B(net134),
    .D(_00268_),
    .Q(\mac_inst.accumulator[20] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _10550_ (.RESET_B(net118),
    .D(net237),
    .Q(\mac_inst.accumulator[21] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _10551_ (.RESET_B(net103),
    .D(_00270_),
    .Q(\mac_inst.accumulator[22] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _10552_ (.RESET_B(net88),
    .D(_00271_),
    .Q(\mac_inst.accumulator[23] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _10553_ (.RESET_B(net73),
    .D(net178),
    .Q(\mac_inst.RDY_get_multiply ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _10554_ (.RESET_B(net58),
    .D(net176),
    .Q(\mac_inst.RDY_get_mac ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _10555_ (.RESET_B(net1490),
    .D(_00274_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _10556_ (.RESET_B(net1500),
    .D(_00275_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _10557_ (.RESET_B(net1499),
    .D(_00276_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _10558_ (.RESET_B(net1497),
    .D(_00277_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _10559_ (.RESET_B(net1489),
    .D(_00278_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _10560_ (.RESET_B(net1497),
    .D(_00279_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _10561_ (.RESET_B(net1489),
    .D(_00280_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _10562_ (.RESET_B(net1500),
    .D(_00281_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_tiehi _10314__28 (.L_HI(net28));
 sg13g2_tiehi _10313__29 (.L_HI(net29));
 sg13g2_tiehi _10312__30 (.L_HI(net30));
 sg13g2_tiehi _10311__31 (.L_HI(net31));
 sg13g2_tiehi _10310__32 (.L_HI(net32));
 sg13g2_tiehi _10281__33 (.L_HI(net33));
 sg13g2_tiehi _10293__34 (.L_HI(net34));
 sg13g2_tiehi _10309__35 (.L_HI(net35));
 sg13g2_tiehi _10294__36 (.L_HI(net36));
 sg13g2_tiehi _10304__37 (.L_HI(net37));
 sg13g2_tiehi _10305__38 (.L_HI(net38));
 sg13g2_tiehi _10306__39 (.L_HI(net39));
 sg13g2_tiehi _10307__40 (.L_HI(net40));
 sg13g2_tiehi _10295__41 (.L_HI(net41));
 sg13g2_tiehi _10530__42 (.L_HI(net42));
 sg13g2_tiehi _10486__43 (.L_HI(net43));
 sg13g2_tiehi _10485__44 (.L_HI(net44));
 sg13g2_tiehi _10529__45 (.L_HI(net45));
 sg13g2_tiehi _10484__46 (.L_HI(net46));
 sg13g2_tiehi _10546__47 (.L_HI(net47));
 sg13g2_tiehi _10483__48 (.L_HI(net48));
 sg13g2_tiehi _10528__49 (.L_HI(net49));
 sg13g2_tiehi _10482__50 (.L_HI(net50));
 sg13g2_tiehi _10481__51 (.L_HI(net51));
 sg13g2_tiehi _10527__52 (.L_HI(net52));
 sg13g2_tiehi _10480__53 (.L_HI(net53));
 sg13g2_tiehi _10545__54 (.L_HI(net54));
 sg13g2_tiehi _10479__55 (.L_HI(net55));
 sg13g2_tiehi _10526__56 (.L_HI(net56));
 sg13g2_tiehi _10478__57 (.L_HI(net57));
 sg13g2_tiehi _10554__58 (.L_HI(net58));
 sg13g2_tiehi _10477__59 (.L_HI(net59));
 sg13g2_tiehi _10525__60 (.L_HI(net60));
 sg13g2_tiehi _10476__61 (.L_HI(net61));
 sg13g2_tiehi _10544__62 (.L_HI(net62));
 sg13g2_tiehi _10475__63 (.L_HI(net63));
 sg13g2_tiehi _10524__64 (.L_HI(net64));
 sg13g2_tiehi _10474__65 (.L_HI(net65));
 sg13g2_tiehi _10473__66 (.L_HI(net66));
 sg13g2_tiehi _10523__67 (.L_HI(net67));
 sg13g2_tiehi _10472__68 (.L_HI(net68));
 sg13g2_tiehi _10543__69 (.L_HI(net69));
 sg13g2_tiehi _10471__70 (.L_HI(net70));
 sg13g2_tiehi _10522__71 (.L_HI(net71));
 sg13g2_tiehi _10470__72 (.L_HI(net72));
 sg13g2_tiehi _10553__73 (.L_HI(net73));
 sg13g2_tiehi _10469__74 (.L_HI(net74));
 sg13g2_tiehi _10521__75 (.L_HI(net75));
 sg13g2_tiehi _10468__76 (.L_HI(net76));
 sg13g2_tiehi _10542__77 (.L_HI(net77));
 sg13g2_tiehi _10467__78 (.L_HI(net78));
 sg13g2_tiehi _10520__79 (.L_HI(net79));
 sg13g2_tiehi _10466__80 (.L_HI(net80));
 sg13g2_tiehi _10465__81 (.L_HI(net81));
 sg13g2_tiehi _10519__82 (.L_HI(net82));
 sg13g2_tiehi _10464__83 (.L_HI(net83));
 sg13g2_tiehi _10541__84 (.L_HI(net84));
 sg13g2_tiehi _10463__85 (.L_HI(net85));
 sg13g2_tiehi _10518__86 (.L_HI(net86));
 sg13g2_tiehi _10462__87 (.L_HI(net87));
 sg13g2_tiehi _10552__88 (.L_HI(net88));
 sg13g2_tiehi _10461__89 (.L_HI(net89));
 sg13g2_tiehi _10517__90 (.L_HI(net90));
 sg13g2_tiehi _10460__91 (.L_HI(net91));
 sg13g2_tiehi _10540__92 (.L_HI(net92));
 sg13g2_tiehi _10459__93 (.L_HI(net93));
 sg13g2_tiehi _10516__94 (.L_HI(net94));
 sg13g2_tiehi _10458__95 (.L_HI(net95));
 sg13g2_tiehi _10457__96 (.L_HI(net96));
 sg13g2_tiehi _10515__97 (.L_HI(net97));
 sg13g2_tiehi _10456__98 (.L_HI(net98));
 sg13g2_tiehi _10539__99 (.L_HI(net99));
 sg13g2_tiehi _10455__100 (.L_HI(net100));
 sg13g2_tiehi _10514__101 (.L_HI(net101));
 sg13g2_tiehi _10454__102 (.L_HI(net102));
 sg13g2_tiehi _10551__103 (.L_HI(net103));
 sg13g2_tiehi _10453__104 (.L_HI(net104));
 sg13g2_tiehi _10513__105 (.L_HI(net105));
 sg13g2_tiehi _10452__106 (.L_HI(net106));
 sg13g2_tiehi _10538__107 (.L_HI(net107));
 sg13g2_tiehi _10451__108 (.L_HI(net108));
 sg13g2_tiehi _10512__109 (.L_HI(net109));
 sg13g2_tiehi _10450__110 (.L_HI(net110));
 sg13g2_tiehi _10449__111 (.L_HI(net111));
 sg13g2_tiehi _10511__112 (.L_HI(net112));
 sg13g2_tiehi _10448__113 (.L_HI(net113));
 sg13g2_tiehi _10537__114 (.L_HI(net114));
 sg13g2_tiehi _10447__115 (.L_HI(net115));
 sg13g2_tiehi _10510__116 (.L_HI(net116));
 sg13g2_tiehi _10446__117 (.L_HI(net117));
 sg13g2_tiehi _10550__118 (.L_HI(net118));
 sg13g2_tiehi _10445__119 (.L_HI(net119));
 sg13g2_tiehi _10509__120 (.L_HI(net120));
 sg13g2_tiehi _10444__121 (.L_HI(net121));
 sg13g2_tiehi _10308__122 (.L_HI(net122));
 sg13g2_tiehi _10536__123 (.L_HI(net123));
 sg13g2_tiehi _10443__124 (.L_HI(net124));
 sg13g2_tiehi _10508__125 (.L_HI(net125));
 sg13g2_tiehi _10442__126 (.L_HI(net126));
 sg13g2_tiehi _10441__127 (.L_HI(net127));
 sg13g2_tiehi _10507__128 (.L_HI(net128));
 sg13g2_tiehi _10440__129 (.L_HI(net129));
 sg13g2_tiehi _10535__130 (.L_HI(net130));
 sg13g2_tiehi _10439__131 (.L_HI(net131));
 sg13g2_tiehi _10506__132 (.L_HI(net132));
 sg13g2_tiehi _10438__133 (.L_HI(net133));
 sg13g2_tiehi _10549__134 (.L_HI(net134));
 sg13g2_tiehi _10437__135 (.L_HI(net135));
 sg13g2_tiehi _10505__136 (.L_HI(net136));
 sg13g2_tiehi _10436__137 (.L_HI(net137));
 sg13g2_tiehi _10435__138 (.L_HI(net138));
 sg13g2_tiehi _10434__139 (.L_HI(net139));
 sg13g2_tiehi _10433__140 (.L_HI(net140));
 sg13g2_tiehi _10432__141 (.L_HI(net141));
 sg13g2_tiehi _10431__142 (.L_HI(net142));
 sg13g2_tiehi _10430__143 (.L_HI(net143));
 sg13g2_tiehi _10429__144 (.L_HI(net144));
 sg13g2_tiehi _10428__145 (.L_HI(net145));
 sg13g2_tiehi _10534__146 (.L_HI(net146));
 sg13g2_tiehi _10427__147 (.L_HI(net147));
 sg13g2_tiehi _10426__148 (.L_HI(net148));
 sg13g2_tiehi _10425__149 (.L_HI(net149));
 sg13g2_tiehi _10493__150 (.L_HI(net150));
 sg13g2_tiehi _10424__151 (.L_HI(net151));
 sg13g2_tiehi _10533__152 (.L_HI(net152));
 sg13g2_tiehi _10423__153 (.L_HI(net153));
 sg13g2_tiehi _10492__154 (.L_HI(net154));
 sg13g2_tiehi _10422__155 (.L_HI(net155));
 sg13g2_tiehi _10548__156 (.L_HI(net156));
 sg13g2_tiehi _10421__157 (.L_HI(net157));
 sg13g2_tiehi _10491__158 (.L_HI(net158));
 sg13g2_tiehi _10420__159 (.L_HI(net159));
 sg13g2_tiehi _10532__160 (.L_HI(net160));
 sg13g2_tiehi _10419__161 (.L_HI(net161));
 sg13g2_tiehi _10490__162 (.L_HI(net162));
 sg13g2_tiehi _10418__163 (.L_HI(net163));
 sg13g2_tiehi _10417__164 (.L_HI(net164));
 sg13g2_tiehi _10489__165 (.L_HI(net165));
 sg13g2_tiehi _10416__166 (.L_HI(net166));
 sg13g2_tiehi _10531__167 (.L_HI(net167));
 sg13g2_tiehi _10415__168 (.L_HI(net168));
 sg13g2_tiehi _10488__169 (.L_HI(net169));
 sg13g2_tiehi _10414__170 (.L_HI(net170));
 sg13g2_tiehi _10547__171 (.L_HI(net171));
 sg13g2_tiehi _10413__172 (.L_HI(net172));
 sg13g2_tiehi _10487__173 (.L_HI(net173));
 sg13g2_tiehi _10412__174 (.L_HI(net174));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_herald_12 (.L_LO(net12));
 sg13g2_tielo tt_um_herald_13 (.L_LO(net13));
 sg13g2_tielo tt_um_herald_14 (.L_LO(net14));
 sg13g2_tielo tt_um_herald_15 (.L_LO(net15));
 sg13g2_tielo tt_um_herald_16 (.L_LO(net16));
 sg13g2_tielo tt_um_herald_17 (.L_LO(net17));
 sg13g2_tielo tt_um_herald_18 (.L_LO(net18));
 sg13g2_tielo tt_um_herald_19 (.L_LO(net19));
 sg13g2_tielo tt_um_herald_20 (.L_LO(net20));
 sg13g2_tielo tt_um_herald_21 (.L_LO(net21));
 sg13g2_tielo tt_um_herald_22 (.L_LO(net22));
 sg13g2_tielo tt_um_herald_23 (.L_LO(net23));
 sg13g2_tielo tt_um_herald_24 (.L_LO(net24));
 sg13g2_tielo tt_um_herald_25 (.L_LO(net25));
 sg13g2_tielo tt_um_herald_26 (.L_LO(net26));
 sg13g2_tiehi _10315__27 (.L_HI(net27));
 sg13g2_buf_8 fanout1019 (.A(_00564_),
    .X(net1019));
 sg13g2_buf_8 fanout1020 (.A(_00552_),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_8 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(_05025_),
    .X(net1023));
 sg13g2_buf_8 fanout1024 (.A(_05025_),
    .X(net1024));
 sg13g2_buf_8 fanout1025 (.A(_05025_),
    .X(net1025));
 sg13g2_buf_8 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_8 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_8 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_8 fanout1029 (.A(_00387_),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(_03936_),
    .X(net1030));
 sg13g2_buf_8 fanout1031 (.A(net1032),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(_00376_),
    .X(net1032));
 sg13g2_buf_8 fanout1033 (.A(net1035),
    .X(net1033));
 sg13g2_buf_1 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_8 fanout1035 (.A(_04850_),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(net1037),
    .X(net1036));
 sg13g2_buf_8 fanout1037 (.A(_04850_),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_8 fanout1039 (.A(net1040),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(_00416_),
    .X(net1040));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_8 fanout1042 (.A(net1043),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(net1044),
    .X(net1043));
 sg13g2_buf_8 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_8 fanout1045 (.A(_00415_),
    .X(net1045));
 sg13g2_buf_8 fanout1046 (.A(net1047),
    .X(net1046));
 sg13g2_buf_8 fanout1047 (.A(_00398_),
    .X(net1047));
 sg13g2_buf_8 fanout1048 (.A(_00397_),
    .X(net1048));
 sg13g2_buf_8 fanout1049 (.A(_04914_),
    .X(net1049));
 sg13g2_buf_8 fanout1050 (.A(net1052),
    .X(net1050));
 sg13g2_buf_1 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_8 fanout1052 (.A(_04897_),
    .X(net1052));
 sg13g2_buf_8 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_8 fanout1054 (.A(_04897_),
    .X(net1054));
 sg13g2_buf_8 fanout1055 (.A(net1058),
    .X(net1055));
 sg13g2_buf_1 fanout1056 (.A(net1058),
    .X(net1056));
 sg13g2_buf_8 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_buf_8 fanout1058 (.A(_04892_),
    .X(net1058));
 sg13g2_buf_8 fanout1059 (.A(net1061),
    .X(net1059));
 sg13g2_buf_1 fanout1060 (.A(net1061),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(_04848_),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(net1063),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(_04848_),
    .X(net1063));
 sg13g2_buf_8 fanout1064 (.A(_04756_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_04756_),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(_03374_),
    .X(net1066));
 sg13g2_buf_8 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_1 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(_01463_),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(net1071),
    .X(net1070));
 sg13g2_buf_8 fanout1071 (.A(_05007_),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(_04983_),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(net1077),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(net1077),
    .X(net1074));
 sg13g2_buf_8 fanout1075 (.A(net1077),
    .X(net1075));
 sg13g2_buf_1 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(_04922_),
    .X(net1077));
 sg13g2_buf_8 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(net1086),
    .X(net1081));
 sg13g2_buf_8 fanout1082 (.A(net1086),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_8 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_8 fanout1086 (.A(net1093),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(net1093),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(net1093),
    .X(net1088));
 sg13g2_buf_8 fanout1089 (.A(net1091),
    .X(net1089));
 sg13g2_buf_1 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_8 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_8 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_buf_8 fanout1093 (.A(_04921_),
    .X(net1093));
 sg13g2_buf_8 fanout1094 (.A(_04912_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_04912_),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_8 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(_04910_),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(_04866_),
    .X(net1100));
 sg13g2_buf_8 fanout1101 (.A(_04859_),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(_04859_),
    .X(net1102));
 sg13g2_buf_8 fanout1103 (.A(_03082_),
    .X(net1103));
 sg13g2_buf_8 fanout1104 (.A(_05006_),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(_05002_),
    .X(net1105));
 sg13g2_buf_8 fanout1106 (.A(_04984_),
    .X(net1106));
 sg13g2_buf_8 fanout1107 (.A(_04908_),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(_04905_),
    .X(net1108));
 sg13g2_buf_8 fanout1109 (.A(_04905_),
    .X(net1109));
 sg13g2_buf_8 fanout1110 (.A(_04869_),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(_04852_),
    .X(net1111));
 sg13g2_buf_8 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(net1116),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1116),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_8 fanout1116 (.A(_04562_),
    .X(net1116));
 sg13g2_buf_8 fanout1117 (.A(_03215_),
    .X(net1117));
 sg13g2_buf_8 fanout1118 (.A(_03081_),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(_00393_),
    .X(net1119));
 sg13g2_buf_1 fanout1120 (.A(_00393_),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_8 fanout1122 (.A(_00392_),
    .X(net1122));
 sg13g2_buf_8 fanout1123 (.A(_00325_),
    .X(net1123));
 sg13g2_buf_8 fanout1124 (.A(_04902_),
    .X(net1124));
 sg13g2_buf_8 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_8 fanout1126 (.A(_04902_),
    .X(net1126));
 sg13g2_buf_8 fanout1127 (.A(_04801_),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(_04801_),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_8 fanout1130 (.A(net1131),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(_04795_),
    .X(net1131));
 sg13g2_buf_8 fanout1132 (.A(net1133),
    .X(net1132));
 sg13g2_buf_8 fanout1133 (.A(_04794_),
    .X(net1133));
 sg13g2_buf_8 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(_04793_),
    .X(net1136));
 sg13g2_buf_8 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(_04792_),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(_04792_),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1144),
    .X(net1141));
 sg13g2_buf_1 fanout1142 (.A(net1144),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(net1144),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(_04770_),
    .X(net1144));
 sg13g2_buf_8 fanout1145 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net1145));
 sg13g2_buf_1 fanout1146 (.A(net530),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_1 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_8 fanout1150 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net522),
    .X(net1151));
 sg13g2_buf_1 fanout1152 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_1 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_8 fanout1156 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .X(net1156));
 sg13g2_buf_8 fanout1157 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .X(net1157));
 sg13g2_buf_1 fanout1158 (.A(net531),
    .X(net1158));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_8 fanout1162 (.A(net558),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_1 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .X(net1166));
 sg13g2_buf_8 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(net515),
    .X(net1168));
 sg13g2_buf_2 fanout1169 (.A(net1171),
    .X(net1169));
 sg13g2_buf_1 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .X(net1172));
 sg13g2_buf_8 fanout1173 (.A(net528),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(net1176),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(net527),
    .X(net1177));
 sg13g2_buf_1 fanout1178 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net1178));
 sg13g2_buf_2 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_2 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_1 fanout1181 (.A(net1183),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_8 fanout1183 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(net1190),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(net1187),
    .X(net1185));
 sg13g2_buf_1 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_8 fanout1187 (.A(net1189),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(net548),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net521),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(net533),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(net1198),
    .X(net1196));
 sg13g2_buf_1 fanout1197 (.A(net1198),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_8 fanout1199 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(net1204),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(net1203),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(net498),
    .X(net1204));
 sg13g2_buf_8 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(net537),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .X(net1207));
 sg13g2_buf_8 fanout1208 (.A(net1213),
    .X(net1208));
 sg13g2_buf_1 fanout1209 (.A(net1213),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1212),
    .X(net1210));
 sg13g2_buf_1 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(net542),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .X(net1215));
 sg13g2_buf_8 fanout1216 (.A(net1218),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(net1222),
    .X(net1219));
 sg13g2_buf_8 fanout1220 (.A(net1222),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_8 fanout1223 (.A(net506),
    .X(net1223));
 sg13g2_buf_8 fanout1224 (.A(net1226),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(net504),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net477),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(net377),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(net1232),
    .X(net1230));
 sg13g2_buf_1 fanout1231 (.A(net1232),
    .X(net1231));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_1 fanout1233 (.A(net524),
    .X(net1233));
 sg13g2_buf_8 fanout1234 (.A(net511),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(net538),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net510),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net1240),
    .X(net1237));
 sg13g2_buf_1 fanout1238 (.A(net1239),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(net1240),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(net540),
    .X(net1240));
 sg13g2_buf_8 fanout1241 (.A(net514),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(net523),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(net499),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net516),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(net513),
    .X(net1245));
 sg13g2_buf_8 fanout1246 (.A(net520),
    .X(net1246));
 sg13g2_buf_8 fanout1247 (.A(net338),
    .X(net1247));
 sg13g2_buf_8 fanout1248 (.A(net518),
    .X(net1248));
 sg13g2_buf_8 fanout1249 (.A(net503),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(net519),
    .X(net1250));
 sg13g2_buf_8 fanout1251 (.A(net507),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(net1253),
    .X(net1252));
 sg13g2_buf_8 fanout1253 (.A(net1254),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net1259),
    .X(net1254));
 sg13g2_buf_8 fanout1255 (.A(net1258),
    .X(net1255));
 sg13g2_buf_8 fanout1256 (.A(net1257),
    .X(net1256));
 sg13g2_buf_1 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_1 fanout1258 (.A(net1259),
    .X(net1258));
 sg13g2_buf_8 fanout1259 (.A(\cordic_inst.cordic_state[7] ),
    .X(net1259));
 sg13g2_buf_8 fanout1260 (.A(net1263),
    .X(net1260));
 sg13g2_buf_1 fanout1261 (.A(net1263),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(net1263),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(net1267),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(net1267),
    .X(net1264));
 sg13g2_buf_1 fanout1265 (.A(net1267),
    .X(net1265));
 sg13g2_buf_8 fanout1266 (.A(net1267),
    .X(net1266));
 sg13g2_buf_8 fanout1267 (.A(net1268),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(\cordic_inst.cordic_state[6] ),
    .X(net1268));
 sg13g2_buf_8 fanout1269 (.A(net1271),
    .X(net1269));
 sg13g2_buf_1 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_8 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_8 fanout1273 (.A(net534),
    .X(net1273));
 sg13g2_buf_8 fanout1274 (.A(net1275),
    .X(net1274));
 sg13g2_buf_8 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_8 fanout1276 (.A(net1281),
    .X(net1276));
 sg13g2_buf_8 fanout1277 (.A(net1280),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(net1280),
    .X(net1278));
 sg13g2_buf_8 fanout1279 (.A(net1280),
    .X(net1279));
 sg13g2_buf_2 fanout1280 (.A(net1281),
    .X(net1280));
 sg13g2_buf_8 fanout1281 (.A(net549),
    .X(net1281));
 sg13g2_buf_8 fanout1282 (.A(net1286),
    .X(net1282));
 sg13g2_buf_8 fanout1283 (.A(net1285),
    .X(net1283));
 sg13g2_buf_8 fanout1284 (.A(net1285),
    .X(net1284));
 sg13g2_buf_8 fanout1285 (.A(net1286),
    .X(net1285));
 sg13g2_buf_8 fanout1286 (.A(net1291),
    .X(net1286));
 sg13g2_buf_8 fanout1287 (.A(net1291),
    .X(net1287));
 sg13g2_buf_8 fanout1288 (.A(net1291),
    .X(net1288));
 sg13g2_buf_8 fanout1289 (.A(net1290),
    .X(net1289));
 sg13g2_buf_8 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_8 fanout1291 (.A(net1292),
    .X(net1291));
 sg13g2_buf_8 fanout1292 (.A(net529),
    .X(net1292));
 sg13g2_buf_8 fanout1293 (.A(net1295),
    .X(net1293));
 sg13g2_buf_8 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_8 fanout1295 (.A(mac_en_mac),
    .X(net1295));
 sg13g2_buf_8 fanout1296 (.A(net1300),
    .X(net1296));
 sg13g2_buf_8 fanout1297 (.A(net1299),
    .X(net1297));
 sg13g2_buf_1 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_8 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_8 fanout1300 (.A(mac_en_multiply),
    .X(net1300));
 sg13g2_buf_8 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_8 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_1 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_8 fanout1304 (.A(net1311),
    .X(net1304));
 sg13g2_buf_8 fanout1305 (.A(net1306),
    .X(net1305));
 sg13g2_buf_8 fanout1306 (.A(net1311),
    .X(net1306));
 sg13g2_buf_8 fanout1307 (.A(net1308),
    .X(net1307));
 sg13g2_buf_1 fanout1308 (.A(net1311),
    .X(net1308));
 sg13g2_buf_8 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_8 fanout1310 (.A(net1311),
    .X(net1310));
 sg13g2_buf_8 fanout1311 (.A(cordic_en_sqrt),
    .X(net1311));
 sg13g2_buf_8 fanout1312 (.A(net1313),
    .X(net1312));
 sg13g2_buf_8 fanout1313 (.A(net1314),
    .X(net1313));
 sg13g2_buf_8 fanout1314 (.A(net1316),
    .X(net1314));
 sg13g2_buf_8 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_8 fanout1316 (.A(cordic_en_atan2),
    .X(net1316));
 sg13g2_buf_8 fanout1317 (.A(cordic_en_sin_cos),
    .X(net1317));
 sg13g2_buf_1 fanout1318 (.A(cordic_en_sin_cos),
    .X(net1318));
 sg13g2_buf_8 fanout1319 (.A(net1321),
    .X(net1319));
 sg13g2_buf_1 fanout1320 (.A(net1321),
    .X(net1320));
 sg13g2_buf_8 fanout1321 (.A(cordic_en_sin_cos),
    .X(net1321));
 sg13g2_buf_8 fanout1322 (.A(net1323),
    .X(net1322));
 sg13g2_buf_8 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_8 fanout1324 (.A(net1325),
    .X(net1324));
 sg13g2_buf_8 fanout1325 (.A(net494),
    .X(net1325));
 sg13g2_buf_8 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_8 fanout1327 (.A(net1328),
    .X(net1327));
 sg13g2_buf_8 fanout1328 (.A(net550),
    .X(net1328));
 sg13g2_buf_8 fanout1329 (.A(net1330),
    .X(net1329));
 sg13g2_buf_8 fanout1330 (.A(net526),
    .X(net1330));
 sg13g2_buf_8 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_8 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_8 fanout1333 (.A(net544),
    .X(net1333));
 sg13g2_buf_8 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_8 fanout1335 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .X(net1335));
 sg13g2_buf_8 fanout1336 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .X(net1336));
 sg13g2_buf_8 fanout1337 (.A(net1341),
    .X(net1337));
 sg13g2_buf_2 fanout1338 (.A(net1341),
    .X(net1338));
 sg13g2_buf_8 fanout1339 (.A(net1340),
    .X(net1339));
 sg13g2_buf_8 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_8 fanout1341 (.A(net556),
    .X(net1341));
 sg13g2_buf_8 fanout1342 (.A(net1347),
    .X(net1342));
 sg13g2_buf_1 fanout1343 (.A(net1347),
    .X(net1343));
 sg13g2_buf_2 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_1 fanout1345 (.A(net1346),
    .X(net1345));
 sg13g2_buf_1 fanout1346 (.A(net1347),
    .X(net1346));
 sg13g2_buf_8 fanout1347 (.A(net546),
    .X(net1347));
 sg13g2_buf_8 fanout1348 (.A(net1351),
    .X(net1348));
 sg13g2_buf_8 fanout1349 (.A(net1350),
    .X(net1349));
 sg13g2_buf_8 fanout1350 (.A(net1351),
    .X(net1350));
 sg13g2_buf_8 fanout1351 (.A(net554),
    .X(net1351));
 sg13g2_buf_8 fanout1352 (.A(net1357),
    .X(net1352));
 sg13g2_buf_8 fanout1353 (.A(net1354),
    .X(net1353));
 sg13g2_buf_8 fanout1354 (.A(net1357),
    .X(net1354));
 sg13g2_buf_8 fanout1355 (.A(net1357),
    .X(net1355));
 sg13g2_buf_1 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_8 fanout1357 (.A(net532),
    .X(net1357));
 sg13g2_buf_8 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_8 fanout1359 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ),
    .X(net1359));
 sg13g2_buf_8 fanout1360 (.A(net1361),
    .X(net1360));
 sg13g2_buf_8 fanout1361 (.A(net1364),
    .X(net1361));
 sg13g2_buf_8 fanout1362 (.A(net1364),
    .X(net1362));
 sg13g2_buf_1 fanout1363 (.A(net1364),
    .X(net1363));
 sg13g2_buf_8 fanout1364 (.A(net512),
    .X(net1364));
 sg13g2_buf_8 fanout1365 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .X(net1365));
 sg13g2_buf_8 fanout1366 (.A(net1371),
    .X(net1366));
 sg13g2_buf_1 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_8 fanout1368 (.A(net1371),
    .X(net1368));
 sg13g2_buf_8 fanout1369 (.A(net1371),
    .X(net1369));
 sg13g2_buf_8 fanout1370 (.A(net1371),
    .X(net1370));
 sg13g2_buf_8 fanout1371 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .X(net1371));
 sg13g2_buf_8 fanout1372 (.A(net1378),
    .X(net1372));
 sg13g2_buf_8 fanout1373 (.A(net1375),
    .X(net1373));
 sg13g2_buf_8 fanout1374 (.A(net1375),
    .X(net1374));
 sg13g2_buf_8 fanout1375 (.A(net1378),
    .X(net1375));
 sg13g2_buf_8 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_8 fanout1377 (.A(net1378),
    .X(net1377));
 sg13g2_buf_8 fanout1378 (.A(net505),
    .X(net1378));
 sg13g2_buf_8 fanout1379 (.A(net1386),
    .X(net1379));
 sg13g2_buf_8 fanout1380 (.A(net1385),
    .X(net1380));
 sg13g2_buf_1 fanout1381 (.A(net1385),
    .X(net1381));
 sg13g2_buf_8 fanout1382 (.A(net1385),
    .X(net1382));
 sg13g2_buf_8 fanout1383 (.A(net1385),
    .X(net1383));
 sg13g2_buf_1 fanout1384 (.A(net1385),
    .X(net1384));
 sg13g2_buf_8 fanout1385 (.A(net1386),
    .X(net1385));
 sg13g2_buf_8 fanout1386 (.A(net551),
    .X(net1386));
 sg13g2_buf_8 fanout1387 (.A(net1393),
    .X(net1387));
 sg13g2_buf_1 fanout1388 (.A(net1393),
    .X(net1388));
 sg13g2_buf_8 fanout1389 (.A(net1393),
    .X(net1389));
 sg13g2_buf_8 fanout1390 (.A(net1392),
    .X(net1390));
 sg13g2_buf_1 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_8 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_8 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_8 fanout1394 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ),
    .X(net1394));
 sg13g2_buf_8 fanout1395 (.A(net1402),
    .X(net1395));
 sg13g2_buf_8 fanout1396 (.A(net1397),
    .X(net1396));
 sg13g2_buf_8 fanout1397 (.A(net1401),
    .X(net1397));
 sg13g2_buf_8 fanout1398 (.A(net1399),
    .X(net1398));
 sg13g2_buf_8 fanout1399 (.A(net1400),
    .X(net1399));
 sg13g2_buf_8 fanout1400 (.A(net1401),
    .X(net1400));
 sg13g2_buf_8 fanout1401 (.A(net1402),
    .X(net1401));
 sg13g2_buf_8 fanout1402 (.A(net535),
    .X(net1402));
 sg13g2_buf_8 fanout1403 (.A(net1404),
    .X(net1403));
 sg13g2_buf_8 fanout1404 (.A(net1405),
    .X(net1404));
 sg13g2_buf_8 fanout1405 (.A(net1408),
    .X(net1405));
 sg13g2_buf_8 fanout1406 (.A(net1407),
    .X(net1406));
 sg13g2_buf_8 fanout1407 (.A(net1408),
    .X(net1407));
 sg13g2_buf_8 fanout1408 (.A(net497),
    .X(net1408));
 sg13g2_buf_8 fanout1409 (.A(net462),
    .X(net1409));
 sg13g2_buf_8 fanout1410 (.A(net1411),
    .X(net1410));
 sg13g2_buf_8 fanout1411 (.A(net555),
    .X(net1411));
 sg13g2_buf_1 fanout1412 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ),
    .X(net1412));
 sg13g2_buf_8 fanout1413 (.A(net1414),
    .X(net1413));
 sg13g2_buf_8 fanout1414 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ),
    .X(net1414));
 sg13g2_buf_8 fanout1415 (.A(net1417),
    .X(net1415));
 sg13g2_buf_8 fanout1416 (.A(net1417),
    .X(net1416));
 sg13g2_buf_8 fanout1417 (.A(net501),
    .X(net1417));
 sg13g2_buf_8 fanout1418 (.A(net1420),
    .X(net1418));
 sg13g2_buf_1 fanout1419 (.A(net1420),
    .X(net1419));
 sg13g2_buf_8 fanout1420 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .X(net1420));
 sg13g2_buf_8 fanout1421 (.A(net1423),
    .X(net1421));
 sg13g2_buf_8 fanout1422 (.A(net1423),
    .X(net1422));
 sg13g2_buf_8 fanout1423 (.A(net541),
    .X(net1423));
 sg13g2_buf_8 fanout1424 (.A(net1427),
    .X(net1424));
 sg13g2_buf_2 fanout1425 (.A(net1427),
    .X(net1425));
 sg13g2_buf_8 fanout1426 (.A(net1427),
    .X(net1426));
 sg13g2_buf_8 fanout1427 (.A(net552),
    .X(net1427));
 sg13g2_buf_8 fanout1428 (.A(net1431),
    .X(net1428));
 sg13g2_buf_2 fanout1429 (.A(net1431),
    .X(net1429));
 sg13g2_buf_8 fanout1430 (.A(net1431),
    .X(net1430));
 sg13g2_buf_8 fanout1431 (.A(net543),
    .X(net1431));
 sg13g2_buf_8 fanout1432 (.A(net1435),
    .X(net1432));
 sg13g2_buf_8 fanout1433 (.A(net1435),
    .X(net1433));
 sg13g2_buf_8 fanout1434 (.A(net1435),
    .X(net1434));
 sg13g2_buf_8 fanout1435 (.A(net539),
    .X(net1435));
 sg13g2_buf_8 fanout1436 (.A(net1440),
    .X(net1436));
 sg13g2_buf_1 fanout1437 (.A(net1440),
    .X(net1437));
 sg13g2_buf_8 fanout1438 (.A(net1440),
    .X(net1438));
 sg13g2_buf_1 fanout1439 (.A(net1440),
    .X(net1439));
 sg13g2_buf_8 fanout1440 (.A(net553),
    .X(net1440));
 sg13g2_buf_8 fanout1441 (.A(net1445),
    .X(net1441));
 sg13g2_buf_2 fanout1442 (.A(net1445),
    .X(net1442));
 sg13g2_buf_8 fanout1443 (.A(net1445),
    .X(net1443));
 sg13g2_buf_8 fanout1444 (.A(net1445),
    .X(net1444));
 sg13g2_buf_8 fanout1445 (.A(net557),
    .X(net1445));
 sg13g2_buf_8 fanout1446 (.A(net1450),
    .X(net1446));
 sg13g2_buf_1 fanout1447 (.A(net1450),
    .X(net1447));
 sg13g2_buf_8 fanout1448 (.A(net1450),
    .X(net1448));
 sg13g2_buf_8 fanout1449 (.A(net1450),
    .X(net1449));
 sg13g2_buf_8 fanout1450 (.A(net547),
    .X(net1450));
 sg13g2_buf_8 fanout1451 (.A(net1452),
    .X(net1451));
 sg13g2_buf_8 fanout1452 (.A(net536),
    .X(net1452));
 sg13g2_buf_8 fanout1453 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .X(net1453));
 sg13g2_buf_8 fanout1454 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .X(net1454));
 sg13g2_buf_8 fanout1455 (.A(net1456),
    .X(net1455));
 sg13g2_buf_8 fanout1456 (.A(net1459),
    .X(net1456));
 sg13g2_buf_8 fanout1457 (.A(net1458),
    .X(net1457));
 sg13g2_buf_8 fanout1458 (.A(net1459),
    .X(net1458));
 sg13g2_buf_8 fanout1459 (.A(net545),
    .X(net1459));
 sg13g2_buf_8 fanout1460 (.A(net1461),
    .X(net1460));
 sg13g2_buf_8 fanout1461 (.A(net525),
    .X(net1461));
 sg13g2_buf_8 fanout1462 (.A(net1463),
    .X(net1462));
 sg13g2_buf_8 fanout1463 (.A(net1464),
    .X(net1463));
 sg13g2_buf_8 fanout1464 (.A(net560),
    .X(net1464));
 sg13g2_buf_8 fanout1465 (.A(net1466),
    .X(net1465));
 sg13g2_buf_8 fanout1466 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ),
    .X(net1466));
 sg13g2_buf_8 fanout1467 (.A(net1468),
    .X(net1467));
 sg13g2_buf_8 fanout1468 (.A(net1469),
    .X(net1468));
 sg13g2_buf_8 fanout1469 (.A(net508),
    .X(net1469));
 sg13g2_buf_8 fanout1470 (.A(net1474),
    .X(net1470));
 sg13g2_buf_8 fanout1471 (.A(net1472),
    .X(net1471));
 sg13g2_buf_8 fanout1472 (.A(net1474),
    .X(net1472));
 sg13g2_buf_8 fanout1473 (.A(net1474),
    .X(net1473));
 sg13g2_buf_8 fanout1474 (.A(net517),
    .X(net1474));
 sg13g2_buf_8 fanout1475 (.A(net201),
    .X(net1475));
 sg13g2_buf_8 fanout1476 (.A(net1477),
    .X(net1476));
 sg13g2_buf_8 fanout1477 (.A(net1481),
    .X(net1477));
 sg13g2_buf_8 fanout1478 (.A(net1481),
    .X(net1478));
 sg13g2_buf_8 fanout1479 (.A(net1480),
    .X(net1479));
 sg13g2_buf_1 fanout1480 (.A(net1481),
    .X(net1480));
 sg13g2_buf_8 fanout1481 (.A(net1488),
    .X(net1481));
 sg13g2_buf_8 fanout1482 (.A(net1483),
    .X(net1482));
 sg13g2_buf_8 fanout1483 (.A(net1484),
    .X(net1483));
 sg13g2_buf_8 fanout1484 (.A(net1488),
    .X(net1484));
 sg13g2_buf_8 fanout1485 (.A(net1488),
    .X(net1485));
 sg13g2_buf_1 fanout1486 (.A(net1487),
    .X(net1486));
 sg13g2_buf_8 fanout1487 (.A(net1488),
    .X(net1487));
 sg13g2_buf_8 fanout1488 (.A(_04800_),
    .X(net1488));
 sg13g2_buf_8 fanout1489 (.A(net1490),
    .X(net1489));
 sg13g2_buf_8 fanout1490 (.A(net1496),
    .X(net1490));
 sg13g2_buf_8 fanout1491 (.A(net1492),
    .X(net1491));
 sg13g2_buf_8 fanout1492 (.A(net1493),
    .X(net1492));
 sg13g2_buf_2 fanout1493 (.A(net1496),
    .X(net1493));
 sg13g2_buf_8 fanout1494 (.A(net1496),
    .X(net1494));
 sg13g2_buf_8 fanout1495 (.A(net1496),
    .X(net1495));
 sg13g2_buf_8 fanout1496 (.A(rst_n),
    .X(net1496));
 sg13g2_buf_8 fanout1497 (.A(net1498),
    .X(net1497));
 sg13g2_buf_8 fanout1498 (.A(net1505),
    .X(net1498));
 sg13g2_buf_8 fanout1499 (.A(net1505),
    .X(net1499));
 sg13g2_buf_8 fanout1500 (.A(net1505),
    .X(net1500));
 sg13g2_buf_8 fanout1501 (.A(net1504),
    .X(net1501));
 sg13g2_buf_8 fanout1502 (.A(net1504),
    .X(net1502));
 sg13g2_buf_8 fanout1503 (.A(net1504),
    .X(net1503));
 sg13g2_buf_8 fanout1504 (.A(net1505),
    .X(net1504));
 sg13g2_buf_8 fanout1505 (.A(rst_n),
    .X(net1505));
 sg13g2_buf_8 fanout1506 (.A(net1509),
    .X(net1506));
 sg13g2_buf_8 fanout1507 (.A(net1509),
    .X(net1507));
 sg13g2_buf_8 fanout1508 (.A(net1509),
    .X(net1508));
 sg13g2_buf_8 fanout1509 (.A(net1522),
    .X(net1509));
 sg13g2_buf_8 fanout1510 (.A(net1513),
    .X(net1510));
 sg13g2_buf_8 fanout1511 (.A(net1513),
    .X(net1511));
 sg13g2_buf_1 fanout1512 (.A(net1513),
    .X(net1512));
 sg13g2_buf_8 fanout1513 (.A(net1522),
    .X(net1513));
 sg13g2_buf_8 fanout1514 (.A(net1515),
    .X(net1514));
 sg13g2_buf_8 fanout1515 (.A(net1522),
    .X(net1515));
 sg13g2_buf_8 fanout1516 (.A(net1520),
    .X(net1516));
 sg13g2_buf_8 fanout1517 (.A(net1519),
    .X(net1517));
 sg13g2_buf_8 fanout1518 (.A(net1520),
    .X(net1518));
 sg13g2_buf_1 fanout1519 (.A(net1520),
    .X(net1519));
 sg13g2_buf_8 fanout1520 (.A(net1521),
    .X(net1520));
 sg13g2_buf_8 fanout1521 (.A(net1522),
    .X(net1521));
 sg13g2_buf_8 fanout1522 (.A(rst_n),
    .X(net1522));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_tielo tt_um_herald_11 (.L_LO(net11));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_1_clk));
 sg13g2_inv_8 clkload5 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_29_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(mac_en_get_mac),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00273_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold3 (.A(mac_en_get_multiply),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00272_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cordic_inst.cordic_state[34] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00112_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac_inst.get_multiply[15] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac_inst.get_multiply[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac_inst.get_multiply[14] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac_inst.get_multiply[4] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac_inst.get_multiply[17] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac_inst.get_multiply[13] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac_inst.get_multiply[12] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac_inst.get_multiply[6] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mac_inst.get_multiply[0] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mac_inst.get_multiply[23] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold17 (.A(\result_reg[16] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00067_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mac_inst.get_multiply[10] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cordic_inst.operation_pending ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold21 (.A(_01460_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac_inst.get_multiply[18] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac_inst.accumulator[20] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold24 (.A(\result_reg[20] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold25 (.A(_00071_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold26 (.A(\result_reg[4] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold27 (.A(\byte_counter[2] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold28 (.A(_00028_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cordic_inst.current_op[2] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mac_inst.accumulator[11] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold31 (.A(_04644_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold32 (.A(_00259_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold33 (.A(\result_reg[19] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold34 (.A(_00070_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold35 (.A(\result_reg[18] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00069_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cmd_reg[6] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold38 (.A(\result_reg[15] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold39 (.A(_00066_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold40 (.A(\result_reg[13] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold41 (.A(_00064_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mac_inst.accumulator[19] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold43 (.A(_00267_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold44 (.A(\result_reg[24] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00110_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cordic_inst.current_op[1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cmd_reg[7] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold48 (.A(\result_reg[25] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold49 (.A(_00111_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mac_inst.accumulator[18] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00266_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold52 (.A(\result_reg[27] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold53 (.A(_00113_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold54 (.A(\result_reg[11] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold55 (.A(_00062_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold56 (.A(\result_reg[21] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold57 (.A(_00072_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold58 (.A(\result_reg[28] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold59 (.A(_00114_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mac_inst.accumulator[13] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold61 (.A(_00261_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mac_inst.accumulator[21] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold63 (.A(_00269_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold64 (.A(\result_reg[30] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00116_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mac_inst.accumulator[14] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold67 (.A(_00262_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mac_inst.accumulator[23] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold69 (.A(\result_reg[1] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00052_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold71 (.A(\result_reg[29] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold72 (.A(_00115_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold73 (.A(\result_reg[17] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00068_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mac_inst.accumulator[12] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold76 (.A(_04651_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00260_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold78 (.A(\result_reg[47] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold79 (.A(_00133_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mac_inst.accumulator[8] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold81 (.A(_04625_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac_inst.get_multiply[9] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold83 (.A(_00233_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold84 (.A(\result_reg[8] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00059_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac_inst.get_multiply[22] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold87 (.A(_04476_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold88 (.A(_00246_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac_inst.accumulator[22] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold90 (.A(_04748_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold91 (.A(\result_reg[46] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold92 (.A(_00132_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mac_inst.accumulator[5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold94 (.A(_04593_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold95 (.A(\result_reg[44] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00130_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac_inst.get_multiply[20] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold98 (.A(_04228_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold99 (.A(_00244_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold100 (.A(\result_reg[33] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00119_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac_inst.get_multiply[21] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold103 (.A(_04353_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold104 (.A(_00245_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold105 (.A(uo_out[4]),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00349_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mac_inst.accumulator[1] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold108 (.A(_04573_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mac_inst.get_multiply[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mac_inst.accumulator[17] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac_inst.get_multiply[19] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold112 (.A(_04104_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold113 (.A(_00243_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mac_inst.get_multiply[16] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold115 (.A(_03705_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold116 (.A(_00240_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold117 (.A(\result_reg[39] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold118 (.A(_00125_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mac_inst.accumulator[16] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold120 (.A(_04695_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold121 (.A(\result_reg[42] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00128_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac_inst.get_multiply[7] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold124 (.A(_00231_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cmd_reg[4] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mac_inst.get_multiply[3] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mac_inst.accumulator[15] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold128 (.A(_00263_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cmd_reg[2] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac_inst.get_multiply[8] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold131 (.A(_00232_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold132 (.A(\result_reg[22] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00073_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold134 (.A(\result_reg[14] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold135 (.A(_00065_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac_inst.get_multiply[2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold137 (.A(uo_out[3]),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold138 (.A(_00344_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold139 (.A(\result_reg[43] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold140 (.A(_00129_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac_inst.accumulator[2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold142 (.A(_04579_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold143 (.A(\result_reg[37] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold144 (.A(_00123_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold145 (.A(uo_out[1]),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold146 (.A(_00334_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cordic_atan2_result[14] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00562_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold149 (.A(\result_reg[35] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold150 (.A(_00121_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold151 (.A(cordic_en_get_sin_cos),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold152 (.A(_01461_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold153 (.A(_01462_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cmd_reg[3] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cmd_reg[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold156 (.A(_04898_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold157 (.A(_00016_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold158 (.A(uo_out[5]),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold159 (.A(_00354_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold160 (.A(\result_reg[31] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold161 (.A(_00117_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold162 (.A(\result_reg[34] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold163 (.A(_00120_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cordic_inst.cordic_state[46] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold165 (.A(_00124_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cmd_reg[5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold167 (.A(uo_out[2]),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00339_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold169 (.A(\result_reg[32] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold170 (.A(_00118_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold171 (.A(\result_reg[12] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00063_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mac_inst.accumulator[7] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold174 (.A(_04614_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cordic_atan2_result[20] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold176 (.A(_00610_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cordic_atan2_result[8] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold178 (.A(\exec_phase[1] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold179 (.A(_04886_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00021_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold181 (.A(\result_reg[45] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold182 (.A(_00131_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold183 (.A(\result_reg[41] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold184 (.A(_00127_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold185 (.A(\result_reg[40] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold186 (.A(_00126_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cordic_atan2_result[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cordic_atan2_result[2] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold189 (.A(uo_out[6]),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold190 (.A(_00359_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold191 (.A(uo_out[0]),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold192 (.A(_00329_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mac_inst.get_multiply[11] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold194 (.A(_03035_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold195 (.A(_00235_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold196 (.A(\result_reg[3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00054_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cordic_atan2_result[12] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold199 (.A(_00539_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold200 (.A(\result_reg[23] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold201 (.A(_00074_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cordic_atan2_result[6] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold203 (.A(_00023_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold204 (.A(_04956_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00014_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cordic_atan2_result[10] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mac_inst.accumulator[10] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold208 (.A(_04643_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold209 (.A(\result_reg[36] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold210 (.A(_00122_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mac_inst.accumulator[4] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold212 (.A(_04592_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mac_inst.accumulator[6] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold214 (.A(_04607_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cordic_atan2_result[21] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold216 (.A(_00617_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold217 (.A(\result_reg[6] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold218 (.A(_00057_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mac_inst.accumulator[3] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold220 (.A(_04585_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cordic_atan2_result[19] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold222 (.A(_00601_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mac_inst.accumulator[0] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cordic_atan2_result[5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold225 (.A(\result_reg[10] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold226 (.A(\cordic_atan2_result[7] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cordic_atan2_result[13] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold228 (.A(_00155_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cordic_atan2_result[16] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold230 (.A(_00578_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cordic_atan2_result[11] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold233 (.A(\result_reg[2] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold234 (.A(_00053_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold235 (.A(\cordic_atan2_result[15] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold236 (.A(_00570_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mac_inst.accumulator[9] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold238 (.A(_04632_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cordic_atan2_result[0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold240 (.A(_00403_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cordic_inst.cordic_state[56] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold242 (.A(_00190_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cordic_inst.current_op[0] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold244 (.A(_04891_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cmd_reg[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold246 (.A(_04847_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold247 (.A(\cordic_atan2_result[22] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00624_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cordic_inst.cordic_state[36] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold250 (.A(\result_reg[7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold251 (.A(\cordic_atan2_result[18] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold252 (.A(_00594_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold253 (.A(\result_reg[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cordic_inst.cordic_state[39] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold255 (.A(wr_prev),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cordic_inst.cordic_state[72] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold257 (.A(_01369_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold258 (.A(cordic_busy),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold259 (.A(_00395_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cordic_atan2_result[1] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold261 (.A(_00424_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cordic_inst.cordic_state[78] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cordic_atan2_result[9] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold264 (.A(_00503_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold266 (.A(_00391_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00134_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold268 (.A(uo_out[7]),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00082_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold270 (.A(\result_reg[9] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold271 (.A(\result_reg[5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold272 (.A(_00056_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold273 (.A(\state[1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cordic_atan2_result[17] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold275 (.A(_00584_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold276 (.A(\byte_counter[1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold277 (.A(_00027_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold278 (.A(\byte_counter[0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold279 (.A(_00026_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cordic_inst.cordic_state[74] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold281 (.A(\cordic_inst.cordic_state[70] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold282 (.A(\state[0] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cordic_atan2_result[23] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00165_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold286 (.A(\cordic_inst.cordic_state[62] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00196_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold288 (.A(\state[2] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cordic_inst.cordic_state[32] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cordic_inst.cordic_state[66] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cordic_inst.cordic_state[41] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cordic_inst.cordic_state[69] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cordic_inst.cordic_state[38] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00172_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold295 (.A(\cordic_inst.cordic_state[65] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold296 (.A(\cmd_reg[0] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold297 (.A(\cordic_inst.cordic_state[71] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cordic_inst.cordic_state[58] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cordic_inst.cordic_state[35] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold300 (.A(\cordic_inst.cordic_state[37] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00171_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cordic_inst.cordic_state[68] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold303 (.A(\exec_phase[2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold304 (.A(_04901_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cordic_inst.cordic_state[40] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cordic_inst.cordic_state[75] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold307 (.A(\cordic_inst.cordic_state[60] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold308 (.A(_01180_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold309 (.A(\cordic_inst.cordic_state[57] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00191_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold311 (.A(\cordic_inst.cordic_state[59] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00193_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cordic_inst.cordic_state[64] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold314 (.A(\cordic_inst.cordic_state[53] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold315 (.A(_00187_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold316 (.A(\cordic_inst.cordic_state[61] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00195_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold318 (.A(\cordic_inst.cordic_state[0] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold319 (.A(_00396_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold320 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold321 (.A(\cordic_inst.cordic_state[63] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold322 (.A(\cordic_inst.cordic_state[54] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold323 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold324 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold325 (.A(\cordic_inst.cordic_state[50] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold326 (.A(\cordic_atan2_result[3] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold327 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cordic_inst.cordic_state[33] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cordic_inst.cordic_state[44] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold330 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold331 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold332 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cordic_inst.cordic_state[42] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold334 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold335 (.A(\cordic_inst.cordic_state[76] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold336 (.A(\cordic_inst.cordic_state[67] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cordic_inst.cordic_state[77] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold338 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold339 (.A(\cordic_inst.cordic_state[48] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold340 (.A(\cordic_inst.cordic_state[52] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold342 (.A(\cordic_inst.cordic_state[49] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold343 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold344 (.A(\cordic_inst.cordic_state[45] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold345 (.A(\cordic_inst.cordic_state[43] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cordic_inst.cordic_state[47] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold347 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold348 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold349 (.A(\cordic_inst.cordic_state[51] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold350 (.A(\cordic_inst.cordic_state[79] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold351 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold352 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold353 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold355 (.A(\cordic_inst.cordic_state[3] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold356 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold358 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold359 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold360 (.A(\cordic_inst.cordic_state[5] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold361 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold362 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold363 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold364 (.A(\cordic_inst.cordic_state[73] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold365 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold366 (.A(\cordic_inst.cordic_state[55] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold367 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold368 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold369 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold370 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold371 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold372 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold373 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold374 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold375 (.A(\cordic_inst.cordic_state[4] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold376 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold377 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold378 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold379 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold381 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold382 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold383 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold385 (.A(\mac_inst.accumulator[4] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold386 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold387 (.A(\cordic_inst.cordic_state[63] ),
    .X(net561));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_fill_2 FILLER_4_637 ();
 sg13g2_fill_1 FILLER_4_639 ();
 sg13g2_decap_8 FILLER_4_646 ();
 sg13g2_decap_8 FILLER_4_653 ();
 sg13g2_fill_2 FILLER_4_660 ();
 sg13g2_fill_1 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_670 ();
 sg13g2_decap_8 FILLER_4_677 ();
 sg13g2_decap_8 FILLER_4_684 ();
 sg13g2_decap_8 FILLER_4_691 ();
 sg13g2_decap_8 FILLER_4_698 ();
 sg13g2_decap_8 FILLER_4_705 ();
 sg13g2_decap_8 FILLER_4_712 ();
 sg13g2_decap_8 FILLER_4_719 ();
 sg13g2_decap_8 FILLER_4_726 ();
 sg13g2_decap_8 FILLER_4_733 ();
 sg13g2_decap_8 FILLER_4_740 ();
 sg13g2_decap_8 FILLER_4_747 ();
 sg13g2_decap_8 FILLER_4_754 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_8 FILLER_4_768 ();
 sg13g2_decap_8 FILLER_4_775 ();
 sg13g2_decap_8 FILLER_4_782 ();
 sg13g2_decap_8 FILLER_4_789 ();
 sg13g2_decap_8 FILLER_4_796 ();
 sg13g2_decap_8 FILLER_4_803 ();
 sg13g2_decap_8 FILLER_4_810 ();
 sg13g2_decap_8 FILLER_4_817 ();
 sg13g2_decap_8 FILLER_4_824 ();
 sg13g2_decap_8 FILLER_4_831 ();
 sg13g2_decap_8 FILLER_4_838 ();
 sg13g2_decap_8 FILLER_4_845 ();
 sg13g2_decap_8 FILLER_4_852 ();
 sg13g2_fill_2 FILLER_4_859 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_4 FILLER_5_56 ();
 sg13g2_fill_1 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_66 ();
 sg13g2_decap_8 FILLER_5_73 ();
 sg13g2_decap_8 FILLER_5_80 ();
 sg13g2_decap_8 FILLER_5_87 ();
 sg13g2_decap_8 FILLER_5_94 ();
 sg13g2_decap_4 FILLER_5_101 ();
 sg13g2_fill_1 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_118 ();
 sg13g2_decap_4 FILLER_5_125 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_decap_8 FILLER_5_148 ();
 sg13g2_decap_4 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_164 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_fill_2 FILLER_5_192 ();
 sg13g2_fill_1 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_220 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_decap_4 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_fill_2 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_decap_8 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_464 ();
 sg13g2_decap_8 FILLER_5_471 ();
 sg13g2_decap_8 FILLER_5_478 ();
 sg13g2_decap_8 FILLER_5_485 ();
 sg13g2_decap_8 FILLER_5_492 ();
 sg13g2_decap_8 FILLER_5_499 ();
 sg13g2_decap_8 FILLER_5_506 ();
 sg13g2_fill_1 FILLER_5_513 ();
 sg13g2_decap_8 FILLER_5_524 ();
 sg13g2_decap_8 FILLER_5_531 ();
 sg13g2_fill_1 FILLER_5_538 ();
 sg13g2_fill_2 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_563 ();
 sg13g2_fill_2 FILLER_5_570 ();
 sg13g2_fill_1 FILLER_5_572 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_fill_1 FILLER_5_594 ();
 sg13g2_decap_4 FILLER_5_608 ();
 sg13g2_fill_2 FILLER_5_612 ();
 sg13g2_decap_8 FILLER_5_619 ();
 sg13g2_decap_8 FILLER_5_626 ();
 sg13g2_fill_2 FILLER_5_633 ();
 sg13g2_fill_1 FILLER_5_635 ();
 sg13g2_decap_4 FILLER_5_656 ();
 sg13g2_fill_2 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_682 ();
 sg13g2_fill_2 FILLER_5_689 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_4 FILLER_5_856 ();
 sg13g2_fill_2 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_30 ();
 sg13g2_fill_1 FILLER_6_37 ();
 sg13g2_fill_1 FILLER_6_51 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_4 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_98 ();
 sg13g2_fill_1 FILLER_6_117 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_189 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_fill_2 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_fill_1 FILLER_6_291 ();
 sg13g2_fill_2 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_311 ();
 sg13g2_decap_4 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_fill_2 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_fill_2 FILLER_6_383 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_fill_2 FILLER_6_413 ();
 sg13g2_fill_1 FILLER_6_415 ();
 sg13g2_fill_1 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_458 ();
 sg13g2_decap_8 FILLER_6_465 ();
 sg13g2_fill_2 FILLER_6_472 ();
 sg13g2_fill_1 FILLER_6_474 ();
 sg13g2_decap_4 FILLER_6_505 ();
 sg13g2_fill_2 FILLER_6_532 ();
 sg13g2_fill_1 FILLER_6_534 ();
 sg13g2_decap_8 FILLER_6_556 ();
 sg13g2_fill_2 FILLER_6_563 ();
 sg13g2_fill_2 FILLER_6_595 ();
 sg13g2_fill_1 FILLER_6_597 ();
 sg13g2_decap_4 FILLER_6_663 ();
 sg13g2_decap_4 FILLER_6_679 ();
 sg13g2_decap_4 FILLER_6_707 ();
 sg13g2_decap_4 FILLER_6_725 ();
 sg13g2_fill_1 FILLER_6_729 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_fill_2 FILLER_6_859 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_20 ();
 sg13g2_decap_8 FILLER_7_30 ();
 sg13g2_decap_4 FILLER_7_37 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_decap_8 FILLER_7_95 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_decap_4 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_131 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_178 ();
 sg13g2_decap_8 FILLER_7_185 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_4 FILLER_7_237 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_259 ();
 sg13g2_fill_2 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_fill_2 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_fill_1 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_2 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_369 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_2 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_7_431 ();
 sg13g2_fill_2 FILLER_7_441 ();
 sg13g2_fill_2 FILLER_7_472 ();
 sg13g2_decap_4 FILLER_7_498 ();
 sg13g2_fill_2 FILLER_7_502 ();
 sg13g2_fill_2 FILLER_7_516 ();
 sg13g2_decap_8 FILLER_7_523 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_fill_1 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_563 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_decap_8 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_600 ();
 sg13g2_fill_2 FILLER_7_607 ();
 sg13g2_fill_2 FILLER_7_614 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_fill_1 FILLER_7_637 ();
 sg13g2_fill_2 FILLER_7_649 ();
 sg13g2_fill_1 FILLER_7_655 ();
 sg13g2_fill_2 FILLER_7_664 ();
 sg13g2_fill_1 FILLER_7_673 ();
 sg13g2_decap_4 FILLER_7_685 ();
 sg13g2_fill_2 FILLER_7_689 ();
 sg13g2_fill_2 FILLER_7_701 ();
 sg13g2_fill_2 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_4 FILLER_7_720 ();
 sg13g2_fill_1 FILLER_7_729 ();
 sg13g2_decap_4 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_decap_8 FILLER_7_758 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_decap_8 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_4 FILLER_7_856 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_22 ();
 sg13g2_decap_8 FILLER_8_27 ();
 sg13g2_fill_1 FILLER_8_34 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_fill_1 FILLER_8_60 ();
 sg13g2_fill_1 FILLER_8_84 ();
 sg13g2_decap_4 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_117 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_4 FILLER_8_228 ();
 sg13g2_fill_2 FILLER_8_232 ();
 sg13g2_fill_2 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_4 FILLER_8_376 ();
 sg13g2_fill_1 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_fill_1 FILLER_8_392 ();
 sg13g2_fill_1 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_fill_2 FILLER_8_433 ();
 sg13g2_decap_8 FILLER_8_443 ();
 sg13g2_fill_2 FILLER_8_450 ();
 sg13g2_decap_8 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_470 ();
 sg13g2_fill_1 FILLER_8_472 ();
 sg13g2_decap_4 FILLER_8_499 ();
 sg13g2_decap_8 FILLER_8_519 ();
 sg13g2_decap_4 FILLER_8_526 ();
 sg13g2_fill_2 FILLER_8_530 ();
 sg13g2_fill_2 FILLER_8_551 ();
 sg13g2_fill_1 FILLER_8_553 ();
 sg13g2_decap_4 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_566 ();
 sg13g2_decap_4 FILLER_8_573 ();
 sg13g2_fill_2 FILLER_8_590 ();
 sg13g2_decap_4 FILLER_8_596 ();
 sg13g2_fill_2 FILLER_8_600 ();
 sg13g2_fill_2 FILLER_8_615 ();
 sg13g2_fill_1 FILLER_8_617 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_fill_2 FILLER_8_637 ();
 sg13g2_fill_1 FILLER_8_639 ();
 sg13g2_fill_2 FILLER_8_655 ();
 sg13g2_fill_1 FILLER_8_657 ();
 sg13g2_decap_4 FILLER_8_662 ();
 sg13g2_fill_1 FILLER_8_666 ();
 sg13g2_decap_4 FILLER_8_679 ();
 sg13g2_fill_2 FILLER_8_683 ();
 sg13g2_fill_1 FILLER_8_698 ();
 sg13g2_decap_4 FILLER_8_740 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_759 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_decap_8 FILLER_8_773 ();
 sg13g2_decap_8 FILLER_8_780 ();
 sg13g2_decap_8 FILLER_8_787 ();
 sg13g2_decap_8 FILLER_8_794 ();
 sg13g2_decap_8 FILLER_8_801 ();
 sg13g2_decap_8 FILLER_8_808 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_822 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_decap_8 FILLER_8_850 ();
 sg13g2_decap_4 FILLER_8_857 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_45 ();
 sg13g2_fill_2 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_fill_2 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_4 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_153 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_256 ();
 sg13g2_decap_4 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_decap_4 FILLER_9_321 ();
 sg13g2_fill_1 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_fill_1 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_fill_1 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_fill_1 FILLER_9_426 ();
 sg13g2_fill_2 FILLER_9_439 ();
 sg13g2_decap_8 FILLER_9_467 ();
 sg13g2_decap_4 FILLER_9_474 ();
 sg13g2_decap_8 FILLER_9_491 ();
 sg13g2_fill_2 FILLER_9_498 ();
 sg13g2_fill_2 FILLER_9_516 ();
 sg13g2_fill_1 FILLER_9_518 ();
 sg13g2_decap_4 FILLER_9_523 ();
 sg13g2_fill_2 FILLER_9_527 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_4 FILLER_9_557 ();
 sg13g2_fill_2 FILLER_9_586 ();
 sg13g2_fill_1 FILLER_9_588 ();
 sg13g2_fill_2 FILLER_9_593 ();
 sg13g2_fill_1 FILLER_9_595 ();
 sg13g2_fill_2 FILLER_9_601 ();
 sg13g2_decap_4 FILLER_9_611 ();
 sg13g2_fill_1 FILLER_9_631 ();
 sg13g2_fill_2 FILLER_9_658 ();
 sg13g2_fill_1 FILLER_9_660 ();
 sg13g2_decap_4 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_fill_1 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_698 ();
 sg13g2_decap_8 FILLER_9_705 ();
 sg13g2_decap_8 FILLER_9_712 ();
 sg13g2_fill_2 FILLER_9_719 ();
 sg13g2_fill_1 FILLER_9_721 ();
 sg13g2_decap_4 FILLER_9_737 ();
 sg13g2_fill_1 FILLER_9_741 ();
 sg13g2_decap_8 FILLER_9_762 ();
 sg13g2_decap_8 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_776 ();
 sg13g2_decap_8 FILLER_9_783 ();
 sg13g2_decap_8 FILLER_9_790 ();
 sg13g2_decap_8 FILLER_9_797 ();
 sg13g2_decap_8 FILLER_9_804 ();
 sg13g2_decap_8 FILLER_9_811 ();
 sg13g2_decap_8 FILLER_9_818 ();
 sg13g2_decap_8 FILLER_9_825 ();
 sg13g2_decap_8 FILLER_9_832 ();
 sg13g2_decap_8 FILLER_9_839 ();
 sg13g2_decap_8 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_853 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_fill_2 FILLER_10_22 ();
 sg13g2_fill_2 FILLER_10_33 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_94 ();
 sg13g2_fill_2 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_150 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_4 FILLER_10_167 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_decap_4 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_fill_1 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_4 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_decap_4 FILLER_10_350 ();
 sg13g2_fill_2 FILLER_10_354 ();
 sg13g2_fill_1 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_fill_1 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_4 FILLER_10_417 ();
 sg13g2_fill_2 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_4 FILLER_10_466 ();
 sg13g2_fill_1 FILLER_10_470 ();
 sg13g2_decap_8 FILLER_10_479 ();
 sg13g2_decap_4 FILLER_10_486 ();
 sg13g2_decap_8 FILLER_10_503 ();
 sg13g2_decap_4 FILLER_10_525 ();
 sg13g2_fill_1 FILLER_10_533 ();
 sg13g2_decap_8 FILLER_10_544 ();
 sg13g2_fill_2 FILLER_10_551 ();
 sg13g2_decap_4 FILLER_10_562 ();
 sg13g2_decap_4 FILLER_10_570 ();
 sg13g2_fill_2 FILLER_10_579 ();
 sg13g2_fill_2 FILLER_10_586 ();
 sg13g2_fill_1 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_597 ();
 sg13g2_fill_1 FILLER_10_604 ();
 sg13g2_decap_8 FILLER_10_626 ();
 sg13g2_decap_4 FILLER_10_633 ();
 sg13g2_fill_1 FILLER_10_637 ();
 sg13g2_fill_1 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_fill_2 FILLER_10_680 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_fill_2 FILLER_10_706 ();
 sg13g2_fill_1 FILLER_10_708 ();
 sg13g2_fill_2 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_32 ();
 sg13g2_fill_1 FILLER_11_34 ();
 sg13g2_decap_8 FILLER_11_38 ();
 sg13g2_decap_4 FILLER_11_45 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_55 ();
 sg13g2_fill_1 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_66 ();
 sg13g2_decap_8 FILLER_11_73 ();
 sg13g2_decap_4 FILLER_11_80 ();
 sg13g2_decap_4 FILLER_11_92 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_4 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_8 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_141 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_4 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_225 ();
 sg13g2_decap_4 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_4 FILLER_11_274 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_decap_4 FILLER_11_283 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_354 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_2 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_410 ();
 sg13g2_fill_2 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_437 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_fill_2 FILLER_11_483 ();
 sg13g2_fill_1 FILLER_11_485 ();
 sg13g2_fill_2 FILLER_11_499 ();
 sg13g2_decap_8 FILLER_11_524 ();
 sg13g2_decap_4 FILLER_11_565 ();
 sg13g2_fill_2 FILLER_11_569 ();
 sg13g2_decap_8 FILLER_11_597 ();
 sg13g2_decap_8 FILLER_11_604 ();
 sg13g2_decap_8 FILLER_11_611 ();
 sg13g2_fill_2 FILLER_11_618 ();
 sg13g2_fill_2 FILLER_11_632 ();
 sg13g2_fill_1 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_652 ();
 sg13g2_fill_1 FILLER_11_659 ();
 sg13g2_fill_2 FILLER_11_684 ();
 sg13g2_decap_4 FILLER_11_707 ();
 sg13g2_fill_1 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_726 ();
 sg13g2_decap_4 FILLER_11_733 ();
 sg13g2_fill_1 FILLER_11_737 ();
 sg13g2_decap_4 FILLER_11_757 ();
 sg13g2_fill_1 FILLER_11_761 ();
 sg13g2_fill_1 FILLER_11_768 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_797 ();
 sg13g2_decap_8 FILLER_11_804 ();
 sg13g2_decap_8 FILLER_11_811 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_8 FILLER_11_825 ();
 sg13g2_decap_8 FILLER_11_832 ();
 sg13g2_decap_8 FILLER_11_839 ();
 sg13g2_decap_8 FILLER_11_846 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_860 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_16 ();
 sg13g2_fill_2 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_fill_2 FILLER_12_33 ();
 sg13g2_decap_8 FILLER_12_59 ();
 sg13g2_decap_4 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_78 ();
 sg13g2_decap_4 FILLER_12_96 ();
 sg13g2_fill_1 FILLER_12_100 ();
 sg13g2_decap_4 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_decap_4 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_decap_4 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_fill_2 FILLER_12_244 ();
 sg13g2_fill_1 FILLER_12_246 ();
 sg13g2_decap_4 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_fill_1 FILLER_12_388 ();
 sg13g2_decap_4 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_fill_1 FILLER_12_421 ();
 sg13g2_decap_4 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_444 ();
 sg13g2_decap_8 FILLER_12_458 ();
 sg13g2_fill_2 FILLER_12_465 ();
 sg13g2_fill_1 FILLER_12_467 ();
 sg13g2_decap_8 FILLER_12_481 ();
 sg13g2_decap_4 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_498 ();
 sg13g2_decap_8 FILLER_12_517 ();
 sg13g2_decap_8 FILLER_12_524 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_4 FILLER_12_550 ();
 sg13g2_decap_4 FILLER_12_562 ();
 sg13g2_decap_4 FILLER_12_578 ();
 sg13g2_fill_1 FILLER_12_582 ();
 sg13g2_decap_8 FILLER_12_604 ();
 sg13g2_fill_2 FILLER_12_611 ();
 sg13g2_decap_4 FILLER_12_629 ();
 sg13g2_fill_2 FILLER_12_633 ();
 sg13g2_fill_2 FILLER_12_640 ();
 sg13g2_fill_1 FILLER_12_642 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_fill_2 FILLER_12_662 ();
 sg13g2_fill_1 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_674 ();
 sg13g2_decap_8 FILLER_12_681 ();
 sg13g2_decap_8 FILLER_12_699 ();
 sg13g2_decap_8 FILLER_12_706 ();
 sg13g2_decap_4 FILLER_12_717 ();
 sg13g2_fill_1 FILLER_12_721 ();
 sg13g2_fill_2 FILLER_12_740 ();
 sg13g2_fill_1 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_748 ();
 sg13g2_fill_2 FILLER_12_755 ();
 sg13g2_fill_2 FILLER_12_778 ();
 sg13g2_decap_8 FILLER_12_801 ();
 sg13g2_decap_8 FILLER_12_808 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_decap_8 FILLER_12_822 ();
 sg13g2_decap_8 FILLER_12_829 ();
 sg13g2_decap_8 FILLER_12_836 ();
 sg13g2_decap_8 FILLER_12_843 ();
 sg13g2_decap_8 FILLER_12_850 ();
 sg13g2_decap_4 FILLER_12_857 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_20 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_decap_4 FILLER_13_53 ();
 sg13g2_fill_2 FILLER_13_57 ();
 sg13g2_decap_4 FILLER_13_80 ();
 sg13g2_fill_2 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_4 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_decap_4 FILLER_13_188 ();
 sg13g2_fill_1 FILLER_13_192 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_239 ();
 sg13g2_fill_2 FILLER_13_253 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_decap_4 FILLER_13_279 ();
 sg13g2_decap_4 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_decap_4 FILLER_13_343 ();
 sg13g2_decap_4 FILLER_13_359 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_393 ();
 sg13g2_fill_1 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_422 ();
 sg13g2_decap_4 FILLER_13_455 ();
 sg13g2_fill_2 FILLER_13_459 ();
 sg13g2_decap_4 FILLER_13_477 ();
 sg13g2_fill_1 FILLER_13_481 ();
 sg13g2_fill_2 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_514 ();
 sg13g2_fill_2 FILLER_13_521 ();
 sg13g2_decap_8 FILLER_13_541 ();
 sg13g2_decap_4 FILLER_13_548 ();
 sg13g2_fill_1 FILLER_13_552 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_4 FILLER_13_586 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_633 ();
 sg13g2_fill_2 FILLER_13_640 ();
 sg13g2_decap_8 FILLER_13_654 ();
 sg13g2_fill_1 FILLER_13_661 ();
 sg13g2_fill_1 FILLER_13_704 ();
 sg13g2_fill_2 FILLER_13_719 ();
 sg13g2_fill_1 FILLER_13_721 ();
 sg13g2_fill_2 FILLER_13_727 ();
 sg13g2_fill_2 FILLER_13_746 ();
 sg13g2_fill_1 FILLER_13_748 ();
 sg13g2_decap_4 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_773 ();
 sg13g2_fill_2 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_825 ();
 sg13g2_decap_8 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_846 ();
 sg13g2_decap_8 FILLER_13_853 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_15 ();
 sg13g2_fill_2 FILLER_14_22 ();
 sg13g2_fill_1 FILLER_14_24 ();
 sg13g2_decap_8 FILLER_14_30 ();
 sg13g2_decap_8 FILLER_14_37 ();
 sg13g2_decap_4 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_99 ();
 sg13g2_decap_4 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_127 ();
 sg13g2_decap_4 FILLER_14_157 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_232 ();
 sg13g2_decap_4 FILLER_14_242 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_decap_4 FILLER_14_261 ();
 sg13g2_fill_2 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_4 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_334 ();
 sg13g2_decap_4 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_373 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_fill_2 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_4 FILLER_14_430 ();
 sg13g2_fill_2 FILLER_14_434 ();
 sg13g2_fill_1 FILLER_14_439 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_fill_2 FILLER_14_452 ();
 sg13g2_fill_1 FILLER_14_454 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_fill_1 FILLER_14_478 ();
 sg13g2_decap_4 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_4 FILLER_14_504 ();
 sg13g2_fill_2 FILLER_14_508 ();
 sg13g2_decap_4 FILLER_14_523 ();
 sg13g2_fill_2 FILLER_14_539 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_fill_2 FILLER_14_551 ();
 sg13g2_decap_4 FILLER_14_558 ();
 sg13g2_fill_2 FILLER_14_562 ();
 sg13g2_decap_4 FILLER_14_577 ();
 sg13g2_fill_1 FILLER_14_581 ();
 sg13g2_decap_4 FILLER_14_600 ();
 sg13g2_fill_2 FILLER_14_604 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_634 ();
 sg13g2_decap_4 FILLER_14_641 ();
 sg13g2_fill_2 FILLER_14_662 ();
 sg13g2_fill_1 FILLER_14_664 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_fill_2 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_fill_2 FILLER_14_710 ();
 sg13g2_decap_4 FILLER_14_725 ();
 sg13g2_decap_4 FILLER_14_746 ();
 sg13g2_decap_4 FILLER_14_757 ();
 sg13g2_fill_1 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_771 ();
 sg13g2_decap_8 FILLER_14_778 ();
 sg13g2_fill_1 FILLER_14_785 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_fill_2 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_4 FILLER_14_856 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_24 ();
 sg13g2_decap_8 FILLER_15_51 ();
 sg13g2_decap_4 FILLER_15_58 ();
 sg13g2_fill_1 FILLER_15_62 ();
 sg13g2_decap_4 FILLER_15_81 ();
 sg13g2_decap_4 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_fill_2 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_4 FILLER_15_156 ();
 sg13g2_fill_1 FILLER_15_160 ();
 sg13g2_decap_4 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_4 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_fill_2 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_decap_4 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_fill_1 FILLER_15_389 ();
 sg13g2_fill_1 FILLER_15_398 ();
 sg13g2_fill_2 FILLER_15_430 ();
 sg13g2_fill_1 FILLER_15_440 ();
 sg13g2_decap_8 FILLER_15_449 ();
 sg13g2_decap_4 FILLER_15_456 ();
 sg13g2_fill_2 FILLER_15_460 ();
 sg13g2_fill_2 FILLER_15_475 ();
 sg13g2_decap_4 FILLER_15_503 ();
 sg13g2_decap_4 FILLER_15_528 ();
 sg13g2_fill_1 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_fill_2 FILLER_15_606 ();
 sg13g2_fill_1 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_624 ();
 sg13g2_decap_8 FILLER_15_631 ();
 sg13g2_fill_2 FILLER_15_638 ();
 sg13g2_decap_4 FILLER_15_661 ();
 sg13g2_fill_2 FILLER_15_665 ();
 sg13g2_decap_4 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_684 ();
 sg13g2_fill_1 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_fill_1 FILLER_15_717 ();
 sg13g2_decap_4 FILLER_15_722 ();
 sg13g2_fill_1 FILLER_15_726 ();
 sg13g2_fill_1 FILLER_15_744 ();
 sg13g2_fill_2 FILLER_15_757 ();
 sg13g2_fill_1 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_fill_1 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_832 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_846 ();
 sg13g2_decap_8 FILLER_15_853 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_57 ();
 sg13g2_decap_4 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_decap_8 FILLER_16_73 ();
 sg13g2_decap_8 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_87 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_1 FILLER_16_117 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_211 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_256 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_2 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_fill_2 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_4 FILLER_16_435 ();
 sg13g2_fill_1 FILLER_16_444 ();
 sg13g2_fill_1 FILLER_16_458 ();
 sg13g2_decap_8 FILLER_16_472 ();
 sg13g2_decap_8 FILLER_16_479 ();
 sg13g2_decap_4 FILLER_16_486 ();
 sg13g2_decap_4 FILLER_16_523 ();
 sg13g2_fill_2 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_547 ();
 sg13g2_decap_8 FILLER_16_554 ();
 sg13g2_fill_2 FILLER_16_561 ();
 sg13g2_decap_4 FILLER_16_576 ();
 sg13g2_fill_1 FILLER_16_580 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_4 FILLER_16_602 ();
 sg13g2_fill_1 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_631 ();
 sg13g2_decap_8 FILLER_16_638 ();
 sg13g2_decap_4 FILLER_16_657 ();
 sg13g2_fill_1 FILLER_16_661 ();
 sg13g2_decap_4 FILLER_16_676 ();
 sg13g2_fill_1 FILLER_16_706 ();
 sg13g2_fill_1 FILLER_16_720 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_fill_2 FILLER_16_754 ();
 sg13g2_fill_1 FILLER_16_756 ();
 sg13g2_decap_4 FILLER_16_762 ();
 sg13g2_fill_2 FILLER_16_771 ();
 sg13g2_fill_2 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_784 ();
 sg13g2_fill_1 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_4 FILLER_16_798 ();
 sg13g2_fill_2 FILLER_16_802 ();
 sg13g2_fill_2 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_9 ();
 sg13g2_fill_2 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_19 ();
 sg13g2_decap_4 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_48 ();
 sg13g2_fill_2 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_decap_4 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_127 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_decap_8 FILLER_17_148 ();
 sg13g2_decap_4 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_decap_4 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_decap_4 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_decap_4 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_295 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_decap_4 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_decap_4 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_4 FILLER_17_421 ();
 sg13g2_decap_8 FILLER_17_446 ();
 sg13g2_decap_4 FILLER_17_453 ();
 sg13g2_fill_2 FILLER_17_457 ();
 sg13g2_decap_8 FILLER_17_471 ();
 sg13g2_decap_8 FILLER_17_478 ();
 sg13g2_decap_4 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_489 ();
 sg13g2_fill_2 FILLER_17_508 ();
 sg13g2_fill_1 FILLER_17_510 ();
 sg13g2_decap_4 FILLER_17_523 ();
 sg13g2_fill_2 FILLER_17_527 ();
 sg13g2_fill_2 FILLER_17_541 ();
 sg13g2_fill_1 FILLER_17_543 ();
 sg13g2_decap_4 FILLER_17_552 ();
 sg13g2_fill_2 FILLER_17_581 ();
 sg13g2_fill_2 FILLER_17_591 ();
 sg13g2_decap_8 FILLER_17_601 ();
 sg13g2_fill_2 FILLER_17_625 ();
 sg13g2_fill_2 FILLER_17_635 ();
 sg13g2_fill_2 FILLER_17_657 ();
 sg13g2_decap_4 FILLER_17_683 ();
 sg13g2_fill_2 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_701 ();
 sg13g2_fill_2 FILLER_17_712 ();
 sg13g2_fill_1 FILLER_17_714 ();
 sg13g2_fill_1 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_4 FILLER_17_739 ();
 sg13g2_fill_2 FILLER_17_743 ();
 sg13g2_fill_1 FILLER_17_772 ();
 sg13g2_decap_4 FILLER_17_793 ();
 sg13g2_fill_2 FILLER_17_797 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_846 ();
 sg13g2_decap_8 FILLER_17_853 ();
 sg13g2_fill_2 FILLER_17_860 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_69 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_decap_4 FILLER_18_101 ();
 sg13g2_decap_4 FILLER_18_113 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_283 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_decap_4 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_4 FILLER_18_422 ();
 sg13g2_fill_2 FILLER_18_438 ();
 sg13g2_fill_1 FILLER_18_440 ();
 sg13g2_decap_8 FILLER_18_449 ();
 sg13g2_decap_4 FILLER_18_456 ();
 sg13g2_fill_2 FILLER_18_472 ();
 sg13g2_decap_4 FILLER_18_482 ();
 sg13g2_fill_2 FILLER_18_486 ();
 sg13g2_decap_8 FILLER_18_496 ();
 sg13g2_decap_4 FILLER_18_503 ();
 sg13g2_fill_2 FILLER_18_507 ();
 sg13g2_decap_4 FILLER_18_526 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_fill_2 FILLER_18_560 ();
 sg13g2_fill_2 FILLER_18_575 ();
 sg13g2_decap_8 FILLER_18_582 ();
 sg13g2_fill_1 FILLER_18_589 ();
 sg13g2_decap_8 FILLER_18_603 ();
 sg13g2_fill_2 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_fill_1 FILLER_18_639 ();
 sg13g2_decap_4 FILLER_18_657 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_fill_2 FILLER_18_689 ();
 sg13g2_fill_2 FILLER_18_707 ();
 sg13g2_fill_1 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_734 ();
 sg13g2_fill_2 FILLER_18_741 ();
 sg13g2_fill_1 FILLER_18_743 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_fill_2 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_fill_2 FILLER_18_799 ();
 sg13g2_fill_1 FILLER_18_801 ();
 sg13g2_decap_4 FILLER_18_807 ();
 sg13g2_fill_1 FILLER_18_811 ();
 sg13g2_fill_1 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_fill_2 FILLER_18_859 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_31 ();
 sg13g2_decap_4 FILLER_19_50 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_127 ();
 sg13g2_decap_4 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_decap_4 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_2 FILLER_19_391 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_419 ();
 sg13g2_fill_1 FILLER_19_421 ();
 sg13g2_decap_4 FILLER_19_444 ();
 sg13g2_fill_2 FILLER_19_448 ();
 sg13g2_fill_2 FILLER_19_463 ();
 sg13g2_fill_1 FILLER_19_465 ();
 sg13g2_decap_8 FILLER_19_502 ();
 sg13g2_fill_1 FILLER_19_509 ();
 sg13g2_fill_2 FILLER_19_523 ();
 sg13g2_fill_1 FILLER_19_525 ();
 sg13g2_decap_4 FILLER_19_531 ();
 sg13g2_fill_1 FILLER_19_535 ();
 sg13g2_decap_4 FILLER_19_553 ();
 sg13g2_fill_2 FILLER_19_580 ();
 sg13g2_fill_1 FILLER_19_582 ();
 sg13g2_decap_4 FILLER_19_591 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_4 FILLER_19_630 ();
 sg13g2_fill_1 FILLER_19_634 ();
 sg13g2_fill_2 FILLER_19_656 ();
 sg13g2_fill_1 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_4 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_4 FILLER_19_720 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_fill_2 FILLER_19_738 ();
 sg13g2_fill_1 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_765 ();
 sg13g2_fill_2 FILLER_19_772 ();
 sg13g2_fill_1 FILLER_19_774 ();
 sg13g2_fill_2 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_790 ();
 sg13g2_decap_4 FILLER_19_803 ();
 sg13g2_fill_1 FILLER_19_807 ();
 sg13g2_decap_4 FILLER_19_821 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_fill_2 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_859 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_8 FILLER_20_31 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_decap_8 FILLER_20_97 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_decap_4 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_decap_8 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_4 FILLER_20_365 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_4 FILLER_20_393 ();
 sg13g2_fill_2 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_4 FILLER_20_450 ();
 sg13g2_fill_2 FILLER_20_454 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_fill_2 FILLER_20_518 ();
 sg13g2_decap_4 FILLER_20_535 ();
 sg13g2_fill_1 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_fill_2 FILLER_20_566 ();
 sg13g2_fill_2 FILLER_20_578 ();
 sg13g2_fill_1 FILLER_20_580 ();
 sg13g2_fill_2 FILLER_20_598 ();
 sg13g2_fill_1 FILLER_20_609 ();
 sg13g2_decap_4 FILLER_20_615 ();
 sg13g2_fill_1 FILLER_20_619 ();
 sg13g2_decap_8 FILLER_20_625 ();
 sg13g2_decap_8 FILLER_20_632 ();
 sg13g2_decap_4 FILLER_20_649 ();
 sg13g2_fill_2 FILLER_20_653 ();
 sg13g2_decap_4 FILLER_20_659 ();
 sg13g2_fill_2 FILLER_20_663 ();
 sg13g2_fill_2 FILLER_20_690 ();
 sg13g2_decap_4 FILLER_20_705 ();
 sg13g2_fill_1 FILLER_20_719 ();
 sg13g2_decap_4 FILLER_20_741 ();
 sg13g2_fill_2 FILLER_20_745 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_795 ();
 sg13g2_fill_2 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_4 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_8 FILLER_21_44 ();
 sg13g2_decap_4 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_118 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_decap_4 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_4 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_364 ();
 sg13g2_decap_4 FILLER_21_390 ();
 sg13g2_fill_1 FILLER_21_394 ();
 sg13g2_decap_4 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_425 ();
 sg13g2_decap_4 FILLER_21_453 ();
 sg13g2_fill_1 FILLER_21_457 ();
 sg13g2_fill_2 FILLER_21_472 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_4 FILLER_21_494 ();
 sg13g2_fill_1 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_516 ();
 sg13g2_decap_8 FILLER_21_526 ();
 sg13g2_decap_4 FILLER_21_533 ();
 sg13g2_decap_4 FILLER_21_550 ();
 sg13g2_fill_1 FILLER_21_554 ();
 sg13g2_decap_4 FILLER_21_559 ();
 sg13g2_fill_1 FILLER_21_563 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_592 ();
 sg13g2_fill_1 FILLER_21_599 ();
 sg13g2_fill_1 FILLER_21_636 ();
 sg13g2_decap_4 FILLER_21_653 ();
 sg13g2_fill_2 FILLER_21_657 ();
 sg13g2_decap_4 FILLER_21_664 ();
 sg13g2_decap_4 FILLER_21_692 ();
 sg13g2_fill_1 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_fill_2 FILLER_21_740 ();
 sg13g2_decap_4 FILLER_21_747 ();
 sg13g2_fill_2 FILLER_21_751 ();
 sg13g2_decap_4 FILLER_21_758 ();
 sg13g2_decap_8 FILLER_21_767 ();
 sg13g2_fill_2 FILLER_21_790 ();
 sg13g2_fill_1 FILLER_21_792 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_fill_2 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_decap_4 FILLER_21_837 ();
 sg13g2_decap_4 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_4 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_4 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_fill_1 FILLER_22_404 ();
 sg13g2_decap_4 FILLER_22_410 ();
 sg13g2_fill_1 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_426 ();
 sg13g2_decap_4 FILLER_22_433 ();
 sg13g2_fill_1 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_447 ();
 sg13g2_decap_8 FILLER_22_454 ();
 sg13g2_fill_1 FILLER_22_480 ();
 sg13g2_decap_4 FILLER_22_489 ();
 sg13g2_fill_1 FILLER_22_493 ();
 sg13g2_fill_2 FILLER_22_512 ();
 sg13g2_decap_8 FILLER_22_527 ();
 sg13g2_fill_1 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_fill_1 FILLER_22_560 ();
 sg13g2_fill_1 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_decap_8 FILLER_22_587 ();
 sg13g2_decap_8 FILLER_22_594 ();
 sg13g2_decap_4 FILLER_22_601 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_fill_2 FILLER_22_618 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_4 FILLER_22_632 ();
 sg13g2_fill_1 FILLER_22_636 ();
 sg13g2_decap_4 FILLER_22_650 ();
 sg13g2_fill_1 FILLER_22_654 ();
 sg13g2_fill_1 FILLER_22_661 ();
 sg13g2_fill_1 FILLER_22_667 ();
 sg13g2_fill_1 FILLER_22_673 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_4 FILLER_22_693 ();
 sg13g2_fill_2 FILLER_22_710 ();
 sg13g2_fill_1 FILLER_22_717 ();
 sg13g2_decap_4 FILLER_22_728 ();
 sg13g2_fill_2 FILLER_22_732 ();
 sg13g2_decap_4 FILLER_22_757 ();
 sg13g2_fill_1 FILLER_22_761 ();
 sg13g2_decap_4 FILLER_22_785 ();
 sg13g2_fill_1 FILLER_22_789 ();
 sg13g2_fill_2 FILLER_22_811 ();
 sg13g2_fill_1 FILLER_22_813 ();
 sg13g2_decap_8 FILLER_22_832 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_decap_8 FILLER_23_61 ();
 sg13g2_decap_8 FILLER_23_68 ();
 sg13g2_fill_2 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_4 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_decap_4 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_4 FILLER_23_319 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_decap_4 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_333 ();
 sg13g2_decap_4 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_4 FILLER_23_402 ();
 sg13g2_fill_2 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_428 ();
 sg13g2_fill_1 FILLER_23_435 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_fill_2 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_fill_2 FILLER_23_483 ();
 sg13g2_fill_2 FILLER_23_514 ();
 sg13g2_fill_1 FILLER_23_520 ();
 sg13g2_decap_4 FILLER_23_526 ();
 sg13g2_fill_2 FILLER_23_530 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_fill_1 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_decap_4 FILLER_23_611 ();
 sg13g2_fill_1 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_4 FILLER_23_637 ();
 sg13g2_fill_2 FILLER_23_655 ();
 sg13g2_fill_2 FILLER_23_667 ();
 sg13g2_fill_1 FILLER_23_669 ();
 sg13g2_decap_4 FILLER_23_685 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_fill_2 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_734 ();
 sg13g2_decap_4 FILLER_23_741 ();
 sg13g2_fill_2 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_773 ();
 sg13g2_fill_1 FILLER_23_780 ();
 sg13g2_fill_2 FILLER_23_789 ();
 sg13g2_fill_1 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_fill_2 FILLER_23_814 ();
 sg13g2_fill_1 FILLER_23_816 ();
 sg13g2_decap_4 FILLER_23_830 ();
 sg13g2_fill_2 FILLER_23_834 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_130 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_decap_8 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_4 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_fill_2 FILLER_24_361 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_403 ();
 sg13g2_fill_1 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_432 ();
 sg13g2_decap_4 FILLER_24_458 ();
 sg13g2_fill_1 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_488 ();
 sg13g2_decap_4 FILLER_24_495 ();
 sg13g2_fill_2 FILLER_24_499 ();
 sg13g2_fill_2 FILLER_24_509 ();
 sg13g2_fill_1 FILLER_24_511 ();
 sg13g2_decap_4 FILLER_24_532 ();
 sg13g2_fill_2 FILLER_24_536 ();
 sg13g2_fill_1 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_566 ();
 sg13g2_decap_4 FILLER_24_588 ();
 sg13g2_fill_1 FILLER_24_592 ();
 sg13g2_fill_2 FILLER_24_608 ();
 sg13g2_fill_1 FILLER_24_610 ();
 sg13g2_fill_2 FILLER_24_624 ();
 sg13g2_fill_1 FILLER_24_626 ();
 sg13g2_decap_4 FILLER_24_653 ();
 sg13g2_fill_2 FILLER_24_657 ();
 sg13g2_decap_8 FILLER_24_663 ();
 sg13g2_fill_2 FILLER_24_670 ();
 sg13g2_decap_4 FILLER_24_677 ();
 sg13g2_fill_2 FILLER_24_681 ();
 sg13g2_decap_4 FILLER_24_697 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_decap_4 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_4 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_fill_1 FILLER_24_789 ();
 sg13g2_fill_1 FILLER_24_794 ();
 sg13g2_decap_4 FILLER_24_803 ();
 sg13g2_fill_2 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_fill_2 FILLER_24_840 ();
 sg13g2_fill_1 FILLER_24_842 ();
 sg13g2_decap_4 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_48 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_decap_4 FILLER_25_76 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_decap_4 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_4 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_4 FILLER_25_390 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_fill_1 FILLER_25_427 ();
 sg13g2_decap_4 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_449 ();
 sg13g2_decap_4 FILLER_25_456 ();
 sg13g2_fill_1 FILLER_25_460 ();
 sg13g2_decap_8 FILLER_25_481 ();
 sg13g2_decap_4 FILLER_25_488 ();
 sg13g2_fill_2 FILLER_25_514 ();
 sg13g2_fill_1 FILLER_25_521 ();
 sg13g2_decap_4 FILLER_25_526 ();
 sg13g2_fill_2 FILLER_25_530 ();
 sg13g2_decap_8 FILLER_25_537 ();
 sg13g2_decap_4 FILLER_25_544 ();
 sg13g2_fill_2 FILLER_25_556 ();
 sg13g2_fill_1 FILLER_25_558 ();
 sg13g2_decap_8 FILLER_25_563 ();
 sg13g2_fill_2 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_580 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_fill_2 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_600 ();
 sg13g2_fill_1 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_decap_4 FILLER_25_655 ();
 sg13g2_fill_1 FILLER_25_659 ();
 sg13g2_fill_1 FILLER_25_689 ();
 sg13g2_fill_1 FILLER_25_707 ();
 sg13g2_decap_4 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_fill_2 FILLER_25_735 ();
 sg13g2_fill_2 FILLER_25_750 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_fill_1 FILLER_25_763 ();
 sg13g2_fill_2 FILLER_25_774 ();
 sg13g2_decap_4 FILLER_25_780 ();
 sg13g2_fill_1 FILLER_25_784 ();
 sg13g2_decap_4 FILLER_25_803 ();
 sg13g2_decap_4 FILLER_25_819 ();
 sg13g2_fill_1 FILLER_25_823 ();
 sg13g2_fill_2 FILLER_25_836 ();
 sg13g2_decap_4 FILLER_25_841 ();
 sg13g2_fill_1 FILLER_25_845 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_decap_8 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_72 ();
 sg13g2_decap_8 FILLER_26_79 ();
 sg13g2_fill_2 FILLER_26_90 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_105 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_4 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_4 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_370 ();
 sg13g2_decap_4 FILLER_26_415 ();
 sg13g2_fill_2 FILLER_26_419 ();
 sg13g2_fill_2 FILLER_26_429 ();
 sg13g2_fill_1 FILLER_26_441 ();
 sg13g2_decap_4 FILLER_26_462 ();
 sg13g2_fill_1 FILLER_26_466 ();
 sg13g2_decap_8 FILLER_26_475 ();
 sg13g2_decap_4 FILLER_26_482 ();
 sg13g2_fill_2 FILLER_26_486 ();
 sg13g2_fill_1 FILLER_26_493 ();
 sg13g2_decap_8 FILLER_26_502 ();
 sg13g2_decap_8 FILLER_26_509 ();
 sg13g2_decap_8 FILLER_26_516 ();
 sg13g2_fill_1 FILLER_26_523 ();
 sg13g2_fill_2 FILLER_26_547 ();
 sg13g2_fill_2 FILLER_26_557 ();
 sg13g2_fill_1 FILLER_26_559 ();
 sg13g2_fill_2 FILLER_26_580 ();
 sg13g2_fill_2 FILLER_26_612 ();
 sg13g2_decap_4 FILLER_26_622 ();
 sg13g2_fill_2 FILLER_26_632 ();
 sg13g2_fill_1 FILLER_26_634 ();
 sg13g2_decap_8 FILLER_26_648 ();
 sg13g2_decap_4 FILLER_26_655 ();
 sg13g2_fill_1 FILLER_26_659 ();
 sg13g2_decap_4 FILLER_26_664 ();
 sg13g2_fill_1 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_fill_1 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_fill_2 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_fill_1 FILLER_26_747 ();
 sg13g2_fill_1 FILLER_26_760 ();
 sg13g2_fill_2 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_fill_2 FILLER_26_779 ();
 sg13g2_fill_1 FILLER_26_781 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_fill_1 FILLER_26_804 ();
 sg13g2_decap_4 FILLER_26_821 ();
 sg13g2_fill_2 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_decap_4 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_4 FILLER_27_158 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_4 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_4 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_398 ();
 sg13g2_fill_2 FILLER_27_412 ();
 sg13g2_fill_1 FILLER_27_414 ();
 sg13g2_decap_4 FILLER_27_440 ();
 sg13g2_fill_1 FILLER_27_444 ();
 sg13g2_decap_8 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_457 ();
 sg13g2_fill_1 FILLER_27_463 ();
 sg13g2_decap_4 FILLER_27_477 ();
 sg13g2_fill_2 FILLER_27_481 ();
 sg13g2_fill_1 FILLER_27_503 ();
 sg13g2_decap_4 FILLER_27_508 ();
 sg13g2_fill_2 FILLER_27_512 ();
 sg13g2_decap_4 FILLER_27_527 ();
 sg13g2_fill_1 FILLER_27_544 ();
 sg13g2_fill_2 FILLER_27_559 ();
 sg13g2_fill_2 FILLER_27_569 ();
 sg13g2_fill_1 FILLER_27_576 ();
 sg13g2_fill_2 FILLER_27_581 ();
 sg13g2_decap_4 FILLER_27_591 ();
 sg13g2_fill_1 FILLER_27_595 ();
 sg13g2_fill_2 FILLER_27_613 ();
 sg13g2_fill_1 FILLER_27_615 ();
 sg13g2_fill_2 FILLER_27_624 ();
 sg13g2_fill_1 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_636 ();
 sg13g2_fill_2 FILLER_27_645 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_decap_8 FILLER_27_652 ();
 sg13g2_fill_2 FILLER_27_659 ();
 sg13g2_decap_4 FILLER_27_678 ();
 sg13g2_fill_2 FILLER_27_682 ();
 sg13g2_fill_2 FILLER_27_711 ();
 sg13g2_fill_1 FILLER_27_713 ();
 sg13g2_decap_4 FILLER_27_738 ();
 sg13g2_decap_8 FILLER_27_773 ();
 sg13g2_fill_1 FILLER_27_780 ();
 sg13g2_decap_4 FILLER_27_794 ();
 sg13g2_decap_4 FILLER_27_803 ();
 sg13g2_fill_1 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_4 FILLER_27_833 ();
 sg13g2_fill_1 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_62 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_404 ();
 sg13g2_fill_2 FILLER_28_411 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_fill_2 FILLER_28_425 ();
 sg13g2_decap_4 FILLER_28_438 ();
 sg13g2_fill_2 FILLER_28_442 ();
 sg13g2_fill_2 FILLER_28_450 ();
 sg13g2_fill_1 FILLER_28_452 ();
 sg13g2_fill_1 FILLER_28_466 ();
 sg13g2_decap_4 FILLER_28_472 ();
 sg13g2_fill_2 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_4 FILLER_28_494 ();
 sg13g2_decap_4 FILLER_28_515 ();
 sg13g2_decap_4 FILLER_28_530 ();
 sg13g2_fill_2 FILLER_28_546 ();
 sg13g2_fill_1 FILLER_28_565 ();
 sg13g2_decap_8 FILLER_28_582 ();
 sg13g2_decap_8 FILLER_28_598 ();
 sg13g2_fill_1 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_663 ();
 sg13g2_decap_4 FILLER_28_710 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_fill_2 FILLER_28_741 ();
 sg13g2_fill_1 FILLER_28_743 ();
 sg13g2_fill_1 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_766 ();
 sg13g2_decap_8 FILLER_28_773 ();
 sg13g2_decap_4 FILLER_28_780 ();
 sg13g2_fill_1 FILLER_28_784 ();
 sg13g2_fill_2 FILLER_28_790 ();
 sg13g2_fill_1 FILLER_28_792 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_fill_1 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_4 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_24 ();
 sg13g2_decap_4 FILLER_29_31 ();
 sg13g2_decap_4 FILLER_29_40 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_80 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_99 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_decap_8 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_131 ();
 sg13g2_decap_4 FILLER_29_138 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_396 ();
 sg13g2_fill_2 FILLER_29_414 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_4 FILLER_29_438 ();
 sg13g2_fill_1 FILLER_29_442 ();
 sg13g2_fill_1 FILLER_29_493 ();
 sg13g2_fill_2 FILLER_29_515 ();
 sg13g2_fill_2 FILLER_29_547 ();
 sg13g2_fill_1 FILLER_29_549 ();
 sg13g2_fill_2 FILLER_29_563 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_fill_2 FILLER_29_592 ();
 sg13g2_decap_4 FILLER_29_598 ();
 sg13g2_fill_1 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_618 ();
 sg13g2_decap_8 FILLER_29_625 ();
 sg13g2_decap_4 FILLER_29_632 ();
 sg13g2_fill_2 FILLER_29_649 ();
 sg13g2_decap_8 FILLER_29_668 ();
 sg13g2_decap_4 FILLER_29_675 ();
 sg13g2_fill_1 FILLER_29_696 ();
 sg13g2_decap_4 FILLER_29_701 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_fill_1 FILLER_29_731 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_753 ();
 sg13g2_fill_2 FILLER_29_766 ();
 sg13g2_fill_1 FILLER_29_768 ();
 sg13g2_decap_4 FILLER_29_777 ();
 sg13g2_fill_1 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_fill_2 FILLER_29_797 ();
 sg13g2_decap_4 FILLER_29_812 ();
 sg13g2_fill_2 FILLER_29_816 ();
 sg13g2_fill_1 FILLER_29_826 ();
 sg13g2_fill_2 FILLER_29_843 ();
 sg13g2_fill_1 FILLER_29_845 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_4 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_decap_4 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_8 FILLER_30_337 ();
 sg13g2_decap_4 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_401 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_decap_4 FILLER_30_418 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_decap_8 FILLER_30_440 ();
 sg13g2_decap_8 FILLER_30_464 ();
 sg13g2_fill_1 FILLER_30_471 ();
 sg13g2_fill_1 FILLER_30_506 ();
 sg13g2_decap_4 FILLER_30_511 ();
 sg13g2_fill_1 FILLER_30_515 ();
 sg13g2_fill_2 FILLER_30_529 ();
 sg13g2_decap_8 FILLER_30_544 ();
 sg13g2_fill_1 FILLER_30_551 ();
 sg13g2_decap_8 FILLER_30_572 ();
 sg13g2_fill_1 FILLER_30_579 ();
 sg13g2_fill_2 FILLER_30_621 ();
 sg13g2_fill_2 FILLER_30_646 ();
 sg13g2_fill_1 FILLER_30_674 ();
 sg13g2_fill_2 FILLER_30_706 ();
 sg13g2_fill_1 FILLER_30_708 ();
 sg13g2_decap_8 FILLER_30_717 ();
 sg13g2_fill_1 FILLER_30_724 ();
 sg13g2_decap_8 FILLER_30_747 ();
 sg13g2_fill_2 FILLER_30_754 ();
 sg13g2_fill_1 FILLER_30_756 ();
 sg13g2_fill_1 FILLER_30_761 ();
 sg13g2_decap_8 FILLER_30_782 ();
 sg13g2_fill_2 FILLER_30_789 ();
 sg13g2_decap_8 FILLER_30_811 ();
 sg13g2_fill_2 FILLER_30_818 ();
 sg13g2_fill_1 FILLER_30_825 ();
 sg13g2_fill_2 FILLER_30_834 ();
 sg13g2_decap_4 FILLER_30_844 ();
 sg13g2_fill_1 FILLER_30_848 ();
 sg13g2_fill_2 FILLER_30_859 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_decap_4 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_33 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_decap_4 FILLER_31_59 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_decap_4 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_114 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_decap_4 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_4 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_decap_4 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_fill_1 FILLER_31_426 ();
 sg13g2_decap_4 FILLER_31_431 ();
 sg13g2_fill_1 FILLER_31_435 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_fill_2 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_464 ();
 sg13g2_fill_2 FILLER_31_481 ();
 sg13g2_fill_2 FILLER_31_496 ();
 sg13g2_fill_1 FILLER_31_498 ();
 sg13g2_fill_2 FILLER_31_525 ();
 sg13g2_decap_4 FILLER_31_551 ();
 sg13g2_fill_1 FILLER_31_555 ();
 sg13g2_fill_2 FILLER_31_583 ();
 sg13g2_fill_1 FILLER_31_585 ();
 sg13g2_decap_4 FILLER_31_603 ();
 sg13g2_fill_1 FILLER_31_607 ();
 sg13g2_fill_2 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_627 ();
 sg13g2_decap_8 FILLER_31_632 ();
 sg13g2_fill_1 FILLER_31_639 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_4 FILLER_31_673 ();
 sg13g2_fill_1 FILLER_31_677 ();
 sg13g2_fill_1 FILLER_31_712 ();
 sg13g2_decap_4 FILLER_31_721 ();
 sg13g2_fill_2 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_751 ();
 sg13g2_decap_4 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_4 FILLER_31_786 ();
 sg13g2_fill_2 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_fill_2 FILLER_31_818 ();
 sg13g2_fill_1 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_824 ();
 sg13g2_decap_4 FILLER_31_836 ();
 sg13g2_fill_1 FILLER_31_840 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_31 ();
 sg13g2_fill_2 FILLER_32_38 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_decap_4 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_99 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_decap_4 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_4 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_294 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_361 ();
 sg13g2_fill_2 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_32_447 ();
 sg13g2_fill_2 FILLER_32_467 ();
 sg13g2_decap_8 FILLER_32_482 ();
 sg13g2_fill_2 FILLER_32_489 ();
 sg13g2_decap_4 FILLER_32_504 ();
 sg13g2_fill_1 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_fill_1 FILLER_32_532 ();
 sg13g2_fill_2 FILLER_32_554 ();
 sg13g2_fill_1 FILLER_32_587 ();
 sg13g2_decap_8 FILLER_32_593 ();
 sg13g2_fill_2 FILLER_32_600 ();
 sg13g2_fill_2 FILLER_32_619 ();
 sg13g2_fill_1 FILLER_32_621 ();
 sg13g2_decap_8 FILLER_32_627 ();
 sg13g2_fill_2 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_fill_2 FILLER_32_675 ();
 sg13g2_fill_1 FILLER_32_677 ();
 sg13g2_decap_4 FILLER_32_691 ();
 sg13g2_fill_1 FILLER_32_695 ();
 sg13g2_fill_2 FILLER_32_700 ();
 sg13g2_fill_1 FILLER_32_702 ();
 sg13g2_decap_4 FILLER_32_734 ();
 sg13g2_decap_4 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_772 ();
 sg13g2_fill_2 FILLER_32_779 ();
 sg13g2_fill_1 FILLER_32_798 ();
 sg13g2_fill_2 FILLER_32_807 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_827 ();
 sg13g2_fill_1 FILLER_32_834 ();
 sg13g2_decap_4 FILLER_32_839 ();
 sg13g2_fill_2 FILLER_32_843 ();
 sg13g2_decap_4 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_61 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_decap_4 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_33_435 ();
 sg13g2_fill_1 FILLER_33_437 ();
 sg13g2_fill_2 FILLER_33_447 ();
 sg13g2_decap_4 FILLER_33_452 ();
 sg13g2_decap_4 FILLER_33_478 ();
 sg13g2_fill_2 FILLER_33_482 ();
 sg13g2_fill_1 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_536 ();
 sg13g2_fill_1 FILLER_33_538 ();
 sg13g2_decap_8 FILLER_33_556 ();
 sg13g2_fill_1 FILLER_33_563 ();
 sg13g2_decap_8 FILLER_33_573 ();
 sg13g2_fill_2 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_592 ();
 sg13g2_decap_4 FILLER_33_607 ();
 sg13g2_fill_1 FILLER_33_611 ();
 sg13g2_fill_2 FILLER_33_616 ();
 sg13g2_fill_1 FILLER_33_618 ();
 sg13g2_fill_2 FILLER_33_634 ();
 sg13g2_fill_1 FILLER_33_636 ();
 sg13g2_decap_8 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_661 ();
 sg13g2_decap_4 FILLER_33_671 ();
 sg13g2_fill_1 FILLER_33_675 ();
 sg13g2_fill_1 FILLER_33_720 ();
 sg13g2_decap_8 FILLER_33_734 ();
 sg13g2_decap_4 FILLER_33_741 ();
 sg13g2_fill_2 FILLER_33_745 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_773 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_fill_2 FILLER_33_807 ();
 sg13g2_fill_1 FILLER_33_809 ();
 sg13g2_fill_2 FILLER_33_818 ();
 sg13g2_fill_1 FILLER_33_820 ();
 sg13g2_fill_2 FILLER_33_829 ();
 sg13g2_fill_1 FILLER_33_831 ();
 sg13g2_fill_1 FILLER_33_845 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_decap_4 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_decap_8 FILLER_34_260 ();
 sg13g2_decap_8 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_531 ();
 sg13g2_decap_4 FILLER_34_551 ();
 sg13g2_fill_1 FILLER_34_555 ();
 sg13g2_fill_1 FILLER_34_564 ();
 sg13g2_fill_2 FILLER_34_589 ();
 sg13g2_fill_1 FILLER_34_591 ();
 sg13g2_decap_8 FILLER_34_604 ();
 sg13g2_fill_2 FILLER_34_611 ();
 sg13g2_fill_1 FILLER_34_613 ();
 sg13g2_decap_8 FILLER_34_622 ();
 sg13g2_fill_2 FILLER_34_629 ();
 sg13g2_fill_1 FILLER_34_631 ();
 sg13g2_decap_8 FILLER_34_648 ();
 sg13g2_fill_2 FILLER_34_655 ();
 sg13g2_fill_2 FILLER_34_680 ();
 sg13g2_fill_1 FILLER_34_682 ();
 sg13g2_decap_8 FILLER_34_702 ();
 sg13g2_fill_2 FILLER_34_709 ();
 sg13g2_decap_4 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_730 ();
 sg13g2_decap_8 FILLER_34_737 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_fill_1 FILLER_34_759 ();
 sg13g2_decap_8 FILLER_34_781 ();
 sg13g2_decap_4 FILLER_34_802 ();
 sg13g2_fill_2 FILLER_34_806 ();
 sg13g2_fill_2 FILLER_34_832 ();
 sg13g2_fill_1 FILLER_34_834 ();
 sg13g2_fill_2 FILLER_34_843 ();
 sg13g2_fill_1 FILLER_34_845 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_75 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_92 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_decap_4 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_160 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_338 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_451 ();
 sg13g2_decap_4 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_484 ();
 sg13g2_fill_1 FILLER_35_503 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_fill_2 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_589 ();
 sg13g2_fill_2 FILLER_35_597 ();
 sg13g2_fill_1 FILLER_35_608 ();
 sg13g2_decap_4 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_622 ();
 sg13g2_fill_2 FILLER_35_650 ();
 sg13g2_decap_4 FILLER_35_657 ();
 sg13g2_fill_2 FILLER_35_661 ();
 sg13g2_fill_2 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_fill_1 FILLER_35_714 ();
 sg13g2_fill_1 FILLER_35_752 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_fill_1 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_4 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_fill_1 FILLER_35_844 ();
 sg13g2_decap_4 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_104 ();
 sg13g2_decap_4 FILLER_36_111 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_decap_4 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_221 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_2 FILLER_36_436 ();
 sg13g2_fill_1 FILLER_36_438 ();
 sg13g2_fill_1 FILLER_36_525 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_fill_2 FILLER_36_571 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_decap_8 FILLER_36_589 ();
 sg13g2_fill_2 FILLER_36_609 ();
 sg13g2_fill_1 FILLER_36_611 ();
 sg13g2_decap_4 FILLER_36_625 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_decap_8 FILLER_36_647 ();
 sg13g2_decap_4 FILLER_36_654 ();
 sg13g2_fill_2 FILLER_36_676 ();
 sg13g2_fill_1 FILLER_36_678 ();
 sg13g2_fill_2 FILLER_36_690 ();
 sg13g2_fill_1 FILLER_36_692 ();
 sg13g2_fill_2 FILLER_36_701 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_fill_2 FILLER_36_731 ();
 sg13g2_fill_1 FILLER_36_738 ();
 sg13g2_decap_4 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_773 ();
 sg13g2_fill_2 FILLER_36_780 ();
 sg13g2_fill_2 FILLER_36_786 ();
 sg13g2_fill_1 FILLER_36_788 ();
 sg13g2_decap_4 FILLER_36_794 ();
 sg13g2_decap_4 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_4 FILLER_36_830 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_73 ();
 sg13g2_fill_2 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_decap_4 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_155 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_4 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_4 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_decap_4 FILLER_37_443 ();
 sg13g2_decap_8 FILLER_37_451 ();
 sg13g2_decap_8 FILLER_37_458 ();
 sg13g2_decap_4 FILLER_37_465 ();
 sg13g2_decap_8 FILLER_37_495 ();
 sg13g2_fill_2 FILLER_37_502 ();
 sg13g2_fill_1 FILLER_37_504 ();
 sg13g2_decap_4 FILLER_37_559 ();
 sg13g2_decap_4 FILLER_37_573 ();
 sg13g2_fill_1 FILLER_37_577 ();
 sg13g2_fill_1 FILLER_37_604 ();
 sg13g2_decap_4 FILLER_37_622 ();
 sg13g2_fill_2 FILLER_37_626 ();
 sg13g2_fill_2 FILLER_37_648 ();
 sg13g2_fill_1 FILLER_37_650 ();
 sg13g2_decap_4 FILLER_37_672 ();
 sg13g2_fill_2 FILLER_37_676 ();
 sg13g2_decap_4 FILLER_37_708 ();
 sg13g2_fill_1 FILLER_37_724 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_fill_2 FILLER_37_756 ();
 sg13g2_fill_2 FILLER_37_762 ();
 sg13g2_decap_4 FILLER_37_772 ();
 sg13g2_fill_2 FILLER_37_776 ();
 sg13g2_decap_4 FILLER_37_800 ();
 sg13g2_fill_1 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_fill_2 FILLER_37_840 ();
 sg13g2_decap_4 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_4 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_45 ();
 sg13g2_decap_8 FILLER_38_52 ();
 sg13g2_decap_8 FILLER_38_59 ();
 sg13g2_decap_8 FILLER_38_69 ();
 sg13g2_decap_8 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_decap_4 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_150 ();
 sg13g2_decap_4 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_decap_4 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_405 ();
 sg13g2_decap_4 FILLER_38_412 ();
 sg13g2_fill_1 FILLER_38_416 ();
 sg13g2_fill_2 FILLER_38_445 ();
 sg13g2_fill_1 FILLER_38_447 ();
 sg13g2_decap_8 FILLER_38_457 ();
 sg13g2_fill_2 FILLER_38_524 ();
 sg13g2_fill_2 FILLER_38_537 ();
 sg13g2_decap_8 FILLER_38_544 ();
 sg13g2_decap_8 FILLER_38_551 ();
 sg13g2_decap_8 FILLER_38_558 ();
 sg13g2_decap_4 FILLER_38_565 ();
 sg13g2_fill_2 FILLER_38_569 ();
 sg13g2_fill_1 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_595 ();
 sg13g2_fill_2 FILLER_38_623 ();
 sg13g2_decap_4 FILLER_38_650 ();
 sg13g2_fill_2 FILLER_38_654 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_decap_8 FILLER_38_671 ();
 sg13g2_fill_2 FILLER_38_682 ();
 sg13g2_fill_1 FILLER_38_684 ();
 sg13g2_decap_4 FILLER_38_703 ();
 sg13g2_decap_4 FILLER_38_720 ();
 sg13g2_fill_2 FILLER_38_724 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_4 FILLER_38_746 ();
 sg13g2_decap_4 FILLER_38_769 ();
 sg13g2_fill_1 FILLER_38_773 ();
 sg13g2_fill_2 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_4 FILLER_38_810 ();
 sg13g2_fill_1 FILLER_38_814 ();
 sg13g2_fill_2 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_4 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_69 ();
 sg13g2_decap_4 FILLER_39_83 ();
 sg13g2_fill_2 FILLER_39_87 ();
 sg13g2_decap_8 FILLER_39_108 ();
 sg13g2_fill_2 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_117 ();
 sg13g2_decap_4 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_207 ();
 sg13g2_fill_2 FILLER_39_230 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_288 ();
 sg13g2_fill_2 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_297 ();
 sg13g2_fill_1 FILLER_39_308 ();
 sg13g2_fill_2 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_2 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_351 ();
 sg13g2_fill_1 FILLER_39_366 ();
 sg13g2_decap_4 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_489 ();
 sg13g2_decap_8 FILLER_39_496 ();
 sg13g2_decap_8 FILLER_39_503 ();
 sg13g2_decap_8 FILLER_39_510 ();
 sg13g2_fill_2 FILLER_39_517 ();
 sg13g2_decap_4 FILLER_39_576 ();
 sg13g2_fill_2 FILLER_39_629 ();
 sg13g2_fill_1 FILLER_39_631 ();
 sg13g2_decap_8 FILLER_39_645 ();
 sg13g2_decap_4 FILLER_39_652 ();
 sg13g2_fill_1 FILLER_39_656 ();
 sg13g2_decap_4 FILLER_39_675 ();
 sg13g2_fill_2 FILLER_39_679 ();
 sg13g2_decap_4 FILLER_39_718 ();
 sg13g2_fill_1 FILLER_39_722 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_4 FILLER_39_756 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_fill_2 FILLER_39_782 ();
 sg13g2_fill_1 FILLER_39_784 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_fill_2 FILLER_39_801 ();
 sg13g2_fill_1 FILLER_39_803 ();
 sg13g2_fill_2 FILLER_39_817 ();
 sg13g2_fill_1 FILLER_39_819 ();
 sg13g2_decap_4 FILLER_39_839 ();
 sg13g2_fill_1 FILLER_39_843 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_4 FILLER_40_53 ();
 sg13g2_fill_2 FILLER_40_57 ();
 sg13g2_fill_2 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_decap_4 FILLER_40_128 ();
 sg13g2_fill_1 FILLER_40_132 ();
 sg13g2_fill_1 FILLER_40_162 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_decap_8 FILLER_40_204 ();
 sg13g2_fill_1 FILLER_40_215 ();
 sg13g2_decap_8 FILLER_40_221 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_2 FILLER_40_276 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_decap_4 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_348 ();
 sg13g2_fill_2 FILLER_40_354 ();
 sg13g2_decap_4 FILLER_40_384 ();
 sg13g2_fill_1 FILLER_40_388 ();
 sg13g2_fill_1 FILLER_40_399 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_decap_4 FILLER_40_449 ();
 sg13g2_fill_1 FILLER_40_453 ();
 sg13g2_decap_8 FILLER_40_458 ();
 sg13g2_fill_2 FILLER_40_465 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_fill_1 FILLER_40_533 ();
 sg13g2_decap_4 FILLER_40_600 ();
 sg13g2_fill_1 FILLER_40_604 ();
 sg13g2_fill_2 FILLER_40_619 ();
 sg13g2_decap_4 FILLER_40_629 ();
 sg13g2_fill_1 FILLER_40_633 ();
 sg13g2_decap_8 FILLER_40_656 ();
 sg13g2_decap_8 FILLER_40_671 ();
 sg13g2_decap_8 FILLER_40_678 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_fill_2 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_713 ();
 sg13g2_decap_8 FILLER_40_750 ();
 sg13g2_fill_1 FILLER_40_757 ();
 sg13g2_fill_1 FILLER_40_762 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_fill_2 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_794 ();
 sg13g2_fill_2 FILLER_40_801 ();
 sg13g2_fill_2 FILLER_40_825 ();
 sg13g2_decap_4 FILLER_40_844 ();
 sg13g2_fill_1 FILLER_40_848 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_28 ();
 sg13g2_decap_4 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_fill_2 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_121 ();
 sg13g2_fill_2 FILLER_41_180 ();
 sg13g2_fill_1 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_203 ();
 sg13g2_decap_4 FILLER_41_233 ();
 sg13g2_fill_2 FILLER_41_243 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_decap_4 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_fill_1 FILLER_41_304 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_fill_2 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_374 ();
 sg13g2_decap_4 FILLER_41_381 ();
 sg13g2_decap_4 FILLER_41_412 ();
 sg13g2_fill_1 FILLER_41_489 ();
 sg13g2_decap_4 FILLER_41_516 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_fill_1 FILLER_41_535 ();
 sg13g2_decap_4 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_4 FILLER_41_654 ();
 sg13g2_fill_2 FILLER_41_658 ();
 sg13g2_decap_4 FILLER_41_669 ();
 sg13g2_fill_1 FILLER_41_673 ();
 sg13g2_decap_4 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_686 ();
 sg13g2_fill_1 FILLER_41_709 ();
 sg13g2_decap_4 FILLER_41_715 ();
 sg13g2_fill_2 FILLER_41_719 ();
 sg13g2_decap_4 FILLER_41_735 ();
 sg13g2_decap_4 FILLER_41_744 ();
 sg13g2_fill_2 FILLER_41_748 ();
 sg13g2_fill_2 FILLER_41_763 ();
 sg13g2_decap_4 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_777 ();
 sg13g2_fill_1 FILLER_41_791 ();
 sg13g2_decap_4 FILLER_41_804 ();
 sg13g2_fill_2 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_fill_1 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_36 ();
 sg13g2_fill_1 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_fill_1 FILLER_42_111 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_133 ();
 sg13g2_decap_4 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_146 ();
 sg13g2_decap_4 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_decap_4 FILLER_42_210 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_fill_1 FILLER_42_241 ();
 sg13g2_fill_2 FILLER_42_314 ();
 sg13g2_fill_2 FILLER_42_336 ();
 sg13g2_fill_2 FILLER_42_346 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_decap_4 FILLER_42_372 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_2 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_fill_2 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_439 ();
 sg13g2_fill_2 FILLER_42_447 ();
 sg13g2_decap_4 FILLER_42_467 ();
 sg13g2_fill_1 FILLER_42_480 ();
 sg13g2_fill_2 FILLER_42_500 ();
 sg13g2_fill_1 FILLER_42_502 ();
 sg13g2_fill_2 FILLER_42_530 ();
 sg13g2_fill_1 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_573 ();
 sg13g2_decap_4 FILLER_42_580 ();
 sg13g2_fill_2 FILLER_42_610 ();
 sg13g2_decap_8 FILLER_42_639 ();
 sg13g2_fill_2 FILLER_42_646 ();
 sg13g2_fill_2 FILLER_42_673 ();
 sg13g2_fill_1 FILLER_42_675 ();
 sg13g2_fill_2 FILLER_42_680 ();
 sg13g2_fill_1 FILLER_42_696 ();
 sg13g2_decap_4 FILLER_42_721 ();
 sg13g2_fill_2 FILLER_42_725 ();
 sg13g2_fill_2 FILLER_42_733 ();
 sg13g2_decap_4 FILLER_42_747 ();
 sg13g2_fill_1 FILLER_42_751 ();
 sg13g2_fill_2 FILLER_42_756 ();
 sg13g2_decap_4 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_fill_2 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_827 ();
 sg13g2_fill_2 FILLER_42_834 ();
 sg13g2_fill_1 FILLER_42_836 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_17 ();
 sg13g2_fill_2 FILLER_43_24 ();
 sg13g2_fill_1 FILLER_43_26 ();
 sg13g2_fill_1 FILLER_43_67 ();
 sg13g2_fill_1 FILLER_43_83 ();
 sg13g2_decap_8 FILLER_43_97 ();
 sg13g2_decap_8 FILLER_43_125 ();
 sg13g2_decap_4 FILLER_43_132 ();
 sg13g2_decap_4 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_2 FILLER_43_154 ();
 sg13g2_fill_1 FILLER_43_156 ();
 sg13g2_decap_8 FILLER_43_162 ();
 sg13g2_fill_2 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_decap_8 FILLER_43_177 ();
 sg13g2_fill_2 FILLER_43_184 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_4 FILLER_43_238 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_decap_4 FILLER_43_256 ();
 sg13g2_fill_2 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_336 ();
 sg13g2_fill_2 FILLER_43_347 ();
 sg13g2_decap_4 FILLER_43_387 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_2 FILLER_43_402 ();
 sg13g2_decap_4 FILLER_43_419 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_43_430 ();
 sg13g2_fill_2 FILLER_43_435 ();
 sg13g2_fill_2 FILLER_43_456 ();
 sg13g2_fill_2 FILLER_43_505 ();
 sg13g2_decap_8 FILLER_43_529 ();
 sg13g2_fill_1 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_542 ();
 sg13g2_decap_4 FILLER_43_549 ();
 sg13g2_fill_2 FILLER_43_553 ();
 sg13g2_fill_1 FILLER_43_606 ();
 sg13g2_fill_2 FILLER_43_635 ();
 sg13g2_fill_1 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_650 ();
 sg13g2_fill_1 FILLER_43_661 ();
 sg13g2_decap_8 FILLER_43_667 ();
 sg13g2_decap_4 FILLER_43_674 ();
 sg13g2_fill_2 FILLER_43_684 ();
 sg13g2_fill_1 FILLER_43_686 ();
 sg13g2_decap_4 FILLER_43_704 ();
 sg13g2_fill_2 FILLER_43_708 ();
 sg13g2_fill_1 FILLER_43_714 ();
 sg13g2_fill_2 FILLER_43_725 ();
 sg13g2_fill_2 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_fill_2 FILLER_43_749 ();
 sg13g2_fill_1 FILLER_43_751 ();
 sg13g2_decap_8 FILLER_43_773 ();
 sg13g2_fill_2 FILLER_43_780 ();
 sg13g2_fill_2 FILLER_43_794 ();
 sg13g2_fill_1 FILLER_43_796 ();
 sg13g2_decap_4 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_decap_4 FILLER_44_113 ();
 sg13g2_fill_1 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_135 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_fill_2 FILLER_44_187 ();
 sg13g2_fill_1 FILLER_44_189 ();
 sg13g2_fill_1 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_4 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_247 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_fill_1 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_342 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_decap_4 FILLER_44_363 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_decap_8 FILLER_44_377 ();
 sg13g2_decap_8 FILLER_44_384 ();
 sg13g2_decap_8 FILLER_44_391 ();
 sg13g2_fill_2 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_400 ();
 sg13g2_decap_4 FILLER_44_417 ();
 sg13g2_fill_2 FILLER_44_421 ();
 sg13g2_decap_8 FILLER_44_442 ();
 sg13g2_decap_8 FILLER_44_449 ();
 sg13g2_fill_1 FILLER_44_456 ();
 sg13g2_decap_8 FILLER_44_474 ();
 sg13g2_fill_1 FILLER_44_481 ();
 sg13g2_decap_8 FILLER_44_499 ();
 sg13g2_decap_8 FILLER_44_506 ();
 sg13g2_fill_2 FILLER_44_513 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_fill_1 FILLER_44_523 ();
 sg13g2_decap_4 FILLER_44_532 ();
 sg13g2_fill_1 FILLER_44_536 ();
 sg13g2_fill_2 FILLER_44_541 ();
 sg13g2_fill_2 FILLER_44_560 ();
 sg13g2_fill_1 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_576 ();
 sg13g2_decap_8 FILLER_44_583 ();
 sg13g2_decap_4 FILLER_44_631 ();
 sg13g2_fill_1 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_fill_2 FILLER_44_683 ();
 sg13g2_decap_4 FILLER_44_696 ();
 sg13g2_fill_2 FILLER_44_700 ();
 sg13g2_fill_2 FILLER_44_738 ();
 sg13g2_fill_1 FILLER_44_740 ();
 sg13g2_decap_4 FILLER_44_762 ();
 sg13g2_decap_8 FILLER_44_771 ();
 sg13g2_decap_4 FILLER_44_778 ();
 sg13g2_decap_4 FILLER_44_794 ();
 sg13g2_fill_2 FILLER_44_798 ();
 sg13g2_fill_2 FILLER_44_804 ();
 sg13g2_decap_4 FILLER_44_822 ();
 sg13g2_fill_2 FILLER_44_826 ();
 sg13g2_fill_2 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_835 ();
 sg13g2_decap_4 FILLER_44_841 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_13 ();
 sg13g2_fill_1 FILLER_45_38 ();
 sg13g2_decap_8 FILLER_45_44 ();
 sg13g2_decap_4 FILLER_45_51 ();
 sg13g2_fill_2 FILLER_45_76 ();
 sg13g2_fill_1 FILLER_45_78 ();
 sg13g2_decap_8 FILLER_45_89 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_2 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_121 ();
 sg13g2_decap_4 FILLER_45_128 ();
 sg13g2_fill_1 FILLER_45_132 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_fill_1 FILLER_45_145 ();
 sg13g2_decap_4 FILLER_45_165 ();
 sg13g2_fill_2 FILLER_45_169 ();
 sg13g2_decap_8 FILLER_45_176 ();
 sg13g2_fill_2 FILLER_45_183 ();
 sg13g2_decap_8 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_204 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_4 FILLER_45_367 ();
 sg13g2_fill_1 FILLER_45_371 ();
 sg13g2_fill_2 FILLER_45_419 ();
 sg13g2_fill_1 FILLER_45_440 ();
 sg13g2_fill_2 FILLER_45_450 ();
 sg13g2_fill_1 FILLER_45_452 ();
 sg13g2_fill_2 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_483 ();
 sg13g2_decap_4 FILLER_45_508 ();
 sg13g2_fill_2 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_569 ();
 sg13g2_fill_2 FILLER_45_610 ();
 sg13g2_fill_1 FILLER_45_612 ();
 sg13g2_decap_4 FILLER_45_627 ();
 sg13g2_fill_1 FILLER_45_631 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_654 ();
 sg13g2_decap_4 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_701 ();
 sg13g2_fill_1 FILLER_45_708 ();
 sg13g2_decap_8 FILLER_45_715 ();
 sg13g2_decap_4 FILLER_45_722 ();
 sg13g2_fill_2 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_decap_8 FILLER_45_783 ();
 sg13g2_decap_4 FILLER_45_790 ();
 sg13g2_fill_1 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_fill_1 FILLER_45_807 ();
 sg13g2_decap_4 FILLER_45_823 ();
 sg13g2_fill_2 FILLER_45_835 ();
 sg13g2_decap_4 FILLER_45_858 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_32 ();
 sg13g2_decap_4 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_92 ();
 sg13g2_decap_4 FILLER_46_145 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_196 ();
 sg13g2_fill_2 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_240 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_4 FILLER_46_259 ();
 sg13g2_decap_4 FILLER_46_267 ();
 sg13g2_fill_2 FILLER_46_313 ();
 sg13g2_fill_1 FILLER_46_342 ();
 sg13g2_fill_2 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_decap_4 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_4 FILLER_46_398 ();
 sg13g2_fill_2 FILLER_46_402 ();
 sg13g2_decap_4 FILLER_46_419 ();
 sg13g2_fill_1 FILLER_46_450 ();
 sg13g2_fill_2 FILLER_46_469 ();
 sg13g2_decap_4 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_512 ();
 sg13g2_decap_8 FILLER_46_542 ();
 sg13g2_fill_2 FILLER_46_549 ();
 sg13g2_fill_1 FILLER_46_551 ();
 sg13g2_decap_4 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_4 FILLER_46_601 ();
 sg13g2_fill_1 FILLER_46_605 ();
 sg13g2_decap_8 FILLER_46_650 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_decap_4 FILLER_46_668 ();
 sg13g2_fill_1 FILLER_46_681 ();
 sg13g2_fill_2 FILLER_46_687 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_718 ();
 sg13g2_fill_1 FILLER_46_720 ();
 sg13g2_decap_8 FILLER_46_736 ();
 sg13g2_decap_4 FILLER_46_743 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_fill_1 FILLER_46_793 ();
 sg13g2_fill_1 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_fill_1 FILLER_46_816 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_4 FILLER_46_836 ();
 sg13g2_fill_2 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_decap_4 FILLER_47_18 ();
 sg13g2_fill_1 FILLER_47_22 ();
 sg13g2_fill_2 FILLER_47_45 ();
 sg13g2_fill_2 FILLER_47_58 ();
 sg13g2_decap_8 FILLER_47_69 ();
 sg13g2_decap_4 FILLER_47_76 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_decap_8 FILLER_47_86 ();
 sg13g2_decap_4 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_97 ();
 sg13g2_decap_4 FILLER_47_117 ();
 sg13g2_fill_2 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_decap_4 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_decap_4 FILLER_47_180 ();
 sg13g2_decap_4 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_243 ();
 sg13g2_fill_1 FILLER_47_250 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_2 FILLER_47_295 ();
 sg13g2_fill_2 FILLER_47_318 ();
 sg13g2_fill_2 FILLER_47_324 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_2 FILLER_47_392 ();
 sg13g2_decap_4 FILLER_47_407 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_fill_2 FILLER_47_455 ();
 sg13g2_fill_2 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_fill_1 FILLER_47_514 ();
 sg13g2_fill_2 FILLER_47_552 ();
 sg13g2_fill_1 FILLER_47_554 ();
 sg13g2_fill_2 FILLER_47_629 ();
 sg13g2_fill_2 FILLER_47_636 ();
 sg13g2_decap_8 FILLER_47_643 ();
 sg13g2_decap_8 FILLER_47_650 ();
 sg13g2_decap_4 FILLER_47_657 ();
 sg13g2_fill_1 FILLER_47_661 ();
 sg13g2_fill_2 FILLER_47_676 ();
 sg13g2_decap_4 FILLER_47_688 ();
 sg13g2_fill_2 FILLER_47_699 ();
 sg13g2_fill_1 FILLER_47_701 ();
 sg13g2_decap_4 FILLER_47_724 ();
 sg13g2_decap_4 FILLER_47_732 ();
 sg13g2_fill_1 FILLER_47_736 ();
 sg13g2_fill_2 FILLER_47_741 ();
 sg13g2_fill_1 FILLER_47_743 ();
 sg13g2_fill_2 FILLER_47_753 ();
 sg13g2_fill_1 FILLER_47_755 ();
 sg13g2_fill_2 FILLER_47_761 ();
 sg13g2_decap_8 FILLER_47_776 ();
 sg13g2_fill_1 FILLER_47_783 ();
 sg13g2_fill_2 FILLER_47_789 ();
 sg13g2_fill_1 FILLER_47_791 ();
 sg13g2_decap_4 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_fill_2 FILLER_47_832 ();
 sg13g2_fill_1 FILLER_47_834 ();
 sg13g2_decap_4 FILLER_47_858 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_108 ();
 sg13g2_decap_4 FILLER_48_122 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_decap_4 FILLER_48_167 ();
 sg13g2_decap_8 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_194 ();
 sg13g2_fill_2 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_203 ();
 sg13g2_fill_2 FILLER_48_213 ();
 sg13g2_decap_8 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_decap_4 FILLER_48_373 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_fill_1 FILLER_48_392 ();
 sg13g2_fill_2 FILLER_48_472 ();
 sg13g2_fill_1 FILLER_48_496 ();
 sg13g2_fill_2 FILLER_48_510 ();
 sg13g2_decap_4 FILLER_48_520 ();
 sg13g2_fill_2 FILLER_48_537 ();
 sg13g2_fill_1 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_584 ();
 sg13g2_fill_1 FILLER_48_586 ();
 sg13g2_decap_8 FILLER_48_591 ();
 sg13g2_decap_8 FILLER_48_607 ();
 sg13g2_fill_1 FILLER_48_633 ();
 sg13g2_fill_2 FILLER_48_654 ();
 sg13g2_fill_1 FILLER_48_656 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_fill_2 FILLER_48_683 ();
 sg13g2_fill_1 FILLER_48_685 ();
 sg13g2_decap_8 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_705 ();
 sg13g2_fill_2 FILLER_48_720 ();
 sg13g2_fill_1 FILLER_48_722 ();
 sg13g2_decap_4 FILLER_48_735 ();
 sg13g2_decap_4 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_776 ();
 sg13g2_decap_4 FILLER_48_783 ();
 sg13g2_fill_1 FILLER_48_823 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_4 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_4 ();
 sg13g2_fill_2 FILLER_49_33 ();
 sg13g2_fill_1 FILLER_49_35 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_72 ();
 sg13g2_decap_4 FILLER_49_79 ();
 sg13g2_fill_1 FILLER_49_83 ();
 sg13g2_decap_8 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_104 ();
 sg13g2_decap_8 FILLER_49_132 ();
 sg13g2_decap_4 FILLER_49_139 ();
 sg13g2_fill_2 FILLER_49_143 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_fill_2 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_fill_2 FILLER_49_242 ();
 sg13g2_fill_2 FILLER_49_257 ();
 sg13g2_fill_1 FILLER_49_259 ();
 sg13g2_fill_2 FILLER_49_270 ();
 sg13g2_fill_2 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_4 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_411 ();
 sg13g2_fill_1 FILLER_49_413 ();
 sg13g2_fill_2 FILLER_49_441 ();
 sg13g2_fill_1 FILLER_49_443 ();
 sg13g2_fill_1 FILLER_49_453 ();
 sg13g2_decap_4 FILLER_49_558 ();
 sg13g2_fill_2 FILLER_49_566 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_fill_2 FILLER_49_578 ();
 sg13g2_fill_2 FILLER_49_612 ();
 sg13g2_fill_1 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_626 ();
 sg13g2_decap_8 FILLER_49_633 ();
 sg13g2_fill_2 FILLER_49_640 ();
 sg13g2_decap_8 FILLER_49_650 ();
 sg13g2_fill_2 FILLER_49_657 ();
 sg13g2_decap_4 FILLER_49_677 ();
 sg13g2_fill_1 FILLER_49_681 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_decap_4 FILLER_49_704 ();
 sg13g2_fill_1 FILLER_49_708 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_4 FILLER_49_740 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_4 FILLER_49_782 ();
 sg13g2_fill_1 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_813 ();
 sg13g2_fill_1 FILLER_49_820 ();
 sg13g2_fill_2 FILLER_49_833 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_43 ();
 sg13g2_decap_4 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_73 ();
 sg13g2_fill_1 FILLER_50_90 ();
 sg13g2_decap_4 FILLER_50_122 ();
 sg13g2_fill_1 FILLER_50_126 ();
 sg13g2_fill_1 FILLER_50_144 ();
 sg13g2_fill_2 FILLER_50_149 ();
 sg13g2_fill_1 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_decap_4 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_171 ();
 sg13g2_decap_4 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_190 ();
 sg13g2_decap_8 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_240 ();
 sg13g2_decap_4 FILLER_50_247 ();
 sg13g2_decap_4 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_fill_1 FILLER_50_281 ();
 sg13g2_decap_4 FILLER_50_320 ();
 sg13g2_fill_1 FILLER_50_332 ();
 sg13g2_decap_8 FILLER_50_355 ();
 sg13g2_decap_8 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_373 ();
 sg13g2_fill_1 FILLER_50_459 ();
 sg13g2_fill_1 FILLER_50_492 ();
 sg13g2_fill_1 FILLER_50_545 ();
 sg13g2_fill_1 FILLER_50_560 ();
 sg13g2_fill_2 FILLER_50_582 ();
 sg13g2_fill_1 FILLER_50_584 ();
 sg13g2_fill_2 FILLER_50_594 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_635 ();
 sg13g2_fill_1 FILLER_50_641 ();
 sg13g2_fill_1 FILLER_50_662 ();
 sg13g2_decap_8 FILLER_50_684 ();
 sg13g2_fill_1 FILLER_50_691 ();
 sg13g2_fill_1 FILLER_50_704 ();
 sg13g2_decap_8 FILLER_50_718 ();
 sg13g2_decap_4 FILLER_50_725 ();
 sg13g2_fill_1 FILLER_50_729 ();
 sg13g2_decap_8 FILLER_50_747 ();
 sg13g2_decap_4 FILLER_50_754 ();
 sg13g2_fill_1 FILLER_50_771 ();
 sg13g2_decap_4 FILLER_50_780 ();
 sg13g2_decap_8 FILLER_50_803 ();
 sg13g2_fill_1 FILLER_50_810 ();
 sg13g2_decap_4 FILLER_50_823 ();
 sg13g2_fill_1 FILLER_50_827 ();
 sg13g2_decap_8 FILLER_50_832 ();
 sg13g2_decap_8 FILLER_50_839 ();
 sg13g2_fill_2 FILLER_50_846 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_4 FILLER_51_68 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_decap_4 FILLER_51_96 ();
 sg13g2_fill_2 FILLER_51_100 ();
 sg13g2_decap_8 FILLER_51_107 ();
 sg13g2_fill_1 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_192 ();
 sg13g2_decap_8 FILLER_51_199 ();
 sg13g2_decap_4 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_decap_8 FILLER_51_246 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_257 ();
 sg13g2_fill_2 FILLER_51_267 ();
 sg13g2_fill_2 FILLER_51_284 ();
 sg13g2_fill_2 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_427 ();
 sg13g2_fill_2 FILLER_51_434 ();
 sg13g2_fill_2 FILLER_51_478 ();
 sg13g2_fill_1 FILLER_51_480 ();
 sg13g2_fill_2 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_521 ();
 sg13g2_fill_2 FILLER_51_536 ();
 sg13g2_fill_1 FILLER_51_564 ();
 sg13g2_fill_2 FILLER_51_570 ();
 sg13g2_fill_1 FILLER_51_572 ();
 sg13g2_fill_2 FILLER_51_597 ();
 sg13g2_fill_1 FILLER_51_599 ();
 sg13g2_decap_8 FILLER_51_628 ();
 sg13g2_fill_2 FILLER_51_635 ();
 sg13g2_decap_8 FILLER_51_653 ();
 sg13g2_decap_4 FILLER_51_660 ();
 sg13g2_fill_2 FILLER_51_664 ();
 sg13g2_decap_4 FILLER_51_679 ();
 sg13g2_decap_8 FILLER_51_689 ();
 sg13g2_fill_2 FILLER_51_713 ();
 sg13g2_fill_1 FILLER_51_715 ();
 sg13g2_decap_4 FILLER_51_728 ();
 sg13g2_fill_1 FILLER_51_732 ();
 sg13g2_decap_8 FILLER_51_759 ();
 sg13g2_decap_4 FILLER_51_766 ();
 sg13g2_decap_4 FILLER_51_775 ();
 sg13g2_fill_2 FILLER_51_779 ();
 sg13g2_fill_1 FILLER_51_786 ();
 sg13g2_decap_8 FILLER_51_799 ();
 sg13g2_fill_2 FILLER_51_806 ();
 sg13g2_fill_1 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_831 ();
 sg13g2_fill_1 FILLER_51_838 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_fill_2 FILLER_52_43 ();
 sg13g2_fill_2 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_58 ();
 sg13g2_decap_8 FILLER_52_64 ();
 sg13g2_decap_8 FILLER_52_71 ();
 sg13g2_decap_8 FILLER_52_94 ();
 sg13g2_decap_8 FILLER_52_101 ();
 sg13g2_fill_2 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_110 ();
 sg13g2_decap_4 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_152 ();
 sg13g2_decap_8 FILLER_52_156 ();
 sg13g2_decap_8 FILLER_52_163 ();
 sg13g2_decap_8 FILLER_52_214 ();
 sg13g2_decap_4 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_225 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_fill_2 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_275 ();
 sg13g2_fill_2 FILLER_52_279 ();
 sg13g2_fill_2 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_295 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_326 ();
 sg13g2_decap_4 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_fill_1 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_410 ();
 sg13g2_fill_1 FILLER_52_416 ();
 sg13g2_fill_1 FILLER_52_430 ();
 sg13g2_decap_4 FILLER_52_444 ();
 sg13g2_fill_2 FILLER_52_501 ();
 sg13g2_decap_8 FILLER_52_511 ();
 sg13g2_fill_2 FILLER_52_546 ();
 sg13g2_fill_1 FILLER_52_548 ();
 sg13g2_decap_4 FILLER_52_585 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_fill_2 FILLER_52_627 ();
 sg13g2_fill_2 FILLER_52_674 ();
 sg13g2_decap_8 FILLER_52_703 ();
 sg13g2_fill_2 FILLER_52_710 ();
 sg13g2_fill_1 FILLER_52_712 ();
 sg13g2_decap_4 FILLER_52_718 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_fill_2 FILLER_52_742 ();
 sg13g2_fill_2 FILLER_52_769 ();
 sg13g2_fill_1 FILLER_52_771 ();
 sg13g2_decap_8 FILLER_52_792 ();
 sg13g2_decap_8 FILLER_52_799 ();
 sg13g2_decap_4 FILLER_52_830 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_4 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_94 ();
 sg13g2_fill_1 FILLER_53_101 ();
 sg13g2_decap_8 FILLER_53_130 ();
 sg13g2_decap_8 FILLER_53_137 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_fill_2 FILLER_53_175 ();
 sg13g2_fill_1 FILLER_53_177 ();
 sg13g2_decap_8 FILLER_53_193 ();
 sg13g2_decap_8 FILLER_53_200 ();
 sg13g2_decap_8 FILLER_53_249 ();
 sg13g2_decap_8 FILLER_53_256 ();
 sg13g2_decap_8 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_decap_8 FILLER_53_292 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_fill_2 FILLER_53_314 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_327 ();
 sg13g2_fill_2 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_fill_2 FILLER_53_367 ();
 sg13g2_decap_4 FILLER_53_382 ();
 sg13g2_fill_2 FILLER_53_386 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_fill_1 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_53_435 ();
 sg13g2_fill_2 FILLER_53_450 ();
 sg13g2_decap_8 FILLER_53_537 ();
 sg13g2_decap_8 FILLER_53_549 ();
 sg13g2_fill_1 FILLER_53_556 ();
 sg13g2_decap_8 FILLER_53_571 ();
 sg13g2_decap_4 FILLER_53_578 ();
 sg13g2_fill_2 FILLER_53_638 ();
 sg13g2_decap_4 FILLER_53_654 ();
 sg13g2_fill_1 FILLER_53_665 ();
 sg13g2_fill_1 FILLER_53_681 ();
 sg13g2_fill_2 FILLER_53_687 ();
 sg13g2_fill_1 FILLER_53_689 ();
 sg13g2_decap_8 FILLER_53_695 ();
 sg13g2_fill_2 FILLER_53_702 ();
 sg13g2_fill_1 FILLER_53_704 ();
 sg13g2_decap_4 FILLER_53_719 ();
 sg13g2_fill_2 FILLER_53_730 ();
 sg13g2_decap_4 FILLER_53_745 ();
 sg13g2_decap_8 FILLER_53_761 ();
 sg13g2_decap_8 FILLER_53_768 ();
 sg13g2_fill_2 FILLER_53_775 ();
 sg13g2_fill_1 FILLER_53_777 ();
 sg13g2_decap_4 FILLER_53_795 ();
 sg13g2_decap_4 FILLER_53_823 ();
 sg13g2_fill_2 FILLER_53_827 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_fill_2 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_decap_4 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_118 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_2 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_decap_4 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_187 ();
 sg13g2_fill_2 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_225 ();
 sg13g2_fill_1 FILLER_54_227 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_fill_1 FILLER_54_245 ();
 sg13g2_decap_4 FILLER_54_267 ();
 sg13g2_fill_2 FILLER_54_271 ();
 sg13g2_fill_2 FILLER_54_294 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_decap_4 FILLER_54_352 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_376 ();
 sg13g2_fill_1 FILLER_54_471 ();
 sg13g2_fill_1 FILLER_54_477 ();
 sg13g2_fill_2 FILLER_54_482 ();
 sg13g2_fill_1 FILLER_54_484 ();
 sg13g2_decap_8 FILLER_54_505 ();
 sg13g2_fill_1 FILLER_54_512 ();
 sg13g2_fill_2 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_527 ();
 sg13g2_decap_4 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_584 ();
 sg13g2_fill_2 FILLER_54_595 ();
 sg13g2_fill_1 FILLER_54_597 ();
 sg13g2_decap_8 FILLER_54_664 ();
 sg13g2_decap_8 FILLER_54_671 ();
 sg13g2_fill_2 FILLER_54_678 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_decap_8 FILLER_54_708 ();
 sg13g2_decap_8 FILLER_54_715 ();
 sg13g2_fill_2 FILLER_54_727 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_fill_2 FILLER_54_743 ();
 sg13g2_fill_2 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_756 ();
 sg13g2_decap_8 FILLER_54_763 ();
 sg13g2_fill_2 FILLER_54_770 ();
 sg13g2_decap_8 FILLER_54_782 ();
 sg13g2_fill_2 FILLER_54_789 ();
 sg13g2_decap_8 FILLER_54_799 ();
 sg13g2_fill_1 FILLER_54_806 ();
 sg13g2_decap_8 FILLER_54_820 ();
 sg13g2_decap_8 FILLER_54_827 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_4 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_fill_2 FILLER_55_27 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_decap_4 FILLER_55_73 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_4 FILLER_55_161 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_decap_4 FILLER_55_180 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_196 ();
 sg13g2_fill_2 FILLER_55_204 ();
 sg13g2_fill_2 FILLER_55_220 ();
 sg13g2_fill_2 FILLER_55_250 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_4 FILLER_55_287 ();
 sg13g2_fill_2 FILLER_55_291 ();
 sg13g2_decap_4 FILLER_55_298 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_decap_4 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_337 ();
 sg13g2_fill_1 FILLER_55_339 ();
 sg13g2_decap_8 FILLER_55_388 ();
 sg13g2_fill_1 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_decap_4 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_55_411 ();
 sg13g2_fill_2 FILLER_55_496 ();
 sg13g2_fill_1 FILLER_55_511 ();
 sg13g2_fill_1 FILLER_55_525 ();
 sg13g2_decap_8 FILLER_55_543 ();
 sg13g2_fill_1 FILLER_55_550 ();
 sg13g2_fill_2 FILLER_55_555 ();
 sg13g2_fill_1 FILLER_55_557 ();
 sg13g2_fill_2 FILLER_55_561 ();
 sg13g2_fill_2 FILLER_55_584 ();
 sg13g2_fill_2 FILLER_55_595 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_625 ();
 sg13g2_fill_1 FILLER_55_639 ();
 sg13g2_decap_8 FILLER_55_663 ();
 sg13g2_fill_2 FILLER_55_670 ();
 sg13g2_decap_8 FILLER_55_685 ();
 sg13g2_fill_1 FILLER_55_692 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_739 ();
 sg13g2_fill_1 FILLER_55_768 ();
 sg13g2_decap_8 FILLER_55_795 ();
 sg13g2_decap_4 FILLER_55_802 ();
 sg13g2_fill_1 FILLER_55_806 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_4 FILLER_55_856 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_4 ();
 sg13g2_decap_8 FILLER_56_9 ();
 sg13g2_fill_2 FILLER_56_16 ();
 sg13g2_decap_8 FILLER_56_62 ();
 sg13g2_fill_2 FILLER_56_69 ();
 sg13g2_fill_1 FILLER_56_71 ();
 sg13g2_decap_4 FILLER_56_80 ();
 sg13g2_fill_2 FILLER_56_84 ();
 sg13g2_fill_1 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_decap_4 FILLER_56_155 ();
 sg13g2_fill_1 FILLER_56_159 ();
 sg13g2_fill_1 FILLER_56_164 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_178 ();
 sg13g2_fill_2 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_decap_8 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_209 ();
 sg13g2_fill_1 FILLER_56_211 ();
 sg13g2_fill_2 FILLER_56_226 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_249 ();
 sg13g2_fill_2 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_decap_8 FILLER_56_304 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_332 ();
 sg13g2_fill_1 FILLER_56_334 ();
 sg13g2_decap_8 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_355 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_2 FILLER_56_419 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_fill_1 FILLER_56_469 ();
 sg13g2_fill_1 FILLER_56_474 ();
 sg13g2_fill_1 FILLER_56_502 ();
 sg13g2_fill_2 FILLER_56_567 ();
 sg13g2_fill_1 FILLER_56_597 ();
 sg13g2_fill_2 FILLER_56_640 ();
 sg13g2_fill_2 FILLER_56_647 ();
 sg13g2_fill_2 FILLER_56_682 ();
 sg13g2_fill_1 FILLER_56_684 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_fill_2 FILLER_56_717 ();
 sg13g2_fill_1 FILLER_56_732 ();
 sg13g2_fill_2 FILLER_56_827 ();
 sg13g2_fill_1 FILLER_56_829 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_38 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_80 ();
 sg13g2_decap_8 FILLER_57_101 ();
 sg13g2_decap_4 FILLER_57_108 ();
 sg13g2_fill_2 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_118 ();
 sg13g2_fill_2 FILLER_57_125 ();
 sg13g2_decap_8 FILLER_57_132 ();
 sg13g2_fill_2 FILLER_57_139 ();
 sg13g2_fill_1 FILLER_57_141 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_1 FILLER_57_184 ();
 sg13g2_decap_4 FILLER_57_189 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_4 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_221 ();
 sg13g2_decap_4 FILLER_57_231 ();
 sg13g2_decap_4 FILLER_57_250 ();
 sg13g2_decap_4 FILLER_57_267 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_decap_4 FILLER_57_286 ();
 sg13g2_fill_2 FILLER_57_290 ();
 sg13g2_decap_4 FILLER_57_317 ();
 sg13g2_fill_2 FILLER_57_321 ();
 sg13g2_fill_1 FILLER_57_330 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_fill_2 FILLER_57_390 ();
 sg13g2_fill_1 FILLER_57_392 ();
 sg13g2_decap_4 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_57_435 ();
 sg13g2_fill_2 FILLER_57_442 ();
 sg13g2_fill_1 FILLER_57_444 ();
 sg13g2_fill_1 FILLER_57_454 ();
 sg13g2_fill_2 FILLER_57_491 ();
 sg13g2_fill_2 FILLER_57_510 ();
 sg13g2_fill_1 FILLER_57_512 ();
 sg13g2_decap_4 FILLER_57_564 ();
 sg13g2_fill_1 FILLER_57_568 ();
 sg13g2_decap_8 FILLER_57_580 ();
 sg13g2_fill_2 FILLER_57_587 ();
 sg13g2_fill_2 FILLER_57_601 ();
 sg13g2_fill_2 FILLER_57_607 ();
 sg13g2_decap_8 FILLER_57_647 ();
 sg13g2_decap_8 FILLER_57_654 ();
 sg13g2_decap_8 FILLER_57_661 ();
 sg13g2_fill_1 FILLER_57_678 ();
 sg13g2_decap_8 FILLER_57_687 ();
 sg13g2_decap_4 FILLER_57_694 ();
 sg13g2_fill_1 FILLER_57_698 ();
 sg13g2_fill_2 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_727 ();
 sg13g2_fill_2 FILLER_57_766 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_fill_2 FILLER_57_785 ();
 sg13g2_fill_1 FILLER_57_801 ();
 sg13g2_fill_1 FILLER_57_821 ();
 sg13g2_fill_2 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_4 ();
 sg13g2_decap_8 FILLER_58_10 ();
 sg13g2_decap_8 FILLER_58_17 ();
 sg13g2_decap_4 FILLER_58_24 ();
 sg13g2_fill_2 FILLER_58_28 ();
 sg13g2_fill_2 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_47 ();
 sg13g2_decap_4 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_60 ();
 sg13g2_decap_8 FILLER_58_72 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_decap_8 FILLER_58_85 ();
 sg13g2_fill_2 FILLER_58_92 ();
 sg13g2_decap_4 FILLER_58_116 ();
 sg13g2_fill_1 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_decap_4 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_143 ();
 sg13g2_decap_4 FILLER_58_159 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_fill_1 FILLER_58_178 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_decap_4 FILLER_58_229 ();
 sg13g2_decap_8 FILLER_58_256 ();
 sg13g2_decap_8 FILLER_58_263 ();
 sg13g2_fill_1 FILLER_58_270 ();
 sg13g2_decap_8 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_299 ();
 sg13g2_fill_1 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_1 FILLER_58_321 ();
 sg13g2_decap_4 FILLER_58_335 ();
 sg13g2_decap_8 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_351 ();
 sg13g2_decap_4 FILLER_58_358 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_2 FILLER_58_367 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_fill_2 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_434 ();
 sg13g2_fill_2 FILLER_58_479 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_fill_2 FILLER_58_554 ();
 sg13g2_fill_1 FILLER_58_556 ();
 sg13g2_decap_8 FILLER_58_561 ();
 sg13g2_fill_2 FILLER_58_568 ();
 sg13g2_fill_1 FILLER_58_570 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_fill_2 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_624 ();
 sg13g2_decap_4 FILLER_58_645 ();
 sg13g2_fill_2 FILLER_58_649 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_fill_2 FILLER_58_711 ();
 sg13g2_fill_1 FILLER_58_713 ();
 sg13g2_fill_2 FILLER_58_720 ();
 sg13g2_decap_8 FILLER_58_732 ();
 sg13g2_decap_8 FILLER_58_739 ();
 sg13g2_fill_2 FILLER_58_746 ();
 sg13g2_fill_2 FILLER_58_775 ();
 sg13g2_fill_1 FILLER_58_796 ();
 sg13g2_fill_1 FILLER_58_818 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_11 ();
 sg13g2_decap_4 FILLER_59_54 ();
 sg13g2_fill_2 FILLER_59_78 ();
 sg13g2_decap_8 FILLER_59_90 ();
 sg13g2_decap_8 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_127 ();
 sg13g2_decap_4 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_4 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_165 ();
 sg13g2_fill_2 FILLER_59_180 ();
 sg13g2_decap_4 FILLER_59_188 ();
 sg13g2_decap_4 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_2 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_254 ();
 sg13g2_decap_4 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_296 ();
 sg13g2_decap_8 FILLER_59_319 ();
 sg13g2_decap_4 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_330 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_420 ();
 sg13g2_decap_8 FILLER_59_449 ();
 sg13g2_fill_2 FILLER_59_456 ();
 sg13g2_fill_1 FILLER_59_458 ();
 sg13g2_decap_8 FILLER_59_476 ();
 sg13g2_fill_2 FILLER_59_483 ();
 sg13g2_fill_1 FILLER_59_485 ();
 sg13g2_decap_4 FILLER_59_499 ();
 sg13g2_fill_1 FILLER_59_503 ();
 sg13g2_fill_1 FILLER_59_517 ();
 sg13g2_decap_4 FILLER_59_522 ();
 sg13g2_decap_8 FILLER_59_579 ();
 sg13g2_fill_2 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_636 ();
 sg13g2_fill_1 FILLER_59_641 ();
 sg13g2_decap_8 FILLER_59_647 ();
 sg13g2_decap_4 FILLER_59_654 ();
 sg13g2_fill_2 FILLER_59_658 ();
 sg13g2_fill_2 FILLER_59_706 ();
 sg13g2_fill_1 FILLER_59_718 ();
 sg13g2_fill_2 FILLER_59_757 ();
 sg13g2_fill_2 FILLER_59_767 ();
 sg13g2_fill_1 FILLER_59_769 ();
 sg13g2_fill_1 FILLER_59_779 ();
 sg13g2_fill_1 FILLER_59_805 ();
 sg13g2_fill_1 FILLER_59_826 ();
 sg13g2_fill_2 FILLER_59_840 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_4 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_82 ();
 sg13g2_decap_8 FILLER_60_87 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_decap_8 FILLER_60_114 ();
 sg13g2_decap_4 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_fill_2 FILLER_60_167 ();
 sg13g2_decap_4 FILLER_60_174 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_4 FILLER_60_203 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_fill_1 FILLER_60_229 ();
 sg13g2_decap_4 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_decap_8 FILLER_60_276 ();
 sg13g2_decap_8 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_326 ();
 sg13g2_fill_2 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_decap_8 FILLER_60_340 ();
 sg13g2_decap_4 FILLER_60_347 ();
 sg13g2_decap_8 FILLER_60_356 ();
 sg13g2_fill_2 FILLER_60_363 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_60_409 ();
 sg13g2_fill_1 FILLER_60_439 ();
 sg13g2_decap_8 FILLER_60_502 ();
 sg13g2_decap_4 FILLER_60_509 ();
 sg13g2_fill_2 FILLER_60_513 ();
 sg13g2_fill_2 FILLER_60_520 ();
 sg13g2_fill_1 FILLER_60_522 ();
 sg13g2_fill_2 FILLER_60_562 ();
 sg13g2_decap_8 FILLER_60_568 ();
 sg13g2_fill_1 FILLER_60_575 ();
 sg13g2_fill_1 FILLER_60_589 ();
 sg13g2_decap_8 FILLER_60_617 ();
 sg13g2_decap_8 FILLER_60_624 ();
 sg13g2_decap_4 FILLER_60_631 ();
 sg13g2_fill_2 FILLER_60_635 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_fill_2 FILLER_60_665 ();
 sg13g2_fill_2 FILLER_60_675 ();
 sg13g2_fill_1 FILLER_60_677 ();
 sg13g2_decap_4 FILLER_60_682 ();
 sg13g2_fill_2 FILLER_60_686 ();
 sg13g2_decap_8 FILLER_60_700 ();
 sg13g2_decap_4 FILLER_60_717 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_726 ();
 sg13g2_decap_4 FILLER_60_737 ();
 sg13g2_fill_1 FILLER_60_741 ();
 sg13g2_decap_8 FILLER_60_746 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_1 FILLER_60_805 ();
 sg13g2_decap_4 FILLER_60_809 ();
 sg13g2_fill_2 FILLER_60_813 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_decap_4 FILLER_61_120 ();
 sg13g2_fill_1 FILLER_61_124 ();
 sg13g2_fill_1 FILLER_61_152 ();
 sg13g2_fill_2 FILLER_61_161 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_decap_4 FILLER_61_170 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_192 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_2 FILLER_61_254 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_decap_4 FILLER_61_300 ();
 sg13g2_fill_2 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_decap_4 FILLER_61_357 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_decap_8 FILLER_61_373 ();
 sg13g2_decap_4 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_430 ();
 sg13g2_fill_2 FILLER_61_439 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_458 ();
 sg13g2_decap_8 FILLER_61_465 ();
 sg13g2_decap_8 FILLER_61_472 ();
 sg13g2_decap_8 FILLER_61_479 ();
 sg13g2_fill_2 FILLER_61_486 ();
 sg13g2_fill_1 FILLER_61_488 ();
 sg13g2_fill_1 FILLER_61_524 ();
 sg13g2_decap_4 FILLER_61_533 ();
 sg13g2_fill_2 FILLER_61_537 ();
 sg13g2_fill_1 FILLER_61_552 ();
 sg13g2_fill_2 FILLER_61_556 ();
 sg13g2_fill_1 FILLER_61_558 ();
 sg13g2_fill_2 FILLER_61_612 ();
 sg13g2_fill_1 FILLER_61_614 ();
 sg13g2_decap_8 FILLER_61_619 ();
 sg13g2_decap_8 FILLER_61_626 ();
 sg13g2_decap_8 FILLER_61_637 ();
 sg13g2_fill_2 FILLER_61_648 ();
 sg13g2_fill_1 FILLER_61_650 ();
 sg13g2_decap_4 FILLER_61_664 ();
 sg13g2_fill_1 FILLER_61_668 ();
 sg13g2_decap_4 FILLER_61_678 ();
 sg13g2_fill_2 FILLER_61_703 ();
 sg13g2_fill_1 FILLER_61_710 ();
 sg13g2_fill_2 FILLER_61_715 ();
 sg13g2_fill_1 FILLER_61_757 ();
 sg13g2_decap_4 FILLER_61_762 ();
 sg13g2_fill_2 FILLER_61_766 ();
 sg13g2_fill_2 FILLER_61_777 ();
 sg13g2_fill_1 FILLER_61_779 ();
 sg13g2_fill_1 FILLER_61_785 ();
 sg13g2_fill_1 FILLER_61_845 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_28 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_decap_8 FILLER_62_87 ();
 sg13g2_decap_8 FILLER_62_94 ();
 sg13g2_decap_4 FILLER_62_101 ();
 sg13g2_decap_4 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_123 ();
 sg13g2_decap_8 FILLER_62_127 ();
 sg13g2_decap_4 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_fill_2 FILLER_62_180 ();
 sg13g2_fill_1 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_195 ();
 sg13g2_fill_2 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_decap_8 FILLER_62_221 ();
 sg13g2_decap_4 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_decap_8 FILLER_62_250 ();
 sg13g2_decap_8 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_264 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_decap_4 FILLER_62_350 ();
 sg13g2_fill_2 FILLER_62_366 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_4 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_392 ();
 sg13g2_decap_4 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_413 ();
 sg13g2_fill_2 FILLER_62_419 ();
 sg13g2_decap_8 FILLER_62_443 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_fill_2 FILLER_62_460 ();
 sg13g2_fill_1 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_484 ();
 sg13g2_decap_4 FILLER_62_491 ();
 sg13g2_fill_1 FILLER_62_500 ();
 sg13g2_fill_1 FILLER_62_514 ();
 sg13g2_decap_4 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_567 ();
 sg13g2_fill_1 FILLER_62_569 ();
 sg13g2_fill_2 FILLER_62_576 ();
 sg13g2_fill_1 FILLER_62_595 ();
 sg13g2_decap_4 FILLER_62_601 ();
 sg13g2_fill_2 FILLER_62_605 ();
 sg13g2_decap_8 FILLER_62_682 ();
 sg13g2_decap_4 FILLER_62_702 ();
 sg13g2_fill_2 FILLER_62_706 ();
 sg13g2_decap_8 FILLER_62_712 ();
 sg13g2_decap_8 FILLER_62_719 ();
 sg13g2_fill_2 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_755 ();
 sg13g2_decap_4 FILLER_62_762 ();
 sg13g2_fill_2 FILLER_62_766 ();
 sg13g2_fill_1 FILLER_62_786 ();
 sg13g2_fill_1 FILLER_62_804 ();
 sg13g2_fill_2 FILLER_62_822 ();
 sg13g2_fill_1 FILLER_62_824 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_2 FILLER_63_45 ();
 sg13g2_decap_8 FILLER_63_60 ();
 sg13g2_decap_8 FILLER_63_67 ();
 sg13g2_fill_2 FILLER_63_94 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_fill_2 FILLER_63_160 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_decap_4 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_220 ();
 sg13g2_decap_4 FILLER_63_227 ();
 sg13g2_decap_4 FILLER_63_254 ();
 sg13g2_decap_8 FILLER_63_271 ();
 sg13g2_decap_8 FILLER_63_278 ();
 sg13g2_decap_8 FILLER_63_285 ();
 sg13g2_decap_8 FILLER_63_292 ();
 sg13g2_decap_8 FILLER_63_299 ();
 sg13g2_decap_4 FILLER_63_306 ();
 sg13g2_fill_2 FILLER_63_310 ();
 sg13g2_decap_8 FILLER_63_341 ();
 sg13g2_decap_4 FILLER_63_370 ();
 sg13g2_decap_4 FILLER_63_423 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_434 ();
 sg13g2_decap_4 FILLER_63_473 ();
 sg13g2_decap_4 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_529 ();
 sg13g2_decap_4 FILLER_63_546 ();
 sg13g2_fill_2 FILLER_63_610 ();
 sg13g2_decap_8 FILLER_63_616 ();
 sg13g2_decap_8 FILLER_63_623 ();
 sg13g2_decap_8 FILLER_63_634 ();
 sg13g2_fill_1 FILLER_63_641 ();
 sg13g2_fill_2 FILLER_63_646 ();
 sg13g2_decap_4 FILLER_63_657 ();
 sg13g2_fill_1 FILLER_63_661 ();
 sg13g2_decap_4 FILLER_63_670 ();
 sg13g2_fill_1 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_710 ();
 sg13g2_decap_4 FILLER_63_740 ();
 sg13g2_fill_1 FILLER_63_744 ();
 sg13g2_decap_8 FILLER_63_755 ();
 sg13g2_fill_2 FILLER_63_815 ();
 sg13g2_fill_2 FILLER_63_827 ();
 sg13g2_fill_2 FILLER_63_843 ();
 sg13g2_fill_1 FILLER_63_845 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_36 ();
 sg13g2_decap_4 FILLER_64_47 ();
 sg13g2_fill_2 FILLER_64_72 ();
 sg13g2_decap_8 FILLER_64_97 ();
 sg13g2_fill_1 FILLER_64_104 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_144 ();
 sg13g2_fill_1 FILLER_64_146 ();
 sg13g2_decap_4 FILLER_64_152 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_decap_4 FILLER_64_161 ();
 sg13g2_fill_2 FILLER_64_165 ();
 sg13g2_decap_8 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_187 ();
 sg13g2_fill_1 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_204 ();
 sg13g2_decap_4 FILLER_64_211 ();
 sg13g2_fill_2 FILLER_64_228 ();
 sg13g2_fill_1 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_282 ();
 sg13g2_decap_4 FILLER_64_293 ();
 sg13g2_fill_2 FILLER_64_297 ();
 sg13g2_decap_8 FILLER_64_304 ();
 sg13g2_decap_8 FILLER_64_311 ();
 sg13g2_decap_4 FILLER_64_318 ();
 sg13g2_decap_8 FILLER_64_332 ();
 sg13g2_decap_8 FILLER_64_339 ();
 sg13g2_decap_4 FILLER_64_346 ();
 sg13g2_decap_4 FILLER_64_387 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_2 FILLER_64_473 ();
 sg13g2_fill_2 FILLER_64_484 ();
 sg13g2_fill_1 FILLER_64_486 ();
 sg13g2_fill_2 FILLER_64_500 ();
 sg13g2_fill_1 FILLER_64_507 ();
 sg13g2_fill_1 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_531 ();
 sg13g2_decap_8 FILLER_64_538 ();
 sg13g2_decap_8 FILLER_64_545 ();
 sg13g2_fill_2 FILLER_64_552 ();
 sg13g2_fill_2 FILLER_64_568 ();
 sg13g2_fill_1 FILLER_64_570 ();
 sg13g2_fill_2 FILLER_64_593 ();
 sg13g2_decap_4 FILLER_64_600 ();
 sg13g2_decap_8 FILLER_64_613 ();
 sg13g2_decap_4 FILLER_64_620 ();
 sg13g2_fill_1 FILLER_64_624 ();
 sg13g2_decap_8 FILLER_64_665 ();
 sg13g2_decap_4 FILLER_64_685 ();
 sg13g2_decap_8 FILLER_64_702 ();
 sg13g2_decap_4 FILLER_64_709 ();
 sg13g2_fill_2 FILLER_64_713 ();
 sg13g2_decap_4 FILLER_64_728 ();
 sg13g2_fill_1 FILLER_64_732 ();
 sg13g2_decap_8 FILLER_64_743 ();
 sg13g2_decap_8 FILLER_64_756 ();
 sg13g2_decap_4 FILLER_64_763 ();
 sg13g2_fill_2 FILLER_64_770 ();
 sg13g2_fill_1 FILLER_64_786 ();
 sg13g2_fill_1 FILLER_64_812 ();
 sg13g2_fill_2 FILLER_64_821 ();
 sg13g2_fill_1 FILLER_65_65 ();
 sg13g2_decap_4 FILLER_65_79 ();
 sg13g2_fill_1 FILLER_65_83 ();
 sg13g2_fill_1 FILLER_65_97 ();
 sg13g2_decap_4 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_127 ();
 sg13g2_fill_2 FILLER_65_148 ();
 sg13g2_fill_1 FILLER_65_150 ();
 sg13g2_fill_1 FILLER_65_182 ();
 sg13g2_decap_4 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_191 ();
 sg13g2_decap_8 FILLER_65_201 ();
 sg13g2_decap_8 FILLER_65_220 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_2 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_236 ();
 sg13g2_decap_4 FILLER_65_254 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_decap_4 FILLER_65_339 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_424 ();
 sg13g2_decap_4 FILLER_65_437 ();
 sg13g2_fill_1 FILLER_65_441 ();
 sg13g2_decap_8 FILLER_65_520 ();
 sg13g2_fill_1 FILLER_65_527 ();
 sg13g2_fill_1 FILLER_65_549 ();
 sg13g2_fill_1 FILLER_65_567 ();
 sg13g2_fill_2 FILLER_65_572 ();
 sg13g2_decap_8 FILLER_65_583 ();
 sg13g2_decap_4 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_642 ();
 sg13g2_decap_8 FILLER_65_664 ();
 sg13g2_decap_8 FILLER_65_671 ();
 sg13g2_decap_8 FILLER_65_678 ();
 sg13g2_fill_1 FILLER_65_705 ();
 sg13g2_fill_2 FILLER_65_711 ();
 sg13g2_fill_2 FILLER_65_717 ();
 sg13g2_fill_1 FILLER_65_747 ();
 sg13g2_fill_2 FILLER_65_754 ();
 sg13g2_fill_1 FILLER_65_810 ();
 sg13g2_fill_1 FILLER_65_820 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_27 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_127 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_decap_8 FILLER_66_162 ();
 sg13g2_decap_4 FILLER_66_169 ();
 sg13g2_fill_2 FILLER_66_178 ();
 sg13g2_decap_8 FILLER_66_184 ();
 sg13g2_fill_1 FILLER_66_191 ();
 sg13g2_decap_8 FILLER_66_205 ();
 sg13g2_fill_2 FILLER_66_217 ();
 sg13g2_fill_2 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_246 ();
 sg13g2_fill_2 FILLER_66_253 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_281 ();
 sg13g2_decap_8 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_300 ();
 sg13g2_fill_1 FILLER_66_302 ();
 sg13g2_decap_8 FILLER_66_332 ();
 sg13g2_decap_4 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_2 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_370 ();
 sg13g2_decap_4 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_66_426 ();
 sg13g2_decap_4 FILLER_66_433 ();
 sg13g2_fill_1 FILLER_66_464 ();
 sg13g2_fill_1 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_503 ();
 sg13g2_decap_4 FILLER_66_510 ();
 sg13g2_decap_4 FILLER_66_554 ();
 sg13g2_fill_1 FILLER_66_558 ();
 sg13g2_fill_1 FILLER_66_572 ();
 sg13g2_decap_4 FILLER_66_578 ();
 sg13g2_fill_1 FILLER_66_582 ();
 sg13g2_decap_4 FILLER_66_587 ();
 sg13g2_decap_4 FILLER_66_605 ();
 sg13g2_fill_2 FILLER_66_618 ();
 sg13g2_decap_8 FILLER_66_624 ();
 sg13g2_fill_1 FILLER_66_631 ();
 sg13g2_decap_8 FILLER_66_683 ();
 sg13g2_fill_2 FILLER_66_690 ();
 sg13g2_fill_1 FILLER_66_692 ();
 sg13g2_decap_8 FILLER_66_710 ();
 sg13g2_fill_2 FILLER_66_798 ();
 sg13g2_fill_1 FILLER_66_800 ();
 sg13g2_fill_1 FILLER_66_828 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_4 ();
 sg13g2_fill_2 FILLER_67_9 ();
 sg13g2_decap_4 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_74 ();
 sg13g2_decap_8 FILLER_67_90 ();
 sg13g2_decap_8 FILLER_67_97 ();
 sg13g2_fill_1 FILLER_67_104 ();
 sg13g2_decap_8 FILLER_67_120 ();
 sg13g2_decap_8 FILLER_67_127 ();
 sg13g2_decap_8 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_145 ();
 sg13g2_decap_4 FILLER_67_156 ();
 sg13g2_fill_2 FILLER_67_160 ();
 sg13g2_decap_8 FILLER_67_183 ();
 sg13g2_decap_8 FILLER_67_190 ();
 sg13g2_fill_2 FILLER_67_217 ();
 sg13g2_fill_1 FILLER_67_219 ();
 sg13g2_decap_8 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_235 ();
 sg13g2_fill_1 FILLER_67_237 ();
 sg13g2_fill_2 FILLER_67_243 ();
 sg13g2_fill_1 FILLER_67_245 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_decap_8 FILLER_67_262 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_fill_2 FILLER_67_316 ();
 sg13g2_fill_1 FILLER_67_318 ();
 sg13g2_decap_4 FILLER_67_344 ();
 sg13g2_fill_1 FILLER_67_348 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_fill_1 FILLER_67_371 ();
 sg13g2_fill_1 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_396 ();
 sg13g2_fill_1 FILLER_67_403 ();
 sg13g2_decap_4 FILLER_67_488 ();
 sg13g2_fill_1 FILLER_67_498 ();
 sg13g2_fill_2 FILLER_67_521 ();
 sg13g2_decap_4 FILLER_67_536 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_fill_2 FILLER_67_574 ();
 sg13g2_fill_1 FILLER_67_576 ();
 sg13g2_fill_2 FILLER_67_604 ();
 sg13g2_fill_1 FILLER_67_606 ();
 sg13g2_fill_2 FILLER_67_634 ();
 sg13g2_fill_1 FILLER_67_636 ();
 sg13g2_decap_8 FILLER_67_653 ();
 sg13g2_decap_8 FILLER_67_660 ();
 sg13g2_decap_4 FILLER_67_667 ();
 sg13g2_fill_2 FILLER_67_689 ();
 sg13g2_fill_1 FILLER_67_691 ();
 sg13g2_fill_1 FILLER_67_705 ();
 sg13g2_fill_2 FILLER_67_712 ();
 sg13g2_fill_1 FILLER_67_714 ();
 sg13g2_decap_4 FILLER_67_719 ();
 sg13g2_fill_1 FILLER_67_723 ();
 sg13g2_decap_8 FILLER_67_743 ();
 sg13g2_decap_4 FILLER_67_750 ();
 sg13g2_decap_4 FILLER_67_779 ();
 sg13g2_decap_8 FILLER_67_796 ();
 sg13g2_fill_2 FILLER_67_803 ();
 sg13g2_fill_1 FILLER_67_805 ();
 sg13g2_fill_1 FILLER_67_833 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_88 ();
 sg13g2_decap_4 FILLER_68_95 ();
 sg13g2_fill_1 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_decap_4 FILLER_68_225 ();
 sg13g2_fill_2 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_271 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_fill_2 FILLER_68_292 ();
 sg13g2_fill_1 FILLER_68_294 ();
 sg13g2_fill_2 FILLER_68_313 ();
 sg13g2_fill_1 FILLER_68_315 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_fill_1 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_344 ();
 sg13g2_fill_1 FILLER_68_351 ();
 sg13g2_fill_1 FILLER_68_357 ();
 sg13g2_fill_2 FILLER_68_363 ();
 sg13g2_fill_1 FILLER_68_426 ();
 sg13g2_fill_2 FILLER_68_436 ();
 sg13g2_fill_2 FILLER_68_470 ();
 sg13g2_fill_2 FILLER_68_584 ();
 sg13g2_decap_8 FILLER_68_592 ();
 sg13g2_decap_8 FILLER_68_599 ();
 sg13g2_decap_8 FILLER_68_610 ();
 sg13g2_decap_8 FILLER_68_617 ();
 sg13g2_decap_8 FILLER_68_624 ();
 sg13g2_fill_2 FILLER_68_631 ();
 sg13g2_fill_1 FILLER_68_633 ();
 sg13g2_decap_4 FILLER_68_647 ();
 sg13g2_fill_1 FILLER_68_651 ();
 sg13g2_fill_1 FILLER_68_665 ();
 sg13g2_decap_4 FILLER_68_670 ();
 sg13g2_fill_2 FILLER_68_695 ();
 sg13g2_fill_2 FILLER_68_702 ();
 sg13g2_decap_4 FILLER_68_718 ();
 sg13g2_fill_2 FILLER_68_756 ();
 sg13g2_fill_2 FILLER_68_771 ();
 sg13g2_fill_2 FILLER_68_813 ();
 sg13g2_fill_1 FILLER_68_833 ();
 sg13g2_fill_2 FILLER_68_843 ();
 sg13g2_fill_1 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_55 ();
 sg13g2_decap_4 FILLER_69_62 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_fill_2 FILLER_69_91 ();
 sg13g2_fill_1 FILLER_69_93 ();
 sg13g2_decap_4 FILLER_69_98 ();
 sg13g2_fill_1 FILLER_69_102 ();
 sg13g2_fill_1 FILLER_69_123 ();
 sg13g2_decap_8 FILLER_69_129 ();
 sg13g2_fill_2 FILLER_69_140 ();
 sg13g2_fill_2 FILLER_69_199 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_2 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_221 ();
 sg13g2_fill_2 FILLER_69_253 ();
 sg13g2_fill_1 FILLER_69_264 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_351 ();
 sg13g2_fill_2 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_436 ();
 sg13g2_fill_2 FILLER_69_443 ();
 sg13g2_fill_1 FILLER_69_445 ();
 sg13g2_decap_4 FILLER_69_456 ();
 sg13g2_fill_1 FILLER_69_460 ();
 sg13g2_fill_2 FILLER_69_465 ();
 sg13g2_fill_1 FILLER_69_467 ();
 sg13g2_fill_2 FILLER_69_499 ();
 sg13g2_fill_2 FILLER_69_510 ();
 sg13g2_decap_4 FILLER_69_562 ();
 sg13g2_fill_1 FILLER_69_566 ();
 sg13g2_fill_1 FILLER_69_600 ();
 sg13g2_fill_1 FILLER_69_628 ();
 sg13g2_decap_8 FILLER_69_642 ();
 sg13g2_fill_2 FILLER_69_649 ();
 sg13g2_fill_1 FILLER_69_663 ();
 sg13g2_fill_2 FILLER_69_684 ();
 sg13g2_fill_2 FILLER_69_696 ();
 sg13g2_decap_8 FILLER_69_726 ();
 sg13g2_fill_1 FILLER_69_733 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_fill_2 FILLER_69_756 ();
 sg13g2_fill_1 FILLER_69_782 ();
 sg13g2_fill_2 FILLER_69_797 ();
 sg13g2_fill_2 FILLER_69_817 ();
 sg13g2_fill_1 FILLER_69_819 ();
 sg13g2_fill_2 FILLER_69_828 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_73 ();
 sg13g2_fill_1 FILLER_70_75 ();
 sg13g2_fill_2 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_87 ();
 sg13g2_decap_8 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_fill_2 FILLER_70_122 ();
 sg13g2_fill_2 FILLER_70_142 ();
 sg13g2_fill_1 FILLER_70_144 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_1 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_219 ();
 sg13g2_decap_4 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_229 ();
 sg13g2_decap_8 FILLER_70_234 ();
 sg13g2_fill_1 FILLER_70_241 ();
 sg13g2_decap_4 FILLER_70_256 ();
 sg13g2_decap_8 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_295 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_327 ();
 sg13g2_fill_1 FILLER_70_329 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_70_478 ();
 sg13g2_fill_2 FILLER_70_489 ();
 sg13g2_fill_1 FILLER_70_491 ();
 sg13g2_fill_2 FILLER_70_501 ();
 sg13g2_fill_1 FILLER_70_503 ();
 sg13g2_decap_4 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_521 ();
 sg13g2_fill_2 FILLER_70_535 ();
 sg13g2_fill_1 FILLER_70_537 ();
 sg13g2_decap_4 FILLER_70_587 ();
 sg13g2_fill_1 FILLER_70_591 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_604 ();
 sg13g2_fill_2 FILLER_70_632 ();
 sg13g2_fill_1 FILLER_70_634 ();
 sg13g2_decap_8 FILLER_70_643 ();
 sg13g2_fill_2 FILLER_70_650 ();
 sg13g2_fill_2 FILLER_70_670 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_fill_2 FILLER_70_695 ();
 sg13g2_fill_1 FILLER_70_697 ();
 sg13g2_fill_2 FILLER_70_713 ();
 sg13g2_fill_1 FILLER_70_715 ();
 sg13g2_fill_1 FILLER_70_725 ();
 sg13g2_decap_4 FILLER_70_772 ();
 sg13g2_fill_2 FILLER_70_789 ();
 sg13g2_fill_1 FILLER_70_836 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_1 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_29 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_fill_2 FILLER_71_59 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_2 FILLER_71_90 ();
 sg13g2_fill_1 FILLER_71_134 ();
 sg13g2_decap_4 FILLER_71_163 ();
 sg13g2_fill_2 FILLER_71_167 ();
 sg13g2_decap_4 FILLER_71_192 ();
 sg13g2_fill_2 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_208 ();
 sg13g2_fill_1 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_decap_4 FILLER_71_267 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_339 ();
 sg13g2_fill_2 FILLER_71_400 ();
 sg13g2_fill_1 FILLER_71_402 ();
 sg13g2_fill_2 FILLER_71_430 ();
 sg13g2_fill_1 FILLER_71_432 ();
 sg13g2_fill_1 FILLER_71_447 ();
 sg13g2_decap_4 FILLER_71_457 ();
 sg13g2_fill_1 FILLER_71_461 ();
 sg13g2_decap_4 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_548 ();
 sg13g2_decap_4 FILLER_71_562 ();
 sg13g2_decap_4 FILLER_71_603 ();
 sg13g2_fill_1 FILLER_71_607 ();
 sg13g2_decap_8 FILLER_71_626 ();
 sg13g2_decap_8 FILLER_71_633 ();
 sg13g2_fill_2 FILLER_71_653 ();
 sg13g2_fill_2 FILLER_71_660 ();
 sg13g2_fill_1 FILLER_71_662 ();
 sg13g2_fill_2 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_679 ();
 sg13g2_fill_2 FILLER_71_689 ();
 sg13g2_fill_2 FILLER_71_732 ();
 sg13g2_fill_1 FILLER_71_734 ();
 sg13g2_fill_1 FILLER_71_747 ();
 sg13g2_fill_1 FILLER_71_784 ();
 sg13g2_fill_2 FILLER_71_832 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_4 ();
 sg13g2_fill_1 FILLER_72_25 ();
 sg13g2_fill_2 FILLER_72_90 ();
 sg13g2_decap_4 FILLER_72_116 ();
 sg13g2_fill_1 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_152 ();
 sg13g2_decap_8 FILLER_72_159 ();
 sg13g2_decap_8 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_248 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_2 FILLER_72_335 ();
 sg13g2_decap_4 FILLER_72_396 ();
 sg13g2_decap_4 FILLER_72_421 ();
 sg13g2_fill_1 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_439 ();
 sg13g2_fill_2 FILLER_72_485 ();
 sg13g2_fill_1 FILLER_72_487 ();
 sg13g2_decap_4 FILLER_72_569 ();
 sg13g2_decap_8 FILLER_72_578 ();
 sg13g2_fill_1 FILLER_72_585 ();
 sg13g2_decap_8 FILLER_72_595 ();
 sg13g2_fill_2 FILLER_72_642 ();
 sg13g2_fill_2 FILLER_72_717 ();
 sg13g2_decap_4 FILLER_72_725 ();
 sg13g2_fill_1 FILLER_72_729 ();
 sg13g2_decap_4 FILLER_72_759 ();
 sg13g2_fill_2 FILLER_72_763 ();
 sg13g2_fill_1 FILLER_72_773 ();
 sg13g2_fill_1 FILLER_72_810 ();
 sg13g2_fill_2 FILLER_72_830 ();
 sg13g2_decap_4 FILLER_72_858 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_4 ();
 sg13g2_fill_1 FILLER_73_24 ();
 sg13g2_fill_2 FILLER_73_39 ();
 sg13g2_decap_4 FILLER_73_123 ();
 sg13g2_decap_4 FILLER_73_160 ();
 sg13g2_fill_1 FILLER_73_172 ();
 sg13g2_decap_4 FILLER_73_197 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_226 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_fill_2 FILLER_73_345 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_368 ();
 sg13g2_decap_4 FILLER_73_378 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_fill_1 FILLER_73_411 ();
 sg13g2_fill_2 FILLER_73_417 ();
 sg13g2_fill_1 FILLER_73_419 ();
 sg13g2_fill_2 FILLER_73_433 ();
 sg13g2_fill_1 FILLER_73_435 ();
 sg13g2_decap_4 FILLER_73_449 ();
 sg13g2_fill_1 FILLER_73_453 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_fill_2 FILLER_73_478 ();
 sg13g2_fill_1 FILLER_73_499 ();
 sg13g2_decap_4 FILLER_73_527 ();
 sg13g2_fill_1 FILLER_73_531 ();
 sg13g2_decap_8 FILLER_73_538 ();
 sg13g2_decap_8 FILLER_73_545 ();
 sg13g2_decap_8 FILLER_73_552 ();
 sg13g2_fill_1 FILLER_73_559 ();
 sg13g2_fill_2 FILLER_73_573 ();
 sg13g2_fill_1 FILLER_73_575 ();
 sg13g2_fill_1 FILLER_73_590 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_fill_2 FILLER_73_647 ();
 sg13g2_fill_1 FILLER_73_649 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_fill_1 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_732 ();
 sg13g2_fill_1 FILLER_73_758 ();
 sg13g2_fill_1 FILLER_73_795 ();
 sg13g2_fill_1 FILLER_73_805 ();
 sg13g2_fill_1 FILLER_73_816 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_85 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_1 FILLER_74_102 ();
 sg13g2_fill_2 FILLER_74_126 ();
 sg13g2_fill_1 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_138 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_fill_1 FILLER_74_199 ();
 sg13g2_fill_2 FILLER_74_254 ();
 sg13g2_fill_2 FILLER_74_265 ();
 sg13g2_fill_1 FILLER_74_267 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_2 FILLER_74_290 ();
 sg13g2_fill_1 FILLER_74_292 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_8 FILLER_74_403 ();
 sg13g2_fill_1 FILLER_74_410 ();
 sg13g2_decap_4 FILLER_74_428 ();
 sg13g2_fill_1 FILLER_74_432 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_fill_2 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_511 ();
 sg13g2_decap_4 FILLER_74_527 ();
 sg13g2_fill_2 FILLER_74_531 ();
 sg13g2_fill_1 FILLER_74_589 ();
 sg13g2_fill_2 FILLER_74_594 ();
 sg13g2_fill_1 FILLER_74_639 ();
 sg13g2_fill_1 FILLER_74_650 ();
 sg13g2_fill_1 FILLER_74_664 ();
 sg13g2_fill_1 FILLER_74_725 ();
 sg13g2_decap_8 FILLER_74_736 ();
 sg13g2_decap_4 FILLER_74_753 ();
 sg13g2_fill_2 FILLER_74_757 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_fill_2 FILLER_74_784 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_decap_4 FILLER_74_834 ();
 sg13g2_fill_2 FILLER_74_838 ();
 sg13g2_fill_2 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_855 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_60 ();
 sg13g2_decap_4 FILLER_75_117 ();
 sg13g2_fill_1 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_149 ();
 sg13g2_fill_1 FILLER_75_151 ();
 sg13g2_fill_2 FILLER_75_209 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_fill_1 FILLER_75_310 ();
 sg13g2_fill_2 FILLER_75_325 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_2 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_370 ();
 sg13g2_fill_1 FILLER_75_372 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_500 ();
 sg13g2_decap_4 FILLER_75_512 ();
 sg13g2_decap_8 FILLER_75_521 ();
 sg13g2_fill_1 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_548 ();
 sg13g2_fill_2 FILLER_75_556 ();
 sg13g2_fill_1 FILLER_75_567 ();
 sg13g2_decap_8 FILLER_75_578 ();
 sg13g2_decap_4 FILLER_75_658 ();
 sg13g2_fill_1 FILLER_75_662 ();
 sg13g2_fill_2 FILLER_75_676 ();
 sg13g2_fill_1 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_701 ();
 sg13g2_fill_1 FILLER_75_708 ();
 sg13g2_decap_4 FILLER_75_713 ();
 sg13g2_fill_2 FILLER_75_717 ();
 sg13g2_decap_4 FILLER_75_747 ();
 sg13g2_fill_1 FILLER_75_751 ();
 sg13g2_fill_1 FILLER_75_780 ();
 sg13g2_fill_2 FILLER_75_821 ();
 sg13g2_fill_1 FILLER_75_823 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_9 ();
 sg13g2_fill_2 FILLER_76_32 ();
 sg13g2_fill_1 FILLER_76_34 ();
 sg13g2_fill_1 FILLER_76_116 ();
 sg13g2_fill_2 FILLER_76_121 ();
 sg13g2_fill_1 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_168 ();
 sg13g2_fill_1 FILLER_76_196 ();
 sg13g2_fill_2 FILLER_76_335 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_fill_2 FILLER_76_369 ();
 sg13g2_fill_1 FILLER_76_392 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_fill_1 FILLER_76_410 ();
 sg13g2_fill_2 FILLER_76_422 ();
 sg13g2_decap_4 FILLER_76_438 ();
 sg13g2_decap_4 FILLER_76_448 ();
 sg13g2_fill_1 FILLER_76_452 ();
 sg13g2_fill_2 FILLER_76_458 ();
 sg13g2_fill_1 FILLER_76_460 ();
 sg13g2_fill_1 FILLER_76_502 ();
 sg13g2_fill_1 FILLER_76_517 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_fill_2 FILLER_76_531 ();
 sg13g2_fill_1 FILLER_76_533 ();
 sg13g2_decap_8 FILLER_76_555 ();
 sg13g2_fill_2 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_fill_1 FILLER_76_628 ();
 sg13g2_decap_4 FILLER_76_669 ();
 sg13g2_fill_1 FILLER_76_673 ();
 sg13g2_decap_4 FILLER_76_687 ();
 sg13g2_fill_1 FILLER_76_691 ();
 sg13g2_fill_2 FILLER_76_739 ();
 sg13g2_fill_1 FILLER_76_741 ();
 sg13g2_fill_1 FILLER_76_752 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_845 ();
 sg13g2_decap_8 FILLER_76_852 ();
 sg13g2_fill_2 FILLER_76_859 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_93 ();
 sg13g2_fill_2 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_163 ();
 sg13g2_fill_1 FILLER_77_200 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_322 ();
 sg13g2_fill_2 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_355 ();
 sg13g2_fill_2 FILLER_77_365 ();
 sg13g2_decap_4 FILLER_77_386 ();
 sg13g2_fill_2 FILLER_77_418 ();
 sg13g2_fill_1 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_435 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_fill_1 FILLER_77_469 ();
 sg13g2_fill_1 FILLER_77_496 ();
 sg13g2_fill_1 FILLER_77_506 ();
 sg13g2_fill_1 FILLER_77_524 ();
 sg13g2_fill_2 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_568 ();
 sg13g2_fill_2 FILLER_77_575 ();
 sg13g2_fill_1 FILLER_77_605 ();
 sg13g2_decap_8 FILLER_77_636 ();
 sg13g2_fill_2 FILLER_77_643 ();
 sg13g2_fill_1 FILLER_77_645 ();
 sg13g2_fill_2 FILLER_77_655 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_fill_1 FILLER_77_701 ();
 sg13g2_decap_4 FILLER_77_730 ();
 sg13g2_fill_1 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_754 ();
 sg13g2_fill_2 FILLER_77_761 ();
 sg13g2_decap_8 FILLER_77_772 ();
 sg13g2_fill_2 FILLER_77_792 ();
 sg13g2_decap_4 FILLER_77_798 ();
 sg13g2_fill_2 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_807 ();
 sg13g2_decap_4 FILLER_77_814 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_decap_4 FILLER_77_824 ();
 sg13g2_fill_1 FILLER_77_828 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_fill_2 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_258 ();
 sg13g2_fill_2 FILLER_78_265 ();
 sg13g2_fill_1 FILLER_78_289 ();
 sg13g2_fill_2 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_366 ();
 sg13g2_fill_1 FILLER_78_387 ();
 sg13g2_fill_1 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_436 ();
 sg13g2_decap_4 FILLER_78_475 ();
 sg13g2_fill_2 FILLER_78_492 ();
 sg13g2_fill_1 FILLER_78_494 ();
 sg13g2_fill_1 FILLER_78_528 ();
 sg13g2_fill_1 FILLER_78_547 ();
 sg13g2_fill_1 FILLER_78_593 ();
 sg13g2_fill_1 FILLER_78_691 ();
 sg13g2_fill_2 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_722 ();
 sg13g2_decap_8 FILLER_78_729 ();
 sg13g2_decap_4 FILLER_78_736 ();
 sg13g2_fill_1 FILLER_78_740 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_decap_8 FILLER_78_776 ();
 sg13g2_decap_8 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_790 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_decap_8 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_8 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_100 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_127 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_fill_1 FILLER_79_366 ();
 sg13g2_fill_2 FILLER_79_379 ();
 sg13g2_fill_1 FILLER_79_381 ();
 sg13g2_decap_4 FILLER_79_428 ();
 sg13g2_fill_2 FILLER_79_432 ();
 sg13g2_decap_4 FILLER_79_467 ();
 sg13g2_fill_2 FILLER_79_471 ();
 sg13g2_decap_4 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_495 ();
 sg13g2_decap_4 FILLER_79_510 ();
 sg13g2_fill_1 FILLER_79_533 ();
 sg13g2_fill_1 FILLER_79_538 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_4 FILLER_79_594 ();
 sg13g2_fill_1 FILLER_79_598 ();
 sg13g2_fill_2 FILLER_79_625 ();
 sg13g2_fill_1 FILLER_79_627 ();
 sg13g2_decap_4 FILLER_79_637 ();
 sg13g2_decap_8 FILLER_79_677 ();
 sg13g2_decap_8 FILLER_79_684 ();
 sg13g2_decap_8 FILLER_79_691 ();
 sg13g2_decap_8 FILLER_79_698 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_fill_1 FILLER_79_712 ();
 sg13g2_decap_8 FILLER_79_722 ();
 sg13g2_decap_8 FILLER_79_729 ();
 sg13g2_decap_4 FILLER_79_736 ();
 sg13g2_fill_1 FILLER_79_740 ();
 sg13g2_decap_4 FILLER_79_750 ();
 sg13g2_fill_2 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_4 FILLER_79_856 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_43 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_216 ();
 sg13g2_fill_2 FILLER_80_223 ();
 sg13g2_fill_1 FILLER_80_225 ();
 sg13g2_fill_1 FILLER_80_241 ();
 sg13g2_fill_1 FILLER_80_251 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_272 ();
 sg13g2_fill_1 FILLER_80_294 ();
 sg13g2_fill_2 FILLER_80_350 ();
 sg13g2_fill_1 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_4 FILLER_80_415 ();
 sg13g2_fill_2 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_fill_2 FILLER_80_456 ();
 sg13g2_fill_1 FILLER_80_458 ();
 sg13g2_decap_4 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_fill_2 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule
